`timescale 1ns/1ps
module add(
    input  [15:0] a,
    input  [15:0] b,
    output  [15:0] o
);
    wire [15:0] x,y,sum;

    assign x=(a[15]==1)?(((a[14:0])==15'b0)?{16'b00000000}:{1'b1,~a[14:0]+1'b1}):({a[15:0]});
    assign y=(b[15]==1)?(((b[14:0])==15'b0)?{16'b00000000}:{1'b1,~b[14:0]+1'b1}):({b[15:0]});//当输入是10000000时转换为00000000参与计算

    assign sum = x + y;

    assign o = (x[15] & y[15])?  {1'b1,~sum[14:0]+1'b1}: //两个负数
                    ( (x[15] || y[15])?(sum[15]?{1'b1,~sum[14:0]+1'b1}:{1'b0,sum[14:0]}): //�?正一�? 
						{1'b0,sum[14:0]} );	// （两个正数）  	

endmodule 
