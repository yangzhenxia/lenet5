# Confidential Information of ARM, Inc.
# Use subject to ARM license.
# Copyright (c) 2022 ARM, Inc.

# ACI Version r1p1

# Reifier 4.0.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;

#name: High Density Single Port Register File RVT RVT Compiler | LOGIC0040LL 40nm Process 0.299um^2 Bit Cell
#version: r1p1
#comment: This is a memory instance
#configuration:  -activity_factor 50 -back_biasing off -bits 144 -bmux off -bus_notation on -check_instname on -diodes on -drive 6 -ema on -frequency 200 -instname sram464x144 -left_bus_delim "[" -mux 2 -mvt "" -name_case upper -power_type otc -prefix "" -pwr_gnd_rename vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -retention on -right_bus_delim "]" -ser none -site_def off -top_layer m5-m10 -words 464 -write_mask off -write_thru off -corners ss_0p99v_0p99v_125c,tt_1p10v_1p10v_125c
MACRO sram464x144
  FOREIGN sram464x144 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 268.38 BY 100.88 ;
  CLASS BLOCK ;
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 134.135 0.0 134.275 0.25 ;
      LAYER M2 ;
      RECT 134.135 0.0 134.275 0.25 ;
      LAYER M3 ;
      RECT 134.135 0.0 134.275 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[5]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.53 0.0 132.67 0.25 ;
      LAYER M2 ;
      RECT 132.53 0.0 132.67 0.25 ;
      LAYER M1 ;
      RECT 132.53 0.0 132.67 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END WEN
  PIN EMA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 136.49 0.0 136.63 0.25 ;
      LAYER M2 ;
      RECT 136.49 0.0 136.63 0.25 ;
      LAYER M3 ;
      RECT 136.49 0.0 136.63 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMA[0]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.11 0.0 132.25 0.25 ;
      LAYER M2 ;
      RECT 132.11 0.0 132.25 0.25 ;
      LAYER M1 ;
      RECT 132.11 0.0 132.25 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[4]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 137.29 0.0 137.43 0.25 ;
      LAYER M2 ;
      RECT 137.29 0.0 137.43 0.25 ;
      LAYER M3 ;
      RECT 137.29 0.0 137.43 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[8]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 128.71 0.0 128.85 0.25 ;
      LAYER M2 ;
      RECT 128.71 0.0 128.85 0.25 ;
      LAYER M1 ;
      RECT 128.71 0.0 128.85 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[1]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 137.57 0.0 137.71 0.25 ;
      LAYER M2 ;
      RECT 137.57 0.0 137.71 0.25 ;
      LAYER M3 ;
      RECT 137.57 0.0 137.71 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[7]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 128.43 0.0 128.57 0.25 ;
      LAYER M2 ;
      RECT 128.43 0.0 128.57 0.25 ;
      LAYER M1 ;
      RECT 128.43 0.0 128.57 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[2]
  PIN EMA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 138.14 0.0 138.28 0.25 ;
      LAYER M2 ;
      RECT 138.14 0.0 138.28 0.25 ;
      LAYER M3 ;
      RECT 138.14 0.0 138.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMA[1]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 126.42 0.0 126.56 0.25 ;
      LAYER M2 ;
      RECT 126.42 0.0 126.56 0.25 ;
      LAYER M1 ;
      RECT 126.42 0.0 126.56 0.25 ;
      LAYER M4 ;
      RECT 126.38 0.0 126.59 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CLK
  PIN EMA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 138.535 0.0 138.675 0.25 ;
      LAYER M2 ;
      RECT 138.535 0.0 138.675 0.25 ;
      LAYER M3 ;
      RECT 138.535 0.0 138.675 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMA[2]
  PIN EMAW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 125.445 0.0 125.585 0.25 ;
      LAYER M2 ;
      RECT 125.445 0.0 125.585 0.25 ;
      LAYER M1 ;
      RECT 125.445 0.0 125.585 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAW[1]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 140.685 0.0 140.825 0.25 ;
      LAYER M2 ;
      RECT 140.685 0.0 140.825 0.25 ;
      LAYER M3 ;
      RECT 140.685 0.0 140.825 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[3]
  PIN EMAW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.63 0.0 124.77 0.25 ;
      LAYER M2 ;
      RECT 124.63 0.0 124.77 0.25 ;
      LAYER M1 ;
      RECT 124.63 0.0 124.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAW[0]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 140.97 0.0 141.11 0.25 ;
      LAYER M2 ;
      RECT 140.97 0.0 141.11 0.25 ;
      LAYER M3 ;
      RECT 140.97 0.0 141.11 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[6]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 121.355 0.0 121.495 0.25 ;
      LAYER M2 ;
      RECT 121.355 0.0 121.495 0.25 ;
      LAYER M1 ;
      RECT 121.355 0.0 121.495 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CEN
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 147.52 0.0 147.66 0.25 ;
      LAYER M2 ;
      RECT 147.52 0.0 147.66 0.25 ;
      LAYER M3 ;
      RECT 147.52 0.0 147.66 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[0]
  PIN RET1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 120.71 0.0 120.85 0.25 ;
      LAYER M2 ;
      RECT 120.71 0.0 120.85 0.25 ;
      LAYER M1 ;
      RECT 120.71 0.0 120.85 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END RET1N
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 148.58 0.0 148.72 0.25 ;
      LAYER M2 ;
      RECT 148.58 0.0 148.72 0.25 ;
      LAYER M3 ;
      RECT 148.58 0.0 148.72 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.66 0.0 119.8 0.25 ;
      LAYER M2 ;
      RECT 119.66 0.0 119.8 0.25 ;
      LAYER M1 ;
      RECT 119.66 0.0 119.8 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[71]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 149.42 0.0 149.56 0.25 ;
      LAYER M2 ;
      RECT 149.42 0.0 149.56 0.25 ;
      LAYER M3 ;
      RECT 149.42 0.0 149.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.82 0.0 118.96 0.25 ;
      LAYER M2 ;
      RECT 118.82 0.0 118.96 0.25 ;
      LAYER M1 ;
      RECT 118.82 0.0 118.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[71]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 149.7 0.0 149.84 0.25 ;
      LAYER M2 ;
      RECT 149.7 0.0 149.84 0.25 ;
      LAYER M3 ;
      RECT 149.7 0.0 149.84 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[73]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.54 0.0 118.68 0.25 ;
      LAYER M2 ;
      RECT 118.54 0.0 118.68 0.25 ;
      LAYER M1 ;
      RECT 118.54 0.0 118.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[70]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 150.47 0.0 150.61 0.25 ;
      LAYER M2 ;
      RECT 150.47 0.0 150.61 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[73]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 117.77 0.0 117.91 0.25 ;
      LAYER M1 ;
      RECT 117.77 0.0 117.91 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[70]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 151.9 0.0 152.04 0.25 ;
      LAYER M2 ;
      RECT 151.9 0.0 152.04 0.25 ;
      LAYER M3 ;
      RECT 151.9 0.0 152.04 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[74]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 116.34 0.0 116.48 0.25 ;
      LAYER M2 ;
      RECT 116.34 0.0 116.48 0.25 ;
      LAYER M1 ;
      RECT 116.34 0.0 116.48 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[69]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 152.74 0.0 152.88 0.25 ;
      LAYER M2 ;
      RECT 152.74 0.0 152.88 0.25 ;
      LAYER M3 ;
      RECT 152.74 0.0 152.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[74]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 115.5 0.0 115.64 0.25 ;
      LAYER M2 ;
      RECT 115.5 0.0 115.64 0.25 ;
      LAYER M1 ;
      RECT 115.5 0.0 115.64 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[69]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 153.02 0.0 153.16 0.25 ;
      LAYER M2 ;
      RECT 153.02 0.0 153.16 0.25 ;
      LAYER M3 ;
      RECT 153.02 0.0 153.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[75]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 115.22 0.0 115.36 0.25 ;
      LAYER M2 ;
      RECT 115.22 0.0 115.36 0.25 ;
      LAYER M1 ;
      RECT 115.22 0.0 115.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[68]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 153.79 0.0 153.93 0.25 ;
      LAYER M2 ;
      RECT 153.79 0.0 153.93 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[75]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 114.45 0.0 114.59 0.25 ;
      LAYER M1 ;
      RECT 114.45 0.0 114.59 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[68]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 155.22 0.0 155.36 0.25 ;
      LAYER M2 ;
      RECT 155.22 0.0 155.36 0.25 ;
      LAYER M3 ;
      RECT 155.22 0.0 155.36 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[76]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 113.02 0.0 113.16 0.25 ;
      LAYER M2 ;
      RECT 113.02 0.0 113.16 0.25 ;
      LAYER M1 ;
      RECT 113.02 0.0 113.16 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[67]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 156.06 0.0 156.2 0.25 ;
      LAYER M2 ;
      RECT 156.06 0.0 156.2 0.25 ;
      LAYER M3 ;
      RECT 156.06 0.0 156.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[76]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.18 0.0 112.32 0.25 ;
      LAYER M2 ;
      RECT 112.18 0.0 112.32 0.25 ;
      LAYER M1 ;
      RECT 112.18 0.0 112.32 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[67]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 156.34 0.0 156.48 0.25 ;
      LAYER M2 ;
      RECT 156.34 0.0 156.48 0.25 ;
      LAYER M3 ;
      RECT 156.34 0.0 156.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[77]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 111.9 0.0 112.04 0.25 ;
      LAYER M2 ;
      RECT 111.9 0.0 112.04 0.25 ;
      LAYER M1 ;
      RECT 111.9 0.0 112.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[66]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 157.11 0.0 157.25 0.25 ;
      LAYER M2 ;
      RECT 157.11 0.0 157.25 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[77]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 111.13 0.0 111.27 0.25 ;
      LAYER M1 ;
      RECT 111.13 0.0 111.27 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[66]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 158.54 0.0 158.68 0.25 ;
      LAYER M2 ;
      RECT 158.54 0.0 158.68 0.25 ;
      LAYER M3 ;
      RECT 158.54 0.0 158.68 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[78]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 109.7 0.0 109.84 0.25 ;
      LAYER M2 ;
      RECT 109.7 0.0 109.84 0.25 ;
      LAYER M1 ;
      RECT 109.7 0.0 109.84 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[65]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 159.38 0.0 159.52 0.25 ;
      LAYER M2 ;
      RECT 159.38 0.0 159.52 0.25 ;
      LAYER M3 ;
      RECT 159.38 0.0 159.52 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[78]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 108.86 0.0 109.0 0.25 ;
      LAYER M2 ;
      RECT 108.86 0.0 109.0 0.25 ;
      LAYER M1 ;
      RECT 108.86 0.0 109.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[65]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 159.66 0.0 159.8 0.25 ;
      LAYER M2 ;
      RECT 159.66 0.0 159.8 0.25 ;
      LAYER M3 ;
      RECT 159.66 0.0 159.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[79]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 108.58 0.0 108.72 0.25 ;
      LAYER M2 ;
      RECT 108.58 0.0 108.72 0.25 ;
      LAYER M1 ;
      RECT 108.58 0.0 108.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[64]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 160.43 0.0 160.57 0.25 ;
      LAYER M2 ;
      RECT 160.43 0.0 160.57 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[79]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 107.81 0.0 107.95 0.25 ;
      LAYER M1 ;
      RECT 107.81 0.0 107.95 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[64]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 161.86 0.0 162.0 0.25 ;
      LAYER M2 ;
      RECT 161.86 0.0 162.0 0.25 ;
      LAYER M3 ;
      RECT 161.86 0.0 162.0 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[80]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.38 0.0 106.52 0.25 ;
      LAYER M2 ;
      RECT 106.38 0.0 106.52 0.25 ;
      LAYER M1 ;
      RECT 106.38 0.0 106.52 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[63]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 162.7 0.0 162.84 0.25 ;
      LAYER M2 ;
      RECT 162.7 0.0 162.84 0.25 ;
      LAYER M3 ;
      RECT 162.7 0.0 162.84 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[80]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.54 0.0 105.68 0.25 ;
      LAYER M2 ;
      RECT 105.54 0.0 105.68 0.25 ;
      LAYER M1 ;
      RECT 105.54 0.0 105.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[63]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 162.98 0.0 163.12 0.25 ;
      LAYER M2 ;
      RECT 162.98 0.0 163.12 0.25 ;
      LAYER M3 ;
      RECT 162.98 0.0 163.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[81]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.26 0.0 105.4 0.25 ;
      LAYER M2 ;
      RECT 105.26 0.0 105.4 0.25 ;
      LAYER M1 ;
      RECT 105.26 0.0 105.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[62]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 163.75 0.0 163.89 0.25 ;
      LAYER M2 ;
      RECT 163.75 0.0 163.89 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[81]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 104.49 0.0 104.63 0.25 ;
      LAYER M1 ;
      RECT 104.49 0.0 104.63 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[62]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 165.18 0.0 165.32 0.25 ;
      LAYER M2 ;
      RECT 165.18 0.0 165.32 0.25 ;
      LAYER M3 ;
      RECT 165.18 0.0 165.32 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[82]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 103.06 0.0 103.2 0.25 ;
      LAYER M2 ;
      RECT 103.06 0.0 103.2 0.25 ;
      LAYER M1 ;
      RECT 103.06 0.0 103.2 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[61]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 166.02 0.0 166.16 0.25 ;
      LAYER M2 ;
      RECT 166.02 0.0 166.16 0.25 ;
      LAYER M3 ;
      RECT 166.02 0.0 166.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[82]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 102.22 0.0 102.36 0.25 ;
      LAYER M2 ;
      RECT 102.22 0.0 102.36 0.25 ;
      LAYER M1 ;
      RECT 102.22 0.0 102.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[61]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 166.3 0.0 166.44 0.25 ;
      LAYER M2 ;
      RECT 166.3 0.0 166.44 0.25 ;
      LAYER M3 ;
      RECT 166.3 0.0 166.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[83]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 101.94 0.0 102.08 0.25 ;
      LAYER M2 ;
      RECT 101.94 0.0 102.08 0.25 ;
      LAYER M1 ;
      RECT 101.94 0.0 102.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[60]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 167.07 0.0 167.21 0.25 ;
      LAYER M2 ;
      RECT 167.07 0.0 167.21 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[83]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 101.17 0.0 101.31 0.25 ;
      LAYER M1 ;
      RECT 101.17 0.0 101.31 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[60]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 168.5 0.0 168.64 0.25 ;
      LAYER M2 ;
      RECT 168.5 0.0 168.64 0.25 ;
      LAYER M3 ;
      RECT 168.5 0.0 168.64 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[84]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 99.74 0.0 99.88 0.25 ;
      LAYER M2 ;
      RECT 99.74 0.0 99.88 0.25 ;
      LAYER M1 ;
      RECT 99.74 0.0 99.88 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[59]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 169.34 0.0 169.48 0.25 ;
      LAYER M2 ;
      RECT 169.34 0.0 169.48 0.25 ;
      LAYER M3 ;
      RECT 169.34 0.0 169.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[84]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.9 0.0 99.04 0.25 ;
      LAYER M2 ;
      RECT 98.9 0.0 99.04 0.25 ;
      LAYER M1 ;
      RECT 98.9 0.0 99.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[59]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 169.62 0.0 169.76 0.25 ;
      LAYER M2 ;
      RECT 169.62 0.0 169.76 0.25 ;
      LAYER M3 ;
      RECT 169.62 0.0 169.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[85]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.62 0.0 98.76 0.25 ;
      LAYER M2 ;
      RECT 98.62 0.0 98.76 0.25 ;
      LAYER M1 ;
      RECT 98.62 0.0 98.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[58]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 170.39 0.0 170.53 0.25 ;
      LAYER M2 ;
      RECT 170.39 0.0 170.53 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[85]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 97.85 0.0 97.99 0.25 ;
      LAYER M1 ;
      RECT 97.85 0.0 97.99 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[58]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 171.82 0.0 171.96 0.25 ;
      LAYER M2 ;
      RECT 171.82 0.0 171.96 0.25 ;
      LAYER M3 ;
      RECT 171.82 0.0 171.96 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[86]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 96.42 0.0 96.56 0.25 ;
      LAYER M2 ;
      RECT 96.42 0.0 96.56 0.25 ;
      LAYER M1 ;
      RECT 96.42 0.0 96.56 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[57]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 172.66 0.0 172.8 0.25 ;
      LAYER M2 ;
      RECT 172.66 0.0 172.8 0.25 ;
      LAYER M3 ;
      RECT 172.66 0.0 172.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[86]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 95.58 0.0 95.72 0.25 ;
      LAYER M2 ;
      RECT 95.58 0.0 95.72 0.25 ;
      LAYER M1 ;
      RECT 95.58 0.0 95.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[57]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 172.94 0.0 173.08 0.25 ;
      LAYER M2 ;
      RECT 172.94 0.0 173.08 0.25 ;
      LAYER M3 ;
      RECT 172.94 0.0 173.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[87]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 95.3 0.0 95.44 0.25 ;
      LAYER M2 ;
      RECT 95.3 0.0 95.44 0.25 ;
      LAYER M1 ;
      RECT 95.3 0.0 95.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[56]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 173.71 0.0 173.85 0.25 ;
      LAYER M2 ;
      RECT 173.71 0.0 173.85 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[87]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 94.53 0.0 94.67 0.25 ;
      LAYER M1 ;
      RECT 94.53 0.0 94.67 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[56]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 175.14 0.0 175.28 0.25 ;
      LAYER M2 ;
      RECT 175.14 0.0 175.28 0.25 ;
      LAYER M3 ;
      RECT 175.14 0.0 175.28 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[88]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.1 0.0 93.24 0.25 ;
      LAYER M2 ;
      RECT 93.1 0.0 93.24 0.25 ;
      LAYER M1 ;
      RECT 93.1 0.0 93.24 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[55]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 175.98 0.0 176.12 0.25 ;
      LAYER M2 ;
      RECT 175.98 0.0 176.12 0.25 ;
      LAYER M3 ;
      RECT 175.98 0.0 176.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[88]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 92.26 0.0 92.4 0.25 ;
      LAYER M2 ;
      RECT 92.26 0.0 92.4 0.25 ;
      LAYER M1 ;
      RECT 92.26 0.0 92.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[55]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 176.26 0.0 176.4 0.25 ;
      LAYER M2 ;
      RECT 176.26 0.0 176.4 0.25 ;
      LAYER M3 ;
      RECT 176.26 0.0 176.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[89]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 91.98 0.0 92.12 0.25 ;
      LAYER M2 ;
      RECT 91.98 0.0 92.12 0.25 ;
      LAYER M1 ;
      RECT 91.98 0.0 92.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[54]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 177.03 0.0 177.17 0.25 ;
      LAYER M2 ;
      RECT 177.03 0.0 177.17 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[89]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 91.21 0.0 91.35 0.25 ;
      LAYER M1 ;
      RECT 91.21 0.0 91.35 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[54]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 178.46 0.0 178.6 0.25 ;
      LAYER M2 ;
      RECT 178.46 0.0 178.6 0.25 ;
      LAYER M3 ;
      RECT 178.46 0.0 178.6 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[90]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 89.78 0.0 89.92 0.25 ;
      LAYER M2 ;
      RECT 89.78 0.0 89.92 0.25 ;
      LAYER M1 ;
      RECT 89.78 0.0 89.92 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[53]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 179.3 0.0 179.44 0.25 ;
      LAYER M2 ;
      RECT 179.3 0.0 179.44 0.25 ;
      LAYER M3 ;
      RECT 179.3 0.0 179.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[90]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.94 0.0 89.08 0.25 ;
      LAYER M2 ;
      RECT 88.94 0.0 89.08 0.25 ;
      LAYER M1 ;
      RECT 88.94 0.0 89.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[53]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 179.58 0.0 179.72 0.25 ;
      LAYER M2 ;
      RECT 179.58 0.0 179.72 0.25 ;
      LAYER M3 ;
      RECT 179.58 0.0 179.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[91]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.66 0.0 88.8 0.25 ;
      LAYER M2 ;
      RECT 88.66 0.0 88.8 0.25 ;
      LAYER M1 ;
      RECT 88.66 0.0 88.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[52]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 180.35 0.0 180.49 0.25 ;
      LAYER M2 ;
      RECT 180.35 0.0 180.49 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[91]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 87.89 0.0 88.03 0.25 ;
      LAYER M1 ;
      RECT 87.89 0.0 88.03 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[52]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 181.78 0.0 181.92 0.25 ;
      LAYER M2 ;
      RECT 181.78 0.0 181.92 0.25 ;
      LAYER M3 ;
      RECT 181.78 0.0 181.92 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[92]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 86.46 0.0 86.6 0.25 ;
      LAYER M2 ;
      RECT 86.46 0.0 86.6 0.25 ;
      LAYER M1 ;
      RECT 86.46 0.0 86.6 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[51]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 182.62 0.0 182.76 0.25 ;
      LAYER M2 ;
      RECT 182.62 0.0 182.76 0.25 ;
      LAYER M3 ;
      RECT 182.62 0.0 182.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[92]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 85.62 0.0 85.76 0.25 ;
      LAYER M2 ;
      RECT 85.62 0.0 85.76 0.25 ;
      LAYER M1 ;
      RECT 85.62 0.0 85.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[51]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 182.9 0.0 183.04 0.25 ;
      LAYER M2 ;
      RECT 182.9 0.0 183.04 0.25 ;
      LAYER M3 ;
      RECT 182.9 0.0 183.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[93]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 85.34 0.0 85.48 0.25 ;
      LAYER M2 ;
      RECT 85.34 0.0 85.48 0.25 ;
      LAYER M1 ;
      RECT 85.34 0.0 85.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[50]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 183.67 0.0 183.81 0.25 ;
      LAYER M2 ;
      RECT 183.67 0.0 183.81 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[93]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 84.57 0.0 84.71 0.25 ;
      LAYER M1 ;
      RECT 84.57 0.0 84.71 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[50]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 185.1 0.0 185.24 0.25 ;
      LAYER M2 ;
      RECT 185.1 0.0 185.24 0.25 ;
      LAYER M3 ;
      RECT 185.1 0.0 185.24 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[94]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 83.14 0.0 83.28 0.25 ;
      LAYER M2 ;
      RECT 83.14 0.0 83.28 0.25 ;
      LAYER M1 ;
      RECT 83.14 0.0 83.28 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[49]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 185.94 0.0 186.08 0.25 ;
      LAYER M2 ;
      RECT 185.94 0.0 186.08 0.25 ;
      LAYER M3 ;
      RECT 185.94 0.0 186.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[94]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 82.3 0.0 82.44 0.25 ;
      LAYER M2 ;
      RECT 82.3 0.0 82.44 0.25 ;
      LAYER M1 ;
      RECT 82.3 0.0 82.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[49]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 186.22 0.0 186.36 0.25 ;
      LAYER M2 ;
      RECT 186.22 0.0 186.36 0.25 ;
      LAYER M3 ;
      RECT 186.22 0.0 186.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[95]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 82.02 0.0 82.16 0.25 ;
      LAYER M2 ;
      RECT 82.02 0.0 82.16 0.25 ;
      LAYER M1 ;
      RECT 82.02 0.0 82.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[48]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 186.99 0.0 187.13 0.25 ;
      LAYER M2 ;
      RECT 186.99 0.0 187.13 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[95]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 81.25 0.0 81.39 0.25 ;
      LAYER M1 ;
      RECT 81.25 0.0 81.39 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[48]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 188.42 0.0 188.56 0.25 ;
      LAYER M2 ;
      RECT 188.42 0.0 188.56 0.25 ;
      LAYER M3 ;
      RECT 188.42 0.0 188.56 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[96]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 79.82 0.0 79.96 0.25 ;
      LAYER M2 ;
      RECT 79.82 0.0 79.96 0.25 ;
      LAYER M1 ;
      RECT 79.82 0.0 79.96 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[47]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 189.26 0.0 189.4 0.25 ;
      LAYER M2 ;
      RECT 189.26 0.0 189.4 0.25 ;
      LAYER M3 ;
      RECT 189.26 0.0 189.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[96]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 78.98 0.0 79.12 0.25 ;
      LAYER M2 ;
      RECT 78.98 0.0 79.12 0.25 ;
      LAYER M1 ;
      RECT 78.98 0.0 79.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[47]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 189.54 0.0 189.68 0.25 ;
      LAYER M2 ;
      RECT 189.54 0.0 189.68 0.25 ;
      LAYER M3 ;
      RECT 189.54 0.0 189.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[97]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 78.7 0.0 78.84 0.25 ;
      LAYER M2 ;
      RECT 78.7 0.0 78.84 0.25 ;
      LAYER M1 ;
      RECT 78.7 0.0 78.84 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[46]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 190.31 0.0 190.45 0.25 ;
      LAYER M2 ;
      RECT 190.31 0.0 190.45 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[97]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 77.93 0.0 78.07 0.25 ;
      LAYER M1 ;
      RECT 77.93 0.0 78.07 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[46]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 191.74 0.0 191.88 0.25 ;
      LAYER M2 ;
      RECT 191.74 0.0 191.88 0.25 ;
      LAYER M3 ;
      RECT 191.74 0.0 191.88 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[98]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.5 0.0 76.64 0.25 ;
      LAYER M2 ;
      RECT 76.5 0.0 76.64 0.25 ;
      LAYER M1 ;
      RECT 76.5 0.0 76.64 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[45]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 192.58 0.0 192.72 0.25 ;
      LAYER M2 ;
      RECT 192.58 0.0 192.72 0.25 ;
      LAYER M3 ;
      RECT 192.58 0.0 192.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[98]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.66 0.0 75.8 0.25 ;
      LAYER M2 ;
      RECT 75.66 0.0 75.8 0.25 ;
      LAYER M1 ;
      RECT 75.66 0.0 75.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[45]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 192.86 0.0 193.0 0.25 ;
      LAYER M2 ;
      RECT 192.86 0.0 193.0 0.25 ;
      LAYER M3 ;
      RECT 192.86 0.0 193.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[99]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.38 0.0 75.52 0.25 ;
      LAYER M2 ;
      RECT 75.38 0.0 75.52 0.25 ;
      LAYER M1 ;
      RECT 75.38 0.0 75.52 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[44]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 193.63 0.0 193.77 0.25 ;
      LAYER M2 ;
      RECT 193.63 0.0 193.77 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[99]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 74.61 0.0 74.75 0.25 ;
      LAYER M1 ;
      RECT 74.61 0.0 74.75 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[44]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 195.06 0.0 195.2 0.25 ;
      LAYER M2 ;
      RECT 195.06 0.0 195.2 0.25 ;
      LAYER M3 ;
      RECT 195.06 0.0 195.2 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[100]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 73.18 0.0 73.32 0.25 ;
      LAYER M2 ;
      RECT 73.18 0.0 73.32 0.25 ;
      LAYER M1 ;
      RECT 73.18 0.0 73.32 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[43]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 195.9 0.0 196.04 0.25 ;
      LAYER M2 ;
      RECT 195.9 0.0 196.04 0.25 ;
      LAYER M3 ;
      RECT 195.9 0.0 196.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[100]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 72.34 0.0 72.48 0.25 ;
      LAYER M2 ;
      RECT 72.34 0.0 72.48 0.25 ;
      LAYER M1 ;
      RECT 72.34 0.0 72.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[43]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 196.18 0.0 196.32 0.25 ;
      LAYER M2 ;
      RECT 196.18 0.0 196.32 0.25 ;
      LAYER M3 ;
      RECT 196.18 0.0 196.32 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[101]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 72.06 0.0 72.2 0.25 ;
      LAYER M2 ;
      RECT 72.06 0.0 72.2 0.25 ;
      LAYER M1 ;
      RECT 72.06 0.0 72.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[42]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 196.95 0.0 197.09 0.25 ;
      LAYER M2 ;
      RECT 196.95 0.0 197.09 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[101]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 71.29 0.0 71.43 0.25 ;
      LAYER M1 ;
      RECT 71.29 0.0 71.43 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[42]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 198.38 0.0 198.52 0.25 ;
      LAYER M2 ;
      RECT 198.38 0.0 198.52 0.25 ;
      LAYER M3 ;
      RECT 198.38 0.0 198.52 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[102]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.86 0.0 70.0 0.25 ;
      LAYER M2 ;
      RECT 69.86 0.0 70.0 0.25 ;
      LAYER M1 ;
      RECT 69.86 0.0 70.0 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[41]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 199.22 0.0 199.36 0.25 ;
      LAYER M2 ;
      RECT 199.22 0.0 199.36 0.25 ;
      LAYER M3 ;
      RECT 199.22 0.0 199.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[102]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.02 0.0 69.16 0.25 ;
      LAYER M2 ;
      RECT 69.02 0.0 69.16 0.25 ;
      LAYER M1 ;
      RECT 69.02 0.0 69.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[41]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 199.5 0.0 199.64 0.25 ;
      LAYER M2 ;
      RECT 199.5 0.0 199.64 0.25 ;
      LAYER M3 ;
      RECT 199.5 0.0 199.64 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[103]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 68.74 0.0 68.88 0.25 ;
      LAYER M2 ;
      RECT 68.74 0.0 68.88 0.25 ;
      LAYER M1 ;
      RECT 68.74 0.0 68.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[40]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 200.27 0.0 200.41 0.25 ;
      LAYER M2 ;
      RECT 200.27 0.0 200.41 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[103]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 67.97 0.0 68.11 0.25 ;
      LAYER M1 ;
      RECT 67.97 0.0 68.11 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[40]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 201.7 0.0 201.84 0.25 ;
      LAYER M2 ;
      RECT 201.7 0.0 201.84 0.25 ;
      LAYER M3 ;
      RECT 201.7 0.0 201.84 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[104]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 66.54 0.0 66.68 0.25 ;
      LAYER M2 ;
      RECT 66.54 0.0 66.68 0.25 ;
      LAYER M1 ;
      RECT 66.54 0.0 66.68 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[39]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 202.54 0.0 202.68 0.25 ;
      LAYER M2 ;
      RECT 202.54 0.0 202.68 0.25 ;
      LAYER M3 ;
      RECT 202.54 0.0 202.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[104]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 65.7 0.0 65.84 0.25 ;
      LAYER M2 ;
      RECT 65.7 0.0 65.84 0.25 ;
      LAYER M1 ;
      RECT 65.7 0.0 65.84 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[39]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 202.82 0.0 202.96 0.25 ;
      LAYER M2 ;
      RECT 202.82 0.0 202.96 0.25 ;
      LAYER M3 ;
      RECT 202.82 0.0 202.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[105]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 65.42 0.0 65.56 0.25 ;
      LAYER M2 ;
      RECT 65.42 0.0 65.56 0.25 ;
      LAYER M1 ;
      RECT 65.42 0.0 65.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[38]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 203.59 0.0 203.73 0.25 ;
      LAYER M2 ;
      RECT 203.59 0.0 203.73 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[105]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 64.65 0.0 64.79 0.25 ;
      LAYER M1 ;
      RECT 64.65 0.0 64.79 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[38]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 205.02 0.0 205.16 0.25 ;
      LAYER M2 ;
      RECT 205.02 0.0 205.16 0.25 ;
      LAYER M3 ;
      RECT 205.02 0.0 205.16 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[106]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.22 0.0 63.36 0.25 ;
      LAYER M2 ;
      RECT 63.22 0.0 63.36 0.25 ;
      LAYER M1 ;
      RECT 63.22 0.0 63.36 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[37]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 205.86 0.0 206.0 0.25 ;
      LAYER M2 ;
      RECT 205.86 0.0 206.0 0.25 ;
      LAYER M3 ;
      RECT 205.86 0.0 206.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[106]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.38 0.0 62.52 0.25 ;
      LAYER M2 ;
      RECT 62.38 0.0 62.52 0.25 ;
      LAYER M1 ;
      RECT 62.38 0.0 62.52 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[37]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 206.14 0.0 206.28 0.25 ;
      LAYER M2 ;
      RECT 206.14 0.0 206.28 0.25 ;
      LAYER M3 ;
      RECT 206.14 0.0 206.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[107]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.1 0.0 62.24 0.25 ;
      LAYER M2 ;
      RECT 62.1 0.0 62.24 0.25 ;
      LAYER M1 ;
      RECT 62.1 0.0 62.24 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[36]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 206.91 0.0 207.05 0.25 ;
      LAYER M2 ;
      RECT 206.91 0.0 207.05 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[107]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 61.33 0.0 61.47 0.25 ;
      LAYER M1 ;
      RECT 61.33 0.0 61.47 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[36]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 208.34 0.0 208.48 0.25 ;
      LAYER M2 ;
      RECT 208.34 0.0 208.48 0.25 ;
      LAYER M3 ;
      RECT 208.34 0.0 208.48 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[108]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 59.9 0.0 60.04 0.25 ;
      LAYER M2 ;
      RECT 59.9 0.0 60.04 0.25 ;
      LAYER M1 ;
      RECT 59.9 0.0 60.04 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[35]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 209.18 0.0 209.32 0.25 ;
      LAYER M2 ;
      RECT 209.18 0.0 209.32 0.25 ;
      LAYER M3 ;
      RECT 209.18 0.0 209.32 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[108]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 59.06 0.0 59.2 0.25 ;
      LAYER M2 ;
      RECT 59.06 0.0 59.2 0.25 ;
      LAYER M1 ;
      RECT 59.06 0.0 59.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[35]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 209.46 0.0 209.6 0.25 ;
      LAYER M2 ;
      RECT 209.46 0.0 209.6 0.25 ;
      LAYER M3 ;
      RECT 209.46 0.0 209.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[109]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 58.78 0.0 58.92 0.25 ;
      LAYER M2 ;
      RECT 58.78 0.0 58.92 0.25 ;
      LAYER M1 ;
      RECT 58.78 0.0 58.92 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[34]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 210.23 0.0 210.37 0.25 ;
      LAYER M2 ;
      RECT 210.23 0.0 210.37 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[109]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 58.01 0.0 58.15 0.25 ;
      LAYER M1 ;
      RECT 58.01 0.0 58.15 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[34]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 211.66 0.0 211.8 0.25 ;
      LAYER M2 ;
      RECT 211.66 0.0 211.8 0.25 ;
      LAYER M3 ;
      RECT 211.66 0.0 211.8 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[110]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.58 0.0 56.72 0.25 ;
      LAYER M2 ;
      RECT 56.58 0.0 56.72 0.25 ;
      LAYER M1 ;
      RECT 56.58 0.0 56.72 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[33]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 212.5 0.0 212.64 0.25 ;
      LAYER M2 ;
      RECT 212.5 0.0 212.64 0.25 ;
      LAYER M3 ;
      RECT 212.5 0.0 212.64 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[110]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 55.74 0.0 55.88 0.25 ;
      LAYER M2 ;
      RECT 55.74 0.0 55.88 0.25 ;
      LAYER M1 ;
      RECT 55.74 0.0 55.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[33]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 212.78 0.0 212.92 0.25 ;
      LAYER M2 ;
      RECT 212.78 0.0 212.92 0.25 ;
      LAYER M3 ;
      RECT 212.78 0.0 212.92 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[111]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 55.46 0.0 55.6 0.25 ;
      LAYER M2 ;
      RECT 55.46 0.0 55.6 0.25 ;
      LAYER M1 ;
      RECT 55.46 0.0 55.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[32]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 213.55 0.0 213.69 0.25 ;
      LAYER M2 ;
      RECT 213.55 0.0 213.69 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[111]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 54.69 0.0 54.83 0.25 ;
      LAYER M1 ;
      RECT 54.69 0.0 54.83 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[32]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 214.98 0.0 215.12 0.25 ;
      LAYER M2 ;
      RECT 214.98 0.0 215.12 0.25 ;
      LAYER M3 ;
      RECT 214.98 0.0 215.12 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[112]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 53.26 0.0 53.4 0.25 ;
      LAYER M2 ;
      RECT 53.26 0.0 53.4 0.25 ;
      LAYER M1 ;
      RECT 53.26 0.0 53.4 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[31]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 215.82 0.0 215.96 0.25 ;
      LAYER M2 ;
      RECT 215.82 0.0 215.96 0.25 ;
      LAYER M3 ;
      RECT 215.82 0.0 215.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[112]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 52.42 0.0 52.56 0.25 ;
      LAYER M2 ;
      RECT 52.42 0.0 52.56 0.25 ;
      LAYER M1 ;
      RECT 52.42 0.0 52.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[31]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 216.1 0.0 216.24 0.25 ;
      LAYER M2 ;
      RECT 216.1 0.0 216.24 0.25 ;
      LAYER M3 ;
      RECT 216.1 0.0 216.24 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[113]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 52.14 0.0 52.28 0.25 ;
      LAYER M2 ;
      RECT 52.14 0.0 52.28 0.25 ;
      LAYER M1 ;
      RECT 52.14 0.0 52.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[30]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 216.87 0.0 217.01 0.25 ;
      LAYER M2 ;
      RECT 216.87 0.0 217.01 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[113]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 51.37 0.0 51.51 0.25 ;
      LAYER M1 ;
      RECT 51.37 0.0 51.51 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[30]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 218.3 0.0 218.44 0.25 ;
      LAYER M2 ;
      RECT 218.3 0.0 218.44 0.25 ;
      LAYER M3 ;
      RECT 218.3 0.0 218.44 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[114]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.94 0.0 50.08 0.25 ;
      LAYER M2 ;
      RECT 49.94 0.0 50.08 0.25 ;
      LAYER M1 ;
      RECT 49.94 0.0 50.08 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[29]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 219.14 0.0 219.28 0.25 ;
      LAYER M2 ;
      RECT 219.14 0.0 219.28 0.25 ;
      LAYER M3 ;
      RECT 219.14 0.0 219.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[114]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.1 0.0 49.24 0.25 ;
      LAYER M2 ;
      RECT 49.1 0.0 49.24 0.25 ;
      LAYER M1 ;
      RECT 49.1 0.0 49.24 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[29]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 219.42 0.0 219.56 0.25 ;
      LAYER M2 ;
      RECT 219.42 0.0 219.56 0.25 ;
      LAYER M3 ;
      RECT 219.42 0.0 219.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[115]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 48.82 0.0 48.96 0.25 ;
      LAYER M2 ;
      RECT 48.82 0.0 48.96 0.25 ;
      LAYER M1 ;
      RECT 48.82 0.0 48.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[28]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 220.19 0.0 220.33 0.25 ;
      LAYER M2 ;
      RECT 220.19 0.0 220.33 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[115]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 48.05 0.0 48.19 0.25 ;
      LAYER M1 ;
      RECT 48.05 0.0 48.19 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[28]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 221.62 0.0 221.76 0.25 ;
      LAYER M2 ;
      RECT 221.62 0.0 221.76 0.25 ;
      LAYER M3 ;
      RECT 221.62 0.0 221.76 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[116]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 46.62 0.0 46.76 0.25 ;
      LAYER M2 ;
      RECT 46.62 0.0 46.76 0.25 ;
      LAYER M1 ;
      RECT 46.62 0.0 46.76 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[27]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 222.46 0.0 222.6 0.25 ;
      LAYER M2 ;
      RECT 222.46 0.0 222.6 0.25 ;
      LAYER M3 ;
      RECT 222.46 0.0 222.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[116]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.78 0.0 45.92 0.25 ;
      LAYER M2 ;
      RECT 45.78 0.0 45.92 0.25 ;
      LAYER M1 ;
      RECT 45.78 0.0 45.92 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[27]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 222.74 0.0 222.88 0.25 ;
      LAYER M2 ;
      RECT 222.74 0.0 222.88 0.25 ;
      LAYER M3 ;
      RECT 222.74 0.0 222.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[117]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.5 0.0 45.64 0.25 ;
      LAYER M2 ;
      RECT 45.5 0.0 45.64 0.25 ;
      LAYER M1 ;
      RECT 45.5 0.0 45.64 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[26]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 223.51 0.0 223.65 0.25 ;
      LAYER M2 ;
      RECT 223.51 0.0 223.65 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[117]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 44.73 0.0 44.87 0.25 ;
      LAYER M1 ;
      RECT 44.73 0.0 44.87 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[26]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 224.94 0.0 225.08 0.25 ;
      LAYER M2 ;
      RECT 224.94 0.0 225.08 0.25 ;
      LAYER M3 ;
      RECT 224.94 0.0 225.08 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[118]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.3 0.0 43.44 0.25 ;
      LAYER M2 ;
      RECT 43.3 0.0 43.44 0.25 ;
      LAYER M1 ;
      RECT 43.3 0.0 43.44 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[25]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 225.78 0.0 225.92 0.25 ;
      LAYER M2 ;
      RECT 225.78 0.0 225.92 0.25 ;
      LAYER M3 ;
      RECT 225.78 0.0 225.92 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[118]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.46 0.0 42.6 0.25 ;
      LAYER M2 ;
      RECT 42.46 0.0 42.6 0.25 ;
      LAYER M1 ;
      RECT 42.46 0.0 42.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[25]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 226.06 0.0 226.2 0.25 ;
      LAYER M2 ;
      RECT 226.06 0.0 226.2 0.25 ;
      LAYER M3 ;
      RECT 226.06 0.0 226.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[119]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.18 0.0 42.32 0.25 ;
      LAYER M2 ;
      RECT 42.18 0.0 42.32 0.25 ;
      LAYER M1 ;
      RECT 42.18 0.0 42.32 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[24]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 226.83 0.0 226.97 0.25 ;
      LAYER M2 ;
      RECT 226.83 0.0 226.97 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[119]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 41.41 0.0 41.55 0.25 ;
      LAYER M1 ;
      RECT 41.41 0.0 41.55 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[24]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 228.26 0.0 228.4 0.25 ;
      LAYER M2 ;
      RECT 228.26 0.0 228.4 0.25 ;
      LAYER M3 ;
      RECT 228.26 0.0 228.4 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[120]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.98 0.0 40.12 0.25 ;
      LAYER M2 ;
      RECT 39.98 0.0 40.12 0.25 ;
      LAYER M1 ;
      RECT 39.98 0.0 40.12 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[23]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 229.1 0.0 229.24 0.25 ;
      LAYER M2 ;
      RECT 229.1 0.0 229.24 0.25 ;
      LAYER M3 ;
      RECT 229.1 0.0 229.24 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[120]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.14 0.0 39.28 0.25 ;
      LAYER M2 ;
      RECT 39.14 0.0 39.28 0.25 ;
      LAYER M1 ;
      RECT 39.14 0.0 39.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[23]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 229.38 0.0 229.52 0.25 ;
      LAYER M2 ;
      RECT 229.38 0.0 229.52 0.25 ;
      LAYER M3 ;
      RECT 229.38 0.0 229.52 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[121]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.86 0.0 39.0 0.25 ;
      LAYER M2 ;
      RECT 38.86 0.0 39.0 0.25 ;
      LAYER M1 ;
      RECT 38.86 0.0 39.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[22]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 230.15 0.0 230.29 0.25 ;
      LAYER M2 ;
      RECT 230.15 0.0 230.29 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[121]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 38.09 0.0 38.23 0.25 ;
      LAYER M1 ;
      RECT 38.09 0.0 38.23 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[22]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 231.58 0.0 231.72 0.25 ;
      LAYER M2 ;
      RECT 231.58 0.0 231.72 0.25 ;
      LAYER M3 ;
      RECT 231.58 0.0 231.72 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[122]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 36.66 0.0 36.8 0.25 ;
      LAYER M2 ;
      RECT 36.66 0.0 36.8 0.25 ;
      LAYER M1 ;
      RECT 36.66 0.0 36.8 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[21]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 232.42 0.0 232.56 0.25 ;
      LAYER M2 ;
      RECT 232.42 0.0 232.56 0.25 ;
      LAYER M3 ;
      RECT 232.42 0.0 232.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[122]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 35.82 0.0 35.96 0.25 ;
      LAYER M2 ;
      RECT 35.82 0.0 35.96 0.25 ;
      LAYER M1 ;
      RECT 35.82 0.0 35.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[21]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 232.7 0.0 232.84 0.25 ;
      LAYER M2 ;
      RECT 232.7 0.0 232.84 0.25 ;
      LAYER M3 ;
      RECT 232.7 0.0 232.84 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[123]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 35.54 0.0 35.68 0.25 ;
      LAYER M2 ;
      RECT 35.54 0.0 35.68 0.25 ;
      LAYER M1 ;
      RECT 35.54 0.0 35.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[20]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 233.47 0.0 233.61 0.25 ;
      LAYER M2 ;
      RECT 233.47 0.0 233.61 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[123]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 34.77 0.0 34.91 0.25 ;
      LAYER M1 ;
      RECT 34.77 0.0 34.91 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[20]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 234.9 0.0 235.04 0.25 ;
      LAYER M2 ;
      RECT 234.9 0.0 235.04 0.25 ;
      LAYER M3 ;
      RECT 234.9 0.0 235.04 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[124]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 33.34 0.0 33.48 0.25 ;
      LAYER M2 ;
      RECT 33.34 0.0 33.48 0.25 ;
      LAYER M1 ;
      RECT 33.34 0.0 33.48 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[19]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 235.74 0.0 235.88 0.25 ;
      LAYER M2 ;
      RECT 235.74 0.0 235.88 0.25 ;
      LAYER M3 ;
      RECT 235.74 0.0 235.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[124]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.5 0.0 32.64 0.25 ;
      LAYER M2 ;
      RECT 32.5 0.0 32.64 0.25 ;
      LAYER M1 ;
      RECT 32.5 0.0 32.64 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[19]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 236.02 0.0 236.16 0.25 ;
      LAYER M2 ;
      RECT 236.02 0.0 236.16 0.25 ;
      LAYER M3 ;
      RECT 236.02 0.0 236.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[125]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.22 0.0 32.36 0.25 ;
      LAYER M2 ;
      RECT 32.22 0.0 32.36 0.25 ;
      LAYER M1 ;
      RECT 32.22 0.0 32.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[18]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 236.79 0.0 236.93 0.25 ;
      LAYER M2 ;
      RECT 236.79 0.0 236.93 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[125]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 31.45 0.0 31.59 0.25 ;
      LAYER M1 ;
      RECT 31.45 0.0 31.59 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[18]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 238.22 0.0 238.36 0.25 ;
      LAYER M2 ;
      RECT 238.22 0.0 238.36 0.25 ;
      LAYER M3 ;
      RECT 238.22 0.0 238.36 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[126]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 30.02 0.0 30.16 0.25 ;
      LAYER M2 ;
      RECT 30.02 0.0 30.16 0.25 ;
      LAYER M1 ;
      RECT 30.02 0.0 30.16 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[17]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 239.06 0.0 239.2 0.25 ;
      LAYER M2 ;
      RECT 239.06 0.0 239.2 0.25 ;
      LAYER M3 ;
      RECT 239.06 0.0 239.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[126]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 29.18 0.0 29.32 0.25 ;
      LAYER M2 ;
      RECT 29.18 0.0 29.32 0.25 ;
      LAYER M1 ;
      RECT 29.18 0.0 29.32 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[17]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 239.34 0.0 239.48 0.25 ;
      LAYER M2 ;
      RECT 239.34 0.0 239.48 0.25 ;
      LAYER M3 ;
      RECT 239.34 0.0 239.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[127]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 28.9 0.0 29.04 0.25 ;
      LAYER M2 ;
      RECT 28.9 0.0 29.04 0.25 ;
      LAYER M1 ;
      RECT 28.9 0.0 29.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[16]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 240.11 0.0 240.25 0.25 ;
      LAYER M2 ;
      RECT 240.11 0.0 240.25 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[127]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 28.13 0.0 28.27 0.25 ;
      LAYER M1 ;
      RECT 28.13 0.0 28.27 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[16]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 241.54 0.0 241.68 0.25 ;
      LAYER M2 ;
      RECT 241.54 0.0 241.68 0.25 ;
      LAYER M3 ;
      RECT 241.54 0.0 241.68 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[128]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.7 0.0 26.84 0.25 ;
      LAYER M2 ;
      RECT 26.7 0.0 26.84 0.25 ;
      LAYER M1 ;
      RECT 26.7 0.0 26.84 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[15]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 242.38 0.0 242.52 0.25 ;
      LAYER M2 ;
      RECT 242.38 0.0 242.52 0.25 ;
      LAYER M3 ;
      RECT 242.38 0.0 242.52 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[128]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.86 0.0 26.0 0.25 ;
      LAYER M2 ;
      RECT 25.86 0.0 26.0 0.25 ;
      LAYER M1 ;
      RECT 25.86 0.0 26.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[15]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 242.66 0.0 242.8 0.25 ;
      LAYER M2 ;
      RECT 242.66 0.0 242.8 0.25 ;
      LAYER M3 ;
      RECT 242.66 0.0 242.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[129]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.58 0.0 25.72 0.25 ;
      LAYER M2 ;
      RECT 25.58 0.0 25.72 0.25 ;
      LAYER M1 ;
      RECT 25.58 0.0 25.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[14]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 243.43 0.0 243.57 0.25 ;
      LAYER M2 ;
      RECT 243.43 0.0 243.57 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[129]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 24.81 0.0 24.95 0.25 ;
      LAYER M1 ;
      RECT 24.81 0.0 24.95 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[14]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 244.86 0.0 245.0 0.25 ;
      LAYER M2 ;
      RECT 244.86 0.0 245.0 0.25 ;
      LAYER M3 ;
      RECT 244.86 0.0 245.0 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[130]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 23.38 0.0 23.52 0.25 ;
      LAYER M2 ;
      RECT 23.38 0.0 23.52 0.25 ;
      LAYER M1 ;
      RECT 23.38 0.0 23.52 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[13]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 245.7 0.0 245.84 0.25 ;
      LAYER M2 ;
      RECT 245.7 0.0 245.84 0.25 ;
      LAYER M3 ;
      RECT 245.7 0.0 245.84 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[130]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 22.54 0.0 22.68 0.25 ;
      LAYER M2 ;
      RECT 22.54 0.0 22.68 0.25 ;
      LAYER M1 ;
      RECT 22.54 0.0 22.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[13]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 245.98 0.0 246.12 0.25 ;
      LAYER M2 ;
      RECT 245.98 0.0 246.12 0.25 ;
      LAYER M3 ;
      RECT 245.98 0.0 246.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[131]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 22.26 0.0 22.4 0.25 ;
      LAYER M2 ;
      RECT 22.26 0.0 22.4 0.25 ;
      LAYER M1 ;
      RECT 22.26 0.0 22.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[12]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 246.75 0.0 246.89 0.25 ;
      LAYER M2 ;
      RECT 246.75 0.0 246.89 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[131]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 21.49 0.0 21.63 0.25 ;
      LAYER M1 ;
      RECT 21.49 0.0 21.63 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[12]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 248.18 0.0 248.32 0.25 ;
      LAYER M2 ;
      RECT 248.18 0.0 248.32 0.25 ;
      LAYER M3 ;
      RECT 248.18 0.0 248.32 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[132]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 20.06 0.0 20.2 0.25 ;
      LAYER M2 ;
      RECT 20.06 0.0 20.2 0.25 ;
      LAYER M1 ;
      RECT 20.06 0.0 20.2 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[11]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 249.02 0.0 249.16 0.25 ;
      LAYER M2 ;
      RECT 249.02 0.0 249.16 0.25 ;
      LAYER M3 ;
      RECT 249.02 0.0 249.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[132]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.22 0.0 19.36 0.25 ;
      LAYER M2 ;
      RECT 19.22 0.0 19.36 0.25 ;
      LAYER M1 ;
      RECT 19.22 0.0 19.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[11]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 249.3 0.0 249.44 0.25 ;
      LAYER M2 ;
      RECT 249.3 0.0 249.44 0.25 ;
      LAYER M3 ;
      RECT 249.3 0.0 249.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[133]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 18.94 0.0 19.08 0.25 ;
      LAYER M2 ;
      RECT 18.94 0.0 19.08 0.25 ;
      LAYER M1 ;
      RECT 18.94 0.0 19.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[10]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 250.07 0.0 250.21 0.25 ;
      LAYER M2 ;
      RECT 250.07 0.0 250.21 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[133]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 18.17 0.0 18.31 0.25 ;
      LAYER M1 ;
      RECT 18.17 0.0 18.31 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[10]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 251.5 0.0 251.64 0.25 ;
      LAYER M2 ;
      RECT 251.5 0.0 251.64 0.25 ;
      LAYER M3 ;
      RECT 251.5 0.0 251.64 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[134]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 16.74 0.0 16.88 0.25 ;
      LAYER M2 ;
      RECT 16.74 0.0 16.88 0.25 ;
      LAYER M1 ;
      RECT 16.74 0.0 16.88 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[9]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 252.34 0.0 252.48 0.25 ;
      LAYER M2 ;
      RECT 252.34 0.0 252.48 0.25 ;
      LAYER M3 ;
      RECT 252.34 0.0 252.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[134]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.9 0.0 16.04 0.25 ;
      LAYER M2 ;
      RECT 15.9 0.0 16.04 0.25 ;
      LAYER M1 ;
      RECT 15.9 0.0 16.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[9]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 252.62 0.0 252.76 0.25 ;
      LAYER M2 ;
      RECT 252.62 0.0 252.76 0.25 ;
      LAYER M3 ;
      RECT 252.62 0.0 252.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[135]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.62 0.0 15.76 0.25 ;
      LAYER M2 ;
      RECT 15.62 0.0 15.76 0.25 ;
      LAYER M1 ;
      RECT 15.62 0.0 15.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[8]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 253.39 0.0 253.53 0.25 ;
      LAYER M2 ;
      RECT 253.39 0.0 253.53 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[135]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 14.85 0.0 14.99 0.25 ;
      LAYER M1 ;
      RECT 14.85 0.0 14.99 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[8]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 254.82 0.0 254.96 0.25 ;
      LAYER M2 ;
      RECT 254.82 0.0 254.96 0.25 ;
      LAYER M3 ;
      RECT 254.82 0.0 254.96 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[136]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.42 0.0 13.56 0.25 ;
      LAYER M2 ;
      RECT 13.42 0.0 13.56 0.25 ;
      LAYER M1 ;
      RECT 13.42 0.0 13.56 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[7]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 255.66 0.0 255.8 0.25 ;
      LAYER M2 ;
      RECT 255.66 0.0 255.8 0.25 ;
      LAYER M3 ;
      RECT 255.66 0.0 255.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[136]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.58 0.0 12.72 0.25 ;
      LAYER M2 ;
      RECT 12.58 0.0 12.72 0.25 ;
      LAYER M1 ;
      RECT 12.58 0.0 12.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[7]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 255.94 0.0 256.08 0.25 ;
      LAYER M2 ;
      RECT 255.94 0.0 256.08 0.25 ;
      LAYER M3 ;
      RECT 255.94 0.0 256.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[137]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.3 0.0 12.44 0.25 ;
      LAYER M2 ;
      RECT 12.3 0.0 12.44 0.25 ;
      LAYER M1 ;
      RECT 12.3 0.0 12.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[6]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 256.71 0.0 256.85 0.25 ;
      LAYER M2 ;
      RECT 256.71 0.0 256.85 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[137]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 11.53 0.0 11.67 0.25 ;
      LAYER M1 ;
      RECT 11.53 0.0 11.67 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[6]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 258.14 0.0 258.28 0.25 ;
      LAYER M2 ;
      RECT 258.14 0.0 258.28 0.25 ;
      LAYER M3 ;
      RECT 258.14 0.0 258.28 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[138]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.1 0.0 10.24 0.25 ;
      LAYER M2 ;
      RECT 10.1 0.0 10.24 0.25 ;
      LAYER M1 ;
      RECT 10.1 0.0 10.24 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[5]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 258.98 0.0 259.12 0.25 ;
      LAYER M2 ;
      RECT 258.98 0.0 259.12 0.25 ;
      LAYER M3 ;
      RECT 258.98 0.0 259.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[138]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.26 0.0 9.4 0.25 ;
      LAYER M2 ;
      RECT 9.26 0.0 9.4 0.25 ;
      LAYER M1 ;
      RECT 9.26 0.0 9.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[5]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 259.26 0.0 259.4 0.25 ;
      LAYER M2 ;
      RECT 259.26 0.0 259.4 0.25 ;
      LAYER M3 ;
      RECT 259.26 0.0 259.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[139]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.98 0.0 9.12 0.25 ;
      LAYER M2 ;
      RECT 8.98 0.0 9.12 0.25 ;
      LAYER M1 ;
      RECT 8.98 0.0 9.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[4]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 260.03 0.0 260.17 0.25 ;
      LAYER M2 ;
      RECT 260.03 0.0 260.17 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[139]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 8.21 0.0 8.35 0.25 ;
      LAYER M1 ;
      RECT 8.21 0.0 8.35 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[4]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 261.46 0.0 261.6 0.25 ;
      LAYER M2 ;
      RECT 261.46 0.0 261.6 0.25 ;
      LAYER M3 ;
      RECT 261.46 0.0 261.6 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[140]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.78 0.0 6.92 0.25 ;
      LAYER M2 ;
      RECT 6.78 0.0 6.92 0.25 ;
      LAYER M1 ;
      RECT 6.78 0.0 6.92 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[3]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 262.3 0.0 262.44 0.25 ;
      LAYER M2 ;
      RECT 262.3 0.0 262.44 0.25 ;
      LAYER M3 ;
      RECT 262.3 0.0 262.44 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[140]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.94 0.0 6.08 0.25 ;
      LAYER M2 ;
      RECT 5.94 0.0 6.08 0.25 ;
      LAYER M1 ;
      RECT 5.94 0.0 6.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[3]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 262.58 0.0 262.72 0.25 ;
      LAYER M2 ;
      RECT 262.58 0.0 262.72 0.25 ;
      LAYER M3 ;
      RECT 262.58 0.0 262.72 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[141]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.66 0.0 5.8 0.25 ;
      LAYER M2 ;
      RECT 5.66 0.0 5.8 0.25 ;
      LAYER M1 ;
      RECT 5.66 0.0 5.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[2]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 263.35 0.0 263.49 0.25 ;
      LAYER M2 ;
      RECT 263.35 0.0 263.49 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[141]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 4.89 0.0 5.03 0.25 ;
      LAYER M1 ;
      RECT 4.89 0.0 5.03 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[2]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 264.78 0.0 264.92 0.25 ;
      LAYER M2 ;
      RECT 264.78 0.0 264.92 0.25 ;
      LAYER M3 ;
      RECT 264.78 0.0 264.92 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[142]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.46 0.0 3.6 0.25 ;
      LAYER M2 ;
      RECT 3.46 0.0 3.6 0.25 ;
      LAYER M1 ;
      RECT 3.46 0.0 3.6 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[1]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 265.62 0.0 265.76 0.25 ;
      LAYER M2 ;
      RECT 265.62 0.0 265.76 0.25 ;
      LAYER M3 ;
      RECT 265.62 0.0 265.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[142]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.62 0.0 2.76 0.25 ;
      LAYER M2 ;
      RECT 2.62 0.0 2.76 0.25 ;
      LAYER M1 ;
      RECT 2.62 0.0 2.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[1]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 265.9 0.0 266.04 0.25 ;
      LAYER M2 ;
      RECT 265.9 0.0 266.04 0.25 ;
      LAYER M3 ;
      RECT 265.9 0.0 266.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[143]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.34 0.0 2.48 0.25 ;
      LAYER M2 ;
      RECT 2.34 0.0 2.48 0.25 ;
      LAYER M1 ;
      RECT 2.34 0.0 2.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[0]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 266.67 0.0 266.81 0.25 ;
      LAYER M2 ;
      RECT 266.67 0.0 266.81 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[143]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 1.57 0.0 1.71 0.25 ;
      LAYER M1 ;
      RECT 1.57 0.0 1.71 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[0]
  PIN VDDPE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.59 0.0 0.7 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 0.995 0.0 1.275 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 4.315 0.0 4.595 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.635 0.0 7.915 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.955 0.0 11.235 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 14.275 0.0 14.555 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.595 0.0 17.875 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.915 0.0 21.195 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 24.235 0.0 24.515 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.555 0.0 27.835 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.875 0.0 31.155 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 34.195 0.0 34.475 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.515 0.0 37.795 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 40.835 0.0 41.115 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.155 0.0 44.435 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.475 0.0 47.755 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.795 0.0 51.075 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 54.115 0.0 54.395 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 57.435 0.0 57.715 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 60.755 0.0 61.035 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.075 0.0 64.355 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.395 0.0 67.675 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.715 0.0 70.995 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.035 0.0 74.315 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 77.355 0.0 77.635 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 80.675 0.0 80.955 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 83.995 0.0 84.275 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.315 0.0 87.595 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.635 0.0 90.915 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 93.955 0.0 94.235 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 97.275 0.0 97.555 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.595 0.0 100.875 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.915 0.0 104.195 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 107.235 0.0 107.515 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 110.555 0.0 110.835 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 113.875 0.0 114.155 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 117.195 0.0 117.475 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.595 0.0 120.705 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 122.375 0.0 122.485 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 124.68 0.0 124.96 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 127.32 0.0 127.53 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.065 0.0 128.215 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.705 0.0 128.935 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 129.415 0.0 129.685 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 131.385 0.0 131.655 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 133.575 0.0 133.785 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 136.5 0.0 136.78 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 137.59 0.0 137.73 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 138.33 0.0 138.48 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 138.69 0.0 138.96 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 141.9 0.0 142.18 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.31 0.0 143.52 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 145.835 0.0 145.975 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 146.765 0.0 146.975 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.675 0.0 147.785 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 150.905 0.0 151.185 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 154.225 0.0 154.505 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 157.545 0.0 157.825 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 160.865 0.0 161.145 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 164.185 0.0 164.465 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 167.505 0.0 167.785 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 170.825 0.0 171.105 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 174.145 0.0 174.425 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.465 0.0 177.745 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 180.785 0.0 181.065 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 184.105 0.0 184.385 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.425 0.0 187.705 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.745 0.0 191.025 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 194.065 0.0 194.345 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 197.385 0.0 197.665 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 200.705 0.0 200.985 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 204.025 0.0 204.305 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.345 0.0 207.625 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 210.665 0.0 210.945 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.985 0.0 214.265 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 217.305 0.0 217.585 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 220.625 0.0 220.905 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 223.945 0.0 224.225 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 227.265 0.0 227.545 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 230.585 0.0 230.865 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 233.905 0.0 234.185 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 237.225 0.0 237.505 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 240.545 0.0 240.825 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 243.865 0.0 244.145 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 247.185 0.0 247.465 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 250.505 0.0 250.785 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 253.825 0.0 254.105 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 257.145 0.0 257.425 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 260.465 0.0 260.745 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 263.785 0.0 264.065 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 267.105 0.0 267.385 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 267.68 0.0 267.79 100.88 ;
      END
    END VDDPE
  PIN VDDCE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.17 0.0 0.28 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 2.405 0.0 2.685 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 5.725 0.0 6.005 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 9.045 0.0 9.325 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.365 0.0 12.645 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.685 0.0 15.965 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.005 0.0 19.285 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 22.325 0.0 22.605 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.645 0.0 25.925 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.965 0.0 29.245 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.285 0.0 32.565 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.605 0.0 35.885 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.925 0.0 39.205 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.245 0.0 42.525 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.565 0.0 45.845 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.885 0.0 49.165 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 52.205 0.0 52.485 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.525 0.0 55.805 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.845 0.0 59.125 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 62.165 0.0 62.445 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 65.485 0.0 65.765 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.805 0.0 69.085 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.125 0.0 72.405 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.445 0.0 75.725 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.765 0.0 79.045 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.085 0.0 82.365 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 85.405 0.0 85.685 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.725 0.0 89.005 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.045 0.0 92.325 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 95.365 0.0 95.645 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.685 0.0 98.965 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 102.005 0.0 102.285 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 105.325 0.0 105.605 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.645 0.0 108.925 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 111.965 0.0 112.245 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 115.285 0.0 115.565 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.605 0.0 118.885 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 121.015 0.0 121.125 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.205 0.0 123.475 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.735 0.0 124.005 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 125.645 0.0 125.905 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 142.51 0.0 142.72 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.315 0.0 144.585 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.925 0.0 145.135 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.255 0.0 147.365 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 149.495 0.0 149.775 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 152.815 0.0 153.095 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.135 0.0 156.415 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 159.455 0.0 159.735 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 162.775 0.0 163.055 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 166.095 0.0 166.375 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 169.415 0.0 169.695 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 172.735 0.0 173.015 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 176.055 0.0 176.335 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 179.375 0.0 179.655 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 182.695 0.0 182.975 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 186.015 0.0 186.295 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 189.335 0.0 189.615 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 192.655 0.0 192.935 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 195.975 0.0 196.255 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.295 0.0 199.575 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 202.615 0.0 202.895 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 205.935 0.0 206.215 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 209.255 0.0 209.535 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 212.575 0.0 212.855 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.895 0.0 216.175 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 219.215 0.0 219.495 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 222.535 0.0 222.815 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.855 0.0 226.135 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.175 0.0 229.455 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.495 0.0 232.775 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.815 0.0 236.095 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.135 0.0 239.415 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.455 0.0 242.735 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 245.775 0.0 246.055 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.095 0.0 249.375 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.415 0.0 252.695 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 255.735 0.0 256.015 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 259.055 0.0 259.335 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.375 0.0 262.655 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 265.695 0.0 265.975 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 268.1 0.0 268.21 100.88 ;
      END
    END VDDCE
  PIN VSSE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.38 0.0 0.49 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 1.915 0.0 2.195 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 5.235 0.0 5.515 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 8.555 0.0 8.835 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 11.875 0.0 12.155 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.195 0.0 15.475 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 18.515 0.0 18.795 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 21.835 0.0 22.115 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.155 0.0 25.435 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.475 0.0 28.755 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 31.795 0.0 32.075 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.115 0.0 35.395 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.435 0.0 38.715 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 41.755 0.0 42.035 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.075 0.0 45.355 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.395 0.0 48.675 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.715 0.0 51.995 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.035 0.0 55.315 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.355 0.0 58.635 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.675 0.0 61.955 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.995 0.0 65.275 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.315 0.0 68.595 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 71.635 0.0 71.915 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.955 0.0 75.235 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.275 0.0 78.555 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.595 0.0 81.875 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.915 0.0 85.195 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.235 0.0 88.515 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 91.555 0.0 91.835 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.875 0.0 95.155 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.195 0.0 98.475 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 101.515 0.0 101.795 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 104.835 0.0 105.115 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.155 0.0 108.435 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 111.475 0.0 111.755 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 114.795 0.0 115.075 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.115 0.0 118.395 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.805 0.0 120.915 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 121.4 0.0 121.55 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 122.04 0.0 122.25 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 124.22 0.0 124.5 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 125.11 0.0 125.32 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 126.73 0.0 127.0 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 130.555 0.0 130.705 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 131.775 0.0 131.885 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 134.305 0.0 134.585 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 136.92 0.0 137.13 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 140.855 0.0 141.005 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 141.38 0.0 141.66 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.03 0.0 143.17 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.66 0.0 143.93 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 146.125 0.0 146.405 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.465 0.0 147.575 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 149.985 0.0 150.265 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 153.305 0.0 153.585 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.625 0.0 156.905 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 159.945 0.0 160.225 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 163.265 0.0 163.545 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 166.585 0.0 166.865 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 169.905 0.0 170.185 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 173.225 0.0 173.505 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 176.545 0.0 176.825 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 179.865 0.0 180.145 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 183.185 0.0 183.465 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 186.505 0.0 186.785 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 189.825 0.0 190.105 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 193.145 0.0 193.425 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.465 0.0 196.745 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.785 0.0 200.065 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 203.105 0.0 203.385 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 206.425 0.0 206.705 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 209.745 0.0 210.025 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.065 0.0 213.345 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 216.385 0.0 216.665 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 219.705 0.0 219.985 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 223.025 0.0 223.305 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 226.345 0.0 226.625 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.665 0.0 229.945 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.985 0.0 233.265 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 236.305 0.0 236.585 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.625 0.0 239.905 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.945 0.0 243.225 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 246.265 0.0 246.545 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.585 0.0 249.865 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.905 0.0 253.185 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 256.225 0.0 256.505 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 259.545 0.0 259.825 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.865 0.0 263.145 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 266.185 0.0 266.465 100.88 ;
      END
    PORT
      LAYER M4 ;
      RECT 267.89 0.0 268.0 100.88 ;
      END
    END VSSE
  OBS
    #otc obstructions
    LAYER M1 DESIGNRULEWIDTH 0.07 ;
    RECT 266.95 0.0 268.38 0.32 ;
    RECT 266.18 0.0 266.53 0.32 ;
    RECT 265.06 0.0 265.48 0.32 ;
    RECT 263.63 0.0 264.64 0.32 ;
    RECT 262.86 0.0 263.21 0.32 ;
    RECT 261.74 0.0 262.16 0.32 ;
    RECT 260.31 0.0 261.32 0.32 ;
    RECT 259.54 0.0 259.89 0.32 ;
    RECT 258.42 0.0 258.84 0.32 ;
    RECT 256.99 0.0 258.0 0.32 ;
    RECT 256.22 0.0 256.57 0.32 ;
    RECT 255.1 0.0 255.52 0.32 ;
    RECT 253.67 0.0 254.68 0.32 ;
    RECT 252.9 0.0 253.25 0.32 ;
    RECT 251.78 0.0 252.2 0.32 ;
    RECT 250.35 0.0 251.36 0.32 ;
    RECT 249.58 0.0 249.93 0.32 ;
    RECT 248.46 0.0 248.88 0.32 ;
    RECT 247.03 0.0 248.04 0.32 ;
    RECT 246.26 0.0 246.61 0.32 ;
    RECT 245.14 0.0 245.56 0.32 ;
    RECT 243.71 0.0 244.72 0.32 ;
    RECT 242.94 0.0 243.29 0.32 ;
    RECT 241.82 0.0 242.24 0.32 ;
    RECT 240.39 0.0 241.4 0.32 ;
    RECT 239.62 0.0 239.97 0.32 ;
    RECT 238.5 0.0 238.92 0.32 ;
    RECT 237.07 0.0 238.08 0.32 ;
    RECT 236.3 0.0 236.65 0.32 ;
    RECT 235.18 0.0 235.6 0.32 ;
    RECT 233.75 0.0 234.76 0.32 ;
    RECT 232.98 0.0 233.33 0.32 ;
    RECT 231.86 0.0 232.28 0.32 ;
    RECT 230.43 0.0 231.44 0.32 ;
    RECT 229.66 0.0 230.01 0.32 ;
    RECT 228.54 0.0 228.96 0.32 ;
    RECT 227.11 0.0 228.12 0.32 ;
    RECT 226.34 0.0 226.69 0.32 ;
    RECT 225.22 0.0 225.64 0.32 ;
    RECT 223.79 0.0 224.8 0.32 ;
    RECT 223.02 0.0 223.37 0.32 ;
    RECT 221.9 0.0 222.32 0.32 ;
    RECT 220.47 0.0 221.48 0.32 ;
    RECT 219.7 0.0 220.05 0.32 ;
    RECT 218.58 0.0 219.0 0.32 ;
    RECT 217.15 0.0 218.16 0.32 ;
    RECT 216.38 0.0 216.73 0.32 ;
    RECT 215.26 0.0 215.68 0.32 ;
    RECT 213.83 0.0 214.84 0.32 ;
    RECT 213.06 0.0 213.41 0.32 ;
    RECT 211.94 0.0 212.36 0.32 ;
    RECT 210.51 0.0 211.52 0.32 ;
    RECT 209.74 0.0 210.09 0.32 ;
    RECT 208.62 0.0 209.04 0.32 ;
    RECT 207.19 0.0 208.2 0.32 ;
    RECT 206.42 0.0 206.77 0.32 ;
    RECT 205.3 0.0 205.72 0.32 ;
    RECT 203.87 0.0 204.88 0.32 ;
    RECT 203.1 0.0 203.45 0.32 ;
    RECT 201.98 0.0 202.4 0.32 ;
    RECT 200.55 0.0 201.56 0.32 ;
    RECT 199.78 0.0 200.13 0.32 ;
    RECT 198.66 0.0 199.08 0.32 ;
    RECT 197.23 0.0 198.24 0.32 ;
    RECT 196.46 0.0 196.81 0.32 ;
    RECT 195.34 0.0 195.76 0.32 ;
    RECT 193.91 0.0 194.92 0.32 ;
    RECT 193.14 0.0 193.49 0.32 ;
    RECT 192.02 0.0 192.44 0.32 ;
    RECT 190.59 0.0 191.6 0.32 ;
    RECT 189.82 0.0 190.17 0.32 ;
    RECT 188.7 0.0 189.12 0.32 ;
    RECT 187.27 0.0 188.28 0.32 ;
    RECT 186.5 0.0 186.85 0.32 ;
    RECT 185.38 0.0 185.8 0.32 ;
    RECT 183.95 0.0 184.96 0.32 ;
    RECT 183.18 0.0 183.53 0.32 ;
    RECT 182.06 0.0 182.48 0.32 ;
    RECT 180.63 0.0 181.64 0.32 ;
    RECT 179.86 0.0 180.21 0.32 ;
    RECT 178.74 0.0 179.16 0.32 ;
    RECT 177.31 0.0 178.32 0.32 ;
    RECT 176.54 0.0 176.89 0.32 ;
    RECT 175.42 0.0 175.84 0.32 ;
    RECT 173.99 0.0 175.0 0.32 ;
    RECT 173.22 0.0 173.57 0.32 ;
    RECT 172.1 0.0 172.52 0.32 ;
    RECT 170.67 0.0 171.68 0.32 ;
    RECT 169.9 0.0 170.25 0.32 ;
    RECT 168.78 0.0 169.2 0.32 ;
    RECT 167.35 0.0 168.36 0.32 ;
    RECT 166.58 0.0 166.93 0.32 ;
    RECT 165.46 0.0 165.88 0.32 ;
    RECT 164.03 0.0 165.04 0.32 ;
    RECT 163.26 0.0 163.61 0.32 ;
    RECT 162.14 0.0 162.56 0.32 ;
    RECT 160.71 0.0 161.72 0.32 ;
    RECT 159.94 0.0 160.29 0.32 ;
    RECT 158.82 0.0 159.24 0.32 ;
    RECT 157.39 0.0 158.4 0.32 ;
    RECT 156.62 0.0 156.97 0.32 ;
    RECT 155.5 0.0 155.92 0.32 ;
    RECT 154.07 0.0 155.08 0.32 ;
    RECT 153.3 0.0 153.65 0.32 ;
    RECT 152.18 0.0 152.6 0.32 ;
    RECT 150.75 0.0 151.76 0.32 ;
    RECT 149.98 0.0 150.33 0.32 ;
    RECT 148.86 0.0 149.28 0.32 ;
    RECT 147.8 0.0 148.44 0.32 ;
    RECT 141.25 0.0 147.38 0.32 ;
    RECT 138.815 0.0 140.545 0.32 ;
    RECT 137.85 0.0 138.0 0.32 ;
    RECT 136.77 0.0 137.15 0.32 ;
    RECT 134.415 0.0 136.35 0.32 ;
    RECT 132.81 0.0 133.995 0.32 ;
    RECT 128.99 0.0 131.97 0.32 ;
    RECT 126.7 0.0 128.29 0.32 ;
    RECT 125.725 0.0 126.28 0.32 ;
    RECT 124.91 0.0 125.305 0.32 ;
    RECT 121.635 0.0 124.49 0.32 ;
    RECT 120.99 0.0 121.215 0.32 ;
    RECT 119.94 0.0 120.57 0.32 ;
    RECT 119.1 0.0 119.52 0.32 ;
    RECT 118.05 0.0 118.4 0.32 ;
    RECT 116.62 0.0 117.63 0.32 ;
    RECT 115.78 0.0 116.2 0.32 ;
    RECT 114.73 0.0 115.08 0.32 ;
    RECT 113.3 0.0 114.31 0.32 ;
    RECT 112.46 0.0 112.88 0.32 ;
    RECT 111.41 0.0 111.76 0.32 ;
    RECT 109.98 0.0 110.99 0.32 ;
    RECT 109.14 0.0 109.56 0.32 ;
    RECT 108.09 0.0 108.44 0.32 ;
    RECT 106.66 0.0 107.67 0.32 ;
    RECT 105.82 0.0 106.24 0.32 ;
    RECT 104.77 0.0 105.12 0.32 ;
    RECT 103.34 0.0 104.35 0.32 ;
    RECT 102.5 0.0 102.92 0.32 ;
    RECT 101.45 0.0 101.8 0.32 ;
    RECT 100.02 0.0 101.03 0.32 ;
    RECT 99.18 0.0 99.6 0.32 ;
    RECT 98.13 0.0 98.48 0.32 ;
    RECT 96.7 0.0 97.71 0.32 ;
    RECT 95.86 0.0 96.28 0.32 ;
    RECT 94.81 0.0 95.16 0.32 ;
    RECT 93.38 0.0 94.39 0.32 ;
    RECT 92.54 0.0 92.96 0.32 ;
    RECT 91.49 0.0 91.84 0.32 ;
    RECT 90.06 0.0 91.07 0.32 ;
    RECT 89.22 0.0 89.64 0.32 ;
    RECT 88.17 0.0 88.52 0.32 ;
    RECT 86.74 0.0 87.75 0.32 ;
    RECT 85.9 0.0 86.32 0.32 ;
    RECT 84.85 0.0 85.2 0.32 ;
    RECT 83.42 0.0 84.43 0.32 ;
    RECT 82.58 0.0 83.0 0.32 ;
    RECT 81.53 0.0 81.88 0.32 ;
    RECT 80.1 0.0 81.11 0.32 ;
    RECT 79.26 0.0 79.68 0.32 ;
    RECT 78.21 0.0 78.56 0.32 ;
    RECT 76.78 0.0 77.79 0.32 ;
    RECT 75.94 0.0 76.36 0.32 ;
    RECT 74.89 0.0 75.24 0.32 ;
    RECT 73.46 0.0 74.47 0.32 ;
    RECT 72.62 0.0 73.04 0.32 ;
    RECT 71.57 0.0 71.92 0.32 ;
    RECT 70.14 0.0 71.15 0.32 ;
    RECT 69.3 0.0 69.72 0.32 ;
    RECT 68.25 0.0 68.6 0.32 ;
    RECT 66.82 0.0 67.83 0.32 ;
    RECT 65.98 0.0 66.4 0.32 ;
    RECT 64.93 0.0 65.28 0.32 ;
    RECT 63.5 0.0 64.51 0.32 ;
    RECT 62.66 0.0 63.08 0.32 ;
    RECT 61.61 0.0 61.96 0.32 ;
    RECT 60.18 0.0 61.19 0.32 ;
    RECT 59.34 0.0 59.76 0.32 ;
    RECT 58.29 0.0 58.64 0.32 ;
    RECT 56.86 0.0 57.87 0.32 ;
    RECT 56.02 0.0 56.44 0.32 ;
    RECT 54.97 0.0 55.32 0.32 ;
    RECT 53.54 0.0 54.55 0.32 ;
    RECT 52.7 0.0 53.12 0.32 ;
    RECT 51.65 0.0 52.0 0.32 ;
    RECT 50.22 0.0 51.23 0.32 ;
    RECT 49.38 0.0 49.8 0.32 ;
    RECT 48.33 0.0 48.68 0.32 ;
    RECT 46.9 0.0 47.91 0.32 ;
    RECT 46.06 0.0 46.48 0.32 ;
    RECT 45.01 0.0 45.36 0.32 ;
    RECT 43.58 0.0 44.59 0.32 ;
    RECT 42.74 0.0 43.16 0.32 ;
    RECT 41.69 0.0 42.04 0.32 ;
    RECT 40.26 0.0 41.27 0.32 ;
    RECT 39.42 0.0 39.84 0.32 ;
    RECT 38.37 0.0 38.72 0.32 ;
    RECT 36.94 0.0 37.95 0.32 ;
    RECT 36.1 0.0 36.52 0.32 ;
    RECT 35.05 0.0 35.4 0.32 ;
    RECT 33.62 0.0 34.63 0.32 ;
    RECT 32.78 0.0 33.2 0.32 ;
    RECT 31.73 0.0 32.08 0.32 ;
    RECT 30.3 0.0 31.31 0.32 ;
    RECT 29.46 0.0 29.88 0.32 ;
    RECT 28.41 0.0 28.76 0.32 ;
    RECT 26.98 0.0 27.99 0.32 ;
    RECT 26.14 0.0 26.56 0.32 ;
    RECT 25.09 0.0 25.44 0.32 ;
    RECT 23.66 0.0 24.67 0.32 ;
    RECT 22.82 0.0 23.24 0.32 ;
    RECT 21.77 0.0 22.12 0.32 ;
    RECT 20.34 0.0 21.35 0.32 ;
    RECT 19.5 0.0 19.92 0.32 ;
    RECT 18.45 0.0 18.8 0.32 ;
    RECT 17.02 0.0 18.03 0.32 ;
    RECT 16.18 0.0 16.6 0.32 ;
    RECT 15.13 0.0 15.48 0.32 ;
    RECT 13.7 0.0 14.71 0.32 ;
    RECT 12.86 0.0 13.28 0.32 ;
    RECT 11.81 0.0 12.16 0.32 ;
    RECT 10.38 0.0 11.39 0.32 ;
    RECT 9.54 0.0 9.96 0.32 ;
    RECT 8.49 0.0 8.84 0.32 ;
    RECT 7.06 0.0 8.07 0.32 ;
    RECT 6.22 0.0 6.64 0.32 ;
    RECT 5.17 0.0 5.52 0.32 ;
    RECT 3.74 0.0 4.75 0.32 ;
    RECT 2.9 0.0 3.32 0.32 ;
    RECT 1.85 0.0 2.2 0.32 ;
    RECT 0.0 0.0 1.43 0.32 ;
    RECT 0.0 0.32 268.38 100.88 ;
    LAYER V1 ;
    RECT 0.0 0.0 268.38 100.88 ;
    LAYER M2 DESIGNRULEWIDTH 0.07 ;
    RECT 266.95 0.0 268.38 0.32 ;
    RECT 266.18 0.0 266.53 0.32 ;
    RECT 265.06 0.0 265.48 0.32 ;
    RECT 263.63 0.0 264.64 0.32 ;
    RECT 262.86 0.0 263.21 0.32 ;
    RECT 261.74 0.0 262.16 0.32 ;
    RECT 260.31 0.0 261.32 0.32 ;
    RECT 259.54 0.0 259.89 0.32 ;
    RECT 258.42 0.0 258.84 0.32 ;
    RECT 256.99 0.0 258.0 0.32 ;
    RECT 256.22 0.0 256.57 0.32 ;
    RECT 255.1 0.0 255.52 0.32 ;
    RECT 253.67 0.0 254.68 0.32 ;
    RECT 252.9 0.0 253.25 0.32 ;
    RECT 251.78 0.0 252.2 0.32 ;
    RECT 250.35 0.0 251.36 0.32 ;
    RECT 249.58 0.0 249.93 0.32 ;
    RECT 248.46 0.0 248.88 0.32 ;
    RECT 247.03 0.0 248.04 0.32 ;
    RECT 246.26 0.0 246.61 0.32 ;
    RECT 245.14 0.0 245.56 0.32 ;
    RECT 243.71 0.0 244.72 0.32 ;
    RECT 242.94 0.0 243.29 0.32 ;
    RECT 241.82 0.0 242.24 0.32 ;
    RECT 240.39 0.0 241.4 0.32 ;
    RECT 239.62 0.0 239.97 0.32 ;
    RECT 238.5 0.0 238.92 0.32 ;
    RECT 237.07 0.0 238.08 0.32 ;
    RECT 236.3 0.0 236.65 0.32 ;
    RECT 235.18 0.0 235.6 0.32 ;
    RECT 233.75 0.0 234.76 0.32 ;
    RECT 232.98 0.0 233.33 0.32 ;
    RECT 231.86 0.0 232.28 0.32 ;
    RECT 230.43 0.0 231.44 0.32 ;
    RECT 229.66 0.0 230.01 0.32 ;
    RECT 228.54 0.0 228.96 0.32 ;
    RECT 227.11 0.0 228.12 0.32 ;
    RECT 226.34 0.0 226.69 0.32 ;
    RECT 225.22 0.0 225.64 0.32 ;
    RECT 223.79 0.0 224.8 0.32 ;
    RECT 223.02 0.0 223.37 0.32 ;
    RECT 221.9 0.0 222.32 0.32 ;
    RECT 220.47 0.0 221.48 0.32 ;
    RECT 219.7 0.0 220.05 0.32 ;
    RECT 218.58 0.0 219.0 0.32 ;
    RECT 217.15 0.0 218.16 0.32 ;
    RECT 216.38 0.0 216.73 0.32 ;
    RECT 215.26 0.0 215.68 0.32 ;
    RECT 213.83 0.0 214.84 0.32 ;
    RECT 213.06 0.0 213.41 0.32 ;
    RECT 211.94 0.0 212.36 0.32 ;
    RECT 210.51 0.0 211.52 0.32 ;
    RECT 209.74 0.0 210.09 0.32 ;
    RECT 208.62 0.0 209.04 0.32 ;
    RECT 207.19 0.0 208.2 0.32 ;
    RECT 206.42 0.0 206.77 0.32 ;
    RECT 205.3 0.0 205.72 0.32 ;
    RECT 203.87 0.0 204.88 0.32 ;
    RECT 203.1 0.0 203.45 0.32 ;
    RECT 201.98 0.0 202.4 0.32 ;
    RECT 200.55 0.0 201.56 0.32 ;
    RECT 199.78 0.0 200.13 0.32 ;
    RECT 198.66 0.0 199.08 0.32 ;
    RECT 197.23 0.0 198.24 0.32 ;
    RECT 196.46 0.0 196.81 0.32 ;
    RECT 195.34 0.0 195.76 0.32 ;
    RECT 193.91 0.0 194.92 0.32 ;
    RECT 193.14 0.0 193.49 0.32 ;
    RECT 192.02 0.0 192.44 0.32 ;
    RECT 190.59 0.0 191.6 0.32 ;
    RECT 189.82 0.0 190.17 0.32 ;
    RECT 188.7 0.0 189.12 0.32 ;
    RECT 187.27 0.0 188.28 0.32 ;
    RECT 186.5 0.0 186.85 0.32 ;
    RECT 185.38 0.0 185.8 0.32 ;
    RECT 183.95 0.0 184.96 0.32 ;
    RECT 183.18 0.0 183.53 0.32 ;
    RECT 182.06 0.0 182.48 0.32 ;
    RECT 180.63 0.0 181.64 0.32 ;
    RECT 179.86 0.0 180.21 0.32 ;
    RECT 178.74 0.0 179.16 0.32 ;
    RECT 177.31 0.0 178.32 0.32 ;
    RECT 176.54 0.0 176.89 0.32 ;
    RECT 175.42 0.0 175.84 0.32 ;
    RECT 173.99 0.0 175.0 0.32 ;
    RECT 173.22 0.0 173.57 0.32 ;
    RECT 172.1 0.0 172.52 0.32 ;
    RECT 170.67 0.0 171.68 0.32 ;
    RECT 169.9 0.0 170.25 0.32 ;
    RECT 168.78 0.0 169.2 0.32 ;
    RECT 167.35 0.0 168.36 0.32 ;
    RECT 166.58 0.0 166.93 0.32 ;
    RECT 165.46 0.0 165.88 0.32 ;
    RECT 164.03 0.0 165.04 0.32 ;
    RECT 163.26 0.0 163.61 0.32 ;
    RECT 162.14 0.0 162.56 0.32 ;
    RECT 160.71 0.0 161.72 0.32 ;
    RECT 159.94 0.0 160.29 0.32 ;
    RECT 158.82 0.0 159.24 0.32 ;
    RECT 157.39 0.0 158.4 0.32 ;
    RECT 156.62 0.0 156.97 0.32 ;
    RECT 155.5 0.0 155.92 0.32 ;
    RECT 154.07 0.0 155.08 0.32 ;
    RECT 153.3 0.0 153.65 0.32 ;
    RECT 152.18 0.0 152.6 0.32 ;
    RECT 150.75 0.0 151.76 0.32 ;
    RECT 149.98 0.0 150.33 0.32 ;
    RECT 148.86 0.0 149.28 0.32 ;
    RECT 147.8 0.0 148.44 0.32 ;
    RECT 141.25 0.0 147.38 0.32 ;
    RECT 138.815 0.0 140.545 0.32 ;
    RECT 137.85 0.0 138.0 0.32 ;
    RECT 136.77 0.0 137.15 0.32 ;
    RECT 134.415 0.0 136.35 0.32 ;
    RECT 132.81 0.0 133.995 0.32 ;
    RECT 128.99 0.0 131.97 0.32 ;
    RECT 126.7 0.0 128.29 0.32 ;
    RECT 125.725 0.0 126.28 0.32 ;
    RECT 124.91 0.0 125.305 0.32 ;
    RECT 121.635 0.0 124.49 0.32 ;
    RECT 120.99 0.0 121.215 0.32 ;
    RECT 119.94 0.0 120.57 0.32 ;
    RECT 119.1 0.0 119.52 0.32 ;
    RECT 118.05 0.0 118.4 0.32 ;
    RECT 116.62 0.0 117.63 0.32 ;
    RECT 115.78 0.0 116.2 0.32 ;
    RECT 114.73 0.0 115.08 0.32 ;
    RECT 113.3 0.0 114.31 0.32 ;
    RECT 112.46 0.0 112.88 0.32 ;
    RECT 111.41 0.0 111.76 0.32 ;
    RECT 109.98 0.0 110.99 0.32 ;
    RECT 109.14 0.0 109.56 0.32 ;
    RECT 108.09 0.0 108.44 0.32 ;
    RECT 106.66 0.0 107.67 0.32 ;
    RECT 105.82 0.0 106.24 0.32 ;
    RECT 104.77 0.0 105.12 0.32 ;
    RECT 103.34 0.0 104.35 0.32 ;
    RECT 102.5 0.0 102.92 0.32 ;
    RECT 101.45 0.0 101.8 0.32 ;
    RECT 100.02 0.0 101.03 0.32 ;
    RECT 99.18 0.0 99.6 0.32 ;
    RECT 98.13 0.0 98.48 0.32 ;
    RECT 96.7 0.0 97.71 0.32 ;
    RECT 95.86 0.0 96.28 0.32 ;
    RECT 94.81 0.0 95.16 0.32 ;
    RECT 93.38 0.0 94.39 0.32 ;
    RECT 92.54 0.0 92.96 0.32 ;
    RECT 91.49 0.0 91.84 0.32 ;
    RECT 90.06 0.0 91.07 0.32 ;
    RECT 89.22 0.0 89.64 0.32 ;
    RECT 88.17 0.0 88.52 0.32 ;
    RECT 86.74 0.0 87.75 0.32 ;
    RECT 85.9 0.0 86.32 0.32 ;
    RECT 84.85 0.0 85.2 0.32 ;
    RECT 83.42 0.0 84.43 0.32 ;
    RECT 82.58 0.0 83.0 0.32 ;
    RECT 81.53 0.0 81.88 0.32 ;
    RECT 80.1 0.0 81.11 0.32 ;
    RECT 79.26 0.0 79.68 0.32 ;
    RECT 78.21 0.0 78.56 0.32 ;
    RECT 76.78 0.0 77.79 0.32 ;
    RECT 75.94 0.0 76.36 0.32 ;
    RECT 74.89 0.0 75.24 0.32 ;
    RECT 73.46 0.0 74.47 0.32 ;
    RECT 72.62 0.0 73.04 0.32 ;
    RECT 71.57 0.0 71.92 0.32 ;
    RECT 70.14 0.0 71.15 0.32 ;
    RECT 69.3 0.0 69.72 0.32 ;
    RECT 68.25 0.0 68.6 0.32 ;
    RECT 66.82 0.0 67.83 0.32 ;
    RECT 65.98 0.0 66.4 0.32 ;
    RECT 64.93 0.0 65.28 0.32 ;
    RECT 63.5 0.0 64.51 0.32 ;
    RECT 62.66 0.0 63.08 0.32 ;
    RECT 61.61 0.0 61.96 0.32 ;
    RECT 60.18 0.0 61.19 0.32 ;
    RECT 59.34 0.0 59.76 0.32 ;
    RECT 58.29 0.0 58.64 0.32 ;
    RECT 56.86 0.0 57.87 0.32 ;
    RECT 56.02 0.0 56.44 0.32 ;
    RECT 54.97 0.0 55.32 0.32 ;
    RECT 53.54 0.0 54.55 0.32 ;
    RECT 52.7 0.0 53.12 0.32 ;
    RECT 51.65 0.0 52.0 0.32 ;
    RECT 50.22 0.0 51.23 0.32 ;
    RECT 49.38 0.0 49.8 0.32 ;
    RECT 48.33 0.0 48.68 0.32 ;
    RECT 46.9 0.0 47.91 0.32 ;
    RECT 46.06 0.0 46.48 0.32 ;
    RECT 45.01 0.0 45.36 0.32 ;
    RECT 43.58 0.0 44.59 0.32 ;
    RECT 42.74 0.0 43.16 0.32 ;
    RECT 41.69 0.0 42.04 0.32 ;
    RECT 40.26 0.0 41.27 0.32 ;
    RECT 39.42 0.0 39.84 0.32 ;
    RECT 38.37 0.0 38.72 0.32 ;
    RECT 36.94 0.0 37.95 0.32 ;
    RECT 36.1 0.0 36.52 0.32 ;
    RECT 35.05 0.0 35.4 0.32 ;
    RECT 33.62 0.0 34.63 0.32 ;
    RECT 32.78 0.0 33.2 0.32 ;
    RECT 31.73 0.0 32.08 0.32 ;
    RECT 30.3 0.0 31.31 0.32 ;
    RECT 29.46 0.0 29.88 0.32 ;
    RECT 28.41 0.0 28.76 0.32 ;
    RECT 26.98 0.0 27.99 0.32 ;
    RECT 26.14 0.0 26.56 0.32 ;
    RECT 25.09 0.0 25.44 0.32 ;
    RECT 23.66 0.0 24.67 0.32 ;
    RECT 22.82 0.0 23.24 0.32 ;
    RECT 21.77 0.0 22.12 0.32 ;
    RECT 20.34 0.0 21.35 0.32 ;
    RECT 19.5 0.0 19.92 0.32 ;
    RECT 18.45 0.0 18.8 0.32 ;
    RECT 17.02 0.0 18.03 0.32 ;
    RECT 16.18 0.0 16.6 0.32 ;
    RECT 15.13 0.0 15.48 0.32 ;
    RECT 13.7 0.0 14.71 0.32 ;
    RECT 12.86 0.0 13.28 0.32 ;
    RECT 11.81 0.0 12.16 0.32 ;
    RECT 10.38 0.0 11.39 0.32 ;
    RECT 9.54 0.0 9.96 0.32 ;
    RECT 8.49 0.0 8.84 0.32 ;
    RECT 7.06 0.0 8.07 0.32 ;
    RECT 6.22 0.0 6.64 0.32 ;
    RECT 5.17 0.0 5.52 0.32 ;
    RECT 3.74 0.0 4.75 0.32 ;
    RECT 2.9 0.0 3.32 0.32 ;
    RECT 1.85 0.0 2.2 0.32 ;
    RECT 0.0 0.0 1.43 0.32 ;
    RECT 0.0 0.32 268.38 100.88 ;
    LAYER V2 ;
    RECT 0.0 0.0 268.38 100.88 ;
    LAYER M3 DESIGNRULEWIDTH 0.07 ;
    RECT 266.18 0.0 268.38 0.32 ;
    RECT 265.06 0.0 265.48 0.32 ;
    RECT 262.86 0.0 264.64 0.32 ;
    RECT 261.74 0.0 262.16 0.32 ;
    RECT 259.54 0.0 261.32 0.32 ;
    RECT 258.42 0.0 258.84 0.32 ;
    RECT 256.22 0.0 258.0 0.32 ;
    RECT 255.1 0.0 255.52 0.32 ;
    RECT 252.9 0.0 254.68 0.32 ;
    RECT 251.78 0.0 252.2 0.32 ;
    RECT 249.58 0.0 251.36 0.32 ;
    RECT 248.46 0.0 248.88 0.32 ;
    RECT 246.26 0.0 248.04 0.32 ;
    RECT 245.14 0.0 245.56 0.32 ;
    RECT 242.94 0.0 244.72 0.32 ;
    RECT 241.82 0.0 242.24 0.32 ;
    RECT 239.62 0.0 241.4 0.32 ;
    RECT 238.5 0.0 238.92 0.32 ;
    RECT 236.3 0.0 238.08 0.32 ;
    RECT 235.18 0.0 235.6 0.32 ;
    RECT 232.98 0.0 234.76 0.32 ;
    RECT 231.86 0.0 232.28 0.32 ;
    RECT 229.66 0.0 231.44 0.32 ;
    RECT 228.54 0.0 228.96 0.32 ;
    RECT 226.34 0.0 228.12 0.32 ;
    RECT 225.22 0.0 225.64 0.32 ;
    RECT 223.02 0.0 224.8 0.32 ;
    RECT 221.9 0.0 222.32 0.32 ;
    RECT 219.7 0.0 221.48 0.32 ;
    RECT 218.58 0.0 219.0 0.32 ;
    RECT 216.38 0.0 218.16 0.32 ;
    RECT 215.26 0.0 215.68 0.32 ;
    RECT 213.06 0.0 214.84 0.32 ;
    RECT 211.94 0.0 212.36 0.32 ;
    RECT 209.74 0.0 211.52 0.32 ;
    RECT 208.62 0.0 209.04 0.32 ;
    RECT 206.42 0.0 208.2 0.32 ;
    RECT 205.3 0.0 205.72 0.32 ;
    RECT 203.1 0.0 204.88 0.32 ;
    RECT 201.98 0.0 202.4 0.32 ;
    RECT 199.78 0.0 201.56 0.32 ;
    RECT 198.66 0.0 199.08 0.32 ;
    RECT 196.46 0.0 198.24 0.32 ;
    RECT 195.34 0.0 195.76 0.32 ;
    RECT 193.14 0.0 194.92 0.32 ;
    RECT 192.02 0.0 192.44 0.32 ;
    RECT 189.82 0.0 191.6 0.32 ;
    RECT 188.7 0.0 189.12 0.32 ;
    RECT 186.5 0.0 188.28 0.32 ;
    RECT 185.38 0.0 185.8 0.32 ;
    RECT 183.18 0.0 184.96 0.32 ;
    RECT 182.06 0.0 182.48 0.32 ;
    RECT 179.86 0.0 181.64 0.32 ;
    RECT 178.74 0.0 179.16 0.32 ;
    RECT 176.54 0.0 178.32 0.32 ;
    RECT 175.42 0.0 175.84 0.32 ;
    RECT 173.22 0.0 175.0 0.32 ;
    RECT 172.1 0.0 172.52 0.32 ;
    RECT 169.9 0.0 171.68 0.32 ;
    RECT 168.78 0.0 169.2 0.32 ;
    RECT 166.58 0.0 168.36 0.32 ;
    RECT 165.46 0.0 165.88 0.32 ;
    RECT 163.26 0.0 165.04 0.32 ;
    RECT 162.14 0.0 162.56 0.32 ;
    RECT 159.94 0.0 161.72 0.32 ;
    RECT 158.82 0.0 159.24 0.32 ;
    RECT 156.62 0.0 158.4 0.32 ;
    RECT 155.5 0.0 155.92 0.32 ;
    RECT 153.3 0.0 155.08 0.32 ;
    RECT 152.18 0.0 152.6 0.32 ;
    RECT 149.98 0.0 151.76 0.32 ;
    RECT 148.86 0.0 149.28 0.32 ;
    RECT 147.8 0.0 148.44 0.32 ;
    RECT 141.25 0.0 147.38 0.32 ;
    RECT 138.815 0.0 140.545 0.32 ;
    RECT 137.85 0.0 138.0 0.32 ;
    RECT 136.77 0.0 137.15 0.32 ;
    RECT 134.415 0.0 136.35 0.32 ;
    RECT 132.81 0.0 133.995 0.32 ;
    RECT 128.99 0.0 131.97 0.32 ;
    RECT 126.7 0.0 128.29 0.32 ;
    RECT 125.725 0.0 126.28 0.32 ;
    RECT 124.91 0.0 125.305 0.32 ;
    RECT 121.635 0.0 124.49 0.32 ;
    RECT 120.99 0.0 121.215 0.32 ;
    RECT 119.94 0.0 120.57 0.32 ;
    RECT 119.1 0.0 119.52 0.32 ;
    RECT 116.62 0.0 118.4 0.32 ;
    RECT 115.78 0.0 116.2 0.32 ;
    RECT 113.3 0.0 115.08 0.32 ;
    RECT 112.46 0.0 112.88 0.32 ;
    RECT 109.98 0.0 111.76 0.32 ;
    RECT 109.14 0.0 109.56 0.32 ;
    RECT 106.66 0.0 108.44 0.32 ;
    RECT 105.82 0.0 106.24 0.32 ;
    RECT 103.34 0.0 105.12 0.32 ;
    RECT 102.5 0.0 102.92 0.32 ;
    RECT 100.02 0.0 101.8 0.32 ;
    RECT 99.18 0.0 99.6 0.32 ;
    RECT 96.7 0.0 98.48 0.32 ;
    RECT 95.86 0.0 96.28 0.32 ;
    RECT 93.38 0.0 95.16 0.32 ;
    RECT 92.54 0.0 92.96 0.32 ;
    RECT 90.06 0.0 91.84 0.32 ;
    RECT 89.22 0.0 89.64 0.32 ;
    RECT 86.74 0.0 88.52 0.32 ;
    RECT 85.9 0.0 86.32 0.32 ;
    RECT 83.42 0.0 85.2 0.32 ;
    RECT 82.58 0.0 83.0 0.32 ;
    RECT 80.1 0.0 81.88 0.32 ;
    RECT 79.26 0.0 79.68 0.32 ;
    RECT 76.78 0.0 78.56 0.32 ;
    RECT 75.94 0.0 76.36 0.32 ;
    RECT 73.46 0.0 75.24 0.32 ;
    RECT 72.62 0.0 73.04 0.32 ;
    RECT 70.14 0.0 71.92 0.32 ;
    RECT 69.3 0.0 69.72 0.32 ;
    RECT 66.82 0.0 68.6 0.32 ;
    RECT 65.98 0.0 66.4 0.32 ;
    RECT 63.5 0.0 65.28 0.32 ;
    RECT 62.66 0.0 63.08 0.32 ;
    RECT 60.18 0.0 61.96 0.32 ;
    RECT 59.34 0.0 59.76 0.32 ;
    RECT 56.86 0.0 58.64 0.32 ;
    RECT 56.02 0.0 56.44 0.32 ;
    RECT 53.54 0.0 55.32 0.32 ;
    RECT 52.7 0.0 53.12 0.32 ;
    RECT 50.22 0.0 52.0 0.32 ;
    RECT 49.38 0.0 49.8 0.32 ;
    RECT 46.9 0.0 48.68 0.32 ;
    RECT 46.06 0.0 46.48 0.32 ;
    RECT 43.58 0.0 45.36 0.32 ;
    RECT 42.74 0.0 43.16 0.32 ;
    RECT 40.26 0.0 42.04 0.32 ;
    RECT 39.42 0.0 39.84 0.32 ;
    RECT 36.94 0.0 38.72 0.32 ;
    RECT 36.1 0.0 36.52 0.32 ;
    RECT 33.62 0.0 35.4 0.32 ;
    RECT 32.78 0.0 33.2 0.32 ;
    RECT 30.3 0.0 32.08 0.32 ;
    RECT 29.46 0.0 29.88 0.32 ;
    RECT 26.98 0.0 28.76 0.32 ;
    RECT 26.14 0.0 26.56 0.32 ;
    RECT 23.66 0.0 25.44 0.32 ;
    RECT 22.82 0.0 23.24 0.32 ;
    RECT 20.34 0.0 22.12 0.32 ;
    RECT 19.5 0.0 19.92 0.32 ;
    RECT 17.02 0.0 18.8 0.32 ;
    RECT 16.18 0.0 16.6 0.32 ;
    RECT 13.7 0.0 15.48 0.32 ;
    RECT 12.86 0.0 13.28 0.32 ;
    RECT 10.38 0.0 12.16 0.32 ;
    RECT 9.54 0.0 9.96 0.32 ;
    RECT 7.06 0.0 8.84 0.32 ;
    RECT 6.22 0.0 6.64 0.32 ;
    RECT 3.74 0.0 5.52 0.32 ;
    RECT 2.9 0.0 3.32 0.32 ;
    RECT 0.0 0.0 2.2 0.32 ;
    RECT 0.0 0.32 268.38 100.88 ;
    LAYER V3 ;
    RECT 0.0 0.0 268.38 100.88 ;
    LAYER V3 ;
    RECT 57.995 0.06 58.065 0.27 ;
    RECT 57.995 0.06 58.065 0.27 ;
    RECT 59.305 0.435 59.585 0.505 ;
    RECT 58.39 0.432 58.6 0.502 ;
    RECT 54.675 0.06 54.745 0.27 ;
    RECT 54.675 0.06 54.745 0.27 ;
    RECT 55.985 0.435 56.265 0.505 ;
    RECT 55.07 0.432 55.28 0.502 ;
    RECT 51.355 0.06 51.425 0.27 ;
    RECT 51.355 0.06 51.425 0.27 ;
    RECT 52.665 0.435 52.945 0.505 ;
    RECT 51.75 0.432 51.96 0.502 ;
    RECT 48.035 0.06 48.105 0.27 ;
    RECT 48.035 0.06 48.105 0.27 ;
    RECT 49.345 0.435 49.625 0.505 ;
    RECT 48.43 0.432 48.64 0.502 ;
    RECT 44.715 0.06 44.785 0.27 ;
    RECT 44.715 0.06 44.785 0.27 ;
    RECT 46.025 0.435 46.305 0.505 ;
    RECT 45.11 0.432 45.32 0.502 ;
    RECT 41.395 0.06 41.465 0.27 ;
    RECT 41.395 0.06 41.465 0.27 ;
    RECT 42.705 0.435 42.985 0.505 ;
    RECT 41.79 0.432 42.0 0.502 ;
    RECT 38.075 0.06 38.145 0.27 ;
    RECT 38.075 0.06 38.145 0.27 ;
    RECT 39.385 0.435 39.665 0.505 ;
    RECT 38.47 0.432 38.68 0.502 ;
    RECT 34.755 0.06 34.825 0.27 ;
    RECT 34.755 0.06 34.825 0.27 ;
    RECT 36.065 0.435 36.345 0.505 ;
    RECT 35.15 0.432 35.36 0.502 ;
    RECT 266.755 0.06 266.825 0.27 ;
    RECT 266.755 0.06 266.825 0.27 ;
    RECT 265.235 0.435 265.515 0.505 ;
    RECT 266.22 0.432 266.43 0.502 ;
    RECT 263.435 0.06 263.505 0.27 ;
    RECT 263.435 0.06 263.505 0.27 ;
    RECT 261.915 0.435 262.195 0.505 ;
    RECT 262.9 0.432 263.11 0.502 ;
    RECT 260.115 0.06 260.185 0.27 ;
    RECT 260.115 0.06 260.185 0.27 ;
    RECT 258.595 0.435 258.875 0.505 ;
    RECT 259.58 0.432 259.79 0.502 ;
    RECT 256.795 0.06 256.865 0.27 ;
    RECT 256.795 0.06 256.865 0.27 ;
    RECT 255.275 0.435 255.555 0.505 ;
    RECT 256.26 0.432 256.47 0.502 ;
    RECT 253.475 0.06 253.545 0.27 ;
    RECT 253.475 0.06 253.545 0.27 ;
    RECT 251.955 0.435 252.235 0.505 ;
    RECT 252.94 0.432 253.15 0.502 ;
    RECT 122.615 0.435 122.855 0.505 ;
    RECT 123.23 0.18 123.98 0.25 ;
    RECT 126.455 0.06 126.525 0.27 ;
    RECT 127.67 0.435 127.92 0.505 ;
    RECT 129.935 0.435 130.2 0.505 ;
    RECT 130.98 0.435 131.23 0.505 ;
    RECT 137.88 0.435 138.13 0.505 ;
    RECT 140.445 0.435 140.715 0.505 ;
    RECT 145.28 0.605 145.35 0.675 ;
    RECT 145.485 0.435 145.695 0.505 ;
    RECT 250.155 0.06 250.225 0.27 ;
    RECT 250.155 0.06 250.225 0.27 ;
    RECT 248.635 0.435 248.915 0.505 ;
    RECT 249.62 0.432 249.83 0.502 ;
    RECT 180.435 0.06 180.505 0.27 ;
    RECT 180.435 0.06 180.505 0.27 ;
    RECT 178.915 0.435 179.195 0.505 ;
    RECT 179.9 0.432 180.11 0.502 ;
    RECT 177.115 0.06 177.185 0.27 ;
    RECT 177.115 0.06 177.185 0.27 ;
    RECT 175.595 0.435 175.875 0.505 ;
    RECT 176.58 0.432 176.79 0.502 ;
    RECT 246.835 0.06 246.905 0.27 ;
    RECT 246.835 0.06 246.905 0.27 ;
    RECT 245.315 0.435 245.595 0.505 ;
    RECT 246.3 0.432 246.51 0.502 ;
    RECT 173.795 0.06 173.865 0.27 ;
    RECT 173.795 0.06 173.865 0.27 ;
    RECT 172.275 0.435 172.555 0.505 ;
    RECT 173.26 0.432 173.47 0.502 ;
    RECT 243.515 0.06 243.585 0.27 ;
    RECT 243.515 0.06 243.585 0.27 ;
    RECT 241.995 0.435 242.275 0.505 ;
    RECT 242.98 0.432 243.19 0.502 ;
    RECT 170.475 0.06 170.545 0.27 ;
    RECT 170.475 0.06 170.545 0.27 ;
    RECT 168.955 0.435 169.235 0.505 ;
    RECT 169.94 0.432 170.15 0.502 ;
    RECT 240.195 0.06 240.265 0.27 ;
    RECT 240.195 0.06 240.265 0.27 ;
    RECT 238.675 0.435 238.955 0.505 ;
    RECT 239.66 0.432 239.87 0.502 ;
    RECT 167.155 0.06 167.225 0.27 ;
    RECT 167.155 0.06 167.225 0.27 ;
    RECT 165.635 0.435 165.915 0.505 ;
    RECT 166.62 0.432 166.83 0.502 ;
    RECT 236.875 0.06 236.945 0.27 ;
    RECT 236.875 0.06 236.945 0.27 ;
    RECT 235.355 0.435 235.635 0.505 ;
    RECT 236.34 0.432 236.55 0.502 ;
    RECT 163.835 0.06 163.905 0.27 ;
    RECT 163.835 0.06 163.905 0.27 ;
    RECT 162.315 0.435 162.595 0.505 ;
    RECT 163.3 0.432 163.51 0.502 ;
    RECT 233.555 0.06 233.625 0.27 ;
    RECT 233.555 0.06 233.625 0.27 ;
    RECT 232.035 0.435 232.315 0.505 ;
    RECT 233.02 0.432 233.23 0.502 ;
    RECT 160.515 0.06 160.585 0.27 ;
    RECT 160.515 0.06 160.585 0.27 ;
    RECT 158.995 0.435 159.275 0.505 ;
    RECT 159.98 0.432 160.19 0.502 ;
    RECT 230.235 0.06 230.305 0.27 ;
    RECT 230.235 0.06 230.305 0.27 ;
    RECT 228.715 0.435 228.995 0.505 ;
    RECT 229.7 0.432 229.91 0.502 ;
    RECT 157.195 0.06 157.265 0.27 ;
    RECT 157.195 0.06 157.265 0.27 ;
    RECT 155.675 0.435 155.955 0.505 ;
    RECT 156.66 0.432 156.87 0.502 ;
    RECT 226.915 0.06 226.985 0.27 ;
    RECT 226.915 0.06 226.985 0.27 ;
    RECT 225.395 0.435 225.675 0.505 ;
    RECT 226.38 0.432 226.59 0.502 ;
    RECT 153.875 0.06 153.945 0.27 ;
    RECT 153.875 0.06 153.945 0.27 ;
    RECT 152.355 0.435 152.635 0.505 ;
    RECT 153.34 0.432 153.55 0.502 ;
    RECT 223.595 0.06 223.665 0.27 ;
    RECT 223.595 0.06 223.665 0.27 ;
    RECT 222.075 0.435 222.355 0.505 ;
    RECT 223.06 0.432 223.27 0.502 ;
    RECT 150.555 0.06 150.625 0.27 ;
    RECT 150.555 0.06 150.625 0.27 ;
    RECT 149.035 0.435 149.315 0.505 ;
    RECT 150.02 0.432 150.23 0.502 ;
    RECT 220.275 0.06 220.345 0.27 ;
    RECT 220.275 0.06 220.345 0.27 ;
    RECT 218.755 0.435 219.035 0.505 ;
    RECT 219.74 0.432 219.95 0.502 ;
    RECT 216.955 0.06 217.025 0.27 ;
    RECT 216.955 0.06 217.025 0.27 ;
    RECT 215.435 0.435 215.715 0.505 ;
    RECT 216.42 0.432 216.63 0.502 ;
    RECT 213.635 0.06 213.705 0.27 ;
    RECT 213.635 0.06 213.705 0.27 ;
    RECT 212.115 0.435 212.395 0.505 ;
    RECT 213.1 0.432 213.31 0.502 ;
    RECT 210.315 0.06 210.385 0.27 ;
    RECT 210.315 0.06 210.385 0.27 ;
    RECT 208.795 0.435 209.075 0.505 ;
    RECT 209.78 0.432 209.99 0.502 ;
    RECT 206.995 0.06 207.065 0.27 ;
    RECT 206.995 0.06 207.065 0.27 ;
    RECT 205.475 0.435 205.755 0.505 ;
    RECT 206.46 0.432 206.67 0.502 ;
    RECT 203.675 0.06 203.745 0.27 ;
    RECT 203.675 0.06 203.745 0.27 ;
    RECT 202.155 0.435 202.435 0.505 ;
    RECT 203.14 0.432 203.35 0.502 ;
    RECT 200.355 0.06 200.425 0.27 ;
    RECT 200.355 0.06 200.425 0.27 ;
    RECT 198.835 0.435 199.115 0.505 ;
    RECT 199.82 0.432 200.03 0.502 ;
    RECT 197.035 0.06 197.105 0.27 ;
    RECT 197.035 0.06 197.105 0.27 ;
    RECT 195.515 0.435 195.795 0.505 ;
    RECT 196.5 0.432 196.71 0.502 ;
    RECT 193.715 0.06 193.785 0.27 ;
    RECT 193.715 0.06 193.785 0.27 ;
    RECT 192.195 0.435 192.475 0.505 ;
    RECT 193.18 0.432 193.39 0.502 ;
    RECT 190.395 0.06 190.465 0.27 ;
    RECT 190.395 0.06 190.465 0.27 ;
    RECT 188.875 0.435 189.155 0.505 ;
    RECT 189.86 0.432 190.07 0.502 ;
    RECT 187.075 0.06 187.145 0.27 ;
    RECT 187.075 0.06 187.145 0.27 ;
    RECT 185.555 0.435 185.835 0.505 ;
    RECT 186.54 0.432 186.75 0.502 ;
    RECT 31.435 0.06 31.505 0.27 ;
    RECT 31.435 0.06 31.505 0.27 ;
    RECT 32.745 0.435 33.025 0.505 ;
    RECT 31.83 0.432 32.04 0.502 ;
    RECT 183.755 0.06 183.825 0.27 ;
    RECT 183.755 0.06 183.825 0.27 ;
    RECT 182.235 0.435 182.515 0.505 ;
    RECT 183.22 0.432 183.43 0.502 ;
    RECT 28.115 0.06 28.185 0.27 ;
    RECT 28.115 0.06 28.185 0.27 ;
    RECT 29.425 0.435 29.705 0.505 ;
    RECT 28.51 0.432 28.72 0.502 ;
    RECT 24.795 0.06 24.865 0.27 ;
    RECT 24.795 0.06 24.865 0.27 ;
    RECT 26.105 0.435 26.385 0.505 ;
    RECT 25.19 0.432 25.4 0.502 ;
    RECT 21.475 0.06 21.545 0.27 ;
    RECT 21.475 0.06 21.545 0.27 ;
    RECT 22.785 0.435 23.065 0.505 ;
    RECT 21.87 0.432 22.08 0.502 ;
    RECT 18.155 0.06 18.225 0.27 ;
    RECT 18.155 0.06 18.225 0.27 ;
    RECT 19.465 0.435 19.745 0.505 ;
    RECT 18.55 0.432 18.76 0.502 ;
    RECT 14.835 0.06 14.905 0.27 ;
    RECT 14.835 0.06 14.905 0.27 ;
    RECT 16.145 0.435 16.425 0.505 ;
    RECT 15.23 0.432 15.44 0.502 ;
    RECT 11.515 0.06 11.585 0.27 ;
    RECT 11.515 0.06 11.585 0.27 ;
    RECT 12.825 0.435 13.105 0.505 ;
    RECT 11.91 0.432 12.12 0.502 ;
    RECT 8.195 0.06 8.265 0.27 ;
    RECT 8.195 0.06 8.265 0.27 ;
    RECT 9.505 0.435 9.785 0.505 ;
    RECT 8.59 0.432 8.8 0.502 ;
    RECT 4.875 0.06 4.945 0.27 ;
    RECT 4.875 0.06 4.945 0.27 ;
    RECT 6.185 0.435 6.465 0.505 ;
    RECT 5.27 0.432 5.48 0.502 ;
    RECT 1.555 0.06 1.625 0.27 ;
    RECT 1.555 0.06 1.625 0.27 ;
    RECT 2.865 0.435 3.145 0.505 ;
    RECT 1.95 0.432 2.16 0.502 ;
    RECT 117.755 0.06 117.825 0.27 ;
    RECT 117.755 0.06 117.825 0.27 ;
    RECT 119.065 0.435 119.345 0.505 ;
    RECT 118.15 0.432 118.36 0.502 ;
    RECT 114.435 0.06 114.505 0.27 ;
    RECT 114.435 0.06 114.505 0.27 ;
    RECT 115.745 0.435 116.025 0.505 ;
    RECT 114.83 0.432 115.04 0.502 ;
    RECT 111.115 0.06 111.185 0.27 ;
    RECT 111.115 0.06 111.185 0.27 ;
    RECT 112.425 0.435 112.705 0.505 ;
    RECT 111.51 0.432 111.72 0.502 ;
    RECT 107.795 0.06 107.865 0.27 ;
    RECT 107.795 0.06 107.865 0.27 ;
    RECT 109.105 0.435 109.385 0.505 ;
    RECT 108.19 0.432 108.4 0.502 ;
    RECT 104.475 0.06 104.545 0.27 ;
    RECT 104.475 0.06 104.545 0.27 ;
    RECT 105.785 0.435 106.065 0.505 ;
    RECT 104.87 0.432 105.08 0.502 ;
    RECT 101.155 0.06 101.225 0.27 ;
    RECT 101.155 0.06 101.225 0.27 ;
    RECT 102.465 0.435 102.745 0.505 ;
    RECT 101.55 0.432 101.76 0.502 ;
    RECT 97.835 0.06 97.905 0.27 ;
    RECT 97.835 0.06 97.905 0.27 ;
    RECT 99.145 0.435 99.425 0.505 ;
    RECT 98.23 0.432 98.44 0.502 ;
    RECT 94.515 0.06 94.585 0.27 ;
    RECT 94.515 0.06 94.585 0.27 ;
    RECT 95.825 0.435 96.105 0.505 ;
    RECT 94.91 0.432 95.12 0.502 ;
    RECT 91.195 0.06 91.265 0.27 ;
    RECT 91.195 0.06 91.265 0.27 ;
    RECT 92.505 0.435 92.785 0.505 ;
    RECT 91.59 0.432 91.8 0.502 ;
    RECT 87.875 0.06 87.945 0.27 ;
    RECT 87.875 0.06 87.945 0.27 ;
    RECT 89.185 0.435 89.465 0.505 ;
    RECT 88.27 0.432 88.48 0.502 ;
    RECT 84.555 0.06 84.625 0.27 ;
    RECT 84.555 0.06 84.625 0.27 ;
    RECT 85.865 0.435 86.145 0.505 ;
    RECT 84.95 0.432 85.16 0.502 ;
    RECT 81.235 0.06 81.305 0.27 ;
    RECT 81.235 0.06 81.305 0.27 ;
    RECT 82.545 0.435 82.825 0.505 ;
    RECT 81.63 0.432 81.84 0.502 ;
    RECT 77.915 0.06 77.985 0.27 ;
    RECT 77.915 0.06 77.985 0.27 ;
    RECT 79.225 0.435 79.505 0.505 ;
    RECT 78.31 0.432 78.52 0.502 ;
    RECT 74.595 0.06 74.665 0.27 ;
    RECT 74.595 0.06 74.665 0.27 ;
    RECT 75.905 0.435 76.185 0.505 ;
    RECT 74.99 0.432 75.2 0.502 ;
    RECT 71.275 0.06 71.345 0.27 ;
    RECT 71.275 0.06 71.345 0.27 ;
    RECT 72.585 0.435 72.865 0.505 ;
    RECT 71.67 0.432 71.88 0.502 ;
    RECT 67.955 0.06 68.025 0.27 ;
    RECT 67.955 0.06 68.025 0.27 ;
    RECT 69.265 0.435 69.545 0.505 ;
    RECT 68.35 0.432 68.56 0.502 ;
    RECT 64.635 0.06 64.705 0.27 ;
    RECT 64.635 0.06 64.705 0.27 ;
    RECT 65.945 0.435 66.225 0.505 ;
    RECT 65.03 0.432 65.24 0.502 ;
    RECT 61.315 0.06 61.385 0.27 ;
    RECT 61.315 0.06 61.385 0.27 ;
    RECT 62.625 0.435 62.905 0.505 ;
    RECT 61.71 0.432 61.92 0.502 ;
    RECT 250.08 36.07 250.29 36.14 ;
    RECT 250.08 36.43 250.29 36.5 ;
    RECT 250.08 36.79 250.29 36.86 ;
    RECT 249.62 36.07 249.83 36.14 ;
    RECT 249.62 36.43 249.83 36.5 ;
    RECT 249.62 36.79 249.83 36.86 ;
    RECT 246.76 36.07 246.97 36.14 ;
    RECT 246.76 36.43 246.97 36.5 ;
    RECT 246.76 36.79 246.97 36.86 ;
    RECT 246.3 36.07 246.51 36.14 ;
    RECT 246.3 36.43 246.51 36.5 ;
    RECT 246.3 36.79 246.51 36.86 ;
    RECT 243.44 36.07 243.65 36.14 ;
    RECT 243.44 36.43 243.65 36.5 ;
    RECT 243.44 36.79 243.65 36.86 ;
    RECT 242.98 36.07 243.19 36.14 ;
    RECT 242.98 36.43 243.19 36.5 ;
    RECT 242.98 36.79 243.19 36.86 ;
    RECT 240.12 36.07 240.33 36.14 ;
    RECT 240.12 36.43 240.33 36.5 ;
    RECT 240.12 36.79 240.33 36.86 ;
    RECT 239.66 36.07 239.87 36.14 ;
    RECT 239.66 36.43 239.87 36.5 ;
    RECT 239.66 36.79 239.87 36.86 ;
    RECT 236.8 36.07 237.01 36.14 ;
    RECT 236.8 36.43 237.01 36.5 ;
    RECT 236.8 36.79 237.01 36.86 ;
    RECT 236.34 36.07 236.55 36.14 ;
    RECT 236.34 36.43 236.55 36.5 ;
    RECT 236.34 36.79 236.55 36.86 ;
    RECT 233.48 36.07 233.69 36.14 ;
    RECT 233.48 36.43 233.69 36.5 ;
    RECT 233.48 36.79 233.69 36.86 ;
    RECT 233.02 36.07 233.23 36.14 ;
    RECT 233.02 36.43 233.23 36.5 ;
    RECT 233.02 36.79 233.23 36.86 ;
    RECT 230.16 36.07 230.37 36.14 ;
    RECT 230.16 36.43 230.37 36.5 ;
    RECT 230.16 36.79 230.37 36.86 ;
    RECT 229.7 36.07 229.91 36.14 ;
    RECT 229.7 36.43 229.91 36.5 ;
    RECT 229.7 36.79 229.91 36.86 ;
    RECT 226.84 36.07 227.05 36.14 ;
    RECT 226.84 36.43 227.05 36.5 ;
    RECT 226.84 36.79 227.05 36.86 ;
    RECT 226.38 36.07 226.59 36.14 ;
    RECT 226.38 36.43 226.59 36.5 ;
    RECT 226.38 36.79 226.59 36.86 ;
    RECT 223.52 36.07 223.73 36.14 ;
    RECT 223.52 36.43 223.73 36.5 ;
    RECT 223.52 36.79 223.73 36.86 ;
    RECT 223.06 36.07 223.27 36.14 ;
    RECT 223.06 36.43 223.27 36.5 ;
    RECT 223.06 36.79 223.27 36.86 ;
    RECT 220.2 36.07 220.41 36.14 ;
    RECT 220.2 36.43 220.41 36.5 ;
    RECT 220.2 36.79 220.41 36.86 ;
    RECT 219.74 36.07 219.95 36.14 ;
    RECT 219.74 36.43 219.95 36.5 ;
    RECT 219.74 36.79 219.95 36.86 ;
    RECT 216.88 36.07 217.09 36.14 ;
    RECT 216.88 36.43 217.09 36.5 ;
    RECT 216.88 36.79 217.09 36.86 ;
    RECT 216.42 36.07 216.63 36.14 ;
    RECT 216.42 36.43 216.63 36.5 ;
    RECT 216.42 36.79 216.63 36.86 ;
    RECT 267.91 36.43 267.98 36.5 ;
    RECT 180.36 36.07 180.57 36.14 ;
    RECT 180.36 36.43 180.57 36.5 ;
    RECT 180.36 36.79 180.57 36.86 ;
    RECT 179.9 36.07 180.11 36.14 ;
    RECT 179.9 36.43 180.11 36.5 ;
    RECT 179.9 36.79 180.11 36.86 ;
    RECT 177.04 36.07 177.25 36.14 ;
    RECT 177.04 36.43 177.25 36.5 ;
    RECT 177.04 36.79 177.25 36.86 ;
    RECT 176.58 36.07 176.79 36.14 ;
    RECT 176.58 36.43 176.79 36.5 ;
    RECT 176.58 36.79 176.79 36.86 ;
    RECT 173.72 36.07 173.93 36.14 ;
    RECT 173.72 36.43 173.93 36.5 ;
    RECT 173.72 36.79 173.93 36.86 ;
    RECT 173.26 36.07 173.47 36.14 ;
    RECT 173.26 36.43 173.47 36.5 ;
    RECT 173.26 36.79 173.47 36.86 ;
    RECT 170.4 36.07 170.61 36.14 ;
    RECT 170.4 36.43 170.61 36.5 ;
    RECT 170.4 36.79 170.61 36.86 ;
    RECT 169.94 36.07 170.15 36.14 ;
    RECT 169.94 36.43 170.15 36.5 ;
    RECT 169.94 36.79 170.15 36.86 ;
    RECT 167.08 36.07 167.29 36.14 ;
    RECT 167.08 36.43 167.29 36.5 ;
    RECT 167.08 36.79 167.29 36.86 ;
    RECT 166.62 36.07 166.83 36.14 ;
    RECT 166.62 36.43 166.83 36.5 ;
    RECT 166.62 36.79 166.83 36.86 ;
    RECT 163.76 36.07 163.97 36.14 ;
    RECT 163.76 36.43 163.97 36.5 ;
    RECT 163.76 36.79 163.97 36.86 ;
    RECT 163.3 36.07 163.51 36.14 ;
    RECT 163.3 36.43 163.51 36.5 ;
    RECT 163.3 36.79 163.51 36.86 ;
    RECT 160.44 36.07 160.65 36.14 ;
    RECT 160.44 36.43 160.65 36.5 ;
    RECT 160.44 36.79 160.65 36.86 ;
    RECT 159.98 36.07 160.19 36.14 ;
    RECT 159.98 36.43 160.19 36.5 ;
    RECT 159.98 36.79 160.19 36.86 ;
    RECT 157.12 36.07 157.33 36.14 ;
    RECT 157.12 36.43 157.33 36.5 ;
    RECT 157.12 36.79 157.33 36.86 ;
    RECT 156.66 36.07 156.87 36.14 ;
    RECT 156.66 36.43 156.87 36.5 ;
    RECT 156.66 36.79 156.87 36.86 ;
    RECT 153.8 36.07 154.01 36.14 ;
    RECT 153.8 36.43 154.01 36.5 ;
    RECT 153.8 36.79 154.01 36.86 ;
    RECT 153.34 36.07 153.55 36.14 ;
    RECT 153.34 36.43 153.55 36.5 ;
    RECT 153.34 36.79 153.55 36.86 ;
    RECT 150.48 36.07 150.69 36.14 ;
    RECT 150.48 36.43 150.69 36.5 ;
    RECT 150.48 36.79 150.69 36.86 ;
    RECT 150.02 36.07 150.23 36.14 ;
    RECT 150.02 36.43 150.23 36.5 ;
    RECT 150.02 36.79 150.23 36.86 ;
    RECT 213.56 36.07 213.77 36.14 ;
    RECT 213.56 36.43 213.77 36.5 ;
    RECT 213.56 36.79 213.77 36.86 ;
    RECT 213.1 36.07 213.31 36.14 ;
    RECT 213.1 36.43 213.31 36.5 ;
    RECT 213.1 36.79 213.31 36.86 ;
    RECT 210.24 36.07 210.45 36.14 ;
    RECT 210.24 36.43 210.45 36.5 ;
    RECT 210.24 36.79 210.45 36.86 ;
    RECT 209.78 36.07 209.99 36.14 ;
    RECT 209.78 36.43 209.99 36.5 ;
    RECT 209.78 36.79 209.99 36.86 ;
    RECT 206.92 36.07 207.13 36.14 ;
    RECT 206.92 36.43 207.13 36.5 ;
    RECT 206.92 36.79 207.13 36.86 ;
    RECT 206.46 36.07 206.67 36.14 ;
    RECT 206.46 36.43 206.67 36.5 ;
    RECT 206.46 36.79 206.67 36.86 ;
    RECT 203.6 36.07 203.81 36.14 ;
    RECT 203.6 36.43 203.81 36.5 ;
    RECT 203.6 36.79 203.81 36.86 ;
    RECT 203.14 36.07 203.35 36.14 ;
    RECT 203.14 36.43 203.35 36.5 ;
    RECT 203.14 36.79 203.35 36.86 ;
    RECT 200.28 36.07 200.49 36.14 ;
    RECT 200.28 36.43 200.49 36.5 ;
    RECT 200.28 36.79 200.49 36.86 ;
    RECT 199.82 36.07 200.03 36.14 ;
    RECT 199.82 36.43 200.03 36.5 ;
    RECT 199.82 36.79 200.03 36.86 ;
    RECT 196.96 36.07 197.17 36.14 ;
    RECT 196.96 36.43 197.17 36.5 ;
    RECT 196.96 36.79 197.17 36.86 ;
    RECT 196.5 36.07 196.71 36.14 ;
    RECT 196.5 36.43 196.71 36.5 ;
    RECT 196.5 36.79 196.71 36.86 ;
    RECT 193.64 36.07 193.85 36.14 ;
    RECT 193.64 36.43 193.85 36.5 ;
    RECT 193.64 36.79 193.85 36.86 ;
    RECT 193.18 36.07 193.39 36.14 ;
    RECT 193.18 36.43 193.39 36.5 ;
    RECT 193.18 36.79 193.39 36.86 ;
    RECT 190.32 36.07 190.53 36.14 ;
    RECT 190.32 36.43 190.53 36.5 ;
    RECT 190.32 36.79 190.53 36.86 ;
    RECT 189.86 36.07 190.07 36.14 ;
    RECT 189.86 36.43 190.07 36.5 ;
    RECT 189.86 36.79 190.07 36.86 ;
    RECT 187.0 36.07 187.21 36.14 ;
    RECT 187.0 36.43 187.21 36.5 ;
    RECT 187.0 36.79 187.21 36.86 ;
    RECT 186.54 36.07 186.75 36.14 ;
    RECT 186.54 36.43 186.75 36.5 ;
    RECT 186.54 36.79 186.75 36.86 ;
    RECT 183.68 36.07 183.89 36.14 ;
    RECT 183.68 36.43 183.89 36.5 ;
    RECT 183.68 36.79 183.89 36.86 ;
    RECT 183.22 36.07 183.43 36.14 ;
    RECT 183.22 36.43 183.43 36.5 ;
    RECT 183.22 36.79 183.43 36.86 ;
    RECT 147.485 36.43 147.555 36.5 ;
    RECT 266.68 36.07 266.89 36.14 ;
    RECT 266.68 36.43 266.89 36.5 ;
    RECT 266.68 36.79 266.89 36.86 ;
    RECT 266.22 36.07 266.43 36.14 ;
    RECT 266.22 36.43 266.43 36.5 ;
    RECT 266.22 36.79 266.43 36.86 ;
    RECT 263.36 36.07 263.57 36.14 ;
    RECT 263.36 36.43 263.57 36.5 ;
    RECT 263.36 36.79 263.57 36.86 ;
    RECT 262.9 36.07 263.11 36.14 ;
    RECT 262.9 36.43 263.11 36.5 ;
    RECT 262.9 36.79 263.11 36.86 ;
    RECT 260.04 36.07 260.25 36.14 ;
    RECT 260.04 36.43 260.25 36.5 ;
    RECT 260.04 36.79 260.25 36.86 ;
    RECT 259.58 36.07 259.79 36.14 ;
    RECT 259.58 36.43 259.79 36.5 ;
    RECT 259.58 36.79 259.79 36.86 ;
    RECT 256.72 36.07 256.93 36.14 ;
    RECT 256.72 36.43 256.93 36.5 ;
    RECT 256.72 36.79 256.93 36.86 ;
    RECT 256.26 36.07 256.47 36.14 ;
    RECT 256.26 36.43 256.47 36.5 ;
    RECT 256.26 36.79 256.47 36.86 ;
    RECT 253.4 36.07 253.61 36.14 ;
    RECT 253.4 36.43 253.61 36.5 ;
    RECT 253.4 36.79 253.61 36.86 ;
    RECT 252.94 36.07 253.15 36.14 ;
    RECT 252.94 36.43 253.15 36.5 ;
    RECT 252.94 36.79 253.15 36.86 ;
    RECT 250.08 75.69 250.29 75.76 ;
    RECT 250.08 76.05 250.29 76.12 ;
    RECT 250.08 76.41 250.29 76.48 ;
    RECT 249.62 75.69 249.83 75.76 ;
    RECT 249.62 76.05 249.83 76.12 ;
    RECT 249.62 76.41 249.83 76.48 ;
    RECT 246.76 75.69 246.97 75.76 ;
    RECT 246.76 76.05 246.97 76.12 ;
    RECT 246.76 76.41 246.97 76.48 ;
    RECT 246.3 75.69 246.51 75.76 ;
    RECT 246.3 76.05 246.51 76.12 ;
    RECT 246.3 76.41 246.51 76.48 ;
    RECT 243.44 75.69 243.65 75.76 ;
    RECT 243.44 76.05 243.65 76.12 ;
    RECT 243.44 76.41 243.65 76.48 ;
    RECT 242.98 75.69 243.19 75.76 ;
    RECT 242.98 76.05 243.19 76.12 ;
    RECT 242.98 76.41 243.19 76.48 ;
    RECT 240.12 75.69 240.33 75.76 ;
    RECT 240.12 76.05 240.33 76.12 ;
    RECT 240.12 76.41 240.33 76.48 ;
    RECT 239.66 75.69 239.87 75.76 ;
    RECT 239.66 76.05 239.87 76.12 ;
    RECT 239.66 76.41 239.87 76.48 ;
    RECT 236.8 75.69 237.01 75.76 ;
    RECT 236.8 76.05 237.01 76.12 ;
    RECT 236.8 76.41 237.01 76.48 ;
    RECT 236.34 75.69 236.55 75.76 ;
    RECT 236.34 76.05 236.55 76.12 ;
    RECT 236.34 76.41 236.55 76.48 ;
    RECT 233.48 75.69 233.69 75.76 ;
    RECT 233.48 76.05 233.69 76.12 ;
    RECT 233.48 76.41 233.69 76.48 ;
    RECT 233.02 75.69 233.23 75.76 ;
    RECT 233.02 76.05 233.23 76.12 ;
    RECT 233.02 76.41 233.23 76.48 ;
    RECT 230.16 75.69 230.37 75.76 ;
    RECT 230.16 76.05 230.37 76.12 ;
    RECT 230.16 76.41 230.37 76.48 ;
    RECT 229.7 75.69 229.91 75.76 ;
    RECT 229.7 76.05 229.91 76.12 ;
    RECT 229.7 76.41 229.91 76.48 ;
    RECT 226.84 75.69 227.05 75.76 ;
    RECT 226.84 76.05 227.05 76.12 ;
    RECT 226.84 76.41 227.05 76.48 ;
    RECT 226.38 75.69 226.59 75.76 ;
    RECT 226.38 76.05 226.59 76.12 ;
    RECT 226.38 76.41 226.59 76.48 ;
    RECT 223.52 75.69 223.73 75.76 ;
    RECT 223.52 76.05 223.73 76.12 ;
    RECT 223.52 76.41 223.73 76.48 ;
    RECT 223.06 75.69 223.27 75.76 ;
    RECT 223.06 76.05 223.27 76.12 ;
    RECT 223.06 76.41 223.27 76.48 ;
    RECT 220.2 75.69 220.41 75.76 ;
    RECT 220.2 76.05 220.41 76.12 ;
    RECT 220.2 76.41 220.41 76.48 ;
    RECT 219.74 75.69 219.95 75.76 ;
    RECT 219.74 76.05 219.95 76.12 ;
    RECT 219.74 76.41 219.95 76.48 ;
    RECT 216.88 75.69 217.09 75.76 ;
    RECT 216.88 76.05 217.09 76.12 ;
    RECT 216.88 76.41 217.09 76.48 ;
    RECT 216.42 75.69 216.63 75.76 ;
    RECT 216.42 76.05 216.63 76.12 ;
    RECT 216.42 76.41 216.63 76.48 ;
    RECT 267.91 76.05 267.98 76.12 ;
    RECT 180.36 75.69 180.57 75.76 ;
    RECT 180.36 76.05 180.57 76.12 ;
    RECT 180.36 76.41 180.57 76.48 ;
    RECT 179.9 75.69 180.11 75.76 ;
    RECT 179.9 76.05 180.11 76.12 ;
    RECT 179.9 76.41 180.11 76.48 ;
    RECT 177.04 75.69 177.25 75.76 ;
    RECT 177.04 76.05 177.25 76.12 ;
    RECT 177.04 76.41 177.25 76.48 ;
    RECT 176.58 75.69 176.79 75.76 ;
    RECT 176.58 76.05 176.79 76.12 ;
    RECT 176.58 76.41 176.79 76.48 ;
    RECT 173.72 75.69 173.93 75.76 ;
    RECT 173.72 76.05 173.93 76.12 ;
    RECT 173.72 76.41 173.93 76.48 ;
    RECT 173.26 75.69 173.47 75.76 ;
    RECT 173.26 76.05 173.47 76.12 ;
    RECT 173.26 76.41 173.47 76.48 ;
    RECT 170.4 75.69 170.61 75.76 ;
    RECT 170.4 76.05 170.61 76.12 ;
    RECT 170.4 76.41 170.61 76.48 ;
    RECT 169.94 75.69 170.15 75.76 ;
    RECT 169.94 76.05 170.15 76.12 ;
    RECT 169.94 76.41 170.15 76.48 ;
    RECT 167.08 75.69 167.29 75.76 ;
    RECT 167.08 76.05 167.29 76.12 ;
    RECT 167.08 76.41 167.29 76.48 ;
    RECT 166.62 75.69 166.83 75.76 ;
    RECT 166.62 76.05 166.83 76.12 ;
    RECT 166.62 76.41 166.83 76.48 ;
    RECT 163.76 75.69 163.97 75.76 ;
    RECT 163.76 76.05 163.97 76.12 ;
    RECT 163.76 76.41 163.97 76.48 ;
    RECT 163.3 75.69 163.51 75.76 ;
    RECT 163.3 76.05 163.51 76.12 ;
    RECT 163.3 76.41 163.51 76.48 ;
    RECT 160.44 75.69 160.65 75.76 ;
    RECT 160.44 76.05 160.65 76.12 ;
    RECT 160.44 76.41 160.65 76.48 ;
    RECT 159.98 75.69 160.19 75.76 ;
    RECT 159.98 76.05 160.19 76.12 ;
    RECT 159.98 76.41 160.19 76.48 ;
    RECT 157.12 75.69 157.33 75.76 ;
    RECT 157.12 76.05 157.33 76.12 ;
    RECT 157.12 76.41 157.33 76.48 ;
    RECT 156.66 75.69 156.87 75.76 ;
    RECT 156.66 76.05 156.87 76.12 ;
    RECT 156.66 76.41 156.87 76.48 ;
    RECT 153.8 75.69 154.01 75.76 ;
    RECT 153.8 76.05 154.01 76.12 ;
    RECT 153.8 76.41 154.01 76.48 ;
    RECT 153.34 75.69 153.55 75.76 ;
    RECT 153.34 76.05 153.55 76.12 ;
    RECT 153.34 76.41 153.55 76.48 ;
    RECT 150.48 75.69 150.69 75.76 ;
    RECT 150.48 76.05 150.69 76.12 ;
    RECT 150.48 76.41 150.69 76.48 ;
    RECT 150.02 75.69 150.23 75.76 ;
    RECT 150.02 76.05 150.23 76.12 ;
    RECT 150.02 76.41 150.23 76.48 ;
    RECT 213.56 75.69 213.77 75.76 ;
    RECT 213.56 76.05 213.77 76.12 ;
    RECT 213.56 76.41 213.77 76.48 ;
    RECT 213.1 75.69 213.31 75.76 ;
    RECT 213.1 76.05 213.31 76.12 ;
    RECT 213.1 76.41 213.31 76.48 ;
    RECT 210.24 75.69 210.45 75.76 ;
    RECT 210.24 76.05 210.45 76.12 ;
    RECT 210.24 76.41 210.45 76.48 ;
    RECT 209.78 75.69 209.99 75.76 ;
    RECT 209.78 76.05 209.99 76.12 ;
    RECT 209.78 76.41 209.99 76.48 ;
    RECT 206.92 75.69 207.13 75.76 ;
    RECT 206.92 76.05 207.13 76.12 ;
    RECT 206.92 76.41 207.13 76.48 ;
    RECT 206.46 75.69 206.67 75.76 ;
    RECT 206.46 76.05 206.67 76.12 ;
    RECT 206.46 76.41 206.67 76.48 ;
    RECT 203.6 75.69 203.81 75.76 ;
    RECT 203.6 76.05 203.81 76.12 ;
    RECT 203.6 76.41 203.81 76.48 ;
    RECT 203.14 75.69 203.35 75.76 ;
    RECT 203.14 76.05 203.35 76.12 ;
    RECT 203.14 76.41 203.35 76.48 ;
    RECT 200.28 75.69 200.49 75.76 ;
    RECT 200.28 76.05 200.49 76.12 ;
    RECT 200.28 76.41 200.49 76.48 ;
    RECT 199.82 75.69 200.03 75.76 ;
    RECT 199.82 76.05 200.03 76.12 ;
    RECT 199.82 76.41 200.03 76.48 ;
    RECT 196.96 75.69 197.17 75.76 ;
    RECT 196.96 76.05 197.17 76.12 ;
    RECT 196.96 76.41 197.17 76.48 ;
    RECT 196.5 75.69 196.71 75.76 ;
    RECT 196.5 76.05 196.71 76.12 ;
    RECT 196.5 76.41 196.71 76.48 ;
    RECT 193.64 75.69 193.85 75.76 ;
    RECT 193.64 76.05 193.85 76.12 ;
    RECT 193.64 76.41 193.85 76.48 ;
    RECT 193.18 75.69 193.39 75.76 ;
    RECT 193.18 76.05 193.39 76.12 ;
    RECT 193.18 76.41 193.39 76.48 ;
    RECT 190.32 75.69 190.53 75.76 ;
    RECT 190.32 76.05 190.53 76.12 ;
    RECT 190.32 76.41 190.53 76.48 ;
    RECT 189.86 75.69 190.07 75.76 ;
    RECT 189.86 76.05 190.07 76.12 ;
    RECT 189.86 76.41 190.07 76.48 ;
    RECT 187.0 75.69 187.21 75.76 ;
    RECT 187.0 76.05 187.21 76.12 ;
    RECT 187.0 76.41 187.21 76.48 ;
    RECT 186.54 75.69 186.75 75.76 ;
    RECT 186.54 76.05 186.75 76.12 ;
    RECT 186.54 76.41 186.75 76.48 ;
    RECT 183.68 75.69 183.89 75.76 ;
    RECT 183.68 76.05 183.89 76.12 ;
    RECT 183.68 76.41 183.89 76.48 ;
    RECT 183.22 75.69 183.43 75.76 ;
    RECT 183.22 76.05 183.43 76.12 ;
    RECT 183.22 76.41 183.43 76.48 ;
    RECT 147.485 76.05 147.555 76.12 ;
    RECT 266.68 75.69 266.89 75.76 ;
    RECT 266.68 76.05 266.89 76.12 ;
    RECT 266.68 76.41 266.89 76.48 ;
    RECT 266.22 75.69 266.43 75.76 ;
    RECT 266.22 76.05 266.43 76.12 ;
    RECT 266.22 76.41 266.43 76.48 ;
    RECT 263.36 75.69 263.57 75.76 ;
    RECT 263.36 76.05 263.57 76.12 ;
    RECT 263.36 76.41 263.57 76.48 ;
    RECT 262.9 75.69 263.11 75.76 ;
    RECT 262.9 76.05 263.11 76.12 ;
    RECT 262.9 76.41 263.11 76.48 ;
    RECT 260.04 75.69 260.25 75.76 ;
    RECT 260.04 76.05 260.25 76.12 ;
    RECT 260.04 76.41 260.25 76.48 ;
    RECT 259.58 75.69 259.79 75.76 ;
    RECT 259.58 76.05 259.79 76.12 ;
    RECT 259.58 76.41 259.79 76.48 ;
    RECT 256.72 75.69 256.93 75.76 ;
    RECT 256.72 76.05 256.93 76.12 ;
    RECT 256.72 76.41 256.93 76.48 ;
    RECT 256.26 75.69 256.47 75.76 ;
    RECT 256.26 76.05 256.47 76.12 ;
    RECT 256.26 76.41 256.47 76.48 ;
    RECT 253.4 75.69 253.61 75.76 ;
    RECT 253.4 76.05 253.61 76.12 ;
    RECT 253.4 76.41 253.61 76.48 ;
    RECT 252.94 75.69 253.15 75.76 ;
    RECT 252.94 76.05 253.15 76.12 ;
    RECT 252.94 76.41 253.15 76.48 ;
    RECT 250.08 74.97 250.29 75.04 ;
    RECT 250.08 75.33 250.29 75.4 ;
    RECT 250.08 75.69 250.29 75.76 ;
    RECT 249.62 74.97 249.83 75.04 ;
    RECT 249.62 75.33 249.83 75.4 ;
    RECT 249.62 75.69 249.83 75.76 ;
    RECT 246.76 74.97 246.97 75.04 ;
    RECT 246.76 75.33 246.97 75.4 ;
    RECT 246.76 75.69 246.97 75.76 ;
    RECT 246.3 74.97 246.51 75.04 ;
    RECT 246.3 75.33 246.51 75.4 ;
    RECT 246.3 75.69 246.51 75.76 ;
    RECT 243.44 74.97 243.65 75.04 ;
    RECT 243.44 75.33 243.65 75.4 ;
    RECT 243.44 75.69 243.65 75.76 ;
    RECT 242.98 74.97 243.19 75.04 ;
    RECT 242.98 75.33 243.19 75.4 ;
    RECT 242.98 75.69 243.19 75.76 ;
    RECT 240.12 74.97 240.33 75.04 ;
    RECT 240.12 75.33 240.33 75.4 ;
    RECT 240.12 75.69 240.33 75.76 ;
    RECT 239.66 74.97 239.87 75.04 ;
    RECT 239.66 75.33 239.87 75.4 ;
    RECT 239.66 75.69 239.87 75.76 ;
    RECT 236.8 74.97 237.01 75.04 ;
    RECT 236.8 75.33 237.01 75.4 ;
    RECT 236.8 75.69 237.01 75.76 ;
    RECT 236.34 74.97 236.55 75.04 ;
    RECT 236.34 75.33 236.55 75.4 ;
    RECT 236.34 75.69 236.55 75.76 ;
    RECT 233.48 74.97 233.69 75.04 ;
    RECT 233.48 75.33 233.69 75.4 ;
    RECT 233.48 75.69 233.69 75.76 ;
    RECT 233.02 74.97 233.23 75.04 ;
    RECT 233.02 75.33 233.23 75.4 ;
    RECT 233.02 75.69 233.23 75.76 ;
    RECT 230.16 74.97 230.37 75.04 ;
    RECT 230.16 75.33 230.37 75.4 ;
    RECT 230.16 75.69 230.37 75.76 ;
    RECT 229.7 74.97 229.91 75.04 ;
    RECT 229.7 75.33 229.91 75.4 ;
    RECT 229.7 75.69 229.91 75.76 ;
    RECT 226.84 74.97 227.05 75.04 ;
    RECT 226.84 75.33 227.05 75.4 ;
    RECT 226.84 75.69 227.05 75.76 ;
    RECT 226.38 74.97 226.59 75.04 ;
    RECT 226.38 75.33 226.59 75.4 ;
    RECT 226.38 75.69 226.59 75.76 ;
    RECT 223.52 74.97 223.73 75.04 ;
    RECT 223.52 75.33 223.73 75.4 ;
    RECT 223.52 75.69 223.73 75.76 ;
    RECT 223.06 74.97 223.27 75.04 ;
    RECT 223.06 75.33 223.27 75.4 ;
    RECT 223.06 75.69 223.27 75.76 ;
    RECT 220.2 74.97 220.41 75.04 ;
    RECT 220.2 75.33 220.41 75.4 ;
    RECT 220.2 75.69 220.41 75.76 ;
    RECT 219.74 74.97 219.95 75.04 ;
    RECT 219.74 75.33 219.95 75.4 ;
    RECT 219.74 75.69 219.95 75.76 ;
    RECT 216.88 74.97 217.09 75.04 ;
    RECT 216.88 75.33 217.09 75.4 ;
    RECT 216.88 75.69 217.09 75.76 ;
    RECT 216.42 74.97 216.63 75.04 ;
    RECT 216.42 75.33 216.63 75.4 ;
    RECT 216.42 75.69 216.63 75.76 ;
    RECT 267.91 75.33 267.98 75.4 ;
    RECT 180.36 74.97 180.57 75.04 ;
    RECT 180.36 75.33 180.57 75.4 ;
    RECT 180.36 75.69 180.57 75.76 ;
    RECT 179.9 74.97 180.11 75.04 ;
    RECT 179.9 75.33 180.11 75.4 ;
    RECT 179.9 75.69 180.11 75.76 ;
    RECT 177.04 74.97 177.25 75.04 ;
    RECT 177.04 75.33 177.25 75.4 ;
    RECT 177.04 75.69 177.25 75.76 ;
    RECT 176.58 74.97 176.79 75.04 ;
    RECT 176.58 75.33 176.79 75.4 ;
    RECT 176.58 75.69 176.79 75.76 ;
    RECT 173.72 74.97 173.93 75.04 ;
    RECT 173.72 75.33 173.93 75.4 ;
    RECT 173.72 75.69 173.93 75.76 ;
    RECT 173.26 74.97 173.47 75.04 ;
    RECT 173.26 75.33 173.47 75.4 ;
    RECT 173.26 75.69 173.47 75.76 ;
    RECT 170.4 74.97 170.61 75.04 ;
    RECT 170.4 75.33 170.61 75.4 ;
    RECT 170.4 75.69 170.61 75.76 ;
    RECT 169.94 74.97 170.15 75.04 ;
    RECT 169.94 75.33 170.15 75.4 ;
    RECT 169.94 75.69 170.15 75.76 ;
    RECT 167.08 74.97 167.29 75.04 ;
    RECT 167.08 75.33 167.29 75.4 ;
    RECT 167.08 75.69 167.29 75.76 ;
    RECT 166.62 74.97 166.83 75.04 ;
    RECT 166.62 75.33 166.83 75.4 ;
    RECT 166.62 75.69 166.83 75.76 ;
    RECT 163.76 74.97 163.97 75.04 ;
    RECT 163.76 75.33 163.97 75.4 ;
    RECT 163.76 75.69 163.97 75.76 ;
    RECT 163.3 74.97 163.51 75.04 ;
    RECT 163.3 75.33 163.51 75.4 ;
    RECT 163.3 75.69 163.51 75.76 ;
    RECT 160.44 74.97 160.65 75.04 ;
    RECT 160.44 75.33 160.65 75.4 ;
    RECT 160.44 75.69 160.65 75.76 ;
    RECT 159.98 74.97 160.19 75.04 ;
    RECT 159.98 75.33 160.19 75.4 ;
    RECT 159.98 75.69 160.19 75.76 ;
    RECT 157.12 74.97 157.33 75.04 ;
    RECT 157.12 75.33 157.33 75.4 ;
    RECT 157.12 75.69 157.33 75.76 ;
    RECT 156.66 74.97 156.87 75.04 ;
    RECT 156.66 75.33 156.87 75.4 ;
    RECT 156.66 75.69 156.87 75.76 ;
    RECT 153.8 74.97 154.01 75.04 ;
    RECT 153.8 75.33 154.01 75.4 ;
    RECT 153.8 75.69 154.01 75.76 ;
    RECT 153.34 74.97 153.55 75.04 ;
    RECT 153.34 75.33 153.55 75.4 ;
    RECT 153.34 75.69 153.55 75.76 ;
    RECT 150.48 74.97 150.69 75.04 ;
    RECT 150.48 75.33 150.69 75.4 ;
    RECT 150.48 75.69 150.69 75.76 ;
    RECT 150.02 74.97 150.23 75.04 ;
    RECT 150.02 75.33 150.23 75.4 ;
    RECT 150.02 75.69 150.23 75.76 ;
    RECT 213.56 74.97 213.77 75.04 ;
    RECT 213.56 75.33 213.77 75.4 ;
    RECT 213.56 75.69 213.77 75.76 ;
    RECT 213.1 74.97 213.31 75.04 ;
    RECT 213.1 75.33 213.31 75.4 ;
    RECT 213.1 75.69 213.31 75.76 ;
    RECT 210.24 74.97 210.45 75.04 ;
    RECT 210.24 75.33 210.45 75.4 ;
    RECT 210.24 75.69 210.45 75.76 ;
    RECT 209.78 74.97 209.99 75.04 ;
    RECT 209.78 75.33 209.99 75.4 ;
    RECT 209.78 75.69 209.99 75.76 ;
    RECT 206.92 74.97 207.13 75.04 ;
    RECT 206.92 75.33 207.13 75.4 ;
    RECT 206.92 75.69 207.13 75.76 ;
    RECT 206.46 74.97 206.67 75.04 ;
    RECT 206.46 75.33 206.67 75.4 ;
    RECT 206.46 75.69 206.67 75.76 ;
    RECT 203.6 74.97 203.81 75.04 ;
    RECT 203.6 75.33 203.81 75.4 ;
    RECT 203.6 75.69 203.81 75.76 ;
    RECT 203.14 74.97 203.35 75.04 ;
    RECT 203.14 75.33 203.35 75.4 ;
    RECT 203.14 75.69 203.35 75.76 ;
    RECT 200.28 74.97 200.49 75.04 ;
    RECT 200.28 75.33 200.49 75.4 ;
    RECT 200.28 75.69 200.49 75.76 ;
    RECT 199.82 74.97 200.03 75.04 ;
    RECT 199.82 75.33 200.03 75.4 ;
    RECT 199.82 75.69 200.03 75.76 ;
    RECT 196.96 74.97 197.17 75.04 ;
    RECT 196.96 75.33 197.17 75.4 ;
    RECT 196.96 75.69 197.17 75.76 ;
    RECT 196.5 74.97 196.71 75.04 ;
    RECT 196.5 75.33 196.71 75.4 ;
    RECT 196.5 75.69 196.71 75.76 ;
    RECT 193.64 74.97 193.85 75.04 ;
    RECT 193.64 75.33 193.85 75.4 ;
    RECT 193.64 75.69 193.85 75.76 ;
    RECT 193.18 74.97 193.39 75.04 ;
    RECT 193.18 75.33 193.39 75.4 ;
    RECT 193.18 75.69 193.39 75.76 ;
    RECT 190.32 74.97 190.53 75.04 ;
    RECT 190.32 75.33 190.53 75.4 ;
    RECT 190.32 75.69 190.53 75.76 ;
    RECT 189.86 74.97 190.07 75.04 ;
    RECT 189.86 75.33 190.07 75.4 ;
    RECT 189.86 75.69 190.07 75.76 ;
    RECT 187.0 74.97 187.21 75.04 ;
    RECT 187.0 75.33 187.21 75.4 ;
    RECT 187.0 75.69 187.21 75.76 ;
    RECT 186.54 74.97 186.75 75.04 ;
    RECT 186.54 75.33 186.75 75.4 ;
    RECT 186.54 75.69 186.75 75.76 ;
    RECT 183.68 74.97 183.89 75.04 ;
    RECT 183.68 75.33 183.89 75.4 ;
    RECT 183.68 75.69 183.89 75.76 ;
    RECT 183.22 74.97 183.43 75.04 ;
    RECT 183.22 75.33 183.43 75.4 ;
    RECT 183.22 75.69 183.43 75.76 ;
    RECT 147.485 75.33 147.555 75.4 ;
    RECT 266.68 74.97 266.89 75.04 ;
    RECT 266.68 75.33 266.89 75.4 ;
    RECT 266.68 75.69 266.89 75.76 ;
    RECT 266.22 74.97 266.43 75.04 ;
    RECT 266.22 75.33 266.43 75.4 ;
    RECT 266.22 75.69 266.43 75.76 ;
    RECT 263.36 74.97 263.57 75.04 ;
    RECT 263.36 75.33 263.57 75.4 ;
    RECT 263.36 75.69 263.57 75.76 ;
    RECT 262.9 74.97 263.11 75.04 ;
    RECT 262.9 75.33 263.11 75.4 ;
    RECT 262.9 75.69 263.11 75.76 ;
    RECT 260.04 74.97 260.25 75.04 ;
    RECT 260.04 75.33 260.25 75.4 ;
    RECT 260.04 75.69 260.25 75.76 ;
    RECT 259.58 74.97 259.79 75.04 ;
    RECT 259.58 75.33 259.79 75.4 ;
    RECT 259.58 75.69 259.79 75.76 ;
    RECT 256.72 74.97 256.93 75.04 ;
    RECT 256.72 75.33 256.93 75.4 ;
    RECT 256.72 75.69 256.93 75.76 ;
    RECT 256.26 74.97 256.47 75.04 ;
    RECT 256.26 75.33 256.47 75.4 ;
    RECT 256.26 75.69 256.47 75.76 ;
    RECT 253.4 74.97 253.61 75.04 ;
    RECT 253.4 75.33 253.61 75.4 ;
    RECT 253.4 75.69 253.61 75.76 ;
    RECT 252.94 74.97 253.15 75.04 ;
    RECT 252.94 75.33 253.15 75.4 ;
    RECT 252.94 75.69 253.15 75.76 ;
    RECT 250.08 74.25 250.29 74.32 ;
    RECT 250.08 74.61 250.29 74.68 ;
    RECT 250.08 74.97 250.29 75.04 ;
    RECT 249.62 74.25 249.83 74.32 ;
    RECT 249.62 74.61 249.83 74.68 ;
    RECT 249.62 74.97 249.83 75.04 ;
    RECT 246.76 74.25 246.97 74.32 ;
    RECT 246.76 74.61 246.97 74.68 ;
    RECT 246.76 74.97 246.97 75.04 ;
    RECT 246.3 74.25 246.51 74.32 ;
    RECT 246.3 74.61 246.51 74.68 ;
    RECT 246.3 74.97 246.51 75.04 ;
    RECT 243.44 74.25 243.65 74.32 ;
    RECT 243.44 74.61 243.65 74.68 ;
    RECT 243.44 74.97 243.65 75.04 ;
    RECT 242.98 74.25 243.19 74.32 ;
    RECT 242.98 74.61 243.19 74.68 ;
    RECT 242.98 74.97 243.19 75.04 ;
    RECT 240.12 74.25 240.33 74.32 ;
    RECT 240.12 74.61 240.33 74.68 ;
    RECT 240.12 74.97 240.33 75.04 ;
    RECT 239.66 74.25 239.87 74.32 ;
    RECT 239.66 74.61 239.87 74.68 ;
    RECT 239.66 74.97 239.87 75.04 ;
    RECT 236.8 74.25 237.01 74.32 ;
    RECT 236.8 74.61 237.01 74.68 ;
    RECT 236.8 74.97 237.01 75.04 ;
    RECT 236.34 74.25 236.55 74.32 ;
    RECT 236.34 74.61 236.55 74.68 ;
    RECT 236.34 74.97 236.55 75.04 ;
    RECT 233.48 74.25 233.69 74.32 ;
    RECT 233.48 74.61 233.69 74.68 ;
    RECT 233.48 74.97 233.69 75.04 ;
    RECT 233.02 74.25 233.23 74.32 ;
    RECT 233.02 74.61 233.23 74.68 ;
    RECT 233.02 74.97 233.23 75.04 ;
    RECT 230.16 74.25 230.37 74.32 ;
    RECT 230.16 74.61 230.37 74.68 ;
    RECT 230.16 74.97 230.37 75.04 ;
    RECT 229.7 74.25 229.91 74.32 ;
    RECT 229.7 74.61 229.91 74.68 ;
    RECT 229.7 74.97 229.91 75.04 ;
    RECT 226.84 74.25 227.05 74.32 ;
    RECT 226.84 74.61 227.05 74.68 ;
    RECT 226.84 74.97 227.05 75.04 ;
    RECT 226.38 74.25 226.59 74.32 ;
    RECT 226.38 74.61 226.59 74.68 ;
    RECT 226.38 74.97 226.59 75.04 ;
    RECT 223.52 74.25 223.73 74.32 ;
    RECT 223.52 74.61 223.73 74.68 ;
    RECT 223.52 74.97 223.73 75.04 ;
    RECT 223.06 74.25 223.27 74.32 ;
    RECT 223.06 74.61 223.27 74.68 ;
    RECT 223.06 74.97 223.27 75.04 ;
    RECT 220.2 74.25 220.41 74.32 ;
    RECT 220.2 74.61 220.41 74.68 ;
    RECT 220.2 74.97 220.41 75.04 ;
    RECT 219.74 74.25 219.95 74.32 ;
    RECT 219.74 74.61 219.95 74.68 ;
    RECT 219.74 74.97 219.95 75.04 ;
    RECT 216.88 74.25 217.09 74.32 ;
    RECT 216.88 74.61 217.09 74.68 ;
    RECT 216.88 74.97 217.09 75.04 ;
    RECT 216.42 74.25 216.63 74.32 ;
    RECT 216.42 74.61 216.63 74.68 ;
    RECT 216.42 74.97 216.63 75.04 ;
    RECT 267.91 74.61 267.98 74.68 ;
    RECT 180.36 74.25 180.57 74.32 ;
    RECT 180.36 74.61 180.57 74.68 ;
    RECT 180.36 74.97 180.57 75.04 ;
    RECT 179.9 74.25 180.11 74.32 ;
    RECT 179.9 74.61 180.11 74.68 ;
    RECT 179.9 74.97 180.11 75.04 ;
    RECT 177.04 74.25 177.25 74.32 ;
    RECT 177.04 74.61 177.25 74.68 ;
    RECT 177.04 74.97 177.25 75.04 ;
    RECT 176.58 74.25 176.79 74.32 ;
    RECT 176.58 74.61 176.79 74.68 ;
    RECT 176.58 74.97 176.79 75.04 ;
    RECT 173.72 74.25 173.93 74.32 ;
    RECT 173.72 74.61 173.93 74.68 ;
    RECT 173.72 74.97 173.93 75.04 ;
    RECT 173.26 74.25 173.47 74.32 ;
    RECT 173.26 74.61 173.47 74.68 ;
    RECT 173.26 74.97 173.47 75.04 ;
    RECT 170.4 74.25 170.61 74.32 ;
    RECT 170.4 74.61 170.61 74.68 ;
    RECT 170.4 74.97 170.61 75.04 ;
    RECT 169.94 74.25 170.15 74.32 ;
    RECT 169.94 74.61 170.15 74.68 ;
    RECT 169.94 74.97 170.15 75.04 ;
    RECT 167.08 74.25 167.29 74.32 ;
    RECT 167.08 74.61 167.29 74.68 ;
    RECT 167.08 74.97 167.29 75.04 ;
    RECT 166.62 74.25 166.83 74.32 ;
    RECT 166.62 74.61 166.83 74.68 ;
    RECT 166.62 74.97 166.83 75.04 ;
    RECT 163.76 74.25 163.97 74.32 ;
    RECT 163.76 74.61 163.97 74.68 ;
    RECT 163.76 74.97 163.97 75.04 ;
    RECT 163.3 74.25 163.51 74.32 ;
    RECT 163.3 74.61 163.51 74.68 ;
    RECT 163.3 74.97 163.51 75.04 ;
    RECT 160.44 74.25 160.65 74.32 ;
    RECT 160.44 74.61 160.65 74.68 ;
    RECT 160.44 74.97 160.65 75.04 ;
    RECT 159.98 74.25 160.19 74.32 ;
    RECT 159.98 74.61 160.19 74.68 ;
    RECT 159.98 74.97 160.19 75.04 ;
    RECT 157.12 74.25 157.33 74.32 ;
    RECT 157.12 74.61 157.33 74.68 ;
    RECT 157.12 74.97 157.33 75.04 ;
    RECT 156.66 74.25 156.87 74.32 ;
    RECT 156.66 74.61 156.87 74.68 ;
    RECT 156.66 74.97 156.87 75.04 ;
    RECT 153.8 74.25 154.01 74.32 ;
    RECT 153.8 74.61 154.01 74.68 ;
    RECT 153.8 74.97 154.01 75.04 ;
    RECT 153.34 74.25 153.55 74.32 ;
    RECT 153.34 74.61 153.55 74.68 ;
    RECT 153.34 74.97 153.55 75.04 ;
    RECT 150.48 74.25 150.69 74.32 ;
    RECT 150.48 74.61 150.69 74.68 ;
    RECT 150.48 74.97 150.69 75.04 ;
    RECT 150.02 74.25 150.23 74.32 ;
    RECT 150.02 74.61 150.23 74.68 ;
    RECT 150.02 74.97 150.23 75.04 ;
    RECT 213.56 74.25 213.77 74.32 ;
    RECT 213.56 74.61 213.77 74.68 ;
    RECT 213.56 74.97 213.77 75.04 ;
    RECT 213.1 74.25 213.31 74.32 ;
    RECT 213.1 74.61 213.31 74.68 ;
    RECT 213.1 74.97 213.31 75.04 ;
    RECT 210.24 74.25 210.45 74.32 ;
    RECT 210.24 74.61 210.45 74.68 ;
    RECT 210.24 74.97 210.45 75.04 ;
    RECT 209.78 74.25 209.99 74.32 ;
    RECT 209.78 74.61 209.99 74.68 ;
    RECT 209.78 74.97 209.99 75.04 ;
    RECT 206.92 74.25 207.13 74.32 ;
    RECT 206.92 74.61 207.13 74.68 ;
    RECT 206.92 74.97 207.13 75.04 ;
    RECT 206.46 74.25 206.67 74.32 ;
    RECT 206.46 74.61 206.67 74.68 ;
    RECT 206.46 74.97 206.67 75.04 ;
    RECT 203.6 74.25 203.81 74.32 ;
    RECT 203.6 74.61 203.81 74.68 ;
    RECT 203.6 74.97 203.81 75.04 ;
    RECT 203.14 74.25 203.35 74.32 ;
    RECT 203.14 74.61 203.35 74.68 ;
    RECT 203.14 74.97 203.35 75.04 ;
    RECT 200.28 74.25 200.49 74.32 ;
    RECT 200.28 74.61 200.49 74.68 ;
    RECT 200.28 74.97 200.49 75.04 ;
    RECT 199.82 74.25 200.03 74.32 ;
    RECT 199.82 74.61 200.03 74.68 ;
    RECT 199.82 74.97 200.03 75.04 ;
    RECT 196.96 74.25 197.17 74.32 ;
    RECT 196.96 74.61 197.17 74.68 ;
    RECT 196.96 74.97 197.17 75.04 ;
    RECT 196.5 74.25 196.71 74.32 ;
    RECT 196.5 74.61 196.71 74.68 ;
    RECT 196.5 74.97 196.71 75.04 ;
    RECT 193.64 74.25 193.85 74.32 ;
    RECT 193.64 74.61 193.85 74.68 ;
    RECT 193.64 74.97 193.85 75.04 ;
    RECT 193.18 74.25 193.39 74.32 ;
    RECT 193.18 74.61 193.39 74.68 ;
    RECT 193.18 74.97 193.39 75.04 ;
    RECT 190.32 74.25 190.53 74.32 ;
    RECT 190.32 74.61 190.53 74.68 ;
    RECT 190.32 74.97 190.53 75.04 ;
    RECT 189.86 74.25 190.07 74.32 ;
    RECT 189.86 74.61 190.07 74.68 ;
    RECT 189.86 74.97 190.07 75.04 ;
    RECT 187.0 74.25 187.21 74.32 ;
    RECT 187.0 74.61 187.21 74.68 ;
    RECT 187.0 74.97 187.21 75.04 ;
    RECT 186.54 74.25 186.75 74.32 ;
    RECT 186.54 74.61 186.75 74.68 ;
    RECT 186.54 74.97 186.75 75.04 ;
    RECT 183.68 74.25 183.89 74.32 ;
    RECT 183.68 74.61 183.89 74.68 ;
    RECT 183.68 74.97 183.89 75.04 ;
    RECT 183.22 74.25 183.43 74.32 ;
    RECT 183.22 74.61 183.43 74.68 ;
    RECT 183.22 74.97 183.43 75.04 ;
    RECT 147.485 74.61 147.555 74.68 ;
    RECT 266.68 74.25 266.89 74.32 ;
    RECT 266.68 74.61 266.89 74.68 ;
    RECT 266.68 74.97 266.89 75.04 ;
    RECT 266.22 74.25 266.43 74.32 ;
    RECT 266.22 74.61 266.43 74.68 ;
    RECT 266.22 74.97 266.43 75.04 ;
    RECT 263.36 74.25 263.57 74.32 ;
    RECT 263.36 74.61 263.57 74.68 ;
    RECT 263.36 74.97 263.57 75.04 ;
    RECT 262.9 74.25 263.11 74.32 ;
    RECT 262.9 74.61 263.11 74.68 ;
    RECT 262.9 74.97 263.11 75.04 ;
    RECT 260.04 74.25 260.25 74.32 ;
    RECT 260.04 74.61 260.25 74.68 ;
    RECT 260.04 74.97 260.25 75.04 ;
    RECT 259.58 74.25 259.79 74.32 ;
    RECT 259.58 74.61 259.79 74.68 ;
    RECT 259.58 74.97 259.79 75.04 ;
    RECT 256.72 74.25 256.93 74.32 ;
    RECT 256.72 74.61 256.93 74.68 ;
    RECT 256.72 74.97 256.93 75.04 ;
    RECT 256.26 74.25 256.47 74.32 ;
    RECT 256.26 74.61 256.47 74.68 ;
    RECT 256.26 74.97 256.47 75.04 ;
    RECT 253.4 74.25 253.61 74.32 ;
    RECT 253.4 74.61 253.61 74.68 ;
    RECT 253.4 74.97 253.61 75.04 ;
    RECT 252.94 74.25 253.15 74.32 ;
    RECT 252.94 74.61 253.15 74.68 ;
    RECT 252.94 74.97 253.15 75.04 ;
    RECT 250.08 73.53 250.29 73.6 ;
    RECT 250.08 73.89 250.29 73.96 ;
    RECT 250.08 74.25 250.29 74.32 ;
    RECT 249.62 73.53 249.83 73.6 ;
    RECT 249.62 73.89 249.83 73.96 ;
    RECT 249.62 74.25 249.83 74.32 ;
    RECT 246.76 73.53 246.97 73.6 ;
    RECT 246.76 73.89 246.97 73.96 ;
    RECT 246.76 74.25 246.97 74.32 ;
    RECT 246.3 73.53 246.51 73.6 ;
    RECT 246.3 73.89 246.51 73.96 ;
    RECT 246.3 74.25 246.51 74.32 ;
    RECT 243.44 73.53 243.65 73.6 ;
    RECT 243.44 73.89 243.65 73.96 ;
    RECT 243.44 74.25 243.65 74.32 ;
    RECT 242.98 73.53 243.19 73.6 ;
    RECT 242.98 73.89 243.19 73.96 ;
    RECT 242.98 74.25 243.19 74.32 ;
    RECT 240.12 73.53 240.33 73.6 ;
    RECT 240.12 73.89 240.33 73.96 ;
    RECT 240.12 74.25 240.33 74.32 ;
    RECT 239.66 73.53 239.87 73.6 ;
    RECT 239.66 73.89 239.87 73.96 ;
    RECT 239.66 74.25 239.87 74.32 ;
    RECT 236.8 73.53 237.01 73.6 ;
    RECT 236.8 73.89 237.01 73.96 ;
    RECT 236.8 74.25 237.01 74.32 ;
    RECT 236.34 73.53 236.55 73.6 ;
    RECT 236.34 73.89 236.55 73.96 ;
    RECT 236.34 74.25 236.55 74.32 ;
    RECT 233.48 73.53 233.69 73.6 ;
    RECT 233.48 73.89 233.69 73.96 ;
    RECT 233.48 74.25 233.69 74.32 ;
    RECT 233.02 73.53 233.23 73.6 ;
    RECT 233.02 73.89 233.23 73.96 ;
    RECT 233.02 74.25 233.23 74.32 ;
    RECT 230.16 73.53 230.37 73.6 ;
    RECT 230.16 73.89 230.37 73.96 ;
    RECT 230.16 74.25 230.37 74.32 ;
    RECT 229.7 73.53 229.91 73.6 ;
    RECT 229.7 73.89 229.91 73.96 ;
    RECT 229.7 74.25 229.91 74.32 ;
    RECT 226.84 73.53 227.05 73.6 ;
    RECT 226.84 73.89 227.05 73.96 ;
    RECT 226.84 74.25 227.05 74.32 ;
    RECT 226.38 73.53 226.59 73.6 ;
    RECT 226.38 73.89 226.59 73.96 ;
    RECT 226.38 74.25 226.59 74.32 ;
    RECT 223.52 73.53 223.73 73.6 ;
    RECT 223.52 73.89 223.73 73.96 ;
    RECT 223.52 74.25 223.73 74.32 ;
    RECT 223.06 73.53 223.27 73.6 ;
    RECT 223.06 73.89 223.27 73.96 ;
    RECT 223.06 74.25 223.27 74.32 ;
    RECT 220.2 73.53 220.41 73.6 ;
    RECT 220.2 73.89 220.41 73.96 ;
    RECT 220.2 74.25 220.41 74.32 ;
    RECT 219.74 73.53 219.95 73.6 ;
    RECT 219.74 73.89 219.95 73.96 ;
    RECT 219.74 74.25 219.95 74.32 ;
    RECT 216.88 73.53 217.09 73.6 ;
    RECT 216.88 73.89 217.09 73.96 ;
    RECT 216.88 74.25 217.09 74.32 ;
    RECT 216.42 73.53 216.63 73.6 ;
    RECT 216.42 73.89 216.63 73.96 ;
    RECT 216.42 74.25 216.63 74.32 ;
    RECT 267.91 73.89 267.98 73.96 ;
    RECT 180.36 73.53 180.57 73.6 ;
    RECT 180.36 73.89 180.57 73.96 ;
    RECT 180.36 74.25 180.57 74.32 ;
    RECT 179.9 73.53 180.11 73.6 ;
    RECT 179.9 73.89 180.11 73.96 ;
    RECT 179.9 74.25 180.11 74.32 ;
    RECT 177.04 73.53 177.25 73.6 ;
    RECT 177.04 73.89 177.25 73.96 ;
    RECT 177.04 74.25 177.25 74.32 ;
    RECT 176.58 73.53 176.79 73.6 ;
    RECT 176.58 73.89 176.79 73.96 ;
    RECT 176.58 74.25 176.79 74.32 ;
    RECT 173.72 73.53 173.93 73.6 ;
    RECT 173.72 73.89 173.93 73.96 ;
    RECT 173.72 74.25 173.93 74.32 ;
    RECT 173.26 73.53 173.47 73.6 ;
    RECT 173.26 73.89 173.47 73.96 ;
    RECT 173.26 74.25 173.47 74.32 ;
    RECT 170.4 73.53 170.61 73.6 ;
    RECT 170.4 73.89 170.61 73.96 ;
    RECT 170.4 74.25 170.61 74.32 ;
    RECT 169.94 73.53 170.15 73.6 ;
    RECT 169.94 73.89 170.15 73.96 ;
    RECT 169.94 74.25 170.15 74.32 ;
    RECT 167.08 73.53 167.29 73.6 ;
    RECT 167.08 73.89 167.29 73.96 ;
    RECT 167.08 74.25 167.29 74.32 ;
    RECT 166.62 73.53 166.83 73.6 ;
    RECT 166.62 73.89 166.83 73.96 ;
    RECT 166.62 74.25 166.83 74.32 ;
    RECT 163.76 73.53 163.97 73.6 ;
    RECT 163.76 73.89 163.97 73.96 ;
    RECT 163.76 74.25 163.97 74.32 ;
    RECT 163.3 73.53 163.51 73.6 ;
    RECT 163.3 73.89 163.51 73.96 ;
    RECT 163.3 74.25 163.51 74.32 ;
    RECT 160.44 73.53 160.65 73.6 ;
    RECT 160.44 73.89 160.65 73.96 ;
    RECT 160.44 74.25 160.65 74.32 ;
    RECT 159.98 73.53 160.19 73.6 ;
    RECT 159.98 73.89 160.19 73.96 ;
    RECT 159.98 74.25 160.19 74.32 ;
    RECT 157.12 73.53 157.33 73.6 ;
    RECT 157.12 73.89 157.33 73.96 ;
    RECT 157.12 74.25 157.33 74.32 ;
    RECT 156.66 73.53 156.87 73.6 ;
    RECT 156.66 73.89 156.87 73.96 ;
    RECT 156.66 74.25 156.87 74.32 ;
    RECT 153.8 73.53 154.01 73.6 ;
    RECT 153.8 73.89 154.01 73.96 ;
    RECT 153.8 74.25 154.01 74.32 ;
    RECT 153.34 73.53 153.55 73.6 ;
    RECT 153.34 73.89 153.55 73.96 ;
    RECT 153.34 74.25 153.55 74.32 ;
    RECT 150.48 73.53 150.69 73.6 ;
    RECT 150.48 73.89 150.69 73.96 ;
    RECT 150.48 74.25 150.69 74.32 ;
    RECT 150.02 73.53 150.23 73.6 ;
    RECT 150.02 73.89 150.23 73.96 ;
    RECT 150.02 74.25 150.23 74.32 ;
    RECT 213.56 73.53 213.77 73.6 ;
    RECT 213.56 73.89 213.77 73.96 ;
    RECT 213.56 74.25 213.77 74.32 ;
    RECT 213.1 73.53 213.31 73.6 ;
    RECT 213.1 73.89 213.31 73.96 ;
    RECT 213.1 74.25 213.31 74.32 ;
    RECT 210.24 73.53 210.45 73.6 ;
    RECT 210.24 73.89 210.45 73.96 ;
    RECT 210.24 74.25 210.45 74.32 ;
    RECT 209.78 73.53 209.99 73.6 ;
    RECT 209.78 73.89 209.99 73.96 ;
    RECT 209.78 74.25 209.99 74.32 ;
    RECT 206.92 73.53 207.13 73.6 ;
    RECT 206.92 73.89 207.13 73.96 ;
    RECT 206.92 74.25 207.13 74.32 ;
    RECT 206.46 73.53 206.67 73.6 ;
    RECT 206.46 73.89 206.67 73.96 ;
    RECT 206.46 74.25 206.67 74.32 ;
    RECT 203.6 73.53 203.81 73.6 ;
    RECT 203.6 73.89 203.81 73.96 ;
    RECT 203.6 74.25 203.81 74.32 ;
    RECT 203.14 73.53 203.35 73.6 ;
    RECT 203.14 73.89 203.35 73.96 ;
    RECT 203.14 74.25 203.35 74.32 ;
    RECT 200.28 73.53 200.49 73.6 ;
    RECT 200.28 73.89 200.49 73.96 ;
    RECT 200.28 74.25 200.49 74.32 ;
    RECT 199.82 73.53 200.03 73.6 ;
    RECT 199.82 73.89 200.03 73.96 ;
    RECT 199.82 74.25 200.03 74.32 ;
    RECT 196.96 73.53 197.17 73.6 ;
    RECT 196.96 73.89 197.17 73.96 ;
    RECT 196.96 74.25 197.17 74.32 ;
    RECT 196.5 73.53 196.71 73.6 ;
    RECT 196.5 73.89 196.71 73.96 ;
    RECT 196.5 74.25 196.71 74.32 ;
    RECT 193.64 73.53 193.85 73.6 ;
    RECT 193.64 73.89 193.85 73.96 ;
    RECT 193.64 74.25 193.85 74.32 ;
    RECT 193.18 73.53 193.39 73.6 ;
    RECT 193.18 73.89 193.39 73.96 ;
    RECT 193.18 74.25 193.39 74.32 ;
    RECT 190.32 73.53 190.53 73.6 ;
    RECT 190.32 73.89 190.53 73.96 ;
    RECT 190.32 74.25 190.53 74.32 ;
    RECT 189.86 73.53 190.07 73.6 ;
    RECT 189.86 73.89 190.07 73.96 ;
    RECT 189.86 74.25 190.07 74.32 ;
    RECT 187.0 73.53 187.21 73.6 ;
    RECT 187.0 73.89 187.21 73.96 ;
    RECT 187.0 74.25 187.21 74.32 ;
    RECT 186.54 73.53 186.75 73.6 ;
    RECT 186.54 73.89 186.75 73.96 ;
    RECT 186.54 74.25 186.75 74.32 ;
    RECT 183.68 73.53 183.89 73.6 ;
    RECT 183.68 73.89 183.89 73.96 ;
    RECT 183.68 74.25 183.89 74.32 ;
    RECT 183.22 73.53 183.43 73.6 ;
    RECT 183.22 73.89 183.43 73.96 ;
    RECT 183.22 74.25 183.43 74.32 ;
    RECT 147.485 73.89 147.555 73.96 ;
    RECT 266.68 73.53 266.89 73.6 ;
    RECT 266.68 73.89 266.89 73.96 ;
    RECT 266.68 74.25 266.89 74.32 ;
    RECT 266.22 73.53 266.43 73.6 ;
    RECT 266.22 73.89 266.43 73.96 ;
    RECT 266.22 74.25 266.43 74.32 ;
    RECT 263.36 73.53 263.57 73.6 ;
    RECT 263.36 73.89 263.57 73.96 ;
    RECT 263.36 74.25 263.57 74.32 ;
    RECT 262.9 73.53 263.11 73.6 ;
    RECT 262.9 73.89 263.11 73.96 ;
    RECT 262.9 74.25 263.11 74.32 ;
    RECT 260.04 73.53 260.25 73.6 ;
    RECT 260.04 73.89 260.25 73.96 ;
    RECT 260.04 74.25 260.25 74.32 ;
    RECT 259.58 73.53 259.79 73.6 ;
    RECT 259.58 73.89 259.79 73.96 ;
    RECT 259.58 74.25 259.79 74.32 ;
    RECT 256.72 73.53 256.93 73.6 ;
    RECT 256.72 73.89 256.93 73.96 ;
    RECT 256.72 74.25 256.93 74.32 ;
    RECT 256.26 73.53 256.47 73.6 ;
    RECT 256.26 73.89 256.47 73.96 ;
    RECT 256.26 74.25 256.47 74.32 ;
    RECT 253.4 73.53 253.61 73.6 ;
    RECT 253.4 73.89 253.61 73.96 ;
    RECT 253.4 74.25 253.61 74.32 ;
    RECT 252.94 73.53 253.15 73.6 ;
    RECT 252.94 73.89 253.15 73.96 ;
    RECT 252.94 74.25 253.15 74.32 ;
    RECT 250.08 72.81 250.29 72.88 ;
    RECT 250.08 73.17 250.29 73.24 ;
    RECT 250.08 73.53 250.29 73.6 ;
    RECT 249.62 72.81 249.83 72.88 ;
    RECT 249.62 73.17 249.83 73.24 ;
    RECT 249.62 73.53 249.83 73.6 ;
    RECT 246.76 72.81 246.97 72.88 ;
    RECT 246.76 73.17 246.97 73.24 ;
    RECT 246.76 73.53 246.97 73.6 ;
    RECT 246.3 72.81 246.51 72.88 ;
    RECT 246.3 73.17 246.51 73.24 ;
    RECT 246.3 73.53 246.51 73.6 ;
    RECT 243.44 72.81 243.65 72.88 ;
    RECT 243.44 73.17 243.65 73.24 ;
    RECT 243.44 73.53 243.65 73.6 ;
    RECT 242.98 72.81 243.19 72.88 ;
    RECT 242.98 73.17 243.19 73.24 ;
    RECT 242.98 73.53 243.19 73.6 ;
    RECT 240.12 72.81 240.33 72.88 ;
    RECT 240.12 73.17 240.33 73.24 ;
    RECT 240.12 73.53 240.33 73.6 ;
    RECT 239.66 72.81 239.87 72.88 ;
    RECT 239.66 73.17 239.87 73.24 ;
    RECT 239.66 73.53 239.87 73.6 ;
    RECT 236.8 72.81 237.01 72.88 ;
    RECT 236.8 73.17 237.01 73.24 ;
    RECT 236.8 73.53 237.01 73.6 ;
    RECT 236.34 72.81 236.55 72.88 ;
    RECT 236.34 73.17 236.55 73.24 ;
    RECT 236.34 73.53 236.55 73.6 ;
    RECT 233.48 72.81 233.69 72.88 ;
    RECT 233.48 73.17 233.69 73.24 ;
    RECT 233.48 73.53 233.69 73.6 ;
    RECT 233.02 72.81 233.23 72.88 ;
    RECT 233.02 73.17 233.23 73.24 ;
    RECT 233.02 73.53 233.23 73.6 ;
    RECT 230.16 72.81 230.37 72.88 ;
    RECT 230.16 73.17 230.37 73.24 ;
    RECT 230.16 73.53 230.37 73.6 ;
    RECT 229.7 72.81 229.91 72.88 ;
    RECT 229.7 73.17 229.91 73.24 ;
    RECT 229.7 73.53 229.91 73.6 ;
    RECT 226.84 72.81 227.05 72.88 ;
    RECT 226.84 73.17 227.05 73.24 ;
    RECT 226.84 73.53 227.05 73.6 ;
    RECT 226.38 72.81 226.59 72.88 ;
    RECT 226.38 73.17 226.59 73.24 ;
    RECT 226.38 73.53 226.59 73.6 ;
    RECT 223.52 72.81 223.73 72.88 ;
    RECT 223.52 73.17 223.73 73.24 ;
    RECT 223.52 73.53 223.73 73.6 ;
    RECT 223.06 72.81 223.27 72.88 ;
    RECT 223.06 73.17 223.27 73.24 ;
    RECT 223.06 73.53 223.27 73.6 ;
    RECT 220.2 72.81 220.41 72.88 ;
    RECT 220.2 73.17 220.41 73.24 ;
    RECT 220.2 73.53 220.41 73.6 ;
    RECT 219.74 72.81 219.95 72.88 ;
    RECT 219.74 73.17 219.95 73.24 ;
    RECT 219.74 73.53 219.95 73.6 ;
    RECT 216.88 72.81 217.09 72.88 ;
    RECT 216.88 73.17 217.09 73.24 ;
    RECT 216.88 73.53 217.09 73.6 ;
    RECT 216.42 72.81 216.63 72.88 ;
    RECT 216.42 73.17 216.63 73.24 ;
    RECT 216.42 73.53 216.63 73.6 ;
    RECT 267.91 73.17 267.98 73.24 ;
    RECT 180.36 72.81 180.57 72.88 ;
    RECT 180.36 73.17 180.57 73.24 ;
    RECT 180.36 73.53 180.57 73.6 ;
    RECT 179.9 72.81 180.11 72.88 ;
    RECT 179.9 73.17 180.11 73.24 ;
    RECT 179.9 73.53 180.11 73.6 ;
    RECT 177.04 72.81 177.25 72.88 ;
    RECT 177.04 73.17 177.25 73.24 ;
    RECT 177.04 73.53 177.25 73.6 ;
    RECT 176.58 72.81 176.79 72.88 ;
    RECT 176.58 73.17 176.79 73.24 ;
    RECT 176.58 73.53 176.79 73.6 ;
    RECT 173.72 72.81 173.93 72.88 ;
    RECT 173.72 73.17 173.93 73.24 ;
    RECT 173.72 73.53 173.93 73.6 ;
    RECT 173.26 72.81 173.47 72.88 ;
    RECT 173.26 73.17 173.47 73.24 ;
    RECT 173.26 73.53 173.47 73.6 ;
    RECT 170.4 72.81 170.61 72.88 ;
    RECT 170.4 73.17 170.61 73.24 ;
    RECT 170.4 73.53 170.61 73.6 ;
    RECT 169.94 72.81 170.15 72.88 ;
    RECT 169.94 73.17 170.15 73.24 ;
    RECT 169.94 73.53 170.15 73.6 ;
    RECT 167.08 72.81 167.29 72.88 ;
    RECT 167.08 73.17 167.29 73.24 ;
    RECT 167.08 73.53 167.29 73.6 ;
    RECT 166.62 72.81 166.83 72.88 ;
    RECT 166.62 73.17 166.83 73.24 ;
    RECT 166.62 73.53 166.83 73.6 ;
    RECT 163.76 72.81 163.97 72.88 ;
    RECT 163.76 73.17 163.97 73.24 ;
    RECT 163.76 73.53 163.97 73.6 ;
    RECT 163.3 72.81 163.51 72.88 ;
    RECT 163.3 73.17 163.51 73.24 ;
    RECT 163.3 73.53 163.51 73.6 ;
    RECT 160.44 72.81 160.65 72.88 ;
    RECT 160.44 73.17 160.65 73.24 ;
    RECT 160.44 73.53 160.65 73.6 ;
    RECT 159.98 72.81 160.19 72.88 ;
    RECT 159.98 73.17 160.19 73.24 ;
    RECT 159.98 73.53 160.19 73.6 ;
    RECT 157.12 72.81 157.33 72.88 ;
    RECT 157.12 73.17 157.33 73.24 ;
    RECT 157.12 73.53 157.33 73.6 ;
    RECT 156.66 72.81 156.87 72.88 ;
    RECT 156.66 73.17 156.87 73.24 ;
    RECT 156.66 73.53 156.87 73.6 ;
    RECT 153.8 72.81 154.01 72.88 ;
    RECT 153.8 73.17 154.01 73.24 ;
    RECT 153.8 73.53 154.01 73.6 ;
    RECT 153.34 72.81 153.55 72.88 ;
    RECT 153.34 73.17 153.55 73.24 ;
    RECT 153.34 73.53 153.55 73.6 ;
    RECT 150.48 72.81 150.69 72.88 ;
    RECT 150.48 73.17 150.69 73.24 ;
    RECT 150.48 73.53 150.69 73.6 ;
    RECT 150.02 72.81 150.23 72.88 ;
    RECT 150.02 73.17 150.23 73.24 ;
    RECT 150.02 73.53 150.23 73.6 ;
    RECT 213.56 72.81 213.77 72.88 ;
    RECT 213.56 73.17 213.77 73.24 ;
    RECT 213.56 73.53 213.77 73.6 ;
    RECT 213.1 72.81 213.31 72.88 ;
    RECT 213.1 73.17 213.31 73.24 ;
    RECT 213.1 73.53 213.31 73.6 ;
    RECT 210.24 72.81 210.45 72.88 ;
    RECT 210.24 73.17 210.45 73.24 ;
    RECT 210.24 73.53 210.45 73.6 ;
    RECT 209.78 72.81 209.99 72.88 ;
    RECT 209.78 73.17 209.99 73.24 ;
    RECT 209.78 73.53 209.99 73.6 ;
    RECT 206.92 72.81 207.13 72.88 ;
    RECT 206.92 73.17 207.13 73.24 ;
    RECT 206.92 73.53 207.13 73.6 ;
    RECT 206.46 72.81 206.67 72.88 ;
    RECT 206.46 73.17 206.67 73.24 ;
    RECT 206.46 73.53 206.67 73.6 ;
    RECT 203.6 72.81 203.81 72.88 ;
    RECT 203.6 73.17 203.81 73.24 ;
    RECT 203.6 73.53 203.81 73.6 ;
    RECT 203.14 72.81 203.35 72.88 ;
    RECT 203.14 73.17 203.35 73.24 ;
    RECT 203.14 73.53 203.35 73.6 ;
    RECT 200.28 72.81 200.49 72.88 ;
    RECT 200.28 73.17 200.49 73.24 ;
    RECT 200.28 73.53 200.49 73.6 ;
    RECT 199.82 72.81 200.03 72.88 ;
    RECT 199.82 73.17 200.03 73.24 ;
    RECT 199.82 73.53 200.03 73.6 ;
    RECT 196.96 72.81 197.17 72.88 ;
    RECT 196.96 73.17 197.17 73.24 ;
    RECT 196.96 73.53 197.17 73.6 ;
    RECT 196.5 72.81 196.71 72.88 ;
    RECT 196.5 73.17 196.71 73.24 ;
    RECT 196.5 73.53 196.71 73.6 ;
    RECT 193.64 72.81 193.85 72.88 ;
    RECT 193.64 73.17 193.85 73.24 ;
    RECT 193.64 73.53 193.85 73.6 ;
    RECT 193.18 72.81 193.39 72.88 ;
    RECT 193.18 73.17 193.39 73.24 ;
    RECT 193.18 73.53 193.39 73.6 ;
    RECT 190.32 72.81 190.53 72.88 ;
    RECT 190.32 73.17 190.53 73.24 ;
    RECT 190.32 73.53 190.53 73.6 ;
    RECT 189.86 72.81 190.07 72.88 ;
    RECT 189.86 73.17 190.07 73.24 ;
    RECT 189.86 73.53 190.07 73.6 ;
    RECT 187.0 72.81 187.21 72.88 ;
    RECT 187.0 73.17 187.21 73.24 ;
    RECT 187.0 73.53 187.21 73.6 ;
    RECT 186.54 72.81 186.75 72.88 ;
    RECT 186.54 73.17 186.75 73.24 ;
    RECT 186.54 73.53 186.75 73.6 ;
    RECT 183.68 72.81 183.89 72.88 ;
    RECT 183.68 73.17 183.89 73.24 ;
    RECT 183.68 73.53 183.89 73.6 ;
    RECT 183.22 72.81 183.43 72.88 ;
    RECT 183.22 73.17 183.43 73.24 ;
    RECT 183.22 73.53 183.43 73.6 ;
    RECT 147.485 73.17 147.555 73.24 ;
    RECT 266.68 72.81 266.89 72.88 ;
    RECT 266.68 73.17 266.89 73.24 ;
    RECT 266.68 73.53 266.89 73.6 ;
    RECT 266.22 72.81 266.43 72.88 ;
    RECT 266.22 73.17 266.43 73.24 ;
    RECT 266.22 73.53 266.43 73.6 ;
    RECT 263.36 72.81 263.57 72.88 ;
    RECT 263.36 73.17 263.57 73.24 ;
    RECT 263.36 73.53 263.57 73.6 ;
    RECT 262.9 72.81 263.11 72.88 ;
    RECT 262.9 73.17 263.11 73.24 ;
    RECT 262.9 73.53 263.11 73.6 ;
    RECT 260.04 72.81 260.25 72.88 ;
    RECT 260.04 73.17 260.25 73.24 ;
    RECT 260.04 73.53 260.25 73.6 ;
    RECT 259.58 72.81 259.79 72.88 ;
    RECT 259.58 73.17 259.79 73.24 ;
    RECT 259.58 73.53 259.79 73.6 ;
    RECT 256.72 72.81 256.93 72.88 ;
    RECT 256.72 73.17 256.93 73.24 ;
    RECT 256.72 73.53 256.93 73.6 ;
    RECT 256.26 72.81 256.47 72.88 ;
    RECT 256.26 73.17 256.47 73.24 ;
    RECT 256.26 73.53 256.47 73.6 ;
    RECT 253.4 72.81 253.61 72.88 ;
    RECT 253.4 73.17 253.61 73.24 ;
    RECT 253.4 73.53 253.61 73.6 ;
    RECT 252.94 72.81 253.15 72.88 ;
    RECT 252.94 73.17 253.15 73.24 ;
    RECT 252.94 73.53 253.15 73.6 ;
    RECT 250.08 20.95 250.29 21.02 ;
    RECT 250.08 21.31 250.29 21.38 ;
    RECT 250.08 21.67 250.29 21.74 ;
    RECT 249.62 20.95 249.83 21.02 ;
    RECT 249.62 21.31 249.83 21.38 ;
    RECT 249.62 21.67 249.83 21.74 ;
    RECT 246.76 20.95 246.97 21.02 ;
    RECT 246.76 21.31 246.97 21.38 ;
    RECT 246.76 21.67 246.97 21.74 ;
    RECT 246.3 20.95 246.51 21.02 ;
    RECT 246.3 21.31 246.51 21.38 ;
    RECT 246.3 21.67 246.51 21.74 ;
    RECT 243.44 20.95 243.65 21.02 ;
    RECT 243.44 21.31 243.65 21.38 ;
    RECT 243.44 21.67 243.65 21.74 ;
    RECT 242.98 20.95 243.19 21.02 ;
    RECT 242.98 21.31 243.19 21.38 ;
    RECT 242.98 21.67 243.19 21.74 ;
    RECT 240.12 20.95 240.33 21.02 ;
    RECT 240.12 21.31 240.33 21.38 ;
    RECT 240.12 21.67 240.33 21.74 ;
    RECT 239.66 20.95 239.87 21.02 ;
    RECT 239.66 21.31 239.87 21.38 ;
    RECT 239.66 21.67 239.87 21.74 ;
    RECT 236.8 20.95 237.01 21.02 ;
    RECT 236.8 21.31 237.01 21.38 ;
    RECT 236.8 21.67 237.01 21.74 ;
    RECT 236.34 20.95 236.55 21.02 ;
    RECT 236.34 21.31 236.55 21.38 ;
    RECT 236.34 21.67 236.55 21.74 ;
    RECT 233.48 20.95 233.69 21.02 ;
    RECT 233.48 21.31 233.69 21.38 ;
    RECT 233.48 21.67 233.69 21.74 ;
    RECT 233.02 20.95 233.23 21.02 ;
    RECT 233.02 21.31 233.23 21.38 ;
    RECT 233.02 21.67 233.23 21.74 ;
    RECT 230.16 20.95 230.37 21.02 ;
    RECT 230.16 21.31 230.37 21.38 ;
    RECT 230.16 21.67 230.37 21.74 ;
    RECT 229.7 20.95 229.91 21.02 ;
    RECT 229.7 21.31 229.91 21.38 ;
    RECT 229.7 21.67 229.91 21.74 ;
    RECT 226.84 20.95 227.05 21.02 ;
    RECT 226.84 21.31 227.05 21.38 ;
    RECT 226.84 21.67 227.05 21.74 ;
    RECT 226.38 20.95 226.59 21.02 ;
    RECT 226.38 21.31 226.59 21.38 ;
    RECT 226.38 21.67 226.59 21.74 ;
    RECT 223.52 20.95 223.73 21.02 ;
    RECT 223.52 21.31 223.73 21.38 ;
    RECT 223.52 21.67 223.73 21.74 ;
    RECT 223.06 20.95 223.27 21.02 ;
    RECT 223.06 21.31 223.27 21.38 ;
    RECT 223.06 21.67 223.27 21.74 ;
    RECT 220.2 20.95 220.41 21.02 ;
    RECT 220.2 21.31 220.41 21.38 ;
    RECT 220.2 21.67 220.41 21.74 ;
    RECT 219.74 20.95 219.95 21.02 ;
    RECT 219.74 21.31 219.95 21.38 ;
    RECT 219.74 21.67 219.95 21.74 ;
    RECT 216.88 20.95 217.09 21.02 ;
    RECT 216.88 21.31 217.09 21.38 ;
    RECT 216.88 21.67 217.09 21.74 ;
    RECT 216.42 20.95 216.63 21.02 ;
    RECT 216.42 21.31 216.63 21.38 ;
    RECT 216.42 21.67 216.63 21.74 ;
    RECT 267.91 21.31 267.98 21.38 ;
    RECT 180.36 20.95 180.57 21.02 ;
    RECT 180.36 21.31 180.57 21.38 ;
    RECT 180.36 21.67 180.57 21.74 ;
    RECT 179.9 20.95 180.11 21.02 ;
    RECT 179.9 21.31 180.11 21.38 ;
    RECT 179.9 21.67 180.11 21.74 ;
    RECT 177.04 20.95 177.25 21.02 ;
    RECT 177.04 21.31 177.25 21.38 ;
    RECT 177.04 21.67 177.25 21.74 ;
    RECT 176.58 20.95 176.79 21.02 ;
    RECT 176.58 21.31 176.79 21.38 ;
    RECT 176.58 21.67 176.79 21.74 ;
    RECT 173.72 20.95 173.93 21.02 ;
    RECT 173.72 21.31 173.93 21.38 ;
    RECT 173.72 21.67 173.93 21.74 ;
    RECT 173.26 20.95 173.47 21.02 ;
    RECT 173.26 21.31 173.47 21.38 ;
    RECT 173.26 21.67 173.47 21.74 ;
    RECT 170.4 20.95 170.61 21.02 ;
    RECT 170.4 21.31 170.61 21.38 ;
    RECT 170.4 21.67 170.61 21.74 ;
    RECT 169.94 20.95 170.15 21.02 ;
    RECT 169.94 21.31 170.15 21.38 ;
    RECT 169.94 21.67 170.15 21.74 ;
    RECT 167.08 20.95 167.29 21.02 ;
    RECT 167.08 21.31 167.29 21.38 ;
    RECT 167.08 21.67 167.29 21.74 ;
    RECT 166.62 20.95 166.83 21.02 ;
    RECT 166.62 21.31 166.83 21.38 ;
    RECT 166.62 21.67 166.83 21.74 ;
    RECT 163.76 20.95 163.97 21.02 ;
    RECT 163.76 21.31 163.97 21.38 ;
    RECT 163.76 21.67 163.97 21.74 ;
    RECT 163.3 20.95 163.51 21.02 ;
    RECT 163.3 21.31 163.51 21.38 ;
    RECT 163.3 21.67 163.51 21.74 ;
    RECT 160.44 20.95 160.65 21.02 ;
    RECT 160.44 21.31 160.65 21.38 ;
    RECT 160.44 21.67 160.65 21.74 ;
    RECT 159.98 20.95 160.19 21.02 ;
    RECT 159.98 21.31 160.19 21.38 ;
    RECT 159.98 21.67 160.19 21.74 ;
    RECT 157.12 20.95 157.33 21.02 ;
    RECT 157.12 21.31 157.33 21.38 ;
    RECT 157.12 21.67 157.33 21.74 ;
    RECT 156.66 20.95 156.87 21.02 ;
    RECT 156.66 21.31 156.87 21.38 ;
    RECT 156.66 21.67 156.87 21.74 ;
    RECT 153.8 20.95 154.01 21.02 ;
    RECT 153.8 21.31 154.01 21.38 ;
    RECT 153.8 21.67 154.01 21.74 ;
    RECT 153.34 20.95 153.55 21.02 ;
    RECT 153.34 21.31 153.55 21.38 ;
    RECT 153.34 21.67 153.55 21.74 ;
    RECT 150.48 20.95 150.69 21.02 ;
    RECT 150.48 21.31 150.69 21.38 ;
    RECT 150.48 21.67 150.69 21.74 ;
    RECT 150.02 20.95 150.23 21.02 ;
    RECT 150.02 21.31 150.23 21.38 ;
    RECT 150.02 21.67 150.23 21.74 ;
    RECT 213.56 20.95 213.77 21.02 ;
    RECT 213.56 21.31 213.77 21.38 ;
    RECT 213.56 21.67 213.77 21.74 ;
    RECT 213.1 20.95 213.31 21.02 ;
    RECT 213.1 21.31 213.31 21.38 ;
    RECT 213.1 21.67 213.31 21.74 ;
    RECT 210.24 20.95 210.45 21.02 ;
    RECT 210.24 21.31 210.45 21.38 ;
    RECT 210.24 21.67 210.45 21.74 ;
    RECT 209.78 20.95 209.99 21.02 ;
    RECT 209.78 21.31 209.99 21.38 ;
    RECT 209.78 21.67 209.99 21.74 ;
    RECT 206.92 20.95 207.13 21.02 ;
    RECT 206.92 21.31 207.13 21.38 ;
    RECT 206.92 21.67 207.13 21.74 ;
    RECT 206.46 20.95 206.67 21.02 ;
    RECT 206.46 21.31 206.67 21.38 ;
    RECT 206.46 21.67 206.67 21.74 ;
    RECT 203.6 20.95 203.81 21.02 ;
    RECT 203.6 21.31 203.81 21.38 ;
    RECT 203.6 21.67 203.81 21.74 ;
    RECT 203.14 20.95 203.35 21.02 ;
    RECT 203.14 21.31 203.35 21.38 ;
    RECT 203.14 21.67 203.35 21.74 ;
    RECT 200.28 20.95 200.49 21.02 ;
    RECT 200.28 21.31 200.49 21.38 ;
    RECT 200.28 21.67 200.49 21.74 ;
    RECT 199.82 20.95 200.03 21.02 ;
    RECT 199.82 21.31 200.03 21.38 ;
    RECT 199.82 21.67 200.03 21.74 ;
    RECT 196.96 20.95 197.17 21.02 ;
    RECT 196.96 21.31 197.17 21.38 ;
    RECT 196.96 21.67 197.17 21.74 ;
    RECT 196.5 20.95 196.71 21.02 ;
    RECT 196.5 21.31 196.71 21.38 ;
    RECT 196.5 21.67 196.71 21.74 ;
    RECT 193.64 20.95 193.85 21.02 ;
    RECT 193.64 21.31 193.85 21.38 ;
    RECT 193.64 21.67 193.85 21.74 ;
    RECT 193.18 20.95 193.39 21.02 ;
    RECT 193.18 21.31 193.39 21.38 ;
    RECT 193.18 21.67 193.39 21.74 ;
    RECT 190.32 20.95 190.53 21.02 ;
    RECT 190.32 21.31 190.53 21.38 ;
    RECT 190.32 21.67 190.53 21.74 ;
    RECT 189.86 20.95 190.07 21.02 ;
    RECT 189.86 21.31 190.07 21.38 ;
    RECT 189.86 21.67 190.07 21.74 ;
    RECT 187.0 20.95 187.21 21.02 ;
    RECT 187.0 21.31 187.21 21.38 ;
    RECT 187.0 21.67 187.21 21.74 ;
    RECT 186.54 20.95 186.75 21.02 ;
    RECT 186.54 21.31 186.75 21.38 ;
    RECT 186.54 21.67 186.75 21.74 ;
    RECT 183.68 20.95 183.89 21.02 ;
    RECT 183.68 21.31 183.89 21.38 ;
    RECT 183.68 21.67 183.89 21.74 ;
    RECT 183.22 20.95 183.43 21.02 ;
    RECT 183.22 21.31 183.43 21.38 ;
    RECT 183.22 21.67 183.43 21.74 ;
    RECT 147.485 21.31 147.555 21.38 ;
    RECT 266.68 20.95 266.89 21.02 ;
    RECT 266.68 21.31 266.89 21.38 ;
    RECT 266.68 21.67 266.89 21.74 ;
    RECT 266.22 20.95 266.43 21.02 ;
    RECT 266.22 21.31 266.43 21.38 ;
    RECT 266.22 21.67 266.43 21.74 ;
    RECT 263.36 20.95 263.57 21.02 ;
    RECT 263.36 21.31 263.57 21.38 ;
    RECT 263.36 21.67 263.57 21.74 ;
    RECT 262.9 20.95 263.11 21.02 ;
    RECT 262.9 21.31 263.11 21.38 ;
    RECT 262.9 21.67 263.11 21.74 ;
    RECT 260.04 20.95 260.25 21.02 ;
    RECT 260.04 21.31 260.25 21.38 ;
    RECT 260.04 21.67 260.25 21.74 ;
    RECT 259.58 20.95 259.79 21.02 ;
    RECT 259.58 21.31 259.79 21.38 ;
    RECT 259.58 21.67 259.79 21.74 ;
    RECT 256.72 20.95 256.93 21.02 ;
    RECT 256.72 21.31 256.93 21.38 ;
    RECT 256.72 21.67 256.93 21.74 ;
    RECT 256.26 20.95 256.47 21.02 ;
    RECT 256.26 21.31 256.47 21.38 ;
    RECT 256.26 21.67 256.47 21.74 ;
    RECT 253.4 20.95 253.61 21.02 ;
    RECT 253.4 21.31 253.61 21.38 ;
    RECT 253.4 21.67 253.61 21.74 ;
    RECT 252.94 20.95 253.15 21.02 ;
    RECT 252.94 21.31 253.15 21.38 ;
    RECT 252.94 21.67 253.15 21.74 ;
    RECT 250.08 20.23 250.29 20.3 ;
    RECT 250.08 20.59 250.29 20.66 ;
    RECT 250.08 20.95 250.29 21.02 ;
    RECT 249.62 20.23 249.83 20.3 ;
    RECT 249.62 20.59 249.83 20.66 ;
    RECT 249.62 20.95 249.83 21.02 ;
    RECT 246.76 20.23 246.97 20.3 ;
    RECT 246.76 20.59 246.97 20.66 ;
    RECT 246.76 20.95 246.97 21.02 ;
    RECT 246.3 20.23 246.51 20.3 ;
    RECT 246.3 20.59 246.51 20.66 ;
    RECT 246.3 20.95 246.51 21.02 ;
    RECT 243.44 20.23 243.65 20.3 ;
    RECT 243.44 20.59 243.65 20.66 ;
    RECT 243.44 20.95 243.65 21.02 ;
    RECT 242.98 20.23 243.19 20.3 ;
    RECT 242.98 20.59 243.19 20.66 ;
    RECT 242.98 20.95 243.19 21.02 ;
    RECT 240.12 20.23 240.33 20.3 ;
    RECT 240.12 20.59 240.33 20.66 ;
    RECT 240.12 20.95 240.33 21.02 ;
    RECT 239.66 20.23 239.87 20.3 ;
    RECT 239.66 20.59 239.87 20.66 ;
    RECT 239.66 20.95 239.87 21.02 ;
    RECT 236.8 20.23 237.01 20.3 ;
    RECT 236.8 20.59 237.01 20.66 ;
    RECT 236.8 20.95 237.01 21.02 ;
    RECT 236.34 20.23 236.55 20.3 ;
    RECT 236.34 20.59 236.55 20.66 ;
    RECT 236.34 20.95 236.55 21.02 ;
    RECT 233.48 20.23 233.69 20.3 ;
    RECT 233.48 20.59 233.69 20.66 ;
    RECT 233.48 20.95 233.69 21.02 ;
    RECT 233.02 20.23 233.23 20.3 ;
    RECT 233.02 20.59 233.23 20.66 ;
    RECT 233.02 20.95 233.23 21.02 ;
    RECT 230.16 20.23 230.37 20.3 ;
    RECT 230.16 20.59 230.37 20.66 ;
    RECT 230.16 20.95 230.37 21.02 ;
    RECT 229.7 20.23 229.91 20.3 ;
    RECT 229.7 20.59 229.91 20.66 ;
    RECT 229.7 20.95 229.91 21.02 ;
    RECT 226.84 20.23 227.05 20.3 ;
    RECT 226.84 20.59 227.05 20.66 ;
    RECT 226.84 20.95 227.05 21.02 ;
    RECT 226.38 20.23 226.59 20.3 ;
    RECT 226.38 20.59 226.59 20.66 ;
    RECT 226.38 20.95 226.59 21.02 ;
    RECT 223.52 20.23 223.73 20.3 ;
    RECT 223.52 20.59 223.73 20.66 ;
    RECT 223.52 20.95 223.73 21.02 ;
    RECT 223.06 20.23 223.27 20.3 ;
    RECT 223.06 20.59 223.27 20.66 ;
    RECT 223.06 20.95 223.27 21.02 ;
    RECT 220.2 20.23 220.41 20.3 ;
    RECT 220.2 20.59 220.41 20.66 ;
    RECT 220.2 20.95 220.41 21.02 ;
    RECT 219.74 20.23 219.95 20.3 ;
    RECT 219.74 20.59 219.95 20.66 ;
    RECT 219.74 20.95 219.95 21.02 ;
    RECT 216.88 20.23 217.09 20.3 ;
    RECT 216.88 20.59 217.09 20.66 ;
    RECT 216.88 20.95 217.09 21.02 ;
    RECT 216.42 20.23 216.63 20.3 ;
    RECT 216.42 20.59 216.63 20.66 ;
    RECT 216.42 20.95 216.63 21.02 ;
    RECT 267.91 20.59 267.98 20.66 ;
    RECT 180.36 20.23 180.57 20.3 ;
    RECT 180.36 20.59 180.57 20.66 ;
    RECT 180.36 20.95 180.57 21.02 ;
    RECT 179.9 20.23 180.11 20.3 ;
    RECT 179.9 20.59 180.11 20.66 ;
    RECT 179.9 20.95 180.11 21.02 ;
    RECT 177.04 20.23 177.25 20.3 ;
    RECT 177.04 20.59 177.25 20.66 ;
    RECT 177.04 20.95 177.25 21.02 ;
    RECT 176.58 20.23 176.79 20.3 ;
    RECT 176.58 20.59 176.79 20.66 ;
    RECT 176.58 20.95 176.79 21.02 ;
    RECT 173.72 20.23 173.93 20.3 ;
    RECT 173.72 20.59 173.93 20.66 ;
    RECT 173.72 20.95 173.93 21.02 ;
    RECT 173.26 20.23 173.47 20.3 ;
    RECT 173.26 20.59 173.47 20.66 ;
    RECT 173.26 20.95 173.47 21.02 ;
    RECT 170.4 20.23 170.61 20.3 ;
    RECT 170.4 20.59 170.61 20.66 ;
    RECT 170.4 20.95 170.61 21.02 ;
    RECT 169.94 20.23 170.15 20.3 ;
    RECT 169.94 20.59 170.15 20.66 ;
    RECT 169.94 20.95 170.15 21.02 ;
    RECT 167.08 20.23 167.29 20.3 ;
    RECT 167.08 20.59 167.29 20.66 ;
    RECT 167.08 20.95 167.29 21.02 ;
    RECT 166.62 20.23 166.83 20.3 ;
    RECT 166.62 20.59 166.83 20.66 ;
    RECT 166.62 20.95 166.83 21.02 ;
    RECT 163.76 20.23 163.97 20.3 ;
    RECT 163.76 20.59 163.97 20.66 ;
    RECT 163.76 20.95 163.97 21.02 ;
    RECT 163.3 20.23 163.51 20.3 ;
    RECT 163.3 20.59 163.51 20.66 ;
    RECT 163.3 20.95 163.51 21.02 ;
    RECT 160.44 20.23 160.65 20.3 ;
    RECT 160.44 20.59 160.65 20.66 ;
    RECT 160.44 20.95 160.65 21.02 ;
    RECT 159.98 20.23 160.19 20.3 ;
    RECT 159.98 20.59 160.19 20.66 ;
    RECT 159.98 20.95 160.19 21.02 ;
    RECT 157.12 20.23 157.33 20.3 ;
    RECT 157.12 20.59 157.33 20.66 ;
    RECT 157.12 20.95 157.33 21.02 ;
    RECT 156.66 20.23 156.87 20.3 ;
    RECT 156.66 20.59 156.87 20.66 ;
    RECT 156.66 20.95 156.87 21.02 ;
    RECT 153.8 20.23 154.01 20.3 ;
    RECT 153.8 20.59 154.01 20.66 ;
    RECT 153.8 20.95 154.01 21.02 ;
    RECT 153.34 20.23 153.55 20.3 ;
    RECT 153.34 20.59 153.55 20.66 ;
    RECT 153.34 20.95 153.55 21.02 ;
    RECT 150.48 20.23 150.69 20.3 ;
    RECT 150.48 20.59 150.69 20.66 ;
    RECT 150.48 20.95 150.69 21.02 ;
    RECT 150.02 20.23 150.23 20.3 ;
    RECT 150.02 20.59 150.23 20.66 ;
    RECT 150.02 20.95 150.23 21.02 ;
    RECT 213.56 20.23 213.77 20.3 ;
    RECT 213.56 20.59 213.77 20.66 ;
    RECT 213.56 20.95 213.77 21.02 ;
    RECT 213.1 20.23 213.31 20.3 ;
    RECT 213.1 20.59 213.31 20.66 ;
    RECT 213.1 20.95 213.31 21.02 ;
    RECT 210.24 20.23 210.45 20.3 ;
    RECT 210.24 20.59 210.45 20.66 ;
    RECT 210.24 20.95 210.45 21.02 ;
    RECT 209.78 20.23 209.99 20.3 ;
    RECT 209.78 20.59 209.99 20.66 ;
    RECT 209.78 20.95 209.99 21.02 ;
    RECT 206.92 20.23 207.13 20.3 ;
    RECT 206.92 20.59 207.13 20.66 ;
    RECT 206.92 20.95 207.13 21.02 ;
    RECT 206.46 20.23 206.67 20.3 ;
    RECT 206.46 20.59 206.67 20.66 ;
    RECT 206.46 20.95 206.67 21.02 ;
    RECT 203.6 20.23 203.81 20.3 ;
    RECT 203.6 20.59 203.81 20.66 ;
    RECT 203.6 20.95 203.81 21.02 ;
    RECT 203.14 20.23 203.35 20.3 ;
    RECT 203.14 20.59 203.35 20.66 ;
    RECT 203.14 20.95 203.35 21.02 ;
    RECT 200.28 20.23 200.49 20.3 ;
    RECT 200.28 20.59 200.49 20.66 ;
    RECT 200.28 20.95 200.49 21.02 ;
    RECT 199.82 20.23 200.03 20.3 ;
    RECT 199.82 20.59 200.03 20.66 ;
    RECT 199.82 20.95 200.03 21.02 ;
    RECT 196.96 20.23 197.17 20.3 ;
    RECT 196.96 20.59 197.17 20.66 ;
    RECT 196.96 20.95 197.17 21.02 ;
    RECT 196.5 20.23 196.71 20.3 ;
    RECT 196.5 20.59 196.71 20.66 ;
    RECT 196.5 20.95 196.71 21.02 ;
    RECT 193.64 20.23 193.85 20.3 ;
    RECT 193.64 20.59 193.85 20.66 ;
    RECT 193.64 20.95 193.85 21.02 ;
    RECT 193.18 20.23 193.39 20.3 ;
    RECT 193.18 20.59 193.39 20.66 ;
    RECT 193.18 20.95 193.39 21.02 ;
    RECT 190.32 20.23 190.53 20.3 ;
    RECT 190.32 20.59 190.53 20.66 ;
    RECT 190.32 20.95 190.53 21.02 ;
    RECT 189.86 20.23 190.07 20.3 ;
    RECT 189.86 20.59 190.07 20.66 ;
    RECT 189.86 20.95 190.07 21.02 ;
    RECT 187.0 20.23 187.21 20.3 ;
    RECT 187.0 20.59 187.21 20.66 ;
    RECT 187.0 20.95 187.21 21.02 ;
    RECT 186.54 20.23 186.75 20.3 ;
    RECT 186.54 20.59 186.75 20.66 ;
    RECT 186.54 20.95 186.75 21.02 ;
    RECT 183.68 20.23 183.89 20.3 ;
    RECT 183.68 20.59 183.89 20.66 ;
    RECT 183.68 20.95 183.89 21.02 ;
    RECT 183.22 20.23 183.43 20.3 ;
    RECT 183.22 20.59 183.43 20.66 ;
    RECT 183.22 20.95 183.43 21.02 ;
    RECT 147.485 20.59 147.555 20.66 ;
    RECT 266.68 20.23 266.89 20.3 ;
    RECT 266.68 20.59 266.89 20.66 ;
    RECT 266.68 20.95 266.89 21.02 ;
    RECT 266.22 20.23 266.43 20.3 ;
    RECT 266.22 20.59 266.43 20.66 ;
    RECT 266.22 20.95 266.43 21.02 ;
    RECT 263.36 20.23 263.57 20.3 ;
    RECT 263.36 20.59 263.57 20.66 ;
    RECT 263.36 20.95 263.57 21.02 ;
    RECT 262.9 20.23 263.11 20.3 ;
    RECT 262.9 20.59 263.11 20.66 ;
    RECT 262.9 20.95 263.11 21.02 ;
    RECT 260.04 20.23 260.25 20.3 ;
    RECT 260.04 20.59 260.25 20.66 ;
    RECT 260.04 20.95 260.25 21.02 ;
    RECT 259.58 20.23 259.79 20.3 ;
    RECT 259.58 20.59 259.79 20.66 ;
    RECT 259.58 20.95 259.79 21.02 ;
    RECT 256.72 20.23 256.93 20.3 ;
    RECT 256.72 20.59 256.93 20.66 ;
    RECT 256.72 20.95 256.93 21.02 ;
    RECT 256.26 20.23 256.47 20.3 ;
    RECT 256.26 20.59 256.47 20.66 ;
    RECT 256.26 20.95 256.47 21.02 ;
    RECT 253.4 20.23 253.61 20.3 ;
    RECT 253.4 20.59 253.61 20.66 ;
    RECT 253.4 20.95 253.61 21.02 ;
    RECT 252.94 20.23 253.15 20.3 ;
    RECT 252.94 20.59 253.15 20.66 ;
    RECT 252.94 20.95 253.15 21.02 ;
    RECT 250.08 19.51 250.29 19.58 ;
    RECT 250.08 19.87 250.29 19.94 ;
    RECT 250.08 20.23 250.29 20.3 ;
    RECT 249.62 19.51 249.83 19.58 ;
    RECT 249.62 19.87 249.83 19.94 ;
    RECT 249.62 20.23 249.83 20.3 ;
    RECT 246.76 19.51 246.97 19.58 ;
    RECT 246.76 19.87 246.97 19.94 ;
    RECT 246.76 20.23 246.97 20.3 ;
    RECT 246.3 19.51 246.51 19.58 ;
    RECT 246.3 19.87 246.51 19.94 ;
    RECT 246.3 20.23 246.51 20.3 ;
    RECT 243.44 19.51 243.65 19.58 ;
    RECT 243.44 19.87 243.65 19.94 ;
    RECT 243.44 20.23 243.65 20.3 ;
    RECT 242.98 19.51 243.19 19.58 ;
    RECT 242.98 19.87 243.19 19.94 ;
    RECT 242.98 20.23 243.19 20.3 ;
    RECT 240.12 19.51 240.33 19.58 ;
    RECT 240.12 19.87 240.33 19.94 ;
    RECT 240.12 20.23 240.33 20.3 ;
    RECT 239.66 19.51 239.87 19.58 ;
    RECT 239.66 19.87 239.87 19.94 ;
    RECT 239.66 20.23 239.87 20.3 ;
    RECT 236.8 19.51 237.01 19.58 ;
    RECT 236.8 19.87 237.01 19.94 ;
    RECT 236.8 20.23 237.01 20.3 ;
    RECT 236.34 19.51 236.55 19.58 ;
    RECT 236.34 19.87 236.55 19.94 ;
    RECT 236.34 20.23 236.55 20.3 ;
    RECT 233.48 19.51 233.69 19.58 ;
    RECT 233.48 19.87 233.69 19.94 ;
    RECT 233.48 20.23 233.69 20.3 ;
    RECT 233.02 19.51 233.23 19.58 ;
    RECT 233.02 19.87 233.23 19.94 ;
    RECT 233.02 20.23 233.23 20.3 ;
    RECT 230.16 19.51 230.37 19.58 ;
    RECT 230.16 19.87 230.37 19.94 ;
    RECT 230.16 20.23 230.37 20.3 ;
    RECT 229.7 19.51 229.91 19.58 ;
    RECT 229.7 19.87 229.91 19.94 ;
    RECT 229.7 20.23 229.91 20.3 ;
    RECT 226.84 19.51 227.05 19.58 ;
    RECT 226.84 19.87 227.05 19.94 ;
    RECT 226.84 20.23 227.05 20.3 ;
    RECT 226.38 19.51 226.59 19.58 ;
    RECT 226.38 19.87 226.59 19.94 ;
    RECT 226.38 20.23 226.59 20.3 ;
    RECT 223.52 19.51 223.73 19.58 ;
    RECT 223.52 19.87 223.73 19.94 ;
    RECT 223.52 20.23 223.73 20.3 ;
    RECT 223.06 19.51 223.27 19.58 ;
    RECT 223.06 19.87 223.27 19.94 ;
    RECT 223.06 20.23 223.27 20.3 ;
    RECT 220.2 19.51 220.41 19.58 ;
    RECT 220.2 19.87 220.41 19.94 ;
    RECT 220.2 20.23 220.41 20.3 ;
    RECT 219.74 19.51 219.95 19.58 ;
    RECT 219.74 19.87 219.95 19.94 ;
    RECT 219.74 20.23 219.95 20.3 ;
    RECT 216.88 19.51 217.09 19.58 ;
    RECT 216.88 19.87 217.09 19.94 ;
    RECT 216.88 20.23 217.09 20.3 ;
    RECT 216.42 19.51 216.63 19.58 ;
    RECT 216.42 19.87 216.63 19.94 ;
    RECT 216.42 20.23 216.63 20.3 ;
    RECT 267.91 19.87 267.98 19.94 ;
    RECT 180.36 19.51 180.57 19.58 ;
    RECT 180.36 19.87 180.57 19.94 ;
    RECT 180.36 20.23 180.57 20.3 ;
    RECT 179.9 19.51 180.11 19.58 ;
    RECT 179.9 19.87 180.11 19.94 ;
    RECT 179.9 20.23 180.11 20.3 ;
    RECT 177.04 19.51 177.25 19.58 ;
    RECT 177.04 19.87 177.25 19.94 ;
    RECT 177.04 20.23 177.25 20.3 ;
    RECT 176.58 19.51 176.79 19.58 ;
    RECT 176.58 19.87 176.79 19.94 ;
    RECT 176.58 20.23 176.79 20.3 ;
    RECT 173.72 19.51 173.93 19.58 ;
    RECT 173.72 19.87 173.93 19.94 ;
    RECT 173.72 20.23 173.93 20.3 ;
    RECT 173.26 19.51 173.47 19.58 ;
    RECT 173.26 19.87 173.47 19.94 ;
    RECT 173.26 20.23 173.47 20.3 ;
    RECT 170.4 19.51 170.61 19.58 ;
    RECT 170.4 19.87 170.61 19.94 ;
    RECT 170.4 20.23 170.61 20.3 ;
    RECT 169.94 19.51 170.15 19.58 ;
    RECT 169.94 19.87 170.15 19.94 ;
    RECT 169.94 20.23 170.15 20.3 ;
    RECT 167.08 19.51 167.29 19.58 ;
    RECT 167.08 19.87 167.29 19.94 ;
    RECT 167.08 20.23 167.29 20.3 ;
    RECT 166.62 19.51 166.83 19.58 ;
    RECT 166.62 19.87 166.83 19.94 ;
    RECT 166.62 20.23 166.83 20.3 ;
    RECT 163.76 19.51 163.97 19.58 ;
    RECT 163.76 19.87 163.97 19.94 ;
    RECT 163.76 20.23 163.97 20.3 ;
    RECT 163.3 19.51 163.51 19.58 ;
    RECT 163.3 19.87 163.51 19.94 ;
    RECT 163.3 20.23 163.51 20.3 ;
    RECT 160.44 19.51 160.65 19.58 ;
    RECT 160.44 19.87 160.65 19.94 ;
    RECT 160.44 20.23 160.65 20.3 ;
    RECT 159.98 19.51 160.19 19.58 ;
    RECT 159.98 19.87 160.19 19.94 ;
    RECT 159.98 20.23 160.19 20.3 ;
    RECT 157.12 19.51 157.33 19.58 ;
    RECT 157.12 19.87 157.33 19.94 ;
    RECT 157.12 20.23 157.33 20.3 ;
    RECT 156.66 19.51 156.87 19.58 ;
    RECT 156.66 19.87 156.87 19.94 ;
    RECT 156.66 20.23 156.87 20.3 ;
    RECT 153.8 19.51 154.01 19.58 ;
    RECT 153.8 19.87 154.01 19.94 ;
    RECT 153.8 20.23 154.01 20.3 ;
    RECT 153.34 19.51 153.55 19.58 ;
    RECT 153.34 19.87 153.55 19.94 ;
    RECT 153.34 20.23 153.55 20.3 ;
    RECT 150.48 19.51 150.69 19.58 ;
    RECT 150.48 19.87 150.69 19.94 ;
    RECT 150.48 20.23 150.69 20.3 ;
    RECT 150.02 19.51 150.23 19.58 ;
    RECT 150.02 19.87 150.23 19.94 ;
    RECT 150.02 20.23 150.23 20.3 ;
    RECT 213.56 19.51 213.77 19.58 ;
    RECT 213.56 19.87 213.77 19.94 ;
    RECT 213.56 20.23 213.77 20.3 ;
    RECT 213.1 19.51 213.31 19.58 ;
    RECT 213.1 19.87 213.31 19.94 ;
    RECT 213.1 20.23 213.31 20.3 ;
    RECT 210.24 19.51 210.45 19.58 ;
    RECT 210.24 19.87 210.45 19.94 ;
    RECT 210.24 20.23 210.45 20.3 ;
    RECT 209.78 19.51 209.99 19.58 ;
    RECT 209.78 19.87 209.99 19.94 ;
    RECT 209.78 20.23 209.99 20.3 ;
    RECT 206.92 19.51 207.13 19.58 ;
    RECT 206.92 19.87 207.13 19.94 ;
    RECT 206.92 20.23 207.13 20.3 ;
    RECT 206.46 19.51 206.67 19.58 ;
    RECT 206.46 19.87 206.67 19.94 ;
    RECT 206.46 20.23 206.67 20.3 ;
    RECT 203.6 19.51 203.81 19.58 ;
    RECT 203.6 19.87 203.81 19.94 ;
    RECT 203.6 20.23 203.81 20.3 ;
    RECT 203.14 19.51 203.35 19.58 ;
    RECT 203.14 19.87 203.35 19.94 ;
    RECT 203.14 20.23 203.35 20.3 ;
    RECT 200.28 19.51 200.49 19.58 ;
    RECT 200.28 19.87 200.49 19.94 ;
    RECT 200.28 20.23 200.49 20.3 ;
    RECT 199.82 19.51 200.03 19.58 ;
    RECT 199.82 19.87 200.03 19.94 ;
    RECT 199.82 20.23 200.03 20.3 ;
    RECT 196.96 19.51 197.17 19.58 ;
    RECT 196.96 19.87 197.17 19.94 ;
    RECT 196.96 20.23 197.17 20.3 ;
    RECT 196.5 19.51 196.71 19.58 ;
    RECT 196.5 19.87 196.71 19.94 ;
    RECT 196.5 20.23 196.71 20.3 ;
    RECT 193.64 19.51 193.85 19.58 ;
    RECT 193.64 19.87 193.85 19.94 ;
    RECT 193.64 20.23 193.85 20.3 ;
    RECT 193.18 19.51 193.39 19.58 ;
    RECT 193.18 19.87 193.39 19.94 ;
    RECT 193.18 20.23 193.39 20.3 ;
    RECT 190.32 19.51 190.53 19.58 ;
    RECT 190.32 19.87 190.53 19.94 ;
    RECT 190.32 20.23 190.53 20.3 ;
    RECT 189.86 19.51 190.07 19.58 ;
    RECT 189.86 19.87 190.07 19.94 ;
    RECT 189.86 20.23 190.07 20.3 ;
    RECT 187.0 19.51 187.21 19.58 ;
    RECT 187.0 19.87 187.21 19.94 ;
    RECT 187.0 20.23 187.21 20.3 ;
    RECT 186.54 19.51 186.75 19.58 ;
    RECT 186.54 19.87 186.75 19.94 ;
    RECT 186.54 20.23 186.75 20.3 ;
    RECT 183.68 19.51 183.89 19.58 ;
    RECT 183.68 19.87 183.89 19.94 ;
    RECT 183.68 20.23 183.89 20.3 ;
    RECT 183.22 19.51 183.43 19.58 ;
    RECT 183.22 19.87 183.43 19.94 ;
    RECT 183.22 20.23 183.43 20.3 ;
    RECT 147.485 19.87 147.555 19.94 ;
    RECT 266.68 19.51 266.89 19.58 ;
    RECT 266.68 19.87 266.89 19.94 ;
    RECT 266.68 20.23 266.89 20.3 ;
    RECT 266.22 19.51 266.43 19.58 ;
    RECT 266.22 19.87 266.43 19.94 ;
    RECT 266.22 20.23 266.43 20.3 ;
    RECT 263.36 19.51 263.57 19.58 ;
    RECT 263.36 19.87 263.57 19.94 ;
    RECT 263.36 20.23 263.57 20.3 ;
    RECT 262.9 19.51 263.11 19.58 ;
    RECT 262.9 19.87 263.11 19.94 ;
    RECT 262.9 20.23 263.11 20.3 ;
    RECT 260.04 19.51 260.25 19.58 ;
    RECT 260.04 19.87 260.25 19.94 ;
    RECT 260.04 20.23 260.25 20.3 ;
    RECT 259.58 19.51 259.79 19.58 ;
    RECT 259.58 19.87 259.79 19.94 ;
    RECT 259.58 20.23 259.79 20.3 ;
    RECT 256.72 19.51 256.93 19.58 ;
    RECT 256.72 19.87 256.93 19.94 ;
    RECT 256.72 20.23 256.93 20.3 ;
    RECT 256.26 19.51 256.47 19.58 ;
    RECT 256.26 19.87 256.47 19.94 ;
    RECT 256.26 20.23 256.47 20.3 ;
    RECT 253.4 19.51 253.61 19.58 ;
    RECT 253.4 19.87 253.61 19.94 ;
    RECT 253.4 20.23 253.61 20.3 ;
    RECT 252.94 19.51 253.15 19.58 ;
    RECT 252.94 19.87 253.15 19.94 ;
    RECT 252.94 20.23 253.15 20.3 ;
    RECT 250.08 35.35 250.29 35.42 ;
    RECT 250.08 35.71 250.29 35.78 ;
    RECT 250.08 36.07 250.29 36.14 ;
    RECT 249.62 35.35 249.83 35.42 ;
    RECT 249.62 35.71 249.83 35.78 ;
    RECT 249.62 36.07 249.83 36.14 ;
    RECT 246.76 35.35 246.97 35.42 ;
    RECT 246.76 35.71 246.97 35.78 ;
    RECT 246.76 36.07 246.97 36.14 ;
    RECT 246.3 35.35 246.51 35.42 ;
    RECT 246.3 35.71 246.51 35.78 ;
    RECT 246.3 36.07 246.51 36.14 ;
    RECT 243.44 35.35 243.65 35.42 ;
    RECT 243.44 35.71 243.65 35.78 ;
    RECT 243.44 36.07 243.65 36.14 ;
    RECT 242.98 35.35 243.19 35.42 ;
    RECT 242.98 35.71 243.19 35.78 ;
    RECT 242.98 36.07 243.19 36.14 ;
    RECT 240.12 35.35 240.33 35.42 ;
    RECT 240.12 35.71 240.33 35.78 ;
    RECT 240.12 36.07 240.33 36.14 ;
    RECT 239.66 35.35 239.87 35.42 ;
    RECT 239.66 35.71 239.87 35.78 ;
    RECT 239.66 36.07 239.87 36.14 ;
    RECT 236.8 35.35 237.01 35.42 ;
    RECT 236.8 35.71 237.01 35.78 ;
    RECT 236.8 36.07 237.01 36.14 ;
    RECT 236.34 35.35 236.55 35.42 ;
    RECT 236.34 35.71 236.55 35.78 ;
    RECT 236.34 36.07 236.55 36.14 ;
    RECT 233.48 35.35 233.69 35.42 ;
    RECT 233.48 35.71 233.69 35.78 ;
    RECT 233.48 36.07 233.69 36.14 ;
    RECT 233.02 35.35 233.23 35.42 ;
    RECT 233.02 35.71 233.23 35.78 ;
    RECT 233.02 36.07 233.23 36.14 ;
    RECT 230.16 35.35 230.37 35.42 ;
    RECT 230.16 35.71 230.37 35.78 ;
    RECT 230.16 36.07 230.37 36.14 ;
    RECT 229.7 35.35 229.91 35.42 ;
    RECT 229.7 35.71 229.91 35.78 ;
    RECT 229.7 36.07 229.91 36.14 ;
    RECT 226.84 35.35 227.05 35.42 ;
    RECT 226.84 35.71 227.05 35.78 ;
    RECT 226.84 36.07 227.05 36.14 ;
    RECT 226.38 35.35 226.59 35.42 ;
    RECT 226.38 35.71 226.59 35.78 ;
    RECT 226.38 36.07 226.59 36.14 ;
    RECT 223.52 35.35 223.73 35.42 ;
    RECT 223.52 35.71 223.73 35.78 ;
    RECT 223.52 36.07 223.73 36.14 ;
    RECT 223.06 35.35 223.27 35.42 ;
    RECT 223.06 35.71 223.27 35.78 ;
    RECT 223.06 36.07 223.27 36.14 ;
    RECT 220.2 35.35 220.41 35.42 ;
    RECT 220.2 35.71 220.41 35.78 ;
    RECT 220.2 36.07 220.41 36.14 ;
    RECT 219.74 35.35 219.95 35.42 ;
    RECT 219.74 35.71 219.95 35.78 ;
    RECT 219.74 36.07 219.95 36.14 ;
    RECT 216.88 35.35 217.09 35.42 ;
    RECT 216.88 35.71 217.09 35.78 ;
    RECT 216.88 36.07 217.09 36.14 ;
    RECT 216.42 35.35 216.63 35.42 ;
    RECT 216.42 35.71 216.63 35.78 ;
    RECT 216.42 36.07 216.63 36.14 ;
    RECT 267.91 35.71 267.98 35.78 ;
    RECT 180.36 35.35 180.57 35.42 ;
    RECT 180.36 35.71 180.57 35.78 ;
    RECT 180.36 36.07 180.57 36.14 ;
    RECT 179.9 35.35 180.11 35.42 ;
    RECT 179.9 35.71 180.11 35.78 ;
    RECT 179.9 36.07 180.11 36.14 ;
    RECT 177.04 35.35 177.25 35.42 ;
    RECT 177.04 35.71 177.25 35.78 ;
    RECT 177.04 36.07 177.25 36.14 ;
    RECT 176.58 35.35 176.79 35.42 ;
    RECT 176.58 35.71 176.79 35.78 ;
    RECT 176.58 36.07 176.79 36.14 ;
    RECT 173.72 35.35 173.93 35.42 ;
    RECT 173.72 35.71 173.93 35.78 ;
    RECT 173.72 36.07 173.93 36.14 ;
    RECT 173.26 35.35 173.47 35.42 ;
    RECT 173.26 35.71 173.47 35.78 ;
    RECT 173.26 36.07 173.47 36.14 ;
    RECT 170.4 35.35 170.61 35.42 ;
    RECT 170.4 35.71 170.61 35.78 ;
    RECT 170.4 36.07 170.61 36.14 ;
    RECT 169.94 35.35 170.15 35.42 ;
    RECT 169.94 35.71 170.15 35.78 ;
    RECT 169.94 36.07 170.15 36.14 ;
    RECT 167.08 35.35 167.29 35.42 ;
    RECT 167.08 35.71 167.29 35.78 ;
    RECT 167.08 36.07 167.29 36.14 ;
    RECT 166.62 35.35 166.83 35.42 ;
    RECT 166.62 35.71 166.83 35.78 ;
    RECT 166.62 36.07 166.83 36.14 ;
    RECT 163.76 35.35 163.97 35.42 ;
    RECT 163.76 35.71 163.97 35.78 ;
    RECT 163.76 36.07 163.97 36.14 ;
    RECT 163.3 35.35 163.51 35.42 ;
    RECT 163.3 35.71 163.51 35.78 ;
    RECT 163.3 36.07 163.51 36.14 ;
    RECT 160.44 35.35 160.65 35.42 ;
    RECT 160.44 35.71 160.65 35.78 ;
    RECT 160.44 36.07 160.65 36.14 ;
    RECT 159.98 35.35 160.19 35.42 ;
    RECT 159.98 35.71 160.19 35.78 ;
    RECT 159.98 36.07 160.19 36.14 ;
    RECT 157.12 35.35 157.33 35.42 ;
    RECT 157.12 35.71 157.33 35.78 ;
    RECT 157.12 36.07 157.33 36.14 ;
    RECT 156.66 35.35 156.87 35.42 ;
    RECT 156.66 35.71 156.87 35.78 ;
    RECT 156.66 36.07 156.87 36.14 ;
    RECT 153.8 35.35 154.01 35.42 ;
    RECT 153.8 35.71 154.01 35.78 ;
    RECT 153.8 36.07 154.01 36.14 ;
    RECT 153.34 35.35 153.55 35.42 ;
    RECT 153.34 35.71 153.55 35.78 ;
    RECT 153.34 36.07 153.55 36.14 ;
    RECT 150.48 35.35 150.69 35.42 ;
    RECT 150.48 35.71 150.69 35.78 ;
    RECT 150.48 36.07 150.69 36.14 ;
    RECT 150.02 35.35 150.23 35.42 ;
    RECT 150.02 35.71 150.23 35.78 ;
    RECT 150.02 36.07 150.23 36.14 ;
    RECT 213.56 35.35 213.77 35.42 ;
    RECT 213.56 35.71 213.77 35.78 ;
    RECT 213.56 36.07 213.77 36.14 ;
    RECT 213.1 35.35 213.31 35.42 ;
    RECT 213.1 35.71 213.31 35.78 ;
    RECT 213.1 36.07 213.31 36.14 ;
    RECT 210.24 35.35 210.45 35.42 ;
    RECT 210.24 35.71 210.45 35.78 ;
    RECT 210.24 36.07 210.45 36.14 ;
    RECT 209.78 35.35 209.99 35.42 ;
    RECT 209.78 35.71 209.99 35.78 ;
    RECT 209.78 36.07 209.99 36.14 ;
    RECT 206.92 35.35 207.13 35.42 ;
    RECT 206.92 35.71 207.13 35.78 ;
    RECT 206.92 36.07 207.13 36.14 ;
    RECT 206.46 35.35 206.67 35.42 ;
    RECT 206.46 35.71 206.67 35.78 ;
    RECT 206.46 36.07 206.67 36.14 ;
    RECT 203.6 35.35 203.81 35.42 ;
    RECT 203.6 35.71 203.81 35.78 ;
    RECT 203.6 36.07 203.81 36.14 ;
    RECT 203.14 35.35 203.35 35.42 ;
    RECT 203.14 35.71 203.35 35.78 ;
    RECT 203.14 36.07 203.35 36.14 ;
    RECT 200.28 35.35 200.49 35.42 ;
    RECT 200.28 35.71 200.49 35.78 ;
    RECT 200.28 36.07 200.49 36.14 ;
    RECT 199.82 35.35 200.03 35.42 ;
    RECT 199.82 35.71 200.03 35.78 ;
    RECT 199.82 36.07 200.03 36.14 ;
    RECT 196.96 35.35 197.17 35.42 ;
    RECT 196.96 35.71 197.17 35.78 ;
    RECT 196.96 36.07 197.17 36.14 ;
    RECT 196.5 35.35 196.71 35.42 ;
    RECT 196.5 35.71 196.71 35.78 ;
    RECT 196.5 36.07 196.71 36.14 ;
    RECT 193.64 35.35 193.85 35.42 ;
    RECT 193.64 35.71 193.85 35.78 ;
    RECT 193.64 36.07 193.85 36.14 ;
    RECT 193.18 35.35 193.39 35.42 ;
    RECT 193.18 35.71 193.39 35.78 ;
    RECT 193.18 36.07 193.39 36.14 ;
    RECT 190.32 35.35 190.53 35.42 ;
    RECT 190.32 35.71 190.53 35.78 ;
    RECT 190.32 36.07 190.53 36.14 ;
    RECT 189.86 35.35 190.07 35.42 ;
    RECT 189.86 35.71 190.07 35.78 ;
    RECT 189.86 36.07 190.07 36.14 ;
    RECT 187.0 35.35 187.21 35.42 ;
    RECT 187.0 35.71 187.21 35.78 ;
    RECT 187.0 36.07 187.21 36.14 ;
    RECT 186.54 35.35 186.75 35.42 ;
    RECT 186.54 35.71 186.75 35.78 ;
    RECT 186.54 36.07 186.75 36.14 ;
    RECT 183.68 35.35 183.89 35.42 ;
    RECT 183.68 35.71 183.89 35.78 ;
    RECT 183.68 36.07 183.89 36.14 ;
    RECT 183.22 35.35 183.43 35.42 ;
    RECT 183.22 35.71 183.43 35.78 ;
    RECT 183.22 36.07 183.43 36.14 ;
    RECT 147.485 35.71 147.555 35.78 ;
    RECT 266.68 35.35 266.89 35.42 ;
    RECT 266.68 35.71 266.89 35.78 ;
    RECT 266.68 36.07 266.89 36.14 ;
    RECT 266.22 35.35 266.43 35.42 ;
    RECT 266.22 35.71 266.43 35.78 ;
    RECT 266.22 36.07 266.43 36.14 ;
    RECT 263.36 35.35 263.57 35.42 ;
    RECT 263.36 35.71 263.57 35.78 ;
    RECT 263.36 36.07 263.57 36.14 ;
    RECT 262.9 35.35 263.11 35.42 ;
    RECT 262.9 35.71 263.11 35.78 ;
    RECT 262.9 36.07 263.11 36.14 ;
    RECT 260.04 35.35 260.25 35.42 ;
    RECT 260.04 35.71 260.25 35.78 ;
    RECT 260.04 36.07 260.25 36.14 ;
    RECT 259.58 35.35 259.79 35.42 ;
    RECT 259.58 35.71 259.79 35.78 ;
    RECT 259.58 36.07 259.79 36.14 ;
    RECT 256.72 35.35 256.93 35.42 ;
    RECT 256.72 35.71 256.93 35.78 ;
    RECT 256.72 36.07 256.93 36.14 ;
    RECT 256.26 35.35 256.47 35.42 ;
    RECT 256.26 35.71 256.47 35.78 ;
    RECT 256.26 36.07 256.47 36.14 ;
    RECT 253.4 35.35 253.61 35.42 ;
    RECT 253.4 35.71 253.61 35.78 ;
    RECT 253.4 36.07 253.61 36.14 ;
    RECT 252.94 35.35 253.15 35.42 ;
    RECT 252.94 35.71 253.15 35.78 ;
    RECT 252.94 36.07 253.15 36.14 ;
    RECT 250.08 18.79 250.29 18.86 ;
    RECT 250.08 19.15 250.29 19.22 ;
    RECT 250.08 19.51 250.29 19.58 ;
    RECT 249.62 18.79 249.83 18.86 ;
    RECT 249.62 19.15 249.83 19.22 ;
    RECT 249.62 19.51 249.83 19.58 ;
    RECT 246.76 18.79 246.97 18.86 ;
    RECT 246.76 19.15 246.97 19.22 ;
    RECT 246.76 19.51 246.97 19.58 ;
    RECT 246.3 18.79 246.51 18.86 ;
    RECT 246.3 19.15 246.51 19.22 ;
    RECT 246.3 19.51 246.51 19.58 ;
    RECT 243.44 18.79 243.65 18.86 ;
    RECT 243.44 19.15 243.65 19.22 ;
    RECT 243.44 19.51 243.65 19.58 ;
    RECT 242.98 18.79 243.19 18.86 ;
    RECT 242.98 19.15 243.19 19.22 ;
    RECT 242.98 19.51 243.19 19.58 ;
    RECT 240.12 18.79 240.33 18.86 ;
    RECT 240.12 19.15 240.33 19.22 ;
    RECT 240.12 19.51 240.33 19.58 ;
    RECT 239.66 18.79 239.87 18.86 ;
    RECT 239.66 19.15 239.87 19.22 ;
    RECT 239.66 19.51 239.87 19.58 ;
    RECT 236.8 18.79 237.01 18.86 ;
    RECT 236.8 19.15 237.01 19.22 ;
    RECT 236.8 19.51 237.01 19.58 ;
    RECT 236.34 18.79 236.55 18.86 ;
    RECT 236.34 19.15 236.55 19.22 ;
    RECT 236.34 19.51 236.55 19.58 ;
    RECT 233.48 18.79 233.69 18.86 ;
    RECT 233.48 19.15 233.69 19.22 ;
    RECT 233.48 19.51 233.69 19.58 ;
    RECT 233.02 18.79 233.23 18.86 ;
    RECT 233.02 19.15 233.23 19.22 ;
    RECT 233.02 19.51 233.23 19.58 ;
    RECT 230.16 18.79 230.37 18.86 ;
    RECT 230.16 19.15 230.37 19.22 ;
    RECT 230.16 19.51 230.37 19.58 ;
    RECT 229.7 18.79 229.91 18.86 ;
    RECT 229.7 19.15 229.91 19.22 ;
    RECT 229.7 19.51 229.91 19.58 ;
    RECT 226.84 18.79 227.05 18.86 ;
    RECT 226.84 19.15 227.05 19.22 ;
    RECT 226.84 19.51 227.05 19.58 ;
    RECT 226.38 18.79 226.59 18.86 ;
    RECT 226.38 19.15 226.59 19.22 ;
    RECT 226.38 19.51 226.59 19.58 ;
    RECT 223.52 18.79 223.73 18.86 ;
    RECT 223.52 19.15 223.73 19.22 ;
    RECT 223.52 19.51 223.73 19.58 ;
    RECT 223.06 18.79 223.27 18.86 ;
    RECT 223.06 19.15 223.27 19.22 ;
    RECT 223.06 19.51 223.27 19.58 ;
    RECT 220.2 18.79 220.41 18.86 ;
    RECT 220.2 19.15 220.41 19.22 ;
    RECT 220.2 19.51 220.41 19.58 ;
    RECT 219.74 18.79 219.95 18.86 ;
    RECT 219.74 19.15 219.95 19.22 ;
    RECT 219.74 19.51 219.95 19.58 ;
    RECT 216.88 18.79 217.09 18.86 ;
    RECT 216.88 19.15 217.09 19.22 ;
    RECT 216.88 19.51 217.09 19.58 ;
    RECT 216.42 18.79 216.63 18.86 ;
    RECT 216.42 19.15 216.63 19.22 ;
    RECT 216.42 19.51 216.63 19.58 ;
    RECT 267.91 19.15 267.98 19.22 ;
    RECT 180.36 18.79 180.57 18.86 ;
    RECT 180.36 19.15 180.57 19.22 ;
    RECT 180.36 19.51 180.57 19.58 ;
    RECT 179.9 18.79 180.11 18.86 ;
    RECT 179.9 19.15 180.11 19.22 ;
    RECT 179.9 19.51 180.11 19.58 ;
    RECT 177.04 18.79 177.25 18.86 ;
    RECT 177.04 19.15 177.25 19.22 ;
    RECT 177.04 19.51 177.25 19.58 ;
    RECT 176.58 18.79 176.79 18.86 ;
    RECT 176.58 19.15 176.79 19.22 ;
    RECT 176.58 19.51 176.79 19.58 ;
    RECT 173.72 18.79 173.93 18.86 ;
    RECT 173.72 19.15 173.93 19.22 ;
    RECT 173.72 19.51 173.93 19.58 ;
    RECT 173.26 18.79 173.47 18.86 ;
    RECT 173.26 19.15 173.47 19.22 ;
    RECT 173.26 19.51 173.47 19.58 ;
    RECT 170.4 18.79 170.61 18.86 ;
    RECT 170.4 19.15 170.61 19.22 ;
    RECT 170.4 19.51 170.61 19.58 ;
    RECT 169.94 18.79 170.15 18.86 ;
    RECT 169.94 19.15 170.15 19.22 ;
    RECT 169.94 19.51 170.15 19.58 ;
    RECT 167.08 18.79 167.29 18.86 ;
    RECT 167.08 19.15 167.29 19.22 ;
    RECT 167.08 19.51 167.29 19.58 ;
    RECT 166.62 18.79 166.83 18.86 ;
    RECT 166.62 19.15 166.83 19.22 ;
    RECT 166.62 19.51 166.83 19.58 ;
    RECT 163.76 18.79 163.97 18.86 ;
    RECT 163.76 19.15 163.97 19.22 ;
    RECT 163.76 19.51 163.97 19.58 ;
    RECT 163.3 18.79 163.51 18.86 ;
    RECT 163.3 19.15 163.51 19.22 ;
    RECT 163.3 19.51 163.51 19.58 ;
    RECT 160.44 18.79 160.65 18.86 ;
    RECT 160.44 19.15 160.65 19.22 ;
    RECT 160.44 19.51 160.65 19.58 ;
    RECT 159.98 18.79 160.19 18.86 ;
    RECT 159.98 19.15 160.19 19.22 ;
    RECT 159.98 19.51 160.19 19.58 ;
    RECT 157.12 18.79 157.33 18.86 ;
    RECT 157.12 19.15 157.33 19.22 ;
    RECT 157.12 19.51 157.33 19.58 ;
    RECT 156.66 18.79 156.87 18.86 ;
    RECT 156.66 19.15 156.87 19.22 ;
    RECT 156.66 19.51 156.87 19.58 ;
    RECT 153.8 18.79 154.01 18.86 ;
    RECT 153.8 19.15 154.01 19.22 ;
    RECT 153.8 19.51 154.01 19.58 ;
    RECT 153.34 18.79 153.55 18.86 ;
    RECT 153.34 19.15 153.55 19.22 ;
    RECT 153.34 19.51 153.55 19.58 ;
    RECT 150.48 18.79 150.69 18.86 ;
    RECT 150.48 19.15 150.69 19.22 ;
    RECT 150.48 19.51 150.69 19.58 ;
    RECT 150.02 18.79 150.23 18.86 ;
    RECT 150.02 19.15 150.23 19.22 ;
    RECT 150.02 19.51 150.23 19.58 ;
    RECT 213.56 18.79 213.77 18.86 ;
    RECT 213.56 19.15 213.77 19.22 ;
    RECT 213.56 19.51 213.77 19.58 ;
    RECT 213.1 18.79 213.31 18.86 ;
    RECT 213.1 19.15 213.31 19.22 ;
    RECT 213.1 19.51 213.31 19.58 ;
    RECT 210.24 18.79 210.45 18.86 ;
    RECT 210.24 19.15 210.45 19.22 ;
    RECT 210.24 19.51 210.45 19.58 ;
    RECT 209.78 18.79 209.99 18.86 ;
    RECT 209.78 19.15 209.99 19.22 ;
    RECT 209.78 19.51 209.99 19.58 ;
    RECT 206.92 18.79 207.13 18.86 ;
    RECT 206.92 19.15 207.13 19.22 ;
    RECT 206.92 19.51 207.13 19.58 ;
    RECT 206.46 18.79 206.67 18.86 ;
    RECT 206.46 19.15 206.67 19.22 ;
    RECT 206.46 19.51 206.67 19.58 ;
    RECT 203.6 18.79 203.81 18.86 ;
    RECT 203.6 19.15 203.81 19.22 ;
    RECT 203.6 19.51 203.81 19.58 ;
    RECT 203.14 18.79 203.35 18.86 ;
    RECT 203.14 19.15 203.35 19.22 ;
    RECT 203.14 19.51 203.35 19.58 ;
    RECT 200.28 18.79 200.49 18.86 ;
    RECT 200.28 19.15 200.49 19.22 ;
    RECT 200.28 19.51 200.49 19.58 ;
    RECT 199.82 18.79 200.03 18.86 ;
    RECT 199.82 19.15 200.03 19.22 ;
    RECT 199.82 19.51 200.03 19.58 ;
    RECT 196.96 18.79 197.17 18.86 ;
    RECT 196.96 19.15 197.17 19.22 ;
    RECT 196.96 19.51 197.17 19.58 ;
    RECT 196.5 18.79 196.71 18.86 ;
    RECT 196.5 19.15 196.71 19.22 ;
    RECT 196.5 19.51 196.71 19.58 ;
    RECT 193.64 18.79 193.85 18.86 ;
    RECT 193.64 19.15 193.85 19.22 ;
    RECT 193.64 19.51 193.85 19.58 ;
    RECT 193.18 18.79 193.39 18.86 ;
    RECT 193.18 19.15 193.39 19.22 ;
    RECT 193.18 19.51 193.39 19.58 ;
    RECT 190.32 18.79 190.53 18.86 ;
    RECT 190.32 19.15 190.53 19.22 ;
    RECT 190.32 19.51 190.53 19.58 ;
    RECT 189.86 18.79 190.07 18.86 ;
    RECT 189.86 19.15 190.07 19.22 ;
    RECT 189.86 19.51 190.07 19.58 ;
    RECT 187.0 18.79 187.21 18.86 ;
    RECT 187.0 19.15 187.21 19.22 ;
    RECT 187.0 19.51 187.21 19.58 ;
    RECT 186.54 18.79 186.75 18.86 ;
    RECT 186.54 19.15 186.75 19.22 ;
    RECT 186.54 19.51 186.75 19.58 ;
    RECT 183.68 18.79 183.89 18.86 ;
    RECT 183.68 19.15 183.89 19.22 ;
    RECT 183.68 19.51 183.89 19.58 ;
    RECT 183.22 18.79 183.43 18.86 ;
    RECT 183.22 19.15 183.43 19.22 ;
    RECT 183.22 19.51 183.43 19.58 ;
    RECT 147.485 19.15 147.555 19.22 ;
    RECT 266.68 18.79 266.89 18.86 ;
    RECT 266.68 19.15 266.89 19.22 ;
    RECT 266.68 19.51 266.89 19.58 ;
    RECT 266.22 18.79 266.43 18.86 ;
    RECT 266.22 19.15 266.43 19.22 ;
    RECT 266.22 19.51 266.43 19.58 ;
    RECT 263.36 18.79 263.57 18.86 ;
    RECT 263.36 19.15 263.57 19.22 ;
    RECT 263.36 19.51 263.57 19.58 ;
    RECT 262.9 18.79 263.11 18.86 ;
    RECT 262.9 19.15 263.11 19.22 ;
    RECT 262.9 19.51 263.11 19.58 ;
    RECT 260.04 18.79 260.25 18.86 ;
    RECT 260.04 19.15 260.25 19.22 ;
    RECT 260.04 19.51 260.25 19.58 ;
    RECT 259.58 18.79 259.79 18.86 ;
    RECT 259.58 19.15 259.79 19.22 ;
    RECT 259.58 19.51 259.79 19.58 ;
    RECT 256.72 18.79 256.93 18.86 ;
    RECT 256.72 19.15 256.93 19.22 ;
    RECT 256.72 19.51 256.93 19.58 ;
    RECT 256.26 18.79 256.47 18.86 ;
    RECT 256.26 19.15 256.47 19.22 ;
    RECT 256.26 19.51 256.47 19.58 ;
    RECT 253.4 18.79 253.61 18.86 ;
    RECT 253.4 19.15 253.61 19.22 ;
    RECT 253.4 19.51 253.61 19.58 ;
    RECT 252.94 18.79 253.15 18.86 ;
    RECT 252.94 19.15 253.15 19.22 ;
    RECT 252.94 19.51 253.15 19.58 ;
    RECT 250.08 34.63 250.29 34.7 ;
    RECT 250.08 34.99 250.29 35.06 ;
    RECT 250.08 35.35 250.29 35.42 ;
    RECT 249.62 34.63 249.83 34.7 ;
    RECT 249.62 34.99 249.83 35.06 ;
    RECT 249.62 35.35 249.83 35.42 ;
    RECT 246.76 34.63 246.97 34.7 ;
    RECT 246.76 34.99 246.97 35.06 ;
    RECT 246.76 35.35 246.97 35.42 ;
    RECT 246.3 34.63 246.51 34.7 ;
    RECT 246.3 34.99 246.51 35.06 ;
    RECT 246.3 35.35 246.51 35.42 ;
    RECT 243.44 34.63 243.65 34.7 ;
    RECT 243.44 34.99 243.65 35.06 ;
    RECT 243.44 35.35 243.65 35.42 ;
    RECT 242.98 34.63 243.19 34.7 ;
    RECT 242.98 34.99 243.19 35.06 ;
    RECT 242.98 35.35 243.19 35.42 ;
    RECT 240.12 34.63 240.33 34.7 ;
    RECT 240.12 34.99 240.33 35.06 ;
    RECT 240.12 35.35 240.33 35.42 ;
    RECT 239.66 34.63 239.87 34.7 ;
    RECT 239.66 34.99 239.87 35.06 ;
    RECT 239.66 35.35 239.87 35.42 ;
    RECT 236.8 34.63 237.01 34.7 ;
    RECT 236.8 34.99 237.01 35.06 ;
    RECT 236.8 35.35 237.01 35.42 ;
    RECT 236.34 34.63 236.55 34.7 ;
    RECT 236.34 34.99 236.55 35.06 ;
    RECT 236.34 35.35 236.55 35.42 ;
    RECT 233.48 34.63 233.69 34.7 ;
    RECT 233.48 34.99 233.69 35.06 ;
    RECT 233.48 35.35 233.69 35.42 ;
    RECT 233.02 34.63 233.23 34.7 ;
    RECT 233.02 34.99 233.23 35.06 ;
    RECT 233.02 35.35 233.23 35.42 ;
    RECT 230.16 34.63 230.37 34.7 ;
    RECT 230.16 34.99 230.37 35.06 ;
    RECT 230.16 35.35 230.37 35.42 ;
    RECT 229.7 34.63 229.91 34.7 ;
    RECT 229.7 34.99 229.91 35.06 ;
    RECT 229.7 35.35 229.91 35.42 ;
    RECT 226.84 34.63 227.05 34.7 ;
    RECT 226.84 34.99 227.05 35.06 ;
    RECT 226.84 35.35 227.05 35.42 ;
    RECT 226.38 34.63 226.59 34.7 ;
    RECT 226.38 34.99 226.59 35.06 ;
    RECT 226.38 35.35 226.59 35.42 ;
    RECT 223.52 34.63 223.73 34.7 ;
    RECT 223.52 34.99 223.73 35.06 ;
    RECT 223.52 35.35 223.73 35.42 ;
    RECT 223.06 34.63 223.27 34.7 ;
    RECT 223.06 34.99 223.27 35.06 ;
    RECT 223.06 35.35 223.27 35.42 ;
    RECT 220.2 34.63 220.41 34.7 ;
    RECT 220.2 34.99 220.41 35.06 ;
    RECT 220.2 35.35 220.41 35.42 ;
    RECT 219.74 34.63 219.95 34.7 ;
    RECT 219.74 34.99 219.95 35.06 ;
    RECT 219.74 35.35 219.95 35.42 ;
    RECT 216.88 34.63 217.09 34.7 ;
    RECT 216.88 34.99 217.09 35.06 ;
    RECT 216.88 35.35 217.09 35.42 ;
    RECT 216.42 34.63 216.63 34.7 ;
    RECT 216.42 34.99 216.63 35.06 ;
    RECT 216.42 35.35 216.63 35.42 ;
    RECT 267.91 34.99 267.98 35.06 ;
    RECT 180.36 34.63 180.57 34.7 ;
    RECT 180.36 34.99 180.57 35.06 ;
    RECT 180.36 35.35 180.57 35.42 ;
    RECT 179.9 34.63 180.11 34.7 ;
    RECT 179.9 34.99 180.11 35.06 ;
    RECT 179.9 35.35 180.11 35.42 ;
    RECT 177.04 34.63 177.25 34.7 ;
    RECT 177.04 34.99 177.25 35.06 ;
    RECT 177.04 35.35 177.25 35.42 ;
    RECT 176.58 34.63 176.79 34.7 ;
    RECT 176.58 34.99 176.79 35.06 ;
    RECT 176.58 35.35 176.79 35.42 ;
    RECT 173.72 34.63 173.93 34.7 ;
    RECT 173.72 34.99 173.93 35.06 ;
    RECT 173.72 35.35 173.93 35.42 ;
    RECT 173.26 34.63 173.47 34.7 ;
    RECT 173.26 34.99 173.47 35.06 ;
    RECT 173.26 35.35 173.47 35.42 ;
    RECT 170.4 34.63 170.61 34.7 ;
    RECT 170.4 34.99 170.61 35.06 ;
    RECT 170.4 35.35 170.61 35.42 ;
    RECT 169.94 34.63 170.15 34.7 ;
    RECT 169.94 34.99 170.15 35.06 ;
    RECT 169.94 35.35 170.15 35.42 ;
    RECT 167.08 34.63 167.29 34.7 ;
    RECT 167.08 34.99 167.29 35.06 ;
    RECT 167.08 35.35 167.29 35.42 ;
    RECT 166.62 34.63 166.83 34.7 ;
    RECT 166.62 34.99 166.83 35.06 ;
    RECT 166.62 35.35 166.83 35.42 ;
    RECT 163.76 34.63 163.97 34.7 ;
    RECT 163.76 34.99 163.97 35.06 ;
    RECT 163.76 35.35 163.97 35.42 ;
    RECT 163.3 34.63 163.51 34.7 ;
    RECT 163.3 34.99 163.51 35.06 ;
    RECT 163.3 35.35 163.51 35.42 ;
    RECT 160.44 34.63 160.65 34.7 ;
    RECT 160.44 34.99 160.65 35.06 ;
    RECT 160.44 35.35 160.65 35.42 ;
    RECT 159.98 34.63 160.19 34.7 ;
    RECT 159.98 34.99 160.19 35.06 ;
    RECT 159.98 35.35 160.19 35.42 ;
    RECT 157.12 34.63 157.33 34.7 ;
    RECT 157.12 34.99 157.33 35.06 ;
    RECT 157.12 35.35 157.33 35.42 ;
    RECT 156.66 34.63 156.87 34.7 ;
    RECT 156.66 34.99 156.87 35.06 ;
    RECT 156.66 35.35 156.87 35.42 ;
    RECT 153.8 34.63 154.01 34.7 ;
    RECT 153.8 34.99 154.01 35.06 ;
    RECT 153.8 35.35 154.01 35.42 ;
    RECT 153.34 34.63 153.55 34.7 ;
    RECT 153.34 34.99 153.55 35.06 ;
    RECT 153.34 35.35 153.55 35.42 ;
    RECT 150.48 34.63 150.69 34.7 ;
    RECT 150.48 34.99 150.69 35.06 ;
    RECT 150.48 35.35 150.69 35.42 ;
    RECT 150.02 34.63 150.23 34.7 ;
    RECT 150.02 34.99 150.23 35.06 ;
    RECT 150.02 35.35 150.23 35.42 ;
    RECT 213.56 34.63 213.77 34.7 ;
    RECT 213.56 34.99 213.77 35.06 ;
    RECT 213.56 35.35 213.77 35.42 ;
    RECT 213.1 34.63 213.31 34.7 ;
    RECT 213.1 34.99 213.31 35.06 ;
    RECT 213.1 35.35 213.31 35.42 ;
    RECT 210.24 34.63 210.45 34.7 ;
    RECT 210.24 34.99 210.45 35.06 ;
    RECT 210.24 35.35 210.45 35.42 ;
    RECT 209.78 34.63 209.99 34.7 ;
    RECT 209.78 34.99 209.99 35.06 ;
    RECT 209.78 35.35 209.99 35.42 ;
    RECT 206.92 34.63 207.13 34.7 ;
    RECT 206.92 34.99 207.13 35.06 ;
    RECT 206.92 35.35 207.13 35.42 ;
    RECT 206.46 34.63 206.67 34.7 ;
    RECT 206.46 34.99 206.67 35.06 ;
    RECT 206.46 35.35 206.67 35.42 ;
    RECT 203.6 34.63 203.81 34.7 ;
    RECT 203.6 34.99 203.81 35.06 ;
    RECT 203.6 35.35 203.81 35.42 ;
    RECT 203.14 34.63 203.35 34.7 ;
    RECT 203.14 34.99 203.35 35.06 ;
    RECT 203.14 35.35 203.35 35.42 ;
    RECT 200.28 34.63 200.49 34.7 ;
    RECT 200.28 34.99 200.49 35.06 ;
    RECT 200.28 35.35 200.49 35.42 ;
    RECT 199.82 34.63 200.03 34.7 ;
    RECT 199.82 34.99 200.03 35.06 ;
    RECT 199.82 35.35 200.03 35.42 ;
    RECT 196.96 34.63 197.17 34.7 ;
    RECT 196.96 34.99 197.17 35.06 ;
    RECT 196.96 35.35 197.17 35.42 ;
    RECT 196.5 34.63 196.71 34.7 ;
    RECT 196.5 34.99 196.71 35.06 ;
    RECT 196.5 35.35 196.71 35.42 ;
    RECT 193.64 34.63 193.85 34.7 ;
    RECT 193.64 34.99 193.85 35.06 ;
    RECT 193.64 35.35 193.85 35.42 ;
    RECT 193.18 34.63 193.39 34.7 ;
    RECT 193.18 34.99 193.39 35.06 ;
    RECT 193.18 35.35 193.39 35.42 ;
    RECT 190.32 34.63 190.53 34.7 ;
    RECT 190.32 34.99 190.53 35.06 ;
    RECT 190.32 35.35 190.53 35.42 ;
    RECT 189.86 34.63 190.07 34.7 ;
    RECT 189.86 34.99 190.07 35.06 ;
    RECT 189.86 35.35 190.07 35.42 ;
    RECT 187.0 34.63 187.21 34.7 ;
    RECT 187.0 34.99 187.21 35.06 ;
    RECT 187.0 35.35 187.21 35.42 ;
    RECT 186.54 34.63 186.75 34.7 ;
    RECT 186.54 34.99 186.75 35.06 ;
    RECT 186.54 35.35 186.75 35.42 ;
    RECT 183.68 34.63 183.89 34.7 ;
    RECT 183.68 34.99 183.89 35.06 ;
    RECT 183.68 35.35 183.89 35.42 ;
    RECT 183.22 34.63 183.43 34.7 ;
    RECT 183.22 34.99 183.43 35.06 ;
    RECT 183.22 35.35 183.43 35.42 ;
    RECT 147.485 34.99 147.555 35.06 ;
    RECT 266.68 34.63 266.89 34.7 ;
    RECT 266.68 34.99 266.89 35.06 ;
    RECT 266.68 35.35 266.89 35.42 ;
    RECT 266.22 34.63 266.43 34.7 ;
    RECT 266.22 34.99 266.43 35.06 ;
    RECT 266.22 35.35 266.43 35.42 ;
    RECT 263.36 34.63 263.57 34.7 ;
    RECT 263.36 34.99 263.57 35.06 ;
    RECT 263.36 35.35 263.57 35.42 ;
    RECT 262.9 34.63 263.11 34.7 ;
    RECT 262.9 34.99 263.11 35.06 ;
    RECT 262.9 35.35 263.11 35.42 ;
    RECT 260.04 34.63 260.25 34.7 ;
    RECT 260.04 34.99 260.25 35.06 ;
    RECT 260.04 35.35 260.25 35.42 ;
    RECT 259.58 34.63 259.79 34.7 ;
    RECT 259.58 34.99 259.79 35.06 ;
    RECT 259.58 35.35 259.79 35.42 ;
    RECT 256.72 34.63 256.93 34.7 ;
    RECT 256.72 34.99 256.93 35.06 ;
    RECT 256.72 35.35 256.93 35.42 ;
    RECT 256.26 34.63 256.47 34.7 ;
    RECT 256.26 34.99 256.47 35.06 ;
    RECT 256.26 35.35 256.47 35.42 ;
    RECT 253.4 34.63 253.61 34.7 ;
    RECT 253.4 34.99 253.61 35.06 ;
    RECT 253.4 35.35 253.61 35.42 ;
    RECT 252.94 34.63 253.15 34.7 ;
    RECT 252.94 34.99 253.15 35.06 ;
    RECT 252.94 35.35 253.15 35.42 ;
    RECT 250.08 18.07 250.29 18.14 ;
    RECT 250.08 18.43 250.29 18.5 ;
    RECT 250.08 18.79 250.29 18.86 ;
    RECT 249.62 18.07 249.83 18.14 ;
    RECT 249.62 18.43 249.83 18.5 ;
    RECT 249.62 18.79 249.83 18.86 ;
    RECT 246.76 18.07 246.97 18.14 ;
    RECT 246.76 18.43 246.97 18.5 ;
    RECT 246.76 18.79 246.97 18.86 ;
    RECT 246.3 18.07 246.51 18.14 ;
    RECT 246.3 18.43 246.51 18.5 ;
    RECT 246.3 18.79 246.51 18.86 ;
    RECT 243.44 18.07 243.65 18.14 ;
    RECT 243.44 18.43 243.65 18.5 ;
    RECT 243.44 18.79 243.65 18.86 ;
    RECT 242.98 18.07 243.19 18.14 ;
    RECT 242.98 18.43 243.19 18.5 ;
    RECT 242.98 18.79 243.19 18.86 ;
    RECT 240.12 18.07 240.33 18.14 ;
    RECT 240.12 18.43 240.33 18.5 ;
    RECT 240.12 18.79 240.33 18.86 ;
    RECT 239.66 18.07 239.87 18.14 ;
    RECT 239.66 18.43 239.87 18.5 ;
    RECT 239.66 18.79 239.87 18.86 ;
    RECT 236.8 18.07 237.01 18.14 ;
    RECT 236.8 18.43 237.01 18.5 ;
    RECT 236.8 18.79 237.01 18.86 ;
    RECT 236.34 18.07 236.55 18.14 ;
    RECT 236.34 18.43 236.55 18.5 ;
    RECT 236.34 18.79 236.55 18.86 ;
    RECT 233.48 18.07 233.69 18.14 ;
    RECT 233.48 18.43 233.69 18.5 ;
    RECT 233.48 18.79 233.69 18.86 ;
    RECT 233.02 18.07 233.23 18.14 ;
    RECT 233.02 18.43 233.23 18.5 ;
    RECT 233.02 18.79 233.23 18.86 ;
    RECT 230.16 18.07 230.37 18.14 ;
    RECT 230.16 18.43 230.37 18.5 ;
    RECT 230.16 18.79 230.37 18.86 ;
    RECT 229.7 18.07 229.91 18.14 ;
    RECT 229.7 18.43 229.91 18.5 ;
    RECT 229.7 18.79 229.91 18.86 ;
    RECT 226.84 18.07 227.05 18.14 ;
    RECT 226.84 18.43 227.05 18.5 ;
    RECT 226.84 18.79 227.05 18.86 ;
    RECT 226.38 18.07 226.59 18.14 ;
    RECT 226.38 18.43 226.59 18.5 ;
    RECT 226.38 18.79 226.59 18.86 ;
    RECT 223.52 18.07 223.73 18.14 ;
    RECT 223.52 18.43 223.73 18.5 ;
    RECT 223.52 18.79 223.73 18.86 ;
    RECT 223.06 18.07 223.27 18.14 ;
    RECT 223.06 18.43 223.27 18.5 ;
    RECT 223.06 18.79 223.27 18.86 ;
    RECT 220.2 18.07 220.41 18.14 ;
    RECT 220.2 18.43 220.41 18.5 ;
    RECT 220.2 18.79 220.41 18.86 ;
    RECT 219.74 18.07 219.95 18.14 ;
    RECT 219.74 18.43 219.95 18.5 ;
    RECT 219.74 18.79 219.95 18.86 ;
    RECT 216.88 18.07 217.09 18.14 ;
    RECT 216.88 18.43 217.09 18.5 ;
    RECT 216.88 18.79 217.09 18.86 ;
    RECT 216.42 18.07 216.63 18.14 ;
    RECT 216.42 18.43 216.63 18.5 ;
    RECT 216.42 18.79 216.63 18.86 ;
    RECT 267.91 18.43 267.98 18.5 ;
    RECT 180.36 18.07 180.57 18.14 ;
    RECT 180.36 18.43 180.57 18.5 ;
    RECT 180.36 18.79 180.57 18.86 ;
    RECT 179.9 18.07 180.11 18.14 ;
    RECT 179.9 18.43 180.11 18.5 ;
    RECT 179.9 18.79 180.11 18.86 ;
    RECT 177.04 18.07 177.25 18.14 ;
    RECT 177.04 18.43 177.25 18.5 ;
    RECT 177.04 18.79 177.25 18.86 ;
    RECT 176.58 18.07 176.79 18.14 ;
    RECT 176.58 18.43 176.79 18.5 ;
    RECT 176.58 18.79 176.79 18.86 ;
    RECT 173.72 18.07 173.93 18.14 ;
    RECT 173.72 18.43 173.93 18.5 ;
    RECT 173.72 18.79 173.93 18.86 ;
    RECT 173.26 18.07 173.47 18.14 ;
    RECT 173.26 18.43 173.47 18.5 ;
    RECT 173.26 18.79 173.47 18.86 ;
    RECT 170.4 18.07 170.61 18.14 ;
    RECT 170.4 18.43 170.61 18.5 ;
    RECT 170.4 18.79 170.61 18.86 ;
    RECT 169.94 18.07 170.15 18.14 ;
    RECT 169.94 18.43 170.15 18.5 ;
    RECT 169.94 18.79 170.15 18.86 ;
    RECT 167.08 18.07 167.29 18.14 ;
    RECT 167.08 18.43 167.29 18.5 ;
    RECT 167.08 18.79 167.29 18.86 ;
    RECT 166.62 18.07 166.83 18.14 ;
    RECT 166.62 18.43 166.83 18.5 ;
    RECT 166.62 18.79 166.83 18.86 ;
    RECT 163.76 18.07 163.97 18.14 ;
    RECT 163.76 18.43 163.97 18.5 ;
    RECT 163.76 18.79 163.97 18.86 ;
    RECT 163.3 18.07 163.51 18.14 ;
    RECT 163.3 18.43 163.51 18.5 ;
    RECT 163.3 18.79 163.51 18.86 ;
    RECT 160.44 18.07 160.65 18.14 ;
    RECT 160.44 18.43 160.65 18.5 ;
    RECT 160.44 18.79 160.65 18.86 ;
    RECT 159.98 18.07 160.19 18.14 ;
    RECT 159.98 18.43 160.19 18.5 ;
    RECT 159.98 18.79 160.19 18.86 ;
    RECT 157.12 18.07 157.33 18.14 ;
    RECT 157.12 18.43 157.33 18.5 ;
    RECT 157.12 18.79 157.33 18.86 ;
    RECT 156.66 18.07 156.87 18.14 ;
    RECT 156.66 18.43 156.87 18.5 ;
    RECT 156.66 18.79 156.87 18.86 ;
    RECT 153.8 18.07 154.01 18.14 ;
    RECT 153.8 18.43 154.01 18.5 ;
    RECT 153.8 18.79 154.01 18.86 ;
    RECT 153.34 18.07 153.55 18.14 ;
    RECT 153.34 18.43 153.55 18.5 ;
    RECT 153.34 18.79 153.55 18.86 ;
    RECT 150.48 18.07 150.69 18.14 ;
    RECT 150.48 18.43 150.69 18.5 ;
    RECT 150.48 18.79 150.69 18.86 ;
    RECT 150.02 18.07 150.23 18.14 ;
    RECT 150.02 18.43 150.23 18.5 ;
    RECT 150.02 18.79 150.23 18.86 ;
    RECT 213.56 18.07 213.77 18.14 ;
    RECT 213.56 18.43 213.77 18.5 ;
    RECT 213.56 18.79 213.77 18.86 ;
    RECT 213.1 18.07 213.31 18.14 ;
    RECT 213.1 18.43 213.31 18.5 ;
    RECT 213.1 18.79 213.31 18.86 ;
    RECT 210.24 18.07 210.45 18.14 ;
    RECT 210.24 18.43 210.45 18.5 ;
    RECT 210.24 18.79 210.45 18.86 ;
    RECT 209.78 18.07 209.99 18.14 ;
    RECT 209.78 18.43 209.99 18.5 ;
    RECT 209.78 18.79 209.99 18.86 ;
    RECT 206.92 18.07 207.13 18.14 ;
    RECT 206.92 18.43 207.13 18.5 ;
    RECT 206.92 18.79 207.13 18.86 ;
    RECT 206.46 18.07 206.67 18.14 ;
    RECT 206.46 18.43 206.67 18.5 ;
    RECT 206.46 18.79 206.67 18.86 ;
    RECT 203.6 18.07 203.81 18.14 ;
    RECT 203.6 18.43 203.81 18.5 ;
    RECT 203.6 18.79 203.81 18.86 ;
    RECT 203.14 18.07 203.35 18.14 ;
    RECT 203.14 18.43 203.35 18.5 ;
    RECT 203.14 18.79 203.35 18.86 ;
    RECT 200.28 18.07 200.49 18.14 ;
    RECT 200.28 18.43 200.49 18.5 ;
    RECT 200.28 18.79 200.49 18.86 ;
    RECT 199.82 18.07 200.03 18.14 ;
    RECT 199.82 18.43 200.03 18.5 ;
    RECT 199.82 18.79 200.03 18.86 ;
    RECT 196.96 18.07 197.17 18.14 ;
    RECT 196.96 18.43 197.17 18.5 ;
    RECT 196.96 18.79 197.17 18.86 ;
    RECT 196.5 18.07 196.71 18.14 ;
    RECT 196.5 18.43 196.71 18.5 ;
    RECT 196.5 18.79 196.71 18.86 ;
    RECT 193.64 18.07 193.85 18.14 ;
    RECT 193.64 18.43 193.85 18.5 ;
    RECT 193.64 18.79 193.85 18.86 ;
    RECT 193.18 18.07 193.39 18.14 ;
    RECT 193.18 18.43 193.39 18.5 ;
    RECT 193.18 18.79 193.39 18.86 ;
    RECT 190.32 18.07 190.53 18.14 ;
    RECT 190.32 18.43 190.53 18.5 ;
    RECT 190.32 18.79 190.53 18.86 ;
    RECT 189.86 18.07 190.07 18.14 ;
    RECT 189.86 18.43 190.07 18.5 ;
    RECT 189.86 18.79 190.07 18.86 ;
    RECT 187.0 18.07 187.21 18.14 ;
    RECT 187.0 18.43 187.21 18.5 ;
    RECT 187.0 18.79 187.21 18.86 ;
    RECT 186.54 18.07 186.75 18.14 ;
    RECT 186.54 18.43 186.75 18.5 ;
    RECT 186.54 18.79 186.75 18.86 ;
    RECT 183.68 18.07 183.89 18.14 ;
    RECT 183.68 18.43 183.89 18.5 ;
    RECT 183.68 18.79 183.89 18.86 ;
    RECT 183.22 18.07 183.43 18.14 ;
    RECT 183.22 18.43 183.43 18.5 ;
    RECT 183.22 18.79 183.43 18.86 ;
    RECT 147.485 18.43 147.555 18.5 ;
    RECT 266.68 18.07 266.89 18.14 ;
    RECT 266.68 18.43 266.89 18.5 ;
    RECT 266.68 18.79 266.89 18.86 ;
    RECT 266.22 18.07 266.43 18.14 ;
    RECT 266.22 18.43 266.43 18.5 ;
    RECT 266.22 18.79 266.43 18.86 ;
    RECT 263.36 18.07 263.57 18.14 ;
    RECT 263.36 18.43 263.57 18.5 ;
    RECT 263.36 18.79 263.57 18.86 ;
    RECT 262.9 18.07 263.11 18.14 ;
    RECT 262.9 18.43 263.11 18.5 ;
    RECT 262.9 18.79 263.11 18.86 ;
    RECT 260.04 18.07 260.25 18.14 ;
    RECT 260.04 18.43 260.25 18.5 ;
    RECT 260.04 18.79 260.25 18.86 ;
    RECT 259.58 18.07 259.79 18.14 ;
    RECT 259.58 18.43 259.79 18.5 ;
    RECT 259.58 18.79 259.79 18.86 ;
    RECT 256.72 18.07 256.93 18.14 ;
    RECT 256.72 18.43 256.93 18.5 ;
    RECT 256.72 18.79 256.93 18.86 ;
    RECT 256.26 18.07 256.47 18.14 ;
    RECT 256.26 18.43 256.47 18.5 ;
    RECT 256.26 18.79 256.47 18.86 ;
    RECT 253.4 18.07 253.61 18.14 ;
    RECT 253.4 18.43 253.61 18.5 ;
    RECT 253.4 18.79 253.61 18.86 ;
    RECT 252.94 18.07 253.15 18.14 ;
    RECT 252.94 18.43 253.15 18.5 ;
    RECT 252.94 18.79 253.15 18.86 ;
    RECT 250.08 33.91 250.29 33.98 ;
    RECT 250.08 34.27 250.29 34.34 ;
    RECT 250.08 34.63 250.29 34.7 ;
    RECT 249.62 33.91 249.83 33.98 ;
    RECT 249.62 34.27 249.83 34.34 ;
    RECT 249.62 34.63 249.83 34.7 ;
    RECT 246.76 33.91 246.97 33.98 ;
    RECT 246.76 34.27 246.97 34.34 ;
    RECT 246.76 34.63 246.97 34.7 ;
    RECT 246.3 33.91 246.51 33.98 ;
    RECT 246.3 34.27 246.51 34.34 ;
    RECT 246.3 34.63 246.51 34.7 ;
    RECT 243.44 33.91 243.65 33.98 ;
    RECT 243.44 34.27 243.65 34.34 ;
    RECT 243.44 34.63 243.65 34.7 ;
    RECT 242.98 33.91 243.19 33.98 ;
    RECT 242.98 34.27 243.19 34.34 ;
    RECT 242.98 34.63 243.19 34.7 ;
    RECT 240.12 33.91 240.33 33.98 ;
    RECT 240.12 34.27 240.33 34.34 ;
    RECT 240.12 34.63 240.33 34.7 ;
    RECT 239.66 33.91 239.87 33.98 ;
    RECT 239.66 34.27 239.87 34.34 ;
    RECT 239.66 34.63 239.87 34.7 ;
    RECT 236.8 33.91 237.01 33.98 ;
    RECT 236.8 34.27 237.01 34.34 ;
    RECT 236.8 34.63 237.01 34.7 ;
    RECT 236.34 33.91 236.55 33.98 ;
    RECT 236.34 34.27 236.55 34.34 ;
    RECT 236.34 34.63 236.55 34.7 ;
    RECT 233.48 33.91 233.69 33.98 ;
    RECT 233.48 34.27 233.69 34.34 ;
    RECT 233.48 34.63 233.69 34.7 ;
    RECT 233.02 33.91 233.23 33.98 ;
    RECT 233.02 34.27 233.23 34.34 ;
    RECT 233.02 34.63 233.23 34.7 ;
    RECT 230.16 33.91 230.37 33.98 ;
    RECT 230.16 34.27 230.37 34.34 ;
    RECT 230.16 34.63 230.37 34.7 ;
    RECT 229.7 33.91 229.91 33.98 ;
    RECT 229.7 34.27 229.91 34.34 ;
    RECT 229.7 34.63 229.91 34.7 ;
    RECT 226.84 33.91 227.05 33.98 ;
    RECT 226.84 34.27 227.05 34.34 ;
    RECT 226.84 34.63 227.05 34.7 ;
    RECT 226.38 33.91 226.59 33.98 ;
    RECT 226.38 34.27 226.59 34.34 ;
    RECT 226.38 34.63 226.59 34.7 ;
    RECT 223.52 33.91 223.73 33.98 ;
    RECT 223.52 34.27 223.73 34.34 ;
    RECT 223.52 34.63 223.73 34.7 ;
    RECT 223.06 33.91 223.27 33.98 ;
    RECT 223.06 34.27 223.27 34.34 ;
    RECT 223.06 34.63 223.27 34.7 ;
    RECT 220.2 33.91 220.41 33.98 ;
    RECT 220.2 34.27 220.41 34.34 ;
    RECT 220.2 34.63 220.41 34.7 ;
    RECT 219.74 33.91 219.95 33.98 ;
    RECT 219.74 34.27 219.95 34.34 ;
    RECT 219.74 34.63 219.95 34.7 ;
    RECT 216.88 33.91 217.09 33.98 ;
    RECT 216.88 34.27 217.09 34.34 ;
    RECT 216.88 34.63 217.09 34.7 ;
    RECT 216.42 33.91 216.63 33.98 ;
    RECT 216.42 34.27 216.63 34.34 ;
    RECT 216.42 34.63 216.63 34.7 ;
    RECT 267.91 34.27 267.98 34.34 ;
    RECT 180.36 33.91 180.57 33.98 ;
    RECT 180.36 34.27 180.57 34.34 ;
    RECT 180.36 34.63 180.57 34.7 ;
    RECT 179.9 33.91 180.11 33.98 ;
    RECT 179.9 34.27 180.11 34.34 ;
    RECT 179.9 34.63 180.11 34.7 ;
    RECT 177.04 33.91 177.25 33.98 ;
    RECT 177.04 34.27 177.25 34.34 ;
    RECT 177.04 34.63 177.25 34.7 ;
    RECT 176.58 33.91 176.79 33.98 ;
    RECT 176.58 34.27 176.79 34.34 ;
    RECT 176.58 34.63 176.79 34.7 ;
    RECT 173.72 33.91 173.93 33.98 ;
    RECT 173.72 34.27 173.93 34.34 ;
    RECT 173.72 34.63 173.93 34.7 ;
    RECT 173.26 33.91 173.47 33.98 ;
    RECT 173.26 34.27 173.47 34.34 ;
    RECT 173.26 34.63 173.47 34.7 ;
    RECT 170.4 33.91 170.61 33.98 ;
    RECT 170.4 34.27 170.61 34.34 ;
    RECT 170.4 34.63 170.61 34.7 ;
    RECT 169.94 33.91 170.15 33.98 ;
    RECT 169.94 34.27 170.15 34.34 ;
    RECT 169.94 34.63 170.15 34.7 ;
    RECT 167.08 33.91 167.29 33.98 ;
    RECT 167.08 34.27 167.29 34.34 ;
    RECT 167.08 34.63 167.29 34.7 ;
    RECT 166.62 33.91 166.83 33.98 ;
    RECT 166.62 34.27 166.83 34.34 ;
    RECT 166.62 34.63 166.83 34.7 ;
    RECT 163.76 33.91 163.97 33.98 ;
    RECT 163.76 34.27 163.97 34.34 ;
    RECT 163.76 34.63 163.97 34.7 ;
    RECT 163.3 33.91 163.51 33.98 ;
    RECT 163.3 34.27 163.51 34.34 ;
    RECT 163.3 34.63 163.51 34.7 ;
    RECT 160.44 33.91 160.65 33.98 ;
    RECT 160.44 34.27 160.65 34.34 ;
    RECT 160.44 34.63 160.65 34.7 ;
    RECT 159.98 33.91 160.19 33.98 ;
    RECT 159.98 34.27 160.19 34.34 ;
    RECT 159.98 34.63 160.19 34.7 ;
    RECT 157.12 33.91 157.33 33.98 ;
    RECT 157.12 34.27 157.33 34.34 ;
    RECT 157.12 34.63 157.33 34.7 ;
    RECT 156.66 33.91 156.87 33.98 ;
    RECT 156.66 34.27 156.87 34.34 ;
    RECT 156.66 34.63 156.87 34.7 ;
    RECT 153.8 33.91 154.01 33.98 ;
    RECT 153.8 34.27 154.01 34.34 ;
    RECT 153.8 34.63 154.01 34.7 ;
    RECT 153.34 33.91 153.55 33.98 ;
    RECT 153.34 34.27 153.55 34.34 ;
    RECT 153.34 34.63 153.55 34.7 ;
    RECT 150.48 33.91 150.69 33.98 ;
    RECT 150.48 34.27 150.69 34.34 ;
    RECT 150.48 34.63 150.69 34.7 ;
    RECT 150.02 33.91 150.23 33.98 ;
    RECT 150.02 34.27 150.23 34.34 ;
    RECT 150.02 34.63 150.23 34.7 ;
    RECT 213.56 33.91 213.77 33.98 ;
    RECT 213.56 34.27 213.77 34.34 ;
    RECT 213.56 34.63 213.77 34.7 ;
    RECT 213.1 33.91 213.31 33.98 ;
    RECT 213.1 34.27 213.31 34.34 ;
    RECT 213.1 34.63 213.31 34.7 ;
    RECT 210.24 33.91 210.45 33.98 ;
    RECT 210.24 34.27 210.45 34.34 ;
    RECT 210.24 34.63 210.45 34.7 ;
    RECT 209.78 33.91 209.99 33.98 ;
    RECT 209.78 34.27 209.99 34.34 ;
    RECT 209.78 34.63 209.99 34.7 ;
    RECT 206.92 33.91 207.13 33.98 ;
    RECT 206.92 34.27 207.13 34.34 ;
    RECT 206.92 34.63 207.13 34.7 ;
    RECT 206.46 33.91 206.67 33.98 ;
    RECT 206.46 34.27 206.67 34.34 ;
    RECT 206.46 34.63 206.67 34.7 ;
    RECT 203.6 33.91 203.81 33.98 ;
    RECT 203.6 34.27 203.81 34.34 ;
    RECT 203.6 34.63 203.81 34.7 ;
    RECT 203.14 33.91 203.35 33.98 ;
    RECT 203.14 34.27 203.35 34.34 ;
    RECT 203.14 34.63 203.35 34.7 ;
    RECT 200.28 33.91 200.49 33.98 ;
    RECT 200.28 34.27 200.49 34.34 ;
    RECT 200.28 34.63 200.49 34.7 ;
    RECT 199.82 33.91 200.03 33.98 ;
    RECT 199.82 34.27 200.03 34.34 ;
    RECT 199.82 34.63 200.03 34.7 ;
    RECT 196.96 33.91 197.17 33.98 ;
    RECT 196.96 34.27 197.17 34.34 ;
    RECT 196.96 34.63 197.17 34.7 ;
    RECT 196.5 33.91 196.71 33.98 ;
    RECT 196.5 34.27 196.71 34.34 ;
    RECT 196.5 34.63 196.71 34.7 ;
    RECT 193.64 33.91 193.85 33.98 ;
    RECT 193.64 34.27 193.85 34.34 ;
    RECT 193.64 34.63 193.85 34.7 ;
    RECT 193.18 33.91 193.39 33.98 ;
    RECT 193.18 34.27 193.39 34.34 ;
    RECT 193.18 34.63 193.39 34.7 ;
    RECT 190.32 33.91 190.53 33.98 ;
    RECT 190.32 34.27 190.53 34.34 ;
    RECT 190.32 34.63 190.53 34.7 ;
    RECT 189.86 33.91 190.07 33.98 ;
    RECT 189.86 34.27 190.07 34.34 ;
    RECT 189.86 34.63 190.07 34.7 ;
    RECT 187.0 33.91 187.21 33.98 ;
    RECT 187.0 34.27 187.21 34.34 ;
    RECT 187.0 34.63 187.21 34.7 ;
    RECT 186.54 33.91 186.75 33.98 ;
    RECT 186.54 34.27 186.75 34.34 ;
    RECT 186.54 34.63 186.75 34.7 ;
    RECT 183.68 33.91 183.89 33.98 ;
    RECT 183.68 34.27 183.89 34.34 ;
    RECT 183.68 34.63 183.89 34.7 ;
    RECT 183.22 33.91 183.43 33.98 ;
    RECT 183.22 34.27 183.43 34.34 ;
    RECT 183.22 34.63 183.43 34.7 ;
    RECT 147.485 34.27 147.555 34.34 ;
    RECT 266.68 33.91 266.89 33.98 ;
    RECT 266.68 34.27 266.89 34.34 ;
    RECT 266.68 34.63 266.89 34.7 ;
    RECT 266.22 33.91 266.43 33.98 ;
    RECT 266.22 34.27 266.43 34.34 ;
    RECT 266.22 34.63 266.43 34.7 ;
    RECT 263.36 33.91 263.57 33.98 ;
    RECT 263.36 34.27 263.57 34.34 ;
    RECT 263.36 34.63 263.57 34.7 ;
    RECT 262.9 33.91 263.11 33.98 ;
    RECT 262.9 34.27 263.11 34.34 ;
    RECT 262.9 34.63 263.11 34.7 ;
    RECT 260.04 33.91 260.25 33.98 ;
    RECT 260.04 34.27 260.25 34.34 ;
    RECT 260.04 34.63 260.25 34.7 ;
    RECT 259.58 33.91 259.79 33.98 ;
    RECT 259.58 34.27 259.79 34.34 ;
    RECT 259.58 34.63 259.79 34.7 ;
    RECT 256.72 33.91 256.93 33.98 ;
    RECT 256.72 34.27 256.93 34.34 ;
    RECT 256.72 34.63 256.93 34.7 ;
    RECT 256.26 33.91 256.47 33.98 ;
    RECT 256.26 34.27 256.47 34.34 ;
    RECT 256.26 34.63 256.47 34.7 ;
    RECT 253.4 33.91 253.61 33.98 ;
    RECT 253.4 34.27 253.61 34.34 ;
    RECT 253.4 34.63 253.61 34.7 ;
    RECT 252.94 33.91 253.15 33.98 ;
    RECT 252.94 34.27 253.15 34.34 ;
    RECT 252.94 34.63 253.15 34.7 ;
    RECT 250.08 17.35 250.29 17.42 ;
    RECT 250.08 17.71 250.29 17.78 ;
    RECT 250.08 18.07 250.29 18.14 ;
    RECT 249.62 17.35 249.83 17.42 ;
    RECT 249.62 17.71 249.83 17.78 ;
    RECT 249.62 18.07 249.83 18.14 ;
    RECT 246.76 17.35 246.97 17.42 ;
    RECT 246.76 17.71 246.97 17.78 ;
    RECT 246.76 18.07 246.97 18.14 ;
    RECT 246.3 17.35 246.51 17.42 ;
    RECT 246.3 17.71 246.51 17.78 ;
    RECT 246.3 18.07 246.51 18.14 ;
    RECT 243.44 17.35 243.65 17.42 ;
    RECT 243.44 17.71 243.65 17.78 ;
    RECT 243.44 18.07 243.65 18.14 ;
    RECT 242.98 17.35 243.19 17.42 ;
    RECT 242.98 17.71 243.19 17.78 ;
    RECT 242.98 18.07 243.19 18.14 ;
    RECT 240.12 17.35 240.33 17.42 ;
    RECT 240.12 17.71 240.33 17.78 ;
    RECT 240.12 18.07 240.33 18.14 ;
    RECT 239.66 17.35 239.87 17.42 ;
    RECT 239.66 17.71 239.87 17.78 ;
    RECT 239.66 18.07 239.87 18.14 ;
    RECT 236.8 17.35 237.01 17.42 ;
    RECT 236.8 17.71 237.01 17.78 ;
    RECT 236.8 18.07 237.01 18.14 ;
    RECT 236.34 17.35 236.55 17.42 ;
    RECT 236.34 17.71 236.55 17.78 ;
    RECT 236.34 18.07 236.55 18.14 ;
    RECT 233.48 17.35 233.69 17.42 ;
    RECT 233.48 17.71 233.69 17.78 ;
    RECT 233.48 18.07 233.69 18.14 ;
    RECT 233.02 17.35 233.23 17.42 ;
    RECT 233.02 17.71 233.23 17.78 ;
    RECT 233.02 18.07 233.23 18.14 ;
    RECT 230.16 17.35 230.37 17.42 ;
    RECT 230.16 17.71 230.37 17.78 ;
    RECT 230.16 18.07 230.37 18.14 ;
    RECT 229.7 17.35 229.91 17.42 ;
    RECT 229.7 17.71 229.91 17.78 ;
    RECT 229.7 18.07 229.91 18.14 ;
    RECT 226.84 17.35 227.05 17.42 ;
    RECT 226.84 17.71 227.05 17.78 ;
    RECT 226.84 18.07 227.05 18.14 ;
    RECT 226.38 17.35 226.59 17.42 ;
    RECT 226.38 17.71 226.59 17.78 ;
    RECT 226.38 18.07 226.59 18.14 ;
    RECT 223.52 17.35 223.73 17.42 ;
    RECT 223.52 17.71 223.73 17.78 ;
    RECT 223.52 18.07 223.73 18.14 ;
    RECT 223.06 17.35 223.27 17.42 ;
    RECT 223.06 17.71 223.27 17.78 ;
    RECT 223.06 18.07 223.27 18.14 ;
    RECT 220.2 17.35 220.41 17.42 ;
    RECT 220.2 17.71 220.41 17.78 ;
    RECT 220.2 18.07 220.41 18.14 ;
    RECT 219.74 17.35 219.95 17.42 ;
    RECT 219.74 17.71 219.95 17.78 ;
    RECT 219.74 18.07 219.95 18.14 ;
    RECT 216.88 17.35 217.09 17.42 ;
    RECT 216.88 17.71 217.09 17.78 ;
    RECT 216.88 18.07 217.09 18.14 ;
    RECT 216.42 17.35 216.63 17.42 ;
    RECT 216.42 17.71 216.63 17.78 ;
    RECT 216.42 18.07 216.63 18.14 ;
    RECT 267.91 17.71 267.98 17.78 ;
    RECT 180.36 17.35 180.57 17.42 ;
    RECT 180.36 17.71 180.57 17.78 ;
    RECT 180.36 18.07 180.57 18.14 ;
    RECT 179.9 17.35 180.11 17.42 ;
    RECT 179.9 17.71 180.11 17.78 ;
    RECT 179.9 18.07 180.11 18.14 ;
    RECT 177.04 17.35 177.25 17.42 ;
    RECT 177.04 17.71 177.25 17.78 ;
    RECT 177.04 18.07 177.25 18.14 ;
    RECT 176.58 17.35 176.79 17.42 ;
    RECT 176.58 17.71 176.79 17.78 ;
    RECT 176.58 18.07 176.79 18.14 ;
    RECT 173.72 17.35 173.93 17.42 ;
    RECT 173.72 17.71 173.93 17.78 ;
    RECT 173.72 18.07 173.93 18.14 ;
    RECT 173.26 17.35 173.47 17.42 ;
    RECT 173.26 17.71 173.47 17.78 ;
    RECT 173.26 18.07 173.47 18.14 ;
    RECT 170.4 17.35 170.61 17.42 ;
    RECT 170.4 17.71 170.61 17.78 ;
    RECT 170.4 18.07 170.61 18.14 ;
    RECT 169.94 17.35 170.15 17.42 ;
    RECT 169.94 17.71 170.15 17.78 ;
    RECT 169.94 18.07 170.15 18.14 ;
    RECT 167.08 17.35 167.29 17.42 ;
    RECT 167.08 17.71 167.29 17.78 ;
    RECT 167.08 18.07 167.29 18.14 ;
    RECT 166.62 17.35 166.83 17.42 ;
    RECT 166.62 17.71 166.83 17.78 ;
    RECT 166.62 18.07 166.83 18.14 ;
    RECT 163.76 17.35 163.97 17.42 ;
    RECT 163.76 17.71 163.97 17.78 ;
    RECT 163.76 18.07 163.97 18.14 ;
    RECT 163.3 17.35 163.51 17.42 ;
    RECT 163.3 17.71 163.51 17.78 ;
    RECT 163.3 18.07 163.51 18.14 ;
    RECT 160.44 17.35 160.65 17.42 ;
    RECT 160.44 17.71 160.65 17.78 ;
    RECT 160.44 18.07 160.65 18.14 ;
    RECT 159.98 17.35 160.19 17.42 ;
    RECT 159.98 17.71 160.19 17.78 ;
    RECT 159.98 18.07 160.19 18.14 ;
    RECT 157.12 17.35 157.33 17.42 ;
    RECT 157.12 17.71 157.33 17.78 ;
    RECT 157.12 18.07 157.33 18.14 ;
    RECT 156.66 17.35 156.87 17.42 ;
    RECT 156.66 17.71 156.87 17.78 ;
    RECT 156.66 18.07 156.87 18.14 ;
    RECT 153.8 17.35 154.01 17.42 ;
    RECT 153.8 17.71 154.01 17.78 ;
    RECT 153.8 18.07 154.01 18.14 ;
    RECT 153.34 17.35 153.55 17.42 ;
    RECT 153.34 17.71 153.55 17.78 ;
    RECT 153.34 18.07 153.55 18.14 ;
    RECT 150.48 17.35 150.69 17.42 ;
    RECT 150.48 17.71 150.69 17.78 ;
    RECT 150.48 18.07 150.69 18.14 ;
    RECT 150.02 17.35 150.23 17.42 ;
    RECT 150.02 17.71 150.23 17.78 ;
    RECT 150.02 18.07 150.23 18.14 ;
    RECT 213.56 17.35 213.77 17.42 ;
    RECT 213.56 17.71 213.77 17.78 ;
    RECT 213.56 18.07 213.77 18.14 ;
    RECT 213.1 17.35 213.31 17.42 ;
    RECT 213.1 17.71 213.31 17.78 ;
    RECT 213.1 18.07 213.31 18.14 ;
    RECT 210.24 17.35 210.45 17.42 ;
    RECT 210.24 17.71 210.45 17.78 ;
    RECT 210.24 18.07 210.45 18.14 ;
    RECT 209.78 17.35 209.99 17.42 ;
    RECT 209.78 17.71 209.99 17.78 ;
    RECT 209.78 18.07 209.99 18.14 ;
    RECT 206.92 17.35 207.13 17.42 ;
    RECT 206.92 17.71 207.13 17.78 ;
    RECT 206.92 18.07 207.13 18.14 ;
    RECT 206.46 17.35 206.67 17.42 ;
    RECT 206.46 17.71 206.67 17.78 ;
    RECT 206.46 18.07 206.67 18.14 ;
    RECT 203.6 17.35 203.81 17.42 ;
    RECT 203.6 17.71 203.81 17.78 ;
    RECT 203.6 18.07 203.81 18.14 ;
    RECT 203.14 17.35 203.35 17.42 ;
    RECT 203.14 17.71 203.35 17.78 ;
    RECT 203.14 18.07 203.35 18.14 ;
    RECT 200.28 17.35 200.49 17.42 ;
    RECT 200.28 17.71 200.49 17.78 ;
    RECT 200.28 18.07 200.49 18.14 ;
    RECT 199.82 17.35 200.03 17.42 ;
    RECT 199.82 17.71 200.03 17.78 ;
    RECT 199.82 18.07 200.03 18.14 ;
    RECT 196.96 17.35 197.17 17.42 ;
    RECT 196.96 17.71 197.17 17.78 ;
    RECT 196.96 18.07 197.17 18.14 ;
    RECT 196.5 17.35 196.71 17.42 ;
    RECT 196.5 17.71 196.71 17.78 ;
    RECT 196.5 18.07 196.71 18.14 ;
    RECT 193.64 17.35 193.85 17.42 ;
    RECT 193.64 17.71 193.85 17.78 ;
    RECT 193.64 18.07 193.85 18.14 ;
    RECT 193.18 17.35 193.39 17.42 ;
    RECT 193.18 17.71 193.39 17.78 ;
    RECT 193.18 18.07 193.39 18.14 ;
    RECT 190.32 17.35 190.53 17.42 ;
    RECT 190.32 17.71 190.53 17.78 ;
    RECT 190.32 18.07 190.53 18.14 ;
    RECT 189.86 17.35 190.07 17.42 ;
    RECT 189.86 17.71 190.07 17.78 ;
    RECT 189.86 18.07 190.07 18.14 ;
    RECT 187.0 17.35 187.21 17.42 ;
    RECT 187.0 17.71 187.21 17.78 ;
    RECT 187.0 18.07 187.21 18.14 ;
    RECT 186.54 17.35 186.75 17.42 ;
    RECT 186.54 17.71 186.75 17.78 ;
    RECT 186.54 18.07 186.75 18.14 ;
    RECT 183.68 17.35 183.89 17.42 ;
    RECT 183.68 17.71 183.89 17.78 ;
    RECT 183.68 18.07 183.89 18.14 ;
    RECT 183.22 17.35 183.43 17.42 ;
    RECT 183.22 17.71 183.43 17.78 ;
    RECT 183.22 18.07 183.43 18.14 ;
    RECT 147.485 17.71 147.555 17.78 ;
    RECT 266.68 17.35 266.89 17.42 ;
    RECT 266.68 17.71 266.89 17.78 ;
    RECT 266.68 18.07 266.89 18.14 ;
    RECT 266.22 17.35 266.43 17.42 ;
    RECT 266.22 17.71 266.43 17.78 ;
    RECT 266.22 18.07 266.43 18.14 ;
    RECT 263.36 17.35 263.57 17.42 ;
    RECT 263.36 17.71 263.57 17.78 ;
    RECT 263.36 18.07 263.57 18.14 ;
    RECT 262.9 17.35 263.11 17.42 ;
    RECT 262.9 17.71 263.11 17.78 ;
    RECT 262.9 18.07 263.11 18.14 ;
    RECT 260.04 17.35 260.25 17.42 ;
    RECT 260.04 17.71 260.25 17.78 ;
    RECT 260.04 18.07 260.25 18.14 ;
    RECT 259.58 17.35 259.79 17.42 ;
    RECT 259.58 17.71 259.79 17.78 ;
    RECT 259.58 18.07 259.79 18.14 ;
    RECT 256.72 17.35 256.93 17.42 ;
    RECT 256.72 17.71 256.93 17.78 ;
    RECT 256.72 18.07 256.93 18.14 ;
    RECT 256.26 17.35 256.47 17.42 ;
    RECT 256.26 17.71 256.47 17.78 ;
    RECT 256.26 18.07 256.47 18.14 ;
    RECT 253.4 17.35 253.61 17.42 ;
    RECT 253.4 17.71 253.61 17.78 ;
    RECT 253.4 18.07 253.61 18.14 ;
    RECT 252.94 17.35 253.15 17.42 ;
    RECT 252.94 17.71 253.15 17.78 ;
    RECT 252.94 18.07 253.15 18.14 ;
    RECT 250.08 33.19 250.29 33.26 ;
    RECT 250.08 33.55 250.29 33.62 ;
    RECT 250.08 33.91 250.29 33.98 ;
    RECT 249.62 33.19 249.83 33.26 ;
    RECT 249.62 33.55 249.83 33.62 ;
    RECT 249.62 33.91 249.83 33.98 ;
    RECT 246.76 33.19 246.97 33.26 ;
    RECT 246.76 33.55 246.97 33.62 ;
    RECT 246.76 33.91 246.97 33.98 ;
    RECT 246.3 33.19 246.51 33.26 ;
    RECT 246.3 33.55 246.51 33.62 ;
    RECT 246.3 33.91 246.51 33.98 ;
    RECT 243.44 33.19 243.65 33.26 ;
    RECT 243.44 33.55 243.65 33.62 ;
    RECT 243.44 33.91 243.65 33.98 ;
    RECT 242.98 33.19 243.19 33.26 ;
    RECT 242.98 33.55 243.19 33.62 ;
    RECT 242.98 33.91 243.19 33.98 ;
    RECT 240.12 33.19 240.33 33.26 ;
    RECT 240.12 33.55 240.33 33.62 ;
    RECT 240.12 33.91 240.33 33.98 ;
    RECT 239.66 33.19 239.87 33.26 ;
    RECT 239.66 33.55 239.87 33.62 ;
    RECT 239.66 33.91 239.87 33.98 ;
    RECT 236.8 33.19 237.01 33.26 ;
    RECT 236.8 33.55 237.01 33.62 ;
    RECT 236.8 33.91 237.01 33.98 ;
    RECT 236.34 33.19 236.55 33.26 ;
    RECT 236.34 33.55 236.55 33.62 ;
    RECT 236.34 33.91 236.55 33.98 ;
    RECT 233.48 33.19 233.69 33.26 ;
    RECT 233.48 33.55 233.69 33.62 ;
    RECT 233.48 33.91 233.69 33.98 ;
    RECT 233.02 33.19 233.23 33.26 ;
    RECT 233.02 33.55 233.23 33.62 ;
    RECT 233.02 33.91 233.23 33.98 ;
    RECT 230.16 33.19 230.37 33.26 ;
    RECT 230.16 33.55 230.37 33.62 ;
    RECT 230.16 33.91 230.37 33.98 ;
    RECT 229.7 33.19 229.91 33.26 ;
    RECT 229.7 33.55 229.91 33.62 ;
    RECT 229.7 33.91 229.91 33.98 ;
    RECT 226.84 33.19 227.05 33.26 ;
    RECT 226.84 33.55 227.05 33.62 ;
    RECT 226.84 33.91 227.05 33.98 ;
    RECT 226.38 33.19 226.59 33.26 ;
    RECT 226.38 33.55 226.59 33.62 ;
    RECT 226.38 33.91 226.59 33.98 ;
    RECT 223.52 33.19 223.73 33.26 ;
    RECT 223.52 33.55 223.73 33.62 ;
    RECT 223.52 33.91 223.73 33.98 ;
    RECT 223.06 33.19 223.27 33.26 ;
    RECT 223.06 33.55 223.27 33.62 ;
    RECT 223.06 33.91 223.27 33.98 ;
    RECT 220.2 33.19 220.41 33.26 ;
    RECT 220.2 33.55 220.41 33.62 ;
    RECT 220.2 33.91 220.41 33.98 ;
    RECT 219.74 33.19 219.95 33.26 ;
    RECT 219.74 33.55 219.95 33.62 ;
    RECT 219.74 33.91 219.95 33.98 ;
    RECT 216.88 33.19 217.09 33.26 ;
    RECT 216.88 33.55 217.09 33.62 ;
    RECT 216.88 33.91 217.09 33.98 ;
    RECT 216.42 33.19 216.63 33.26 ;
    RECT 216.42 33.55 216.63 33.62 ;
    RECT 216.42 33.91 216.63 33.98 ;
    RECT 267.91 33.55 267.98 33.62 ;
    RECT 180.36 33.19 180.57 33.26 ;
    RECT 180.36 33.55 180.57 33.62 ;
    RECT 180.36 33.91 180.57 33.98 ;
    RECT 179.9 33.19 180.11 33.26 ;
    RECT 179.9 33.55 180.11 33.62 ;
    RECT 179.9 33.91 180.11 33.98 ;
    RECT 177.04 33.19 177.25 33.26 ;
    RECT 177.04 33.55 177.25 33.62 ;
    RECT 177.04 33.91 177.25 33.98 ;
    RECT 176.58 33.19 176.79 33.26 ;
    RECT 176.58 33.55 176.79 33.62 ;
    RECT 176.58 33.91 176.79 33.98 ;
    RECT 173.72 33.19 173.93 33.26 ;
    RECT 173.72 33.55 173.93 33.62 ;
    RECT 173.72 33.91 173.93 33.98 ;
    RECT 173.26 33.19 173.47 33.26 ;
    RECT 173.26 33.55 173.47 33.62 ;
    RECT 173.26 33.91 173.47 33.98 ;
    RECT 170.4 33.19 170.61 33.26 ;
    RECT 170.4 33.55 170.61 33.62 ;
    RECT 170.4 33.91 170.61 33.98 ;
    RECT 169.94 33.19 170.15 33.26 ;
    RECT 169.94 33.55 170.15 33.62 ;
    RECT 169.94 33.91 170.15 33.98 ;
    RECT 167.08 33.19 167.29 33.26 ;
    RECT 167.08 33.55 167.29 33.62 ;
    RECT 167.08 33.91 167.29 33.98 ;
    RECT 166.62 33.19 166.83 33.26 ;
    RECT 166.62 33.55 166.83 33.62 ;
    RECT 166.62 33.91 166.83 33.98 ;
    RECT 163.76 33.19 163.97 33.26 ;
    RECT 163.76 33.55 163.97 33.62 ;
    RECT 163.76 33.91 163.97 33.98 ;
    RECT 163.3 33.19 163.51 33.26 ;
    RECT 163.3 33.55 163.51 33.62 ;
    RECT 163.3 33.91 163.51 33.98 ;
    RECT 160.44 33.19 160.65 33.26 ;
    RECT 160.44 33.55 160.65 33.62 ;
    RECT 160.44 33.91 160.65 33.98 ;
    RECT 159.98 33.19 160.19 33.26 ;
    RECT 159.98 33.55 160.19 33.62 ;
    RECT 159.98 33.91 160.19 33.98 ;
    RECT 157.12 33.19 157.33 33.26 ;
    RECT 157.12 33.55 157.33 33.62 ;
    RECT 157.12 33.91 157.33 33.98 ;
    RECT 156.66 33.19 156.87 33.26 ;
    RECT 156.66 33.55 156.87 33.62 ;
    RECT 156.66 33.91 156.87 33.98 ;
    RECT 153.8 33.19 154.01 33.26 ;
    RECT 153.8 33.55 154.01 33.62 ;
    RECT 153.8 33.91 154.01 33.98 ;
    RECT 153.34 33.19 153.55 33.26 ;
    RECT 153.34 33.55 153.55 33.62 ;
    RECT 153.34 33.91 153.55 33.98 ;
    RECT 150.48 33.19 150.69 33.26 ;
    RECT 150.48 33.55 150.69 33.62 ;
    RECT 150.48 33.91 150.69 33.98 ;
    RECT 150.02 33.19 150.23 33.26 ;
    RECT 150.02 33.55 150.23 33.62 ;
    RECT 150.02 33.91 150.23 33.98 ;
    RECT 213.56 33.19 213.77 33.26 ;
    RECT 213.56 33.55 213.77 33.62 ;
    RECT 213.56 33.91 213.77 33.98 ;
    RECT 213.1 33.19 213.31 33.26 ;
    RECT 213.1 33.55 213.31 33.62 ;
    RECT 213.1 33.91 213.31 33.98 ;
    RECT 210.24 33.19 210.45 33.26 ;
    RECT 210.24 33.55 210.45 33.62 ;
    RECT 210.24 33.91 210.45 33.98 ;
    RECT 209.78 33.19 209.99 33.26 ;
    RECT 209.78 33.55 209.99 33.62 ;
    RECT 209.78 33.91 209.99 33.98 ;
    RECT 206.92 33.19 207.13 33.26 ;
    RECT 206.92 33.55 207.13 33.62 ;
    RECT 206.92 33.91 207.13 33.98 ;
    RECT 206.46 33.19 206.67 33.26 ;
    RECT 206.46 33.55 206.67 33.62 ;
    RECT 206.46 33.91 206.67 33.98 ;
    RECT 203.6 33.19 203.81 33.26 ;
    RECT 203.6 33.55 203.81 33.62 ;
    RECT 203.6 33.91 203.81 33.98 ;
    RECT 203.14 33.19 203.35 33.26 ;
    RECT 203.14 33.55 203.35 33.62 ;
    RECT 203.14 33.91 203.35 33.98 ;
    RECT 200.28 33.19 200.49 33.26 ;
    RECT 200.28 33.55 200.49 33.62 ;
    RECT 200.28 33.91 200.49 33.98 ;
    RECT 199.82 33.19 200.03 33.26 ;
    RECT 199.82 33.55 200.03 33.62 ;
    RECT 199.82 33.91 200.03 33.98 ;
    RECT 196.96 33.19 197.17 33.26 ;
    RECT 196.96 33.55 197.17 33.62 ;
    RECT 196.96 33.91 197.17 33.98 ;
    RECT 196.5 33.19 196.71 33.26 ;
    RECT 196.5 33.55 196.71 33.62 ;
    RECT 196.5 33.91 196.71 33.98 ;
    RECT 193.64 33.19 193.85 33.26 ;
    RECT 193.64 33.55 193.85 33.62 ;
    RECT 193.64 33.91 193.85 33.98 ;
    RECT 193.18 33.19 193.39 33.26 ;
    RECT 193.18 33.55 193.39 33.62 ;
    RECT 193.18 33.91 193.39 33.98 ;
    RECT 190.32 33.19 190.53 33.26 ;
    RECT 190.32 33.55 190.53 33.62 ;
    RECT 190.32 33.91 190.53 33.98 ;
    RECT 189.86 33.19 190.07 33.26 ;
    RECT 189.86 33.55 190.07 33.62 ;
    RECT 189.86 33.91 190.07 33.98 ;
    RECT 187.0 33.19 187.21 33.26 ;
    RECT 187.0 33.55 187.21 33.62 ;
    RECT 187.0 33.91 187.21 33.98 ;
    RECT 186.54 33.19 186.75 33.26 ;
    RECT 186.54 33.55 186.75 33.62 ;
    RECT 186.54 33.91 186.75 33.98 ;
    RECT 183.68 33.19 183.89 33.26 ;
    RECT 183.68 33.55 183.89 33.62 ;
    RECT 183.68 33.91 183.89 33.98 ;
    RECT 183.22 33.19 183.43 33.26 ;
    RECT 183.22 33.55 183.43 33.62 ;
    RECT 183.22 33.91 183.43 33.98 ;
    RECT 147.485 33.55 147.555 33.62 ;
    RECT 266.68 33.19 266.89 33.26 ;
    RECT 266.68 33.55 266.89 33.62 ;
    RECT 266.68 33.91 266.89 33.98 ;
    RECT 266.22 33.19 266.43 33.26 ;
    RECT 266.22 33.55 266.43 33.62 ;
    RECT 266.22 33.91 266.43 33.98 ;
    RECT 263.36 33.19 263.57 33.26 ;
    RECT 263.36 33.55 263.57 33.62 ;
    RECT 263.36 33.91 263.57 33.98 ;
    RECT 262.9 33.19 263.11 33.26 ;
    RECT 262.9 33.55 263.11 33.62 ;
    RECT 262.9 33.91 263.11 33.98 ;
    RECT 260.04 33.19 260.25 33.26 ;
    RECT 260.04 33.55 260.25 33.62 ;
    RECT 260.04 33.91 260.25 33.98 ;
    RECT 259.58 33.19 259.79 33.26 ;
    RECT 259.58 33.55 259.79 33.62 ;
    RECT 259.58 33.91 259.79 33.98 ;
    RECT 256.72 33.19 256.93 33.26 ;
    RECT 256.72 33.55 256.93 33.62 ;
    RECT 256.72 33.91 256.93 33.98 ;
    RECT 256.26 33.19 256.47 33.26 ;
    RECT 256.26 33.55 256.47 33.62 ;
    RECT 256.26 33.91 256.47 33.98 ;
    RECT 253.4 33.19 253.61 33.26 ;
    RECT 253.4 33.55 253.61 33.62 ;
    RECT 253.4 33.91 253.61 33.98 ;
    RECT 252.94 33.19 253.15 33.26 ;
    RECT 252.94 33.55 253.15 33.62 ;
    RECT 252.94 33.91 253.15 33.98 ;
    RECT 250.08 16.63 250.29 16.7 ;
    RECT 250.08 16.99 250.29 17.06 ;
    RECT 250.08 17.35 250.29 17.42 ;
    RECT 249.62 16.63 249.83 16.7 ;
    RECT 249.62 16.99 249.83 17.06 ;
    RECT 249.62 17.35 249.83 17.42 ;
    RECT 246.76 16.63 246.97 16.7 ;
    RECT 246.76 16.99 246.97 17.06 ;
    RECT 246.76 17.35 246.97 17.42 ;
    RECT 246.3 16.63 246.51 16.7 ;
    RECT 246.3 16.99 246.51 17.06 ;
    RECT 246.3 17.35 246.51 17.42 ;
    RECT 243.44 16.63 243.65 16.7 ;
    RECT 243.44 16.99 243.65 17.06 ;
    RECT 243.44 17.35 243.65 17.42 ;
    RECT 242.98 16.63 243.19 16.7 ;
    RECT 242.98 16.99 243.19 17.06 ;
    RECT 242.98 17.35 243.19 17.42 ;
    RECT 240.12 16.63 240.33 16.7 ;
    RECT 240.12 16.99 240.33 17.06 ;
    RECT 240.12 17.35 240.33 17.42 ;
    RECT 239.66 16.63 239.87 16.7 ;
    RECT 239.66 16.99 239.87 17.06 ;
    RECT 239.66 17.35 239.87 17.42 ;
    RECT 236.8 16.63 237.01 16.7 ;
    RECT 236.8 16.99 237.01 17.06 ;
    RECT 236.8 17.35 237.01 17.42 ;
    RECT 236.34 16.63 236.55 16.7 ;
    RECT 236.34 16.99 236.55 17.06 ;
    RECT 236.34 17.35 236.55 17.42 ;
    RECT 233.48 16.63 233.69 16.7 ;
    RECT 233.48 16.99 233.69 17.06 ;
    RECT 233.48 17.35 233.69 17.42 ;
    RECT 233.02 16.63 233.23 16.7 ;
    RECT 233.02 16.99 233.23 17.06 ;
    RECT 233.02 17.35 233.23 17.42 ;
    RECT 230.16 16.63 230.37 16.7 ;
    RECT 230.16 16.99 230.37 17.06 ;
    RECT 230.16 17.35 230.37 17.42 ;
    RECT 229.7 16.63 229.91 16.7 ;
    RECT 229.7 16.99 229.91 17.06 ;
    RECT 229.7 17.35 229.91 17.42 ;
    RECT 226.84 16.63 227.05 16.7 ;
    RECT 226.84 16.99 227.05 17.06 ;
    RECT 226.84 17.35 227.05 17.42 ;
    RECT 226.38 16.63 226.59 16.7 ;
    RECT 226.38 16.99 226.59 17.06 ;
    RECT 226.38 17.35 226.59 17.42 ;
    RECT 223.52 16.63 223.73 16.7 ;
    RECT 223.52 16.99 223.73 17.06 ;
    RECT 223.52 17.35 223.73 17.42 ;
    RECT 223.06 16.63 223.27 16.7 ;
    RECT 223.06 16.99 223.27 17.06 ;
    RECT 223.06 17.35 223.27 17.42 ;
    RECT 220.2 16.63 220.41 16.7 ;
    RECT 220.2 16.99 220.41 17.06 ;
    RECT 220.2 17.35 220.41 17.42 ;
    RECT 219.74 16.63 219.95 16.7 ;
    RECT 219.74 16.99 219.95 17.06 ;
    RECT 219.74 17.35 219.95 17.42 ;
    RECT 216.88 16.63 217.09 16.7 ;
    RECT 216.88 16.99 217.09 17.06 ;
    RECT 216.88 17.35 217.09 17.42 ;
    RECT 216.42 16.63 216.63 16.7 ;
    RECT 216.42 16.99 216.63 17.06 ;
    RECT 216.42 17.35 216.63 17.42 ;
    RECT 267.91 16.99 267.98 17.06 ;
    RECT 180.36 16.63 180.57 16.7 ;
    RECT 180.36 16.99 180.57 17.06 ;
    RECT 180.36 17.35 180.57 17.42 ;
    RECT 179.9 16.63 180.11 16.7 ;
    RECT 179.9 16.99 180.11 17.06 ;
    RECT 179.9 17.35 180.11 17.42 ;
    RECT 177.04 16.63 177.25 16.7 ;
    RECT 177.04 16.99 177.25 17.06 ;
    RECT 177.04 17.35 177.25 17.42 ;
    RECT 176.58 16.63 176.79 16.7 ;
    RECT 176.58 16.99 176.79 17.06 ;
    RECT 176.58 17.35 176.79 17.42 ;
    RECT 173.72 16.63 173.93 16.7 ;
    RECT 173.72 16.99 173.93 17.06 ;
    RECT 173.72 17.35 173.93 17.42 ;
    RECT 173.26 16.63 173.47 16.7 ;
    RECT 173.26 16.99 173.47 17.06 ;
    RECT 173.26 17.35 173.47 17.42 ;
    RECT 170.4 16.63 170.61 16.7 ;
    RECT 170.4 16.99 170.61 17.06 ;
    RECT 170.4 17.35 170.61 17.42 ;
    RECT 169.94 16.63 170.15 16.7 ;
    RECT 169.94 16.99 170.15 17.06 ;
    RECT 169.94 17.35 170.15 17.42 ;
    RECT 167.08 16.63 167.29 16.7 ;
    RECT 167.08 16.99 167.29 17.06 ;
    RECT 167.08 17.35 167.29 17.42 ;
    RECT 166.62 16.63 166.83 16.7 ;
    RECT 166.62 16.99 166.83 17.06 ;
    RECT 166.62 17.35 166.83 17.42 ;
    RECT 163.76 16.63 163.97 16.7 ;
    RECT 163.76 16.99 163.97 17.06 ;
    RECT 163.76 17.35 163.97 17.42 ;
    RECT 163.3 16.63 163.51 16.7 ;
    RECT 163.3 16.99 163.51 17.06 ;
    RECT 163.3 17.35 163.51 17.42 ;
    RECT 160.44 16.63 160.65 16.7 ;
    RECT 160.44 16.99 160.65 17.06 ;
    RECT 160.44 17.35 160.65 17.42 ;
    RECT 159.98 16.63 160.19 16.7 ;
    RECT 159.98 16.99 160.19 17.06 ;
    RECT 159.98 17.35 160.19 17.42 ;
    RECT 157.12 16.63 157.33 16.7 ;
    RECT 157.12 16.99 157.33 17.06 ;
    RECT 157.12 17.35 157.33 17.42 ;
    RECT 156.66 16.63 156.87 16.7 ;
    RECT 156.66 16.99 156.87 17.06 ;
    RECT 156.66 17.35 156.87 17.42 ;
    RECT 153.8 16.63 154.01 16.7 ;
    RECT 153.8 16.99 154.01 17.06 ;
    RECT 153.8 17.35 154.01 17.42 ;
    RECT 153.34 16.63 153.55 16.7 ;
    RECT 153.34 16.99 153.55 17.06 ;
    RECT 153.34 17.35 153.55 17.42 ;
    RECT 150.48 16.63 150.69 16.7 ;
    RECT 150.48 16.99 150.69 17.06 ;
    RECT 150.48 17.35 150.69 17.42 ;
    RECT 150.02 16.63 150.23 16.7 ;
    RECT 150.02 16.99 150.23 17.06 ;
    RECT 150.02 17.35 150.23 17.42 ;
    RECT 213.56 16.63 213.77 16.7 ;
    RECT 213.56 16.99 213.77 17.06 ;
    RECT 213.56 17.35 213.77 17.42 ;
    RECT 213.1 16.63 213.31 16.7 ;
    RECT 213.1 16.99 213.31 17.06 ;
    RECT 213.1 17.35 213.31 17.42 ;
    RECT 210.24 16.63 210.45 16.7 ;
    RECT 210.24 16.99 210.45 17.06 ;
    RECT 210.24 17.35 210.45 17.42 ;
    RECT 209.78 16.63 209.99 16.7 ;
    RECT 209.78 16.99 209.99 17.06 ;
    RECT 209.78 17.35 209.99 17.42 ;
    RECT 206.92 16.63 207.13 16.7 ;
    RECT 206.92 16.99 207.13 17.06 ;
    RECT 206.92 17.35 207.13 17.42 ;
    RECT 206.46 16.63 206.67 16.7 ;
    RECT 206.46 16.99 206.67 17.06 ;
    RECT 206.46 17.35 206.67 17.42 ;
    RECT 203.6 16.63 203.81 16.7 ;
    RECT 203.6 16.99 203.81 17.06 ;
    RECT 203.6 17.35 203.81 17.42 ;
    RECT 203.14 16.63 203.35 16.7 ;
    RECT 203.14 16.99 203.35 17.06 ;
    RECT 203.14 17.35 203.35 17.42 ;
    RECT 200.28 16.63 200.49 16.7 ;
    RECT 200.28 16.99 200.49 17.06 ;
    RECT 200.28 17.35 200.49 17.42 ;
    RECT 199.82 16.63 200.03 16.7 ;
    RECT 199.82 16.99 200.03 17.06 ;
    RECT 199.82 17.35 200.03 17.42 ;
    RECT 196.96 16.63 197.17 16.7 ;
    RECT 196.96 16.99 197.17 17.06 ;
    RECT 196.96 17.35 197.17 17.42 ;
    RECT 196.5 16.63 196.71 16.7 ;
    RECT 196.5 16.99 196.71 17.06 ;
    RECT 196.5 17.35 196.71 17.42 ;
    RECT 193.64 16.63 193.85 16.7 ;
    RECT 193.64 16.99 193.85 17.06 ;
    RECT 193.64 17.35 193.85 17.42 ;
    RECT 193.18 16.63 193.39 16.7 ;
    RECT 193.18 16.99 193.39 17.06 ;
    RECT 193.18 17.35 193.39 17.42 ;
    RECT 190.32 16.63 190.53 16.7 ;
    RECT 190.32 16.99 190.53 17.06 ;
    RECT 190.32 17.35 190.53 17.42 ;
    RECT 189.86 16.63 190.07 16.7 ;
    RECT 189.86 16.99 190.07 17.06 ;
    RECT 189.86 17.35 190.07 17.42 ;
    RECT 187.0 16.63 187.21 16.7 ;
    RECT 187.0 16.99 187.21 17.06 ;
    RECT 187.0 17.35 187.21 17.42 ;
    RECT 186.54 16.63 186.75 16.7 ;
    RECT 186.54 16.99 186.75 17.06 ;
    RECT 186.54 17.35 186.75 17.42 ;
    RECT 183.68 16.63 183.89 16.7 ;
    RECT 183.68 16.99 183.89 17.06 ;
    RECT 183.68 17.35 183.89 17.42 ;
    RECT 183.22 16.63 183.43 16.7 ;
    RECT 183.22 16.99 183.43 17.06 ;
    RECT 183.22 17.35 183.43 17.42 ;
    RECT 147.485 16.99 147.555 17.06 ;
    RECT 266.68 16.63 266.89 16.7 ;
    RECT 266.68 16.99 266.89 17.06 ;
    RECT 266.68 17.35 266.89 17.42 ;
    RECT 266.22 16.63 266.43 16.7 ;
    RECT 266.22 16.99 266.43 17.06 ;
    RECT 266.22 17.35 266.43 17.42 ;
    RECT 263.36 16.63 263.57 16.7 ;
    RECT 263.36 16.99 263.57 17.06 ;
    RECT 263.36 17.35 263.57 17.42 ;
    RECT 262.9 16.63 263.11 16.7 ;
    RECT 262.9 16.99 263.11 17.06 ;
    RECT 262.9 17.35 263.11 17.42 ;
    RECT 260.04 16.63 260.25 16.7 ;
    RECT 260.04 16.99 260.25 17.06 ;
    RECT 260.04 17.35 260.25 17.42 ;
    RECT 259.58 16.63 259.79 16.7 ;
    RECT 259.58 16.99 259.79 17.06 ;
    RECT 259.58 17.35 259.79 17.42 ;
    RECT 256.72 16.63 256.93 16.7 ;
    RECT 256.72 16.99 256.93 17.06 ;
    RECT 256.72 17.35 256.93 17.42 ;
    RECT 256.26 16.63 256.47 16.7 ;
    RECT 256.26 16.99 256.47 17.06 ;
    RECT 256.26 17.35 256.47 17.42 ;
    RECT 253.4 16.63 253.61 16.7 ;
    RECT 253.4 16.99 253.61 17.06 ;
    RECT 253.4 17.35 253.61 17.42 ;
    RECT 252.94 16.63 253.15 16.7 ;
    RECT 252.94 16.99 253.15 17.06 ;
    RECT 252.94 17.35 253.15 17.42 ;
    RECT 250.08 32.47 250.29 32.54 ;
    RECT 250.08 32.83 250.29 32.9 ;
    RECT 250.08 33.19 250.29 33.26 ;
    RECT 249.62 32.47 249.83 32.54 ;
    RECT 249.62 32.83 249.83 32.9 ;
    RECT 249.62 33.19 249.83 33.26 ;
    RECT 246.76 32.47 246.97 32.54 ;
    RECT 246.76 32.83 246.97 32.9 ;
    RECT 246.76 33.19 246.97 33.26 ;
    RECT 246.3 32.47 246.51 32.54 ;
    RECT 246.3 32.83 246.51 32.9 ;
    RECT 246.3 33.19 246.51 33.26 ;
    RECT 243.44 32.47 243.65 32.54 ;
    RECT 243.44 32.83 243.65 32.9 ;
    RECT 243.44 33.19 243.65 33.26 ;
    RECT 242.98 32.47 243.19 32.54 ;
    RECT 242.98 32.83 243.19 32.9 ;
    RECT 242.98 33.19 243.19 33.26 ;
    RECT 240.12 32.47 240.33 32.54 ;
    RECT 240.12 32.83 240.33 32.9 ;
    RECT 240.12 33.19 240.33 33.26 ;
    RECT 239.66 32.47 239.87 32.54 ;
    RECT 239.66 32.83 239.87 32.9 ;
    RECT 239.66 33.19 239.87 33.26 ;
    RECT 236.8 32.47 237.01 32.54 ;
    RECT 236.8 32.83 237.01 32.9 ;
    RECT 236.8 33.19 237.01 33.26 ;
    RECT 236.34 32.47 236.55 32.54 ;
    RECT 236.34 32.83 236.55 32.9 ;
    RECT 236.34 33.19 236.55 33.26 ;
    RECT 233.48 32.47 233.69 32.54 ;
    RECT 233.48 32.83 233.69 32.9 ;
    RECT 233.48 33.19 233.69 33.26 ;
    RECT 233.02 32.47 233.23 32.54 ;
    RECT 233.02 32.83 233.23 32.9 ;
    RECT 233.02 33.19 233.23 33.26 ;
    RECT 230.16 32.47 230.37 32.54 ;
    RECT 230.16 32.83 230.37 32.9 ;
    RECT 230.16 33.19 230.37 33.26 ;
    RECT 229.7 32.47 229.91 32.54 ;
    RECT 229.7 32.83 229.91 32.9 ;
    RECT 229.7 33.19 229.91 33.26 ;
    RECT 226.84 32.47 227.05 32.54 ;
    RECT 226.84 32.83 227.05 32.9 ;
    RECT 226.84 33.19 227.05 33.26 ;
    RECT 226.38 32.47 226.59 32.54 ;
    RECT 226.38 32.83 226.59 32.9 ;
    RECT 226.38 33.19 226.59 33.26 ;
    RECT 223.52 32.47 223.73 32.54 ;
    RECT 223.52 32.83 223.73 32.9 ;
    RECT 223.52 33.19 223.73 33.26 ;
    RECT 223.06 32.47 223.27 32.54 ;
    RECT 223.06 32.83 223.27 32.9 ;
    RECT 223.06 33.19 223.27 33.26 ;
    RECT 220.2 32.47 220.41 32.54 ;
    RECT 220.2 32.83 220.41 32.9 ;
    RECT 220.2 33.19 220.41 33.26 ;
    RECT 219.74 32.47 219.95 32.54 ;
    RECT 219.74 32.83 219.95 32.9 ;
    RECT 219.74 33.19 219.95 33.26 ;
    RECT 216.88 32.47 217.09 32.54 ;
    RECT 216.88 32.83 217.09 32.9 ;
    RECT 216.88 33.19 217.09 33.26 ;
    RECT 216.42 32.47 216.63 32.54 ;
    RECT 216.42 32.83 216.63 32.9 ;
    RECT 216.42 33.19 216.63 33.26 ;
    RECT 267.91 32.83 267.98 32.9 ;
    RECT 180.36 32.47 180.57 32.54 ;
    RECT 180.36 32.83 180.57 32.9 ;
    RECT 180.36 33.19 180.57 33.26 ;
    RECT 179.9 32.47 180.11 32.54 ;
    RECT 179.9 32.83 180.11 32.9 ;
    RECT 179.9 33.19 180.11 33.26 ;
    RECT 177.04 32.47 177.25 32.54 ;
    RECT 177.04 32.83 177.25 32.9 ;
    RECT 177.04 33.19 177.25 33.26 ;
    RECT 176.58 32.47 176.79 32.54 ;
    RECT 176.58 32.83 176.79 32.9 ;
    RECT 176.58 33.19 176.79 33.26 ;
    RECT 173.72 32.47 173.93 32.54 ;
    RECT 173.72 32.83 173.93 32.9 ;
    RECT 173.72 33.19 173.93 33.26 ;
    RECT 173.26 32.47 173.47 32.54 ;
    RECT 173.26 32.83 173.47 32.9 ;
    RECT 173.26 33.19 173.47 33.26 ;
    RECT 170.4 32.47 170.61 32.54 ;
    RECT 170.4 32.83 170.61 32.9 ;
    RECT 170.4 33.19 170.61 33.26 ;
    RECT 169.94 32.47 170.15 32.54 ;
    RECT 169.94 32.83 170.15 32.9 ;
    RECT 169.94 33.19 170.15 33.26 ;
    RECT 167.08 32.47 167.29 32.54 ;
    RECT 167.08 32.83 167.29 32.9 ;
    RECT 167.08 33.19 167.29 33.26 ;
    RECT 166.62 32.47 166.83 32.54 ;
    RECT 166.62 32.83 166.83 32.9 ;
    RECT 166.62 33.19 166.83 33.26 ;
    RECT 163.76 32.47 163.97 32.54 ;
    RECT 163.76 32.83 163.97 32.9 ;
    RECT 163.76 33.19 163.97 33.26 ;
    RECT 163.3 32.47 163.51 32.54 ;
    RECT 163.3 32.83 163.51 32.9 ;
    RECT 163.3 33.19 163.51 33.26 ;
    RECT 160.44 32.47 160.65 32.54 ;
    RECT 160.44 32.83 160.65 32.9 ;
    RECT 160.44 33.19 160.65 33.26 ;
    RECT 159.98 32.47 160.19 32.54 ;
    RECT 159.98 32.83 160.19 32.9 ;
    RECT 159.98 33.19 160.19 33.26 ;
    RECT 157.12 32.47 157.33 32.54 ;
    RECT 157.12 32.83 157.33 32.9 ;
    RECT 157.12 33.19 157.33 33.26 ;
    RECT 156.66 32.47 156.87 32.54 ;
    RECT 156.66 32.83 156.87 32.9 ;
    RECT 156.66 33.19 156.87 33.26 ;
    RECT 153.8 32.47 154.01 32.54 ;
    RECT 153.8 32.83 154.01 32.9 ;
    RECT 153.8 33.19 154.01 33.26 ;
    RECT 153.34 32.47 153.55 32.54 ;
    RECT 153.34 32.83 153.55 32.9 ;
    RECT 153.34 33.19 153.55 33.26 ;
    RECT 150.48 32.47 150.69 32.54 ;
    RECT 150.48 32.83 150.69 32.9 ;
    RECT 150.48 33.19 150.69 33.26 ;
    RECT 150.02 32.47 150.23 32.54 ;
    RECT 150.02 32.83 150.23 32.9 ;
    RECT 150.02 33.19 150.23 33.26 ;
    RECT 213.56 32.47 213.77 32.54 ;
    RECT 213.56 32.83 213.77 32.9 ;
    RECT 213.56 33.19 213.77 33.26 ;
    RECT 213.1 32.47 213.31 32.54 ;
    RECT 213.1 32.83 213.31 32.9 ;
    RECT 213.1 33.19 213.31 33.26 ;
    RECT 210.24 32.47 210.45 32.54 ;
    RECT 210.24 32.83 210.45 32.9 ;
    RECT 210.24 33.19 210.45 33.26 ;
    RECT 209.78 32.47 209.99 32.54 ;
    RECT 209.78 32.83 209.99 32.9 ;
    RECT 209.78 33.19 209.99 33.26 ;
    RECT 206.92 32.47 207.13 32.54 ;
    RECT 206.92 32.83 207.13 32.9 ;
    RECT 206.92 33.19 207.13 33.26 ;
    RECT 206.46 32.47 206.67 32.54 ;
    RECT 206.46 32.83 206.67 32.9 ;
    RECT 206.46 33.19 206.67 33.26 ;
    RECT 203.6 32.47 203.81 32.54 ;
    RECT 203.6 32.83 203.81 32.9 ;
    RECT 203.6 33.19 203.81 33.26 ;
    RECT 203.14 32.47 203.35 32.54 ;
    RECT 203.14 32.83 203.35 32.9 ;
    RECT 203.14 33.19 203.35 33.26 ;
    RECT 200.28 32.47 200.49 32.54 ;
    RECT 200.28 32.83 200.49 32.9 ;
    RECT 200.28 33.19 200.49 33.26 ;
    RECT 199.82 32.47 200.03 32.54 ;
    RECT 199.82 32.83 200.03 32.9 ;
    RECT 199.82 33.19 200.03 33.26 ;
    RECT 196.96 32.47 197.17 32.54 ;
    RECT 196.96 32.83 197.17 32.9 ;
    RECT 196.96 33.19 197.17 33.26 ;
    RECT 196.5 32.47 196.71 32.54 ;
    RECT 196.5 32.83 196.71 32.9 ;
    RECT 196.5 33.19 196.71 33.26 ;
    RECT 193.64 32.47 193.85 32.54 ;
    RECT 193.64 32.83 193.85 32.9 ;
    RECT 193.64 33.19 193.85 33.26 ;
    RECT 193.18 32.47 193.39 32.54 ;
    RECT 193.18 32.83 193.39 32.9 ;
    RECT 193.18 33.19 193.39 33.26 ;
    RECT 190.32 32.47 190.53 32.54 ;
    RECT 190.32 32.83 190.53 32.9 ;
    RECT 190.32 33.19 190.53 33.26 ;
    RECT 189.86 32.47 190.07 32.54 ;
    RECT 189.86 32.83 190.07 32.9 ;
    RECT 189.86 33.19 190.07 33.26 ;
    RECT 187.0 32.47 187.21 32.54 ;
    RECT 187.0 32.83 187.21 32.9 ;
    RECT 187.0 33.19 187.21 33.26 ;
    RECT 186.54 32.47 186.75 32.54 ;
    RECT 186.54 32.83 186.75 32.9 ;
    RECT 186.54 33.19 186.75 33.26 ;
    RECT 183.68 32.47 183.89 32.54 ;
    RECT 183.68 32.83 183.89 32.9 ;
    RECT 183.68 33.19 183.89 33.26 ;
    RECT 183.22 32.47 183.43 32.54 ;
    RECT 183.22 32.83 183.43 32.9 ;
    RECT 183.22 33.19 183.43 33.26 ;
    RECT 147.485 32.83 147.555 32.9 ;
    RECT 266.68 32.47 266.89 32.54 ;
    RECT 266.68 32.83 266.89 32.9 ;
    RECT 266.68 33.19 266.89 33.26 ;
    RECT 266.22 32.47 266.43 32.54 ;
    RECT 266.22 32.83 266.43 32.9 ;
    RECT 266.22 33.19 266.43 33.26 ;
    RECT 263.36 32.47 263.57 32.54 ;
    RECT 263.36 32.83 263.57 32.9 ;
    RECT 263.36 33.19 263.57 33.26 ;
    RECT 262.9 32.47 263.11 32.54 ;
    RECT 262.9 32.83 263.11 32.9 ;
    RECT 262.9 33.19 263.11 33.26 ;
    RECT 260.04 32.47 260.25 32.54 ;
    RECT 260.04 32.83 260.25 32.9 ;
    RECT 260.04 33.19 260.25 33.26 ;
    RECT 259.58 32.47 259.79 32.54 ;
    RECT 259.58 32.83 259.79 32.9 ;
    RECT 259.58 33.19 259.79 33.26 ;
    RECT 256.72 32.47 256.93 32.54 ;
    RECT 256.72 32.83 256.93 32.9 ;
    RECT 256.72 33.19 256.93 33.26 ;
    RECT 256.26 32.47 256.47 32.54 ;
    RECT 256.26 32.83 256.47 32.9 ;
    RECT 256.26 33.19 256.47 33.26 ;
    RECT 253.4 32.47 253.61 32.54 ;
    RECT 253.4 32.83 253.61 32.9 ;
    RECT 253.4 33.19 253.61 33.26 ;
    RECT 252.94 32.47 253.15 32.54 ;
    RECT 252.94 32.83 253.15 32.9 ;
    RECT 252.94 33.19 253.15 33.26 ;
    RECT 250.08 72.09 250.29 72.16 ;
    RECT 250.08 72.45 250.29 72.52 ;
    RECT 250.08 72.81 250.29 72.88 ;
    RECT 249.62 72.09 249.83 72.16 ;
    RECT 249.62 72.45 249.83 72.52 ;
    RECT 249.62 72.81 249.83 72.88 ;
    RECT 246.76 72.09 246.97 72.16 ;
    RECT 246.76 72.45 246.97 72.52 ;
    RECT 246.76 72.81 246.97 72.88 ;
    RECT 246.3 72.09 246.51 72.16 ;
    RECT 246.3 72.45 246.51 72.52 ;
    RECT 246.3 72.81 246.51 72.88 ;
    RECT 243.44 72.09 243.65 72.16 ;
    RECT 243.44 72.45 243.65 72.52 ;
    RECT 243.44 72.81 243.65 72.88 ;
    RECT 242.98 72.09 243.19 72.16 ;
    RECT 242.98 72.45 243.19 72.52 ;
    RECT 242.98 72.81 243.19 72.88 ;
    RECT 240.12 72.09 240.33 72.16 ;
    RECT 240.12 72.45 240.33 72.52 ;
    RECT 240.12 72.81 240.33 72.88 ;
    RECT 239.66 72.09 239.87 72.16 ;
    RECT 239.66 72.45 239.87 72.52 ;
    RECT 239.66 72.81 239.87 72.88 ;
    RECT 236.8 72.09 237.01 72.16 ;
    RECT 236.8 72.45 237.01 72.52 ;
    RECT 236.8 72.81 237.01 72.88 ;
    RECT 236.34 72.09 236.55 72.16 ;
    RECT 236.34 72.45 236.55 72.52 ;
    RECT 236.34 72.81 236.55 72.88 ;
    RECT 233.48 72.09 233.69 72.16 ;
    RECT 233.48 72.45 233.69 72.52 ;
    RECT 233.48 72.81 233.69 72.88 ;
    RECT 233.02 72.09 233.23 72.16 ;
    RECT 233.02 72.45 233.23 72.52 ;
    RECT 233.02 72.81 233.23 72.88 ;
    RECT 230.16 72.09 230.37 72.16 ;
    RECT 230.16 72.45 230.37 72.52 ;
    RECT 230.16 72.81 230.37 72.88 ;
    RECT 229.7 72.09 229.91 72.16 ;
    RECT 229.7 72.45 229.91 72.52 ;
    RECT 229.7 72.81 229.91 72.88 ;
    RECT 226.84 72.09 227.05 72.16 ;
    RECT 226.84 72.45 227.05 72.52 ;
    RECT 226.84 72.81 227.05 72.88 ;
    RECT 226.38 72.09 226.59 72.16 ;
    RECT 226.38 72.45 226.59 72.52 ;
    RECT 226.38 72.81 226.59 72.88 ;
    RECT 223.52 72.09 223.73 72.16 ;
    RECT 223.52 72.45 223.73 72.52 ;
    RECT 223.52 72.81 223.73 72.88 ;
    RECT 223.06 72.09 223.27 72.16 ;
    RECT 223.06 72.45 223.27 72.52 ;
    RECT 223.06 72.81 223.27 72.88 ;
    RECT 220.2 72.09 220.41 72.16 ;
    RECT 220.2 72.45 220.41 72.52 ;
    RECT 220.2 72.81 220.41 72.88 ;
    RECT 219.74 72.09 219.95 72.16 ;
    RECT 219.74 72.45 219.95 72.52 ;
    RECT 219.74 72.81 219.95 72.88 ;
    RECT 216.88 72.09 217.09 72.16 ;
    RECT 216.88 72.45 217.09 72.52 ;
    RECT 216.88 72.81 217.09 72.88 ;
    RECT 216.42 72.09 216.63 72.16 ;
    RECT 216.42 72.45 216.63 72.52 ;
    RECT 216.42 72.81 216.63 72.88 ;
    RECT 267.91 72.45 267.98 72.52 ;
    RECT 180.36 72.09 180.57 72.16 ;
    RECT 180.36 72.45 180.57 72.52 ;
    RECT 180.36 72.81 180.57 72.88 ;
    RECT 179.9 72.09 180.11 72.16 ;
    RECT 179.9 72.45 180.11 72.52 ;
    RECT 179.9 72.81 180.11 72.88 ;
    RECT 177.04 72.09 177.25 72.16 ;
    RECT 177.04 72.45 177.25 72.52 ;
    RECT 177.04 72.81 177.25 72.88 ;
    RECT 176.58 72.09 176.79 72.16 ;
    RECT 176.58 72.45 176.79 72.52 ;
    RECT 176.58 72.81 176.79 72.88 ;
    RECT 173.72 72.09 173.93 72.16 ;
    RECT 173.72 72.45 173.93 72.52 ;
    RECT 173.72 72.81 173.93 72.88 ;
    RECT 173.26 72.09 173.47 72.16 ;
    RECT 173.26 72.45 173.47 72.52 ;
    RECT 173.26 72.81 173.47 72.88 ;
    RECT 170.4 72.09 170.61 72.16 ;
    RECT 170.4 72.45 170.61 72.52 ;
    RECT 170.4 72.81 170.61 72.88 ;
    RECT 169.94 72.09 170.15 72.16 ;
    RECT 169.94 72.45 170.15 72.52 ;
    RECT 169.94 72.81 170.15 72.88 ;
    RECT 167.08 72.09 167.29 72.16 ;
    RECT 167.08 72.45 167.29 72.52 ;
    RECT 167.08 72.81 167.29 72.88 ;
    RECT 166.62 72.09 166.83 72.16 ;
    RECT 166.62 72.45 166.83 72.52 ;
    RECT 166.62 72.81 166.83 72.88 ;
    RECT 163.76 72.09 163.97 72.16 ;
    RECT 163.76 72.45 163.97 72.52 ;
    RECT 163.76 72.81 163.97 72.88 ;
    RECT 163.3 72.09 163.51 72.16 ;
    RECT 163.3 72.45 163.51 72.52 ;
    RECT 163.3 72.81 163.51 72.88 ;
    RECT 160.44 72.09 160.65 72.16 ;
    RECT 160.44 72.45 160.65 72.52 ;
    RECT 160.44 72.81 160.65 72.88 ;
    RECT 159.98 72.09 160.19 72.16 ;
    RECT 159.98 72.45 160.19 72.52 ;
    RECT 159.98 72.81 160.19 72.88 ;
    RECT 157.12 72.09 157.33 72.16 ;
    RECT 157.12 72.45 157.33 72.52 ;
    RECT 157.12 72.81 157.33 72.88 ;
    RECT 156.66 72.09 156.87 72.16 ;
    RECT 156.66 72.45 156.87 72.52 ;
    RECT 156.66 72.81 156.87 72.88 ;
    RECT 153.8 72.09 154.01 72.16 ;
    RECT 153.8 72.45 154.01 72.52 ;
    RECT 153.8 72.81 154.01 72.88 ;
    RECT 153.34 72.09 153.55 72.16 ;
    RECT 153.34 72.45 153.55 72.52 ;
    RECT 153.34 72.81 153.55 72.88 ;
    RECT 150.48 72.09 150.69 72.16 ;
    RECT 150.48 72.45 150.69 72.52 ;
    RECT 150.48 72.81 150.69 72.88 ;
    RECT 150.02 72.09 150.23 72.16 ;
    RECT 150.02 72.45 150.23 72.52 ;
    RECT 150.02 72.81 150.23 72.88 ;
    RECT 213.56 72.09 213.77 72.16 ;
    RECT 213.56 72.45 213.77 72.52 ;
    RECT 213.56 72.81 213.77 72.88 ;
    RECT 213.1 72.09 213.31 72.16 ;
    RECT 213.1 72.45 213.31 72.52 ;
    RECT 213.1 72.81 213.31 72.88 ;
    RECT 210.24 72.09 210.45 72.16 ;
    RECT 210.24 72.45 210.45 72.52 ;
    RECT 210.24 72.81 210.45 72.88 ;
    RECT 209.78 72.09 209.99 72.16 ;
    RECT 209.78 72.45 209.99 72.52 ;
    RECT 209.78 72.81 209.99 72.88 ;
    RECT 206.92 72.09 207.13 72.16 ;
    RECT 206.92 72.45 207.13 72.52 ;
    RECT 206.92 72.81 207.13 72.88 ;
    RECT 206.46 72.09 206.67 72.16 ;
    RECT 206.46 72.45 206.67 72.52 ;
    RECT 206.46 72.81 206.67 72.88 ;
    RECT 203.6 72.09 203.81 72.16 ;
    RECT 203.6 72.45 203.81 72.52 ;
    RECT 203.6 72.81 203.81 72.88 ;
    RECT 203.14 72.09 203.35 72.16 ;
    RECT 203.14 72.45 203.35 72.52 ;
    RECT 203.14 72.81 203.35 72.88 ;
    RECT 200.28 72.09 200.49 72.16 ;
    RECT 200.28 72.45 200.49 72.52 ;
    RECT 200.28 72.81 200.49 72.88 ;
    RECT 199.82 72.09 200.03 72.16 ;
    RECT 199.82 72.45 200.03 72.52 ;
    RECT 199.82 72.81 200.03 72.88 ;
    RECT 196.96 72.09 197.17 72.16 ;
    RECT 196.96 72.45 197.17 72.52 ;
    RECT 196.96 72.81 197.17 72.88 ;
    RECT 196.5 72.09 196.71 72.16 ;
    RECT 196.5 72.45 196.71 72.52 ;
    RECT 196.5 72.81 196.71 72.88 ;
    RECT 193.64 72.09 193.85 72.16 ;
    RECT 193.64 72.45 193.85 72.52 ;
    RECT 193.64 72.81 193.85 72.88 ;
    RECT 193.18 72.09 193.39 72.16 ;
    RECT 193.18 72.45 193.39 72.52 ;
    RECT 193.18 72.81 193.39 72.88 ;
    RECT 190.32 72.09 190.53 72.16 ;
    RECT 190.32 72.45 190.53 72.52 ;
    RECT 190.32 72.81 190.53 72.88 ;
    RECT 189.86 72.09 190.07 72.16 ;
    RECT 189.86 72.45 190.07 72.52 ;
    RECT 189.86 72.81 190.07 72.88 ;
    RECT 187.0 72.09 187.21 72.16 ;
    RECT 187.0 72.45 187.21 72.52 ;
    RECT 187.0 72.81 187.21 72.88 ;
    RECT 186.54 72.09 186.75 72.16 ;
    RECT 186.54 72.45 186.75 72.52 ;
    RECT 186.54 72.81 186.75 72.88 ;
    RECT 183.68 72.09 183.89 72.16 ;
    RECT 183.68 72.45 183.89 72.52 ;
    RECT 183.68 72.81 183.89 72.88 ;
    RECT 183.22 72.09 183.43 72.16 ;
    RECT 183.22 72.45 183.43 72.52 ;
    RECT 183.22 72.81 183.43 72.88 ;
    RECT 147.485 72.45 147.555 72.52 ;
    RECT 266.68 72.09 266.89 72.16 ;
    RECT 266.68 72.45 266.89 72.52 ;
    RECT 266.68 72.81 266.89 72.88 ;
    RECT 266.22 72.09 266.43 72.16 ;
    RECT 266.22 72.45 266.43 72.52 ;
    RECT 266.22 72.81 266.43 72.88 ;
    RECT 263.36 72.09 263.57 72.16 ;
    RECT 263.36 72.45 263.57 72.52 ;
    RECT 263.36 72.81 263.57 72.88 ;
    RECT 262.9 72.09 263.11 72.16 ;
    RECT 262.9 72.45 263.11 72.52 ;
    RECT 262.9 72.81 263.11 72.88 ;
    RECT 260.04 72.09 260.25 72.16 ;
    RECT 260.04 72.45 260.25 72.52 ;
    RECT 260.04 72.81 260.25 72.88 ;
    RECT 259.58 72.09 259.79 72.16 ;
    RECT 259.58 72.45 259.79 72.52 ;
    RECT 259.58 72.81 259.79 72.88 ;
    RECT 256.72 72.09 256.93 72.16 ;
    RECT 256.72 72.45 256.93 72.52 ;
    RECT 256.72 72.81 256.93 72.88 ;
    RECT 256.26 72.09 256.47 72.16 ;
    RECT 256.26 72.45 256.47 72.52 ;
    RECT 256.26 72.81 256.47 72.88 ;
    RECT 253.4 72.09 253.61 72.16 ;
    RECT 253.4 72.45 253.61 72.52 ;
    RECT 253.4 72.81 253.61 72.88 ;
    RECT 252.94 72.09 253.15 72.16 ;
    RECT 252.94 72.45 253.15 72.52 ;
    RECT 252.94 72.81 253.15 72.88 ;
    RECT 250.08 15.91 250.29 15.98 ;
    RECT 250.08 16.27 250.29 16.34 ;
    RECT 250.08 16.63 250.29 16.7 ;
    RECT 249.62 15.91 249.83 15.98 ;
    RECT 249.62 16.27 249.83 16.34 ;
    RECT 249.62 16.63 249.83 16.7 ;
    RECT 246.76 15.91 246.97 15.98 ;
    RECT 246.76 16.27 246.97 16.34 ;
    RECT 246.76 16.63 246.97 16.7 ;
    RECT 246.3 15.91 246.51 15.98 ;
    RECT 246.3 16.27 246.51 16.34 ;
    RECT 246.3 16.63 246.51 16.7 ;
    RECT 243.44 15.91 243.65 15.98 ;
    RECT 243.44 16.27 243.65 16.34 ;
    RECT 243.44 16.63 243.65 16.7 ;
    RECT 242.98 15.91 243.19 15.98 ;
    RECT 242.98 16.27 243.19 16.34 ;
    RECT 242.98 16.63 243.19 16.7 ;
    RECT 240.12 15.91 240.33 15.98 ;
    RECT 240.12 16.27 240.33 16.34 ;
    RECT 240.12 16.63 240.33 16.7 ;
    RECT 239.66 15.91 239.87 15.98 ;
    RECT 239.66 16.27 239.87 16.34 ;
    RECT 239.66 16.63 239.87 16.7 ;
    RECT 236.8 15.91 237.01 15.98 ;
    RECT 236.8 16.27 237.01 16.34 ;
    RECT 236.8 16.63 237.01 16.7 ;
    RECT 236.34 15.91 236.55 15.98 ;
    RECT 236.34 16.27 236.55 16.34 ;
    RECT 236.34 16.63 236.55 16.7 ;
    RECT 233.48 15.91 233.69 15.98 ;
    RECT 233.48 16.27 233.69 16.34 ;
    RECT 233.48 16.63 233.69 16.7 ;
    RECT 233.02 15.91 233.23 15.98 ;
    RECT 233.02 16.27 233.23 16.34 ;
    RECT 233.02 16.63 233.23 16.7 ;
    RECT 230.16 15.91 230.37 15.98 ;
    RECT 230.16 16.27 230.37 16.34 ;
    RECT 230.16 16.63 230.37 16.7 ;
    RECT 229.7 15.91 229.91 15.98 ;
    RECT 229.7 16.27 229.91 16.34 ;
    RECT 229.7 16.63 229.91 16.7 ;
    RECT 226.84 15.91 227.05 15.98 ;
    RECT 226.84 16.27 227.05 16.34 ;
    RECT 226.84 16.63 227.05 16.7 ;
    RECT 226.38 15.91 226.59 15.98 ;
    RECT 226.38 16.27 226.59 16.34 ;
    RECT 226.38 16.63 226.59 16.7 ;
    RECT 223.52 15.91 223.73 15.98 ;
    RECT 223.52 16.27 223.73 16.34 ;
    RECT 223.52 16.63 223.73 16.7 ;
    RECT 223.06 15.91 223.27 15.98 ;
    RECT 223.06 16.27 223.27 16.34 ;
    RECT 223.06 16.63 223.27 16.7 ;
    RECT 220.2 15.91 220.41 15.98 ;
    RECT 220.2 16.27 220.41 16.34 ;
    RECT 220.2 16.63 220.41 16.7 ;
    RECT 219.74 15.91 219.95 15.98 ;
    RECT 219.74 16.27 219.95 16.34 ;
    RECT 219.74 16.63 219.95 16.7 ;
    RECT 216.88 15.91 217.09 15.98 ;
    RECT 216.88 16.27 217.09 16.34 ;
    RECT 216.88 16.63 217.09 16.7 ;
    RECT 216.42 15.91 216.63 15.98 ;
    RECT 216.42 16.27 216.63 16.34 ;
    RECT 216.42 16.63 216.63 16.7 ;
    RECT 267.91 16.27 267.98 16.34 ;
    RECT 180.36 15.91 180.57 15.98 ;
    RECT 180.36 16.27 180.57 16.34 ;
    RECT 180.36 16.63 180.57 16.7 ;
    RECT 179.9 15.91 180.11 15.98 ;
    RECT 179.9 16.27 180.11 16.34 ;
    RECT 179.9 16.63 180.11 16.7 ;
    RECT 177.04 15.91 177.25 15.98 ;
    RECT 177.04 16.27 177.25 16.34 ;
    RECT 177.04 16.63 177.25 16.7 ;
    RECT 176.58 15.91 176.79 15.98 ;
    RECT 176.58 16.27 176.79 16.34 ;
    RECT 176.58 16.63 176.79 16.7 ;
    RECT 173.72 15.91 173.93 15.98 ;
    RECT 173.72 16.27 173.93 16.34 ;
    RECT 173.72 16.63 173.93 16.7 ;
    RECT 173.26 15.91 173.47 15.98 ;
    RECT 173.26 16.27 173.47 16.34 ;
    RECT 173.26 16.63 173.47 16.7 ;
    RECT 170.4 15.91 170.61 15.98 ;
    RECT 170.4 16.27 170.61 16.34 ;
    RECT 170.4 16.63 170.61 16.7 ;
    RECT 169.94 15.91 170.15 15.98 ;
    RECT 169.94 16.27 170.15 16.34 ;
    RECT 169.94 16.63 170.15 16.7 ;
    RECT 167.08 15.91 167.29 15.98 ;
    RECT 167.08 16.27 167.29 16.34 ;
    RECT 167.08 16.63 167.29 16.7 ;
    RECT 166.62 15.91 166.83 15.98 ;
    RECT 166.62 16.27 166.83 16.34 ;
    RECT 166.62 16.63 166.83 16.7 ;
    RECT 163.76 15.91 163.97 15.98 ;
    RECT 163.76 16.27 163.97 16.34 ;
    RECT 163.76 16.63 163.97 16.7 ;
    RECT 163.3 15.91 163.51 15.98 ;
    RECT 163.3 16.27 163.51 16.34 ;
    RECT 163.3 16.63 163.51 16.7 ;
    RECT 160.44 15.91 160.65 15.98 ;
    RECT 160.44 16.27 160.65 16.34 ;
    RECT 160.44 16.63 160.65 16.7 ;
    RECT 159.98 15.91 160.19 15.98 ;
    RECT 159.98 16.27 160.19 16.34 ;
    RECT 159.98 16.63 160.19 16.7 ;
    RECT 157.12 15.91 157.33 15.98 ;
    RECT 157.12 16.27 157.33 16.34 ;
    RECT 157.12 16.63 157.33 16.7 ;
    RECT 156.66 15.91 156.87 15.98 ;
    RECT 156.66 16.27 156.87 16.34 ;
    RECT 156.66 16.63 156.87 16.7 ;
    RECT 153.8 15.91 154.01 15.98 ;
    RECT 153.8 16.27 154.01 16.34 ;
    RECT 153.8 16.63 154.01 16.7 ;
    RECT 153.34 15.91 153.55 15.98 ;
    RECT 153.34 16.27 153.55 16.34 ;
    RECT 153.34 16.63 153.55 16.7 ;
    RECT 150.48 15.91 150.69 15.98 ;
    RECT 150.48 16.27 150.69 16.34 ;
    RECT 150.48 16.63 150.69 16.7 ;
    RECT 150.02 15.91 150.23 15.98 ;
    RECT 150.02 16.27 150.23 16.34 ;
    RECT 150.02 16.63 150.23 16.7 ;
    RECT 213.56 15.91 213.77 15.98 ;
    RECT 213.56 16.27 213.77 16.34 ;
    RECT 213.56 16.63 213.77 16.7 ;
    RECT 213.1 15.91 213.31 15.98 ;
    RECT 213.1 16.27 213.31 16.34 ;
    RECT 213.1 16.63 213.31 16.7 ;
    RECT 210.24 15.91 210.45 15.98 ;
    RECT 210.24 16.27 210.45 16.34 ;
    RECT 210.24 16.63 210.45 16.7 ;
    RECT 209.78 15.91 209.99 15.98 ;
    RECT 209.78 16.27 209.99 16.34 ;
    RECT 209.78 16.63 209.99 16.7 ;
    RECT 206.92 15.91 207.13 15.98 ;
    RECT 206.92 16.27 207.13 16.34 ;
    RECT 206.92 16.63 207.13 16.7 ;
    RECT 206.46 15.91 206.67 15.98 ;
    RECT 206.46 16.27 206.67 16.34 ;
    RECT 206.46 16.63 206.67 16.7 ;
    RECT 203.6 15.91 203.81 15.98 ;
    RECT 203.6 16.27 203.81 16.34 ;
    RECT 203.6 16.63 203.81 16.7 ;
    RECT 203.14 15.91 203.35 15.98 ;
    RECT 203.14 16.27 203.35 16.34 ;
    RECT 203.14 16.63 203.35 16.7 ;
    RECT 200.28 15.91 200.49 15.98 ;
    RECT 200.28 16.27 200.49 16.34 ;
    RECT 200.28 16.63 200.49 16.7 ;
    RECT 199.82 15.91 200.03 15.98 ;
    RECT 199.82 16.27 200.03 16.34 ;
    RECT 199.82 16.63 200.03 16.7 ;
    RECT 196.96 15.91 197.17 15.98 ;
    RECT 196.96 16.27 197.17 16.34 ;
    RECT 196.96 16.63 197.17 16.7 ;
    RECT 196.5 15.91 196.71 15.98 ;
    RECT 196.5 16.27 196.71 16.34 ;
    RECT 196.5 16.63 196.71 16.7 ;
    RECT 193.64 15.91 193.85 15.98 ;
    RECT 193.64 16.27 193.85 16.34 ;
    RECT 193.64 16.63 193.85 16.7 ;
    RECT 193.18 15.91 193.39 15.98 ;
    RECT 193.18 16.27 193.39 16.34 ;
    RECT 193.18 16.63 193.39 16.7 ;
    RECT 190.32 15.91 190.53 15.98 ;
    RECT 190.32 16.27 190.53 16.34 ;
    RECT 190.32 16.63 190.53 16.7 ;
    RECT 189.86 15.91 190.07 15.98 ;
    RECT 189.86 16.27 190.07 16.34 ;
    RECT 189.86 16.63 190.07 16.7 ;
    RECT 187.0 15.91 187.21 15.98 ;
    RECT 187.0 16.27 187.21 16.34 ;
    RECT 187.0 16.63 187.21 16.7 ;
    RECT 186.54 15.91 186.75 15.98 ;
    RECT 186.54 16.27 186.75 16.34 ;
    RECT 186.54 16.63 186.75 16.7 ;
    RECT 183.68 15.91 183.89 15.98 ;
    RECT 183.68 16.27 183.89 16.34 ;
    RECT 183.68 16.63 183.89 16.7 ;
    RECT 183.22 15.91 183.43 15.98 ;
    RECT 183.22 16.27 183.43 16.34 ;
    RECT 183.22 16.63 183.43 16.7 ;
    RECT 147.485 16.27 147.555 16.34 ;
    RECT 266.68 15.91 266.89 15.98 ;
    RECT 266.68 16.27 266.89 16.34 ;
    RECT 266.68 16.63 266.89 16.7 ;
    RECT 266.22 15.91 266.43 15.98 ;
    RECT 266.22 16.27 266.43 16.34 ;
    RECT 266.22 16.63 266.43 16.7 ;
    RECT 263.36 15.91 263.57 15.98 ;
    RECT 263.36 16.27 263.57 16.34 ;
    RECT 263.36 16.63 263.57 16.7 ;
    RECT 262.9 15.91 263.11 15.98 ;
    RECT 262.9 16.27 263.11 16.34 ;
    RECT 262.9 16.63 263.11 16.7 ;
    RECT 260.04 15.91 260.25 15.98 ;
    RECT 260.04 16.27 260.25 16.34 ;
    RECT 260.04 16.63 260.25 16.7 ;
    RECT 259.58 15.91 259.79 15.98 ;
    RECT 259.58 16.27 259.79 16.34 ;
    RECT 259.58 16.63 259.79 16.7 ;
    RECT 256.72 15.91 256.93 15.98 ;
    RECT 256.72 16.27 256.93 16.34 ;
    RECT 256.72 16.63 256.93 16.7 ;
    RECT 256.26 15.91 256.47 15.98 ;
    RECT 256.26 16.27 256.47 16.34 ;
    RECT 256.26 16.63 256.47 16.7 ;
    RECT 253.4 15.91 253.61 15.98 ;
    RECT 253.4 16.27 253.61 16.34 ;
    RECT 253.4 16.63 253.61 16.7 ;
    RECT 252.94 15.91 253.15 15.98 ;
    RECT 252.94 16.27 253.15 16.34 ;
    RECT 252.94 16.63 253.15 16.7 ;
    RECT 250.08 31.75 250.29 31.82 ;
    RECT 250.08 32.11 250.29 32.18 ;
    RECT 250.08 32.47 250.29 32.54 ;
    RECT 249.62 31.75 249.83 31.82 ;
    RECT 249.62 32.11 249.83 32.18 ;
    RECT 249.62 32.47 249.83 32.54 ;
    RECT 246.76 31.75 246.97 31.82 ;
    RECT 246.76 32.11 246.97 32.18 ;
    RECT 246.76 32.47 246.97 32.54 ;
    RECT 246.3 31.75 246.51 31.82 ;
    RECT 246.3 32.11 246.51 32.18 ;
    RECT 246.3 32.47 246.51 32.54 ;
    RECT 243.44 31.75 243.65 31.82 ;
    RECT 243.44 32.11 243.65 32.18 ;
    RECT 243.44 32.47 243.65 32.54 ;
    RECT 242.98 31.75 243.19 31.82 ;
    RECT 242.98 32.11 243.19 32.18 ;
    RECT 242.98 32.47 243.19 32.54 ;
    RECT 240.12 31.75 240.33 31.82 ;
    RECT 240.12 32.11 240.33 32.18 ;
    RECT 240.12 32.47 240.33 32.54 ;
    RECT 239.66 31.75 239.87 31.82 ;
    RECT 239.66 32.11 239.87 32.18 ;
    RECT 239.66 32.47 239.87 32.54 ;
    RECT 236.8 31.75 237.01 31.82 ;
    RECT 236.8 32.11 237.01 32.18 ;
    RECT 236.8 32.47 237.01 32.54 ;
    RECT 236.34 31.75 236.55 31.82 ;
    RECT 236.34 32.11 236.55 32.18 ;
    RECT 236.34 32.47 236.55 32.54 ;
    RECT 233.48 31.75 233.69 31.82 ;
    RECT 233.48 32.11 233.69 32.18 ;
    RECT 233.48 32.47 233.69 32.54 ;
    RECT 233.02 31.75 233.23 31.82 ;
    RECT 233.02 32.11 233.23 32.18 ;
    RECT 233.02 32.47 233.23 32.54 ;
    RECT 230.16 31.75 230.37 31.82 ;
    RECT 230.16 32.11 230.37 32.18 ;
    RECT 230.16 32.47 230.37 32.54 ;
    RECT 229.7 31.75 229.91 31.82 ;
    RECT 229.7 32.11 229.91 32.18 ;
    RECT 229.7 32.47 229.91 32.54 ;
    RECT 226.84 31.75 227.05 31.82 ;
    RECT 226.84 32.11 227.05 32.18 ;
    RECT 226.84 32.47 227.05 32.54 ;
    RECT 226.38 31.75 226.59 31.82 ;
    RECT 226.38 32.11 226.59 32.18 ;
    RECT 226.38 32.47 226.59 32.54 ;
    RECT 223.52 31.75 223.73 31.82 ;
    RECT 223.52 32.11 223.73 32.18 ;
    RECT 223.52 32.47 223.73 32.54 ;
    RECT 223.06 31.75 223.27 31.82 ;
    RECT 223.06 32.11 223.27 32.18 ;
    RECT 223.06 32.47 223.27 32.54 ;
    RECT 220.2 31.75 220.41 31.82 ;
    RECT 220.2 32.11 220.41 32.18 ;
    RECT 220.2 32.47 220.41 32.54 ;
    RECT 219.74 31.75 219.95 31.82 ;
    RECT 219.74 32.11 219.95 32.18 ;
    RECT 219.74 32.47 219.95 32.54 ;
    RECT 216.88 31.75 217.09 31.82 ;
    RECT 216.88 32.11 217.09 32.18 ;
    RECT 216.88 32.47 217.09 32.54 ;
    RECT 216.42 31.75 216.63 31.82 ;
    RECT 216.42 32.11 216.63 32.18 ;
    RECT 216.42 32.47 216.63 32.54 ;
    RECT 267.91 32.11 267.98 32.18 ;
    RECT 180.36 31.75 180.57 31.82 ;
    RECT 180.36 32.11 180.57 32.18 ;
    RECT 180.36 32.47 180.57 32.54 ;
    RECT 179.9 31.75 180.11 31.82 ;
    RECT 179.9 32.11 180.11 32.18 ;
    RECT 179.9 32.47 180.11 32.54 ;
    RECT 177.04 31.75 177.25 31.82 ;
    RECT 177.04 32.11 177.25 32.18 ;
    RECT 177.04 32.47 177.25 32.54 ;
    RECT 176.58 31.75 176.79 31.82 ;
    RECT 176.58 32.11 176.79 32.18 ;
    RECT 176.58 32.47 176.79 32.54 ;
    RECT 173.72 31.75 173.93 31.82 ;
    RECT 173.72 32.11 173.93 32.18 ;
    RECT 173.72 32.47 173.93 32.54 ;
    RECT 173.26 31.75 173.47 31.82 ;
    RECT 173.26 32.11 173.47 32.18 ;
    RECT 173.26 32.47 173.47 32.54 ;
    RECT 170.4 31.75 170.61 31.82 ;
    RECT 170.4 32.11 170.61 32.18 ;
    RECT 170.4 32.47 170.61 32.54 ;
    RECT 169.94 31.75 170.15 31.82 ;
    RECT 169.94 32.11 170.15 32.18 ;
    RECT 169.94 32.47 170.15 32.54 ;
    RECT 167.08 31.75 167.29 31.82 ;
    RECT 167.08 32.11 167.29 32.18 ;
    RECT 167.08 32.47 167.29 32.54 ;
    RECT 166.62 31.75 166.83 31.82 ;
    RECT 166.62 32.11 166.83 32.18 ;
    RECT 166.62 32.47 166.83 32.54 ;
    RECT 163.76 31.75 163.97 31.82 ;
    RECT 163.76 32.11 163.97 32.18 ;
    RECT 163.76 32.47 163.97 32.54 ;
    RECT 163.3 31.75 163.51 31.82 ;
    RECT 163.3 32.11 163.51 32.18 ;
    RECT 163.3 32.47 163.51 32.54 ;
    RECT 160.44 31.75 160.65 31.82 ;
    RECT 160.44 32.11 160.65 32.18 ;
    RECT 160.44 32.47 160.65 32.54 ;
    RECT 159.98 31.75 160.19 31.82 ;
    RECT 159.98 32.11 160.19 32.18 ;
    RECT 159.98 32.47 160.19 32.54 ;
    RECT 157.12 31.75 157.33 31.82 ;
    RECT 157.12 32.11 157.33 32.18 ;
    RECT 157.12 32.47 157.33 32.54 ;
    RECT 156.66 31.75 156.87 31.82 ;
    RECT 156.66 32.11 156.87 32.18 ;
    RECT 156.66 32.47 156.87 32.54 ;
    RECT 153.8 31.75 154.01 31.82 ;
    RECT 153.8 32.11 154.01 32.18 ;
    RECT 153.8 32.47 154.01 32.54 ;
    RECT 153.34 31.75 153.55 31.82 ;
    RECT 153.34 32.11 153.55 32.18 ;
    RECT 153.34 32.47 153.55 32.54 ;
    RECT 150.48 31.75 150.69 31.82 ;
    RECT 150.48 32.11 150.69 32.18 ;
    RECT 150.48 32.47 150.69 32.54 ;
    RECT 150.02 31.75 150.23 31.82 ;
    RECT 150.02 32.11 150.23 32.18 ;
    RECT 150.02 32.47 150.23 32.54 ;
    RECT 213.56 31.75 213.77 31.82 ;
    RECT 213.56 32.11 213.77 32.18 ;
    RECT 213.56 32.47 213.77 32.54 ;
    RECT 213.1 31.75 213.31 31.82 ;
    RECT 213.1 32.11 213.31 32.18 ;
    RECT 213.1 32.47 213.31 32.54 ;
    RECT 210.24 31.75 210.45 31.82 ;
    RECT 210.24 32.11 210.45 32.18 ;
    RECT 210.24 32.47 210.45 32.54 ;
    RECT 209.78 31.75 209.99 31.82 ;
    RECT 209.78 32.11 209.99 32.18 ;
    RECT 209.78 32.47 209.99 32.54 ;
    RECT 206.92 31.75 207.13 31.82 ;
    RECT 206.92 32.11 207.13 32.18 ;
    RECT 206.92 32.47 207.13 32.54 ;
    RECT 206.46 31.75 206.67 31.82 ;
    RECT 206.46 32.11 206.67 32.18 ;
    RECT 206.46 32.47 206.67 32.54 ;
    RECT 203.6 31.75 203.81 31.82 ;
    RECT 203.6 32.11 203.81 32.18 ;
    RECT 203.6 32.47 203.81 32.54 ;
    RECT 203.14 31.75 203.35 31.82 ;
    RECT 203.14 32.11 203.35 32.18 ;
    RECT 203.14 32.47 203.35 32.54 ;
    RECT 200.28 31.75 200.49 31.82 ;
    RECT 200.28 32.11 200.49 32.18 ;
    RECT 200.28 32.47 200.49 32.54 ;
    RECT 199.82 31.75 200.03 31.82 ;
    RECT 199.82 32.11 200.03 32.18 ;
    RECT 199.82 32.47 200.03 32.54 ;
    RECT 196.96 31.75 197.17 31.82 ;
    RECT 196.96 32.11 197.17 32.18 ;
    RECT 196.96 32.47 197.17 32.54 ;
    RECT 196.5 31.75 196.71 31.82 ;
    RECT 196.5 32.11 196.71 32.18 ;
    RECT 196.5 32.47 196.71 32.54 ;
    RECT 193.64 31.75 193.85 31.82 ;
    RECT 193.64 32.11 193.85 32.18 ;
    RECT 193.64 32.47 193.85 32.54 ;
    RECT 193.18 31.75 193.39 31.82 ;
    RECT 193.18 32.11 193.39 32.18 ;
    RECT 193.18 32.47 193.39 32.54 ;
    RECT 190.32 31.75 190.53 31.82 ;
    RECT 190.32 32.11 190.53 32.18 ;
    RECT 190.32 32.47 190.53 32.54 ;
    RECT 189.86 31.75 190.07 31.82 ;
    RECT 189.86 32.11 190.07 32.18 ;
    RECT 189.86 32.47 190.07 32.54 ;
    RECT 187.0 31.75 187.21 31.82 ;
    RECT 187.0 32.11 187.21 32.18 ;
    RECT 187.0 32.47 187.21 32.54 ;
    RECT 186.54 31.75 186.75 31.82 ;
    RECT 186.54 32.11 186.75 32.18 ;
    RECT 186.54 32.47 186.75 32.54 ;
    RECT 183.68 31.75 183.89 31.82 ;
    RECT 183.68 32.11 183.89 32.18 ;
    RECT 183.68 32.47 183.89 32.54 ;
    RECT 183.22 31.75 183.43 31.82 ;
    RECT 183.22 32.11 183.43 32.18 ;
    RECT 183.22 32.47 183.43 32.54 ;
    RECT 147.485 32.11 147.555 32.18 ;
    RECT 266.68 31.75 266.89 31.82 ;
    RECT 266.68 32.11 266.89 32.18 ;
    RECT 266.68 32.47 266.89 32.54 ;
    RECT 266.22 31.75 266.43 31.82 ;
    RECT 266.22 32.11 266.43 32.18 ;
    RECT 266.22 32.47 266.43 32.54 ;
    RECT 263.36 31.75 263.57 31.82 ;
    RECT 263.36 32.11 263.57 32.18 ;
    RECT 263.36 32.47 263.57 32.54 ;
    RECT 262.9 31.75 263.11 31.82 ;
    RECT 262.9 32.11 263.11 32.18 ;
    RECT 262.9 32.47 263.11 32.54 ;
    RECT 260.04 31.75 260.25 31.82 ;
    RECT 260.04 32.11 260.25 32.18 ;
    RECT 260.04 32.47 260.25 32.54 ;
    RECT 259.58 31.75 259.79 31.82 ;
    RECT 259.58 32.11 259.79 32.18 ;
    RECT 259.58 32.47 259.79 32.54 ;
    RECT 256.72 31.75 256.93 31.82 ;
    RECT 256.72 32.11 256.93 32.18 ;
    RECT 256.72 32.47 256.93 32.54 ;
    RECT 256.26 31.75 256.47 31.82 ;
    RECT 256.26 32.11 256.47 32.18 ;
    RECT 256.26 32.47 256.47 32.54 ;
    RECT 253.4 31.75 253.61 31.82 ;
    RECT 253.4 32.11 253.61 32.18 ;
    RECT 253.4 32.47 253.61 32.54 ;
    RECT 252.94 31.75 253.15 31.82 ;
    RECT 252.94 32.11 253.15 32.18 ;
    RECT 252.94 32.47 253.15 32.54 ;
    RECT 250.08 71.37 250.29 71.44 ;
    RECT 250.08 71.73 250.29 71.8 ;
    RECT 250.08 72.09 250.29 72.16 ;
    RECT 249.62 71.37 249.83 71.44 ;
    RECT 249.62 71.73 249.83 71.8 ;
    RECT 249.62 72.09 249.83 72.16 ;
    RECT 246.76 71.37 246.97 71.44 ;
    RECT 246.76 71.73 246.97 71.8 ;
    RECT 246.76 72.09 246.97 72.16 ;
    RECT 246.3 71.37 246.51 71.44 ;
    RECT 246.3 71.73 246.51 71.8 ;
    RECT 246.3 72.09 246.51 72.16 ;
    RECT 243.44 71.37 243.65 71.44 ;
    RECT 243.44 71.73 243.65 71.8 ;
    RECT 243.44 72.09 243.65 72.16 ;
    RECT 242.98 71.37 243.19 71.44 ;
    RECT 242.98 71.73 243.19 71.8 ;
    RECT 242.98 72.09 243.19 72.16 ;
    RECT 240.12 71.37 240.33 71.44 ;
    RECT 240.12 71.73 240.33 71.8 ;
    RECT 240.12 72.09 240.33 72.16 ;
    RECT 239.66 71.37 239.87 71.44 ;
    RECT 239.66 71.73 239.87 71.8 ;
    RECT 239.66 72.09 239.87 72.16 ;
    RECT 236.8 71.37 237.01 71.44 ;
    RECT 236.8 71.73 237.01 71.8 ;
    RECT 236.8 72.09 237.01 72.16 ;
    RECT 236.34 71.37 236.55 71.44 ;
    RECT 236.34 71.73 236.55 71.8 ;
    RECT 236.34 72.09 236.55 72.16 ;
    RECT 233.48 71.37 233.69 71.44 ;
    RECT 233.48 71.73 233.69 71.8 ;
    RECT 233.48 72.09 233.69 72.16 ;
    RECT 233.02 71.37 233.23 71.44 ;
    RECT 233.02 71.73 233.23 71.8 ;
    RECT 233.02 72.09 233.23 72.16 ;
    RECT 230.16 71.37 230.37 71.44 ;
    RECT 230.16 71.73 230.37 71.8 ;
    RECT 230.16 72.09 230.37 72.16 ;
    RECT 229.7 71.37 229.91 71.44 ;
    RECT 229.7 71.73 229.91 71.8 ;
    RECT 229.7 72.09 229.91 72.16 ;
    RECT 226.84 71.37 227.05 71.44 ;
    RECT 226.84 71.73 227.05 71.8 ;
    RECT 226.84 72.09 227.05 72.16 ;
    RECT 226.38 71.37 226.59 71.44 ;
    RECT 226.38 71.73 226.59 71.8 ;
    RECT 226.38 72.09 226.59 72.16 ;
    RECT 223.52 71.37 223.73 71.44 ;
    RECT 223.52 71.73 223.73 71.8 ;
    RECT 223.52 72.09 223.73 72.16 ;
    RECT 223.06 71.37 223.27 71.44 ;
    RECT 223.06 71.73 223.27 71.8 ;
    RECT 223.06 72.09 223.27 72.16 ;
    RECT 220.2 71.37 220.41 71.44 ;
    RECT 220.2 71.73 220.41 71.8 ;
    RECT 220.2 72.09 220.41 72.16 ;
    RECT 219.74 71.37 219.95 71.44 ;
    RECT 219.74 71.73 219.95 71.8 ;
    RECT 219.74 72.09 219.95 72.16 ;
    RECT 216.88 71.37 217.09 71.44 ;
    RECT 216.88 71.73 217.09 71.8 ;
    RECT 216.88 72.09 217.09 72.16 ;
    RECT 216.42 71.37 216.63 71.44 ;
    RECT 216.42 71.73 216.63 71.8 ;
    RECT 216.42 72.09 216.63 72.16 ;
    RECT 267.91 71.73 267.98 71.8 ;
    RECT 180.36 71.37 180.57 71.44 ;
    RECT 180.36 71.73 180.57 71.8 ;
    RECT 180.36 72.09 180.57 72.16 ;
    RECT 179.9 71.37 180.11 71.44 ;
    RECT 179.9 71.73 180.11 71.8 ;
    RECT 179.9 72.09 180.11 72.16 ;
    RECT 177.04 71.37 177.25 71.44 ;
    RECT 177.04 71.73 177.25 71.8 ;
    RECT 177.04 72.09 177.25 72.16 ;
    RECT 176.58 71.37 176.79 71.44 ;
    RECT 176.58 71.73 176.79 71.8 ;
    RECT 176.58 72.09 176.79 72.16 ;
    RECT 173.72 71.37 173.93 71.44 ;
    RECT 173.72 71.73 173.93 71.8 ;
    RECT 173.72 72.09 173.93 72.16 ;
    RECT 173.26 71.37 173.47 71.44 ;
    RECT 173.26 71.73 173.47 71.8 ;
    RECT 173.26 72.09 173.47 72.16 ;
    RECT 170.4 71.37 170.61 71.44 ;
    RECT 170.4 71.73 170.61 71.8 ;
    RECT 170.4 72.09 170.61 72.16 ;
    RECT 169.94 71.37 170.15 71.44 ;
    RECT 169.94 71.73 170.15 71.8 ;
    RECT 169.94 72.09 170.15 72.16 ;
    RECT 167.08 71.37 167.29 71.44 ;
    RECT 167.08 71.73 167.29 71.8 ;
    RECT 167.08 72.09 167.29 72.16 ;
    RECT 166.62 71.37 166.83 71.44 ;
    RECT 166.62 71.73 166.83 71.8 ;
    RECT 166.62 72.09 166.83 72.16 ;
    RECT 163.76 71.37 163.97 71.44 ;
    RECT 163.76 71.73 163.97 71.8 ;
    RECT 163.76 72.09 163.97 72.16 ;
    RECT 163.3 71.37 163.51 71.44 ;
    RECT 163.3 71.73 163.51 71.8 ;
    RECT 163.3 72.09 163.51 72.16 ;
    RECT 160.44 71.37 160.65 71.44 ;
    RECT 160.44 71.73 160.65 71.8 ;
    RECT 160.44 72.09 160.65 72.16 ;
    RECT 159.98 71.37 160.19 71.44 ;
    RECT 159.98 71.73 160.19 71.8 ;
    RECT 159.98 72.09 160.19 72.16 ;
    RECT 157.12 71.37 157.33 71.44 ;
    RECT 157.12 71.73 157.33 71.8 ;
    RECT 157.12 72.09 157.33 72.16 ;
    RECT 156.66 71.37 156.87 71.44 ;
    RECT 156.66 71.73 156.87 71.8 ;
    RECT 156.66 72.09 156.87 72.16 ;
    RECT 153.8 71.37 154.01 71.44 ;
    RECT 153.8 71.73 154.01 71.8 ;
    RECT 153.8 72.09 154.01 72.16 ;
    RECT 153.34 71.37 153.55 71.44 ;
    RECT 153.34 71.73 153.55 71.8 ;
    RECT 153.34 72.09 153.55 72.16 ;
    RECT 150.48 71.37 150.69 71.44 ;
    RECT 150.48 71.73 150.69 71.8 ;
    RECT 150.48 72.09 150.69 72.16 ;
    RECT 150.02 71.37 150.23 71.44 ;
    RECT 150.02 71.73 150.23 71.8 ;
    RECT 150.02 72.09 150.23 72.16 ;
    RECT 213.56 71.37 213.77 71.44 ;
    RECT 213.56 71.73 213.77 71.8 ;
    RECT 213.56 72.09 213.77 72.16 ;
    RECT 213.1 71.37 213.31 71.44 ;
    RECT 213.1 71.73 213.31 71.8 ;
    RECT 213.1 72.09 213.31 72.16 ;
    RECT 210.24 71.37 210.45 71.44 ;
    RECT 210.24 71.73 210.45 71.8 ;
    RECT 210.24 72.09 210.45 72.16 ;
    RECT 209.78 71.37 209.99 71.44 ;
    RECT 209.78 71.73 209.99 71.8 ;
    RECT 209.78 72.09 209.99 72.16 ;
    RECT 206.92 71.37 207.13 71.44 ;
    RECT 206.92 71.73 207.13 71.8 ;
    RECT 206.92 72.09 207.13 72.16 ;
    RECT 206.46 71.37 206.67 71.44 ;
    RECT 206.46 71.73 206.67 71.8 ;
    RECT 206.46 72.09 206.67 72.16 ;
    RECT 203.6 71.37 203.81 71.44 ;
    RECT 203.6 71.73 203.81 71.8 ;
    RECT 203.6 72.09 203.81 72.16 ;
    RECT 203.14 71.37 203.35 71.44 ;
    RECT 203.14 71.73 203.35 71.8 ;
    RECT 203.14 72.09 203.35 72.16 ;
    RECT 200.28 71.37 200.49 71.44 ;
    RECT 200.28 71.73 200.49 71.8 ;
    RECT 200.28 72.09 200.49 72.16 ;
    RECT 199.82 71.37 200.03 71.44 ;
    RECT 199.82 71.73 200.03 71.8 ;
    RECT 199.82 72.09 200.03 72.16 ;
    RECT 196.96 71.37 197.17 71.44 ;
    RECT 196.96 71.73 197.17 71.8 ;
    RECT 196.96 72.09 197.17 72.16 ;
    RECT 196.5 71.37 196.71 71.44 ;
    RECT 196.5 71.73 196.71 71.8 ;
    RECT 196.5 72.09 196.71 72.16 ;
    RECT 193.64 71.37 193.85 71.44 ;
    RECT 193.64 71.73 193.85 71.8 ;
    RECT 193.64 72.09 193.85 72.16 ;
    RECT 193.18 71.37 193.39 71.44 ;
    RECT 193.18 71.73 193.39 71.8 ;
    RECT 193.18 72.09 193.39 72.16 ;
    RECT 190.32 71.37 190.53 71.44 ;
    RECT 190.32 71.73 190.53 71.8 ;
    RECT 190.32 72.09 190.53 72.16 ;
    RECT 189.86 71.37 190.07 71.44 ;
    RECT 189.86 71.73 190.07 71.8 ;
    RECT 189.86 72.09 190.07 72.16 ;
    RECT 187.0 71.37 187.21 71.44 ;
    RECT 187.0 71.73 187.21 71.8 ;
    RECT 187.0 72.09 187.21 72.16 ;
    RECT 186.54 71.37 186.75 71.44 ;
    RECT 186.54 71.73 186.75 71.8 ;
    RECT 186.54 72.09 186.75 72.16 ;
    RECT 183.68 71.37 183.89 71.44 ;
    RECT 183.68 71.73 183.89 71.8 ;
    RECT 183.68 72.09 183.89 72.16 ;
    RECT 183.22 71.37 183.43 71.44 ;
    RECT 183.22 71.73 183.43 71.8 ;
    RECT 183.22 72.09 183.43 72.16 ;
    RECT 147.485 71.73 147.555 71.8 ;
    RECT 266.68 71.37 266.89 71.44 ;
    RECT 266.68 71.73 266.89 71.8 ;
    RECT 266.68 72.09 266.89 72.16 ;
    RECT 266.22 71.37 266.43 71.44 ;
    RECT 266.22 71.73 266.43 71.8 ;
    RECT 266.22 72.09 266.43 72.16 ;
    RECT 263.36 71.37 263.57 71.44 ;
    RECT 263.36 71.73 263.57 71.8 ;
    RECT 263.36 72.09 263.57 72.16 ;
    RECT 262.9 71.37 263.11 71.44 ;
    RECT 262.9 71.73 263.11 71.8 ;
    RECT 262.9 72.09 263.11 72.16 ;
    RECT 260.04 71.37 260.25 71.44 ;
    RECT 260.04 71.73 260.25 71.8 ;
    RECT 260.04 72.09 260.25 72.16 ;
    RECT 259.58 71.37 259.79 71.44 ;
    RECT 259.58 71.73 259.79 71.8 ;
    RECT 259.58 72.09 259.79 72.16 ;
    RECT 256.72 71.37 256.93 71.44 ;
    RECT 256.72 71.73 256.93 71.8 ;
    RECT 256.72 72.09 256.93 72.16 ;
    RECT 256.26 71.37 256.47 71.44 ;
    RECT 256.26 71.73 256.47 71.8 ;
    RECT 256.26 72.09 256.47 72.16 ;
    RECT 253.4 71.37 253.61 71.44 ;
    RECT 253.4 71.73 253.61 71.8 ;
    RECT 253.4 72.09 253.61 72.16 ;
    RECT 252.94 71.37 253.15 71.44 ;
    RECT 252.94 71.73 253.15 71.8 ;
    RECT 252.94 72.09 253.15 72.16 ;
    RECT 250.08 15.19 250.29 15.26 ;
    RECT 250.08 15.55 250.29 15.62 ;
    RECT 250.08 15.91 250.29 15.98 ;
    RECT 249.62 15.19 249.83 15.26 ;
    RECT 249.62 15.55 249.83 15.62 ;
    RECT 249.62 15.91 249.83 15.98 ;
    RECT 246.76 15.19 246.97 15.26 ;
    RECT 246.76 15.55 246.97 15.62 ;
    RECT 246.76 15.91 246.97 15.98 ;
    RECT 246.3 15.19 246.51 15.26 ;
    RECT 246.3 15.55 246.51 15.62 ;
    RECT 246.3 15.91 246.51 15.98 ;
    RECT 243.44 15.19 243.65 15.26 ;
    RECT 243.44 15.55 243.65 15.62 ;
    RECT 243.44 15.91 243.65 15.98 ;
    RECT 242.98 15.19 243.19 15.26 ;
    RECT 242.98 15.55 243.19 15.62 ;
    RECT 242.98 15.91 243.19 15.98 ;
    RECT 240.12 15.19 240.33 15.26 ;
    RECT 240.12 15.55 240.33 15.62 ;
    RECT 240.12 15.91 240.33 15.98 ;
    RECT 239.66 15.19 239.87 15.26 ;
    RECT 239.66 15.55 239.87 15.62 ;
    RECT 239.66 15.91 239.87 15.98 ;
    RECT 236.8 15.19 237.01 15.26 ;
    RECT 236.8 15.55 237.01 15.62 ;
    RECT 236.8 15.91 237.01 15.98 ;
    RECT 236.34 15.19 236.55 15.26 ;
    RECT 236.34 15.55 236.55 15.62 ;
    RECT 236.34 15.91 236.55 15.98 ;
    RECT 233.48 15.19 233.69 15.26 ;
    RECT 233.48 15.55 233.69 15.62 ;
    RECT 233.48 15.91 233.69 15.98 ;
    RECT 233.02 15.19 233.23 15.26 ;
    RECT 233.02 15.55 233.23 15.62 ;
    RECT 233.02 15.91 233.23 15.98 ;
    RECT 230.16 15.19 230.37 15.26 ;
    RECT 230.16 15.55 230.37 15.62 ;
    RECT 230.16 15.91 230.37 15.98 ;
    RECT 229.7 15.19 229.91 15.26 ;
    RECT 229.7 15.55 229.91 15.62 ;
    RECT 229.7 15.91 229.91 15.98 ;
    RECT 226.84 15.19 227.05 15.26 ;
    RECT 226.84 15.55 227.05 15.62 ;
    RECT 226.84 15.91 227.05 15.98 ;
    RECT 226.38 15.19 226.59 15.26 ;
    RECT 226.38 15.55 226.59 15.62 ;
    RECT 226.38 15.91 226.59 15.98 ;
    RECT 223.52 15.19 223.73 15.26 ;
    RECT 223.52 15.55 223.73 15.62 ;
    RECT 223.52 15.91 223.73 15.98 ;
    RECT 223.06 15.19 223.27 15.26 ;
    RECT 223.06 15.55 223.27 15.62 ;
    RECT 223.06 15.91 223.27 15.98 ;
    RECT 220.2 15.19 220.41 15.26 ;
    RECT 220.2 15.55 220.41 15.62 ;
    RECT 220.2 15.91 220.41 15.98 ;
    RECT 219.74 15.19 219.95 15.26 ;
    RECT 219.74 15.55 219.95 15.62 ;
    RECT 219.74 15.91 219.95 15.98 ;
    RECT 216.88 15.19 217.09 15.26 ;
    RECT 216.88 15.55 217.09 15.62 ;
    RECT 216.88 15.91 217.09 15.98 ;
    RECT 216.42 15.19 216.63 15.26 ;
    RECT 216.42 15.55 216.63 15.62 ;
    RECT 216.42 15.91 216.63 15.98 ;
    RECT 267.91 15.55 267.98 15.62 ;
    RECT 180.36 15.19 180.57 15.26 ;
    RECT 180.36 15.55 180.57 15.62 ;
    RECT 180.36 15.91 180.57 15.98 ;
    RECT 179.9 15.19 180.11 15.26 ;
    RECT 179.9 15.55 180.11 15.62 ;
    RECT 179.9 15.91 180.11 15.98 ;
    RECT 177.04 15.19 177.25 15.26 ;
    RECT 177.04 15.55 177.25 15.62 ;
    RECT 177.04 15.91 177.25 15.98 ;
    RECT 176.58 15.19 176.79 15.26 ;
    RECT 176.58 15.55 176.79 15.62 ;
    RECT 176.58 15.91 176.79 15.98 ;
    RECT 173.72 15.19 173.93 15.26 ;
    RECT 173.72 15.55 173.93 15.62 ;
    RECT 173.72 15.91 173.93 15.98 ;
    RECT 173.26 15.19 173.47 15.26 ;
    RECT 173.26 15.55 173.47 15.62 ;
    RECT 173.26 15.91 173.47 15.98 ;
    RECT 170.4 15.19 170.61 15.26 ;
    RECT 170.4 15.55 170.61 15.62 ;
    RECT 170.4 15.91 170.61 15.98 ;
    RECT 169.94 15.19 170.15 15.26 ;
    RECT 169.94 15.55 170.15 15.62 ;
    RECT 169.94 15.91 170.15 15.98 ;
    RECT 167.08 15.19 167.29 15.26 ;
    RECT 167.08 15.55 167.29 15.62 ;
    RECT 167.08 15.91 167.29 15.98 ;
    RECT 166.62 15.19 166.83 15.26 ;
    RECT 166.62 15.55 166.83 15.62 ;
    RECT 166.62 15.91 166.83 15.98 ;
    RECT 163.76 15.19 163.97 15.26 ;
    RECT 163.76 15.55 163.97 15.62 ;
    RECT 163.76 15.91 163.97 15.98 ;
    RECT 163.3 15.19 163.51 15.26 ;
    RECT 163.3 15.55 163.51 15.62 ;
    RECT 163.3 15.91 163.51 15.98 ;
    RECT 160.44 15.19 160.65 15.26 ;
    RECT 160.44 15.55 160.65 15.62 ;
    RECT 160.44 15.91 160.65 15.98 ;
    RECT 159.98 15.19 160.19 15.26 ;
    RECT 159.98 15.55 160.19 15.62 ;
    RECT 159.98 15.91 160.19 15.98 ;
    RECT 157.12 15.19 157.33 15.26 ;
    RECT 157.12 15.55 157.33 15.62 ;
    RECT 157.12 15.91 157.33 15.98 ;
    RECT 156.66 15.19 156.87 15.26 ;
    RECT 156.66 15.55 156.87 15.62 ;
    RECT 156.66 15.91 156.87 15.98 ;
    RECT 153.8 15.19 154.01 15.26 ;
    RECT 153.8 15.55 154.01 15.62 ;
    RECT 153.8 15.91 154.01 15.98 ;
    RECT 153.34 15.19 153.55 15.26 ;
    RECT 153.34 15.55 153.55 15.62 ;
    RECT 153.34 15.91 153.55 15.98 ;
    RECT 150.48 15.19 150.69 15.26 ;
    RECT 150.48 15.55 150.69 15.62 ;
    RECT 150.48 15.91 150.69 15.98 ;
    RECT 150.02 15.19 150.23 15.26 ;
    RECT 150.02 15.55 150.23 15.62 ;
    RECT 150.02 15.91 150.23 15.98 ;
    RECT 213.56 15.19 213.77 15.26 ;
    RECT 213.56 15.55 213.77 15.62 ;
    RECT 213.56 15.91 213.77 15.98 ;
    RECT 213.1 15.19 213.31 15.26 ;
    RECT 213.1 15.55 213.31 15.62 ;
    RECT 213.1 15.91 213.31 15.98 ;
    RECT 210.24 15.19 210.45 15.26 ;
    RECT 210.24 15.55 210.45 15.62 ;
    RECT 210.24 15.91 210.45 15.98 ;
    RECT 209.78 15.19 209.99 15.26 ;
    RECT 209.78 15.55 209.99 15.62 ;
    RECT 209.78 15.91 209.99 15.98 ;
    RECT 206.92 15.19 207.13 15.26 ;
    RECT 206.92 15.55 207.13 15.62 ;
    RECT 206.92 15.91 207.13 15.98 ;
    RECT 206.46 15.19 206.67 15.26 ;
    RECT 206.46 15.55 206.67 15.62 ;
    RECT 206.46 15.91 206.67 15.98 ;
    RECT 203.6 15.19 203.81 15.26 ;
    RECT 203.6 15.55 203.81 15.62 ;
    RECT 203.6 15.91 203.81 15.98 ;
    RECT 203.14 15.19 203.35 15.26 ;
    RECT 203.14 15.55 203.35 15.62 ;
    RECT 203.14 15.91 203.35 15.98 ;
    RECT 200.28 15.19 200.49 15.26 ;
    RECT 200.28 15.55 200.49 15.62 ;
    RECT 200.28 15.91 200.49 15.98 ;
    RECT 199.82 15.19 200.03 15.26 ;
    RECT 199.82 15.55 200.03 15.62 ;
    RECT 199.82 15.91 200.03 15.98 ;
    RECT 196.96 15.19 197.17 15.26 ;
    RECT 196.96 15.55 197.17 15.62 ;
    RECT 196.96 15.91 197.17 15.98 ;
    RECT 196.5 15.19 196.71 15.26 ;
    RECT 196.5 15.55 196.71 15.62 ;
    RECT 196.5 15.91 196.71 15.98 ;
    RECT 193.64 15.19 193.85 15.26 ;
    RECT 193.64 15.55 193.85 15.62 ;
    RECT 193.64 15.91 193.85 15.98 ;
    RECT 193.18 15.19 193.39 15.26 ;
    RECT 193.18 15.55 193.39 15.62 ;
    RECT 193.18 15.91 193.39 15.98 ;
    RECT 190.32 15.19 190.53 15.26 ;
    RECT 190.32 15.55 190.53 15.62 ;
    RECT 190.32 15.91 190.53 15.98 ;
    RECT 189.86 15.19 190.07 15.26 ;
    RECT 189.86 15.55 190.07 15.62 ;
    RECT 189.86 15.91 190.07 15.98 ;
    RECT 187.0 15.19 187.21 15.26 ;
    RECT 187.0 15.55 187.21 15.62 ;
    RECT 187.0 15.91 187.21 15.98 ;
    RECT 186.54 15.19 186.75 15.26 ;
    RECT 186.54 15.55 186.75 15.62 ;
    RECT 186.54 15.91 186.75 15.98 ;
    RECT 183.68 15.19 183.89 15.26 ;
    RECT 183.68 15.55 183.89 15.62 ;
    RECT 183.68 15.91 183.89 15.98 ;
    RECT 183.22 15.19 183.43 15.26 ;
    RECT 183.22 15.55 183.43 15.62 ;
    RECT 183.22 15.91 183.43 15.98 ;
    RECT 147.485 15.55 147.555 15.62 ;
    RECT 266.68 15.19 266.89 15.26 ;
    RECT 266.68 15.55 266.89 15.62 ;
    RECT 266.68 15.91 266.89 15.98 ;
    RECT 266.22 15.19 266.43 15.26 ;
    RECT 266.22 15.55 266.43 15.62 ;
    RECT 266.22 15.91 266.43 15.98 ;
    RECT 263.36 15.19 263.57 15.26 ;
    RECT 263.36 15.55 263.57 15.62 ;
    RECT 263.36 15.91 263.57 15.98 ;
    RECT 262.9 15.19 263.11 15.26 ;
    RECT 262.9 15.55 263.11 15.62 ;
    RECT 262.9 15.91 263.11 15.98 ;
    RECT 260.04 15.19 260.25 15.26 ;
    RECT 260.04 15.55 260.25 15.62 ;
    RECT 260.04 15.91 260.25 15.98 ;
    RECT 259.58 15.19 259.79 15.26 ;
    RECT 259.58 15.55 259.79 15.62 ;
    RECT 259.58 15.91 259.79 15.98 ;
    RECT 256.72 15.19 256.93 15.26 ;
    RECT 256.72 15.55 256.93 15.62 ;
    RECT 256.72 15.91 256.93 15.98 ;
    RECT 256.26 15.19 256.47 15.26 ;
    RECT 256.26 15.55 256.47 15.62 ;
    RECT 256.26 15.91 256.47 15.98 ;
    RECT 253.4 15.19 253.61 15.26 ;
    RECT 253.4 15.55 253.61 15.62 ;
    RECT 253.4 15.91 253.61 15.98 ;
    RECT 252.94 15.19 253.15 15.26 ;
    RECT 252.94 15.55 253.15 15.62 ;
    RECT 252.94 15.91 253.15 15.98 ;
    RECT 250.08 31.03 250.29 31.1 ;
    RECT 250.08 31.39 250.29 31.46 ;
    RECT 250.08 31.75 250.29 31.82 ;
    RECT 249.62 31.03 249.83 31.1 ;
    RECT 249.62 31.39 249.83 31.46 ;
    RECT 249.62 31.75 249.83 31.82 ;
    RECT 246.76 31.03 246.97 31.1 ;
    RECT 246.76 31.39 246.97 31.46 ;
    RECT 246.76 31.75 246.97 31.82 ;
    RECT 246.3 31.03 246.51 31.1 ;
    RECT 246.3 31.39 246.51 31.46 ;
    RECT 246.3 31.75 246.51 31.82 ;
    RECT 243.44 31.03 243.65 31.1 ;
    RECT 243.44 31.39 243.65 31.46 ;
    RECT 243.44 31.75 243.65 31.82 ;
    RECT 242.98 31.03 243.19 31.1 ;
    RECT 242.98 31.39 243.19 31.46 ;
    RECT 242.98 31.75 243.19 31.82 ;
    RECT 240.12 31.03 240.33 31.1 ;
    RECT 240.12 31.39 240.33 31.46 ;
    RECT 240.12 31.75 240.33 31.82 ;
    RECT 239.66 31.03 239.87 31.1 ;
    RECT 239.66 31.39 239.87 31.46 ;
    RECT 239.66 31.75 239.87 31.82 ;
    RECT 236.8 31.03 237.01 31.1 ;
    RECT 236.8 31.39 237.01 31.46 ;
    RECT 236.8 31.75 237.01 31.82 ;
    RECT 236.34 31.03 236.55 31.1 ;
    RECT 236.34 31.39 236.55 31.46 ;
    RECT 236.34 31.75 236.55 31.82 ;
    RECT 233.48 31.03 233.69 31.1 ;
    RECT 233.48 31.39 233.69 31.46 ;
    RECT 233.48 31.75 233.69 31.82 ;
    RECT 233.02 31.03 233.23 31.1 ;
    RECT 233.02 31.39 233.23 31.46 ;
    RECT 233.02 31.75 233.23 31.82 ;
    RECT 230.16 31.03 230.37 31.1 ;
    RECT 230.16 31.39 230.37 31.46 ;
    RECT 230.16 31.75 230.37 31.82 ;
    RECT 229.7 31.03 229.91 31.1 ;
    RECT 229.7 31.39 229.91 31.46 ;
    RECT 229.7 31.75 229.91 31.82 ;
    RECT 226.84 31.03 227.05 31.1 ;
    RECT 226.84 31.39 227.05 31.46 ;
    RECT 226.84 31.75 227.05 31.82 ;
    RECT 226.38 31.03 226.59 31.1 ;
    RECT 226.38 31.39 226.59 31.46 ;
    RECT 226.38 31.75 226.59 31.82 ;
    RECT 223.52 31.03 223.73 31.1 ;
    RECT 223.52 31.39 223.73 31.46 ;
    RECT 223.52 31.75 223.73 31.82 ;
    RECT 223.06 31.03 223.27 31.1 ;
    RECT 223.06 31.39 223.27 31.46 ;
    RECT 223.06 31.75 223.27 31.82 ;
    RECT 220.2 31.03 220.41 31.1 ;
    RECT 220.2 31.39 220.41 31.46 ;
    RECT 220.2 31.75 220.41 31.82 ;
    RECT 219.74 31.03 219.95 31.1 ;
    RECT 219.74 31.39 219.95 31.46 ;
    RECT 219.74 31.75 219.95 31.82 ;
    RECT 216.88 31.03 217.09 31.1 ;
    RECT 216.88 31.39 217.09 31.46 ;
    RECT 216.88 31.75 217.09 31.82 ;
    RECT 216.42 31.03 216.63 31.1 ;
    RECT 216.42 31.39 216.63 31.46 ;
    RECT 216.42 31.75 216.63 31.82 ;
    RECT 267.91 31.39 267.98 31.46 ;
    RECT 180.36 31.03 180.57 31.1 ;
    RECT 180.36 31.39 180.57 31.46 ;
    RECT 180.36 31.75 180.57 31.82 ;
    RECT 179.9 31.03 180.11 31.1 ;
    RECT 179.9 31.39 180.11 31.46 ;
    RECT 179.9 31.75 180.11 31.82 ;
    RECT 177.04 31.03 177.25 31.1 ;
    RECT 177.04 31.39 177.25 31.46 ;
    RECT 177.04 31.75 177.25 31.82 ;
    RECT 176.58 31.03 176.79 31.1 ;
    RECT 176.58 31.39 176.79 31.46 ;
    RECT 176.58 31.75 176.79 31.82 ;
    RECT 173.72 31.03 173.93 31.1 ;
    RECT 173.72 31.39 173.93 31.46 ;
    RECT 173.72 31.75 173.93 31.82 ;
    RECT 173.26 31.03 173.47 31.1 ;
    RECT 173.26 31.39 173.47 31.46 ;
    RECT 173.26 31.75 173.47 31.82 ;
    RECT 170.4 31.03 170.61 31.1 ;
    RECT 170.4 31.39 170.61 31.46 ;
    RECT 170.4 31.75 170.61 31.82 ;
    RECT 169.94 31.03 170.15 31.1 ;
    RECT 169.94 31.39 170.15 31.46 ;
    RECT 169.94 31.75 170.15 31.82 ;
    RECT 167.08 31.03 167.29 31.1 ;
    RECT 167.08 31.39 167.29 31.46 ;
    RECT 167.08 31.75 167.29 31.82 ;
    RECT 166.62 31.03 166.83 31.1 ;
    RECT 166.62 31.39 166.83 31.46 ;
    RECT 166.62 31.75 166.83 31.82 ;
    RECT 163.76 31.03 163.97 31.1 ;
    RECT 163.76 31.39 163.97 31.46 ;
    RECT 163.76 31.75 163.97 31.82 ;
    RECT 163.3 31.03 163.51 31.1 ;
    RECT 163.3 31.39 163.51 31.46 ;
    RECT 163.3 31.75 163.51 31.82 ;
    RECT 160.44 31.03 160.65 31.1 ;
    RECT 160.44 31.39 160.65 31.46 ;
    RECT 160.44 31.75 160.65 31.82 ;
    RECT 159.98 31.03 160.19 31.1 ;
    RECT 159.98 31.39 160.19 31.46 ;
    RECT 159.98 31.75 160.19 31.82 ;
    RECT 157.12 31.03 157.33 31.1 ;
    RECT 157.12 31.39 157.33 31.46 ;
    RECT 157.12 31.75 157.33 31.82 ;
    RECT 156.66 31.03 156.87 31.1 ;
    RECT 156.66 31.39 156.87 31.46 ;
    RECT 156.66 31.75 156.87 31.82 ;
    RECT 153.8 31.03 154.01 31.1 ;
    RECT 153.8 31.39 154.01 31.46 ;
    RECT 153.8 31.75 154.01 31.82 ;
    RECT 153.34 31.03 153.55 31.1 ;
    RECT 153.34 31.39 153.55 31.46 ;
    RECT 153.34 31.75 153.55 31.82 ;
    RECT 150.48 31.03 150.69 31.1 ;
    RECT 150.48 31.39 150.69 31.46 ;
    RECT 150.48 31.75 150.69 31.82 ;
    RECT 150.02 31.03 150.23 31.1 ;
    RECT 150.02 31.39 150.23 31.46 ;
    RECT 150.02 31.75 150.23 31.82 ;
    RECT 213.56 31.03 213.77 31.1 ;
    RECT 213.56 31.39 213.77 31.46 ;
    RECT 213.56 31.75 213.77 31.82 ;
    RECT 213.1 31.03 213.31 31.1 ;
    RECT 213.1 31.39 213.31 31.46 ;
    RECT 213.1 31.75 213.31 31.82 ;
    RECT 210.24 31.03 210.45 31.1 ;
    RECT 210.24 31.39 210.45 31.46 ;
    RECT 210.24 31.75 210.45 31.82 ;
    RECT 209.78 31.03 209.99 31.1 ;
    RECT 209.78 31.39 209.99 31.46 ;
    RECT 209.78 31.75 209.99 31.82 ;
    RECT 206.92 31.03 207.13 31.1 ;
    RECT 206.92 31.39 207.13 31.46 ;
    RECT 206.92 31.75 207.13 31.82 ;
    RECT 206.46 31.03 206.67 31.1 ;
    RECT 206.46 31.39 206.67 31.46 ;
    RECT 206.46 31.75 206.67 31.82 ;
    RECT 203.6 31.03 203.81 31.1 ;
    RECT 203.6 31.39 203.81 31.46 ;
    RECT 203.6 31.75 203.81 31.82 ;
    RECT 203.14 31.03 203.35 31.1 ;
    RECT 203.14 31.39 203.35 31.46 ;
    RECT 203.14 31.75 203.35 31.82 ;
    RECT 200.28 31.03 200.49 31.1 ;
    RECT 200.28 31.39 200.49 31.46 ;
    RECT 200.28 31.75 200.49 31.82 ;
    RECT 199.82 31.03 200.03 31.1 ;
    RECT 199.82 31.39 200.03 31.46 ;
    RECT 199.82 31.75 200.03 31.82 ;
    RECT 196.96 31.03 197.17 31.1 ;
    RECT 196.96 31.39 197.17 31.46 ;
    RECT 196.96 31.75 197.17 31.82 ;
    RECT 196.5 31.03 196.71 31.1 ;
    RECT 196.5 31.39 196.71 31.46 ;
    RECT 196.5 31.75 196.71 31.82 ;
    RECT 193.64 31.03 193.85 31.1 ;
    RECT 193.64 31.39 193.85 31.46 ;
    RECT 193.64 31.75 193.85 31.82 ;
    RECT 193.18 31.03 193.39 31.1 ;
    RECT 193.18 31.39 193.39 31.46 ;
    RECT 193.18 31.75 193.39 31.82 ;
    RECT 190.32 31.03 190.53 31.1 ;
    RECT 190.32 31.39 190.53 31.46 ;
    RECT 190.32 31.75 190.53 31.82 ;
    RECT 189.86 31.03 190.07 31.1 ;
    RECT 189.86 31.39 190.07 31.46 ;
    RECT 189.86 31.75 190.07 31.82 ;
    RECT 187.0 31.03 187.21 31.1 ;
    RECT 187.0 31.39 187.21 31.46 ;
    RECT 187.0 31.75 187.21 31.82 ;
    RECT 186.54 31.03 186.75 31.1 ;
    RECT 186.54 31.39 186.75 31.46 ;
    RECT 186.54 31.75 186.75 31.82 ;
    RECT 183.68 31.03 183.89 31.1 ;
    RECT 183.68 31.39 183.89 31.46 ;
    RECT 183.68 31.75 183.89 31.82 ;
    RECT 183.22 31.03 183.43 31.1 ;
    RECT 183.22 31.39 183.43 31.46 ;
    RECT 183.22 31.75 183.43 31.82 ;
    RECT 147.485 31.39 147.555 31.46 ;
    RECT 266.68 31.03 266.89 31.1 ;
    RECT 266.68 31.39 266.89 31.46 ;
    RECT 266.68 31.75 266.89 31.82 ;
    RECT 266.22 31.03 266.43 31.1 ;
    RECT 266.22 31.39 266.43 31.46 ;
    RECT 266.22 31.75 266.43 31.82 ;
    RECT 263.36 31.03 263.57 31.1 ;
    RECT 263.36 31.39 263.57 31.46 ;
    RECT 263.36 31.75 263.57 31.82 ;
    RECT 262.9 31.03 263.11 31.1 ;
    RECT 262.9 31.39 263.11 31.46 ;
    RECT 262.9 31.75 263.11 31.82 ;
    RECT 260.04 31.03 260.25 31.1 ;
    RECT 260.04 31.39 260.25 31.46 ;
    RECT 260.04 31.75 260.25 31.82 ;
    RECT 259.58 31.03 259.79 31.1 ;
    RECT 259.58 31.39 259.79 31.46 ;
    RECT 259.58 31.75 259.79 31.82 ;
    RECT 256.72 31.03 256.93 31.1 ;
    RECT 256.72 31.39 256.93 31.46 ;
    RECT 256.72 31.75 256.93 31.82 ;
    RECT 256.26 31.03 256.47 31.1 ;
    RECT 256.26 31.39 256.47 31.46 ;
    RECT 256.26 31.75 256.47 31.82 ;
    RECT 253.4 31.03 253.61 31.1 ;
    RECT 253.4 31.39 253.61 31.46 ;
    RECT 253.4 31.75 253.61 31.82 ;
    RECT 252.94 31.03 253.15 31.1 ;
    RECT 252.94 31.39 253.15 31.46 ;
    RECT 252.94 31.75 253.15 31.82 ;
    RECT 250.08 70.65 250.29 70.72 ;
    RECT 250.08 71.01 250.29 71.08 ;
    RECT 250.08 71.37 250.29 71.44 ;
    RECT 249.62 70.65 249.83 70.72 ;
    RECT 249.62 71.01 249.83 71.08 ;
    RECT 249.62 71.37 249.83 71.44 ;
    RECT 246.76 70.65 246.97 70.72 ;
    RECT 246.76 71.01 246.97 71.08 ;
    RECT 246.76 71.37 246.97 71.44 ;
    RECT 246.3 70.65 246.51 70.72 ;
    RECT 246.3 71.01 246.51 71.08 ;
    RECT 246.3 71.37 246.51 71.44 ;
    RECT 243.44 70.65 243.65 70.72 ;
    RECT 243.44 71.01 243.65 71.08 ;
    RECT 243.44 71.37 243.65 71.44 ;
    RECT 242.98 70.65 243.19 70.72 ;
    RECT 242.98 71.01 243.19 71.08 ;
    RECT 242.98 71.37 243.19 71.44 ;
    RECT 240.12 70.65 240.33 70.72 ;
    RECT 240.12 71.01 240.33 71.08 ;
    RECT 240.12 71.37 240.33 71.44 ;
    RECT 239.66 70.65 239.87 70.72 ;
    RECT 239.66 71.01 239.87 71.08 ;
    RECT 239.66 71.37 239.87 71.44 ;
    RECT 236.8 70.65 237.01 70.72 ;
    RECT 236.8 71.01 237.01 71.08 ;
    RECT 236.8 71.37 237.01 71.44 ;
    RECT 236.34 70.65 236.55 70.72 ;
    RECT 236.34 71.01 236.55 71.08 ;
    RECT 236.34 71.37 236.55 71.44 ;
    RECT 233.48 70.65 233.69 70.72 ;
    RECT 233.48 71.01 233.69 71.08 ;
    RECT 233.48 71.37 233.69 71.44 ;
    RECT 233.02 70.65 233.23 70.72 ;
    RECT 233.02 71.01 233.23 71.08 ;
    RECT 233.02 71.37 233.23 71.44 ;
    RECT 230.16 70.65 230.37 70.72 ;
    RECT 230.16 71.01 230.37 71.08 ;
    RECT 230.16 71.37 230.37 71.44 ;
    RECT 229.7 70.65 229.91 70.72 ;
    RECT 229.7 71.01 229.91 71.08 ;
    RECT 229.7 71.37 229.91 71.44 ;
    RECT 226.84 70.65 227.05 70.72 ;
    RECT 226.84 71.01 227.05 71.08 ;
    RECT 226.84 71.37 227.05 71.44 ;
    RECT 226.38 70.65 226.59 70.72 ;
    RECT 226.38 71.01 226.59 71.08 ;
    RECT 226.38 71.37 226.59 71.44 ;
    RECT 223.52 70.65 223.73 70.72 ;
    RECT 223.52 71.01 223.73 71.08 ;
    RECT 223.52 71.37 223.73 71.44 ;
    RECT 223.06 70.65 223.27 70.72 ;
    RECT 223.06 71.01 223.27 71.08 ;
    RECT 223.06 71.37 223.27 71.44 ;
    RECT 220.2 70.65 220.41 70.72 ;
    RECT 220.2 71.01 220.41 71.08 ;
    RECT 220.2 71.37 220.41 71.44 ;
    RECT 219.74 70.65 219.95 70.72 ;
    RECT 219.74 71.01 219.95 71.08 ;
    RECT 219.74 71.37 219.95 71.44 ;
    RECT 216.88 70.65 217.09 70.72 ;
    RECT 216.88 71.01 217.09 71.08 ;
    RECT 216.88 71.37 217.09 71.44 ;
    RECT 216.42 70.65 216.63 70.72 ;
    RECT 216.42 71.01 216.63 71.08 ;
    RECT 216.42 71.37 216.63 71.44 ;
    RECT 267.91 71.01 267.98 71.08 ;
    RECT 180.36 70.65 180.57 70.72 ;
    RECT 180.36 71.01 180.57 71.08 ;
    RECT 180.36 71.37 180.57 71.44 ;
    RECT 179.9 70.65 180.11 70.72 ;
    RECT 179.9 71.01 180.11 71.08 ;
    RECT 179.9 71.37 180.11 71.44 ;
    RECT 177.04 70.65 177.25 70.72 ;
    RECT 177.04 71.01 177.25 71.08 ;
    RECT 177.04 71.37 177.25 71.44 ;
    RECT 176.58 70.65 176.79 70.72 ;
    RECT 176.58 71.01 176.79 71.08 ;
    RECT 176.58 71.37 176.79 71.44 ;
    RECT 173.72 70.65 173.93 70.72 ;
    RECT 173.72 71.01 173.93 71.08 ;
    RECT 173.72 71.37 173.93 71.44 ;
    RECT 173.26 70.65 173.47 70.72 ;
    RECT 173.26 71.01 173.47 71.08 ;
    RECT 173.26 71.37 173.47 71.44 ;
    RECT 170.4 70.65 170.61 70.72 ;
    RECT 170.4 71.01 170.61 71.08 ;
    RECT 170.4 71.37 170.61 71.44 ;
    RECT 169.94 70.65 170.15 70.72 ;
    RECT 169.94 71.01 170.15 71.08 ;
    RECT 169.94 71.37 170.15 71.44 ;
    RECT 167.08 70.65 167.29 70.72 ;
    RECT 167.08 71.01 167.29 71.08 ;
    RECT 167.08 71.37 167.29 71.44 ;
    RECT 166.62 70.65 166.83 70.72 ;
    RECT 166.62 71.01 166.83 71.08 ;
    RECT 166.62 71.37 166.83 71.44 ;
    RECT 163.76 70.65 163.97 70.72 ;
    RECT 163.76 71.01 163.97 71.08 ;
    RECT 163.76 71.37 163.97 71.44 ;
    RECT 163.3 70.65 163.51 70.72 ;
    RECT 163.3 71.01 163.51 71.08 ;
    RECT 163.3 71.37 163.51 71.44 ;
    RECT 160.44 70.65 160.65 70.72 ;
    RECT 160.44 71.01 160.65 71.08 ;
    RECT 160.44 71.37 160.65 71.44 ;
    RECT 159.98 70.65 160.19 70.72 ;
    RECT 159.98 71.01 160.19 71.08 ;
    RECT 159.98 71.37 160.19 71.44 ;
    RECT 157.12 70.65 157.33 70.72 ;
    RECT 157.12 71.01 157.33 71.08 ;
    RECT 157.12 71.37 157.33 71.44 ;
    RECT 156.66 70.65 156.87 70.72 ;
    RECT 156.66 71.01 156.87 71.08 ;
    RECT 156.66 71.37 156.87 71.44 ;
    RECT 153.8 70.65 154.01 70.72 ;
    RECT 153.8 71.01 154.01 71.08 ;
    RECT 153.8 71.37 154.01 71.44 ;
    RECT 153.34 70.65 153.55 70.72 ;
    RECT 153.34 71.01 153.55 71.08 ;
    RECT 153.34 71.37 153.55 71.44 ;
    RECT 150.48 70.65 150.69 70.72 ;
    RECT 150.48 71.01 150.69 71.08 ;
    RECT 150.48 71.37 150.69 71.44 ;
    RECT 150.02 70.65 150.23 70.72 ;
    RECT 150.02 71.01 150.23 71.08 ;
    RECT 150.02 71.37 150.23 71.44 ;
    RECT 213.56 70.65 213.77 70.72 ;
    RECT 213.56 71.01 213.77 71.08 ;
    RECT 213.56 71.37 213.77 71.44 ;
    RECT 213.1 70.65 213.31 70.72 ;
    RECT 213.1 71.01 213.31 71.08 ;
    RECT 213.1 71.37 213.31 71.44 ;
    RECT 210.24 70.65 210.45 70.72 ;
    RECT 210.24 71.01 210.45 71.08 ;
    RECT 210.24 71.37 210.45 71.44 ;
    RECT 209.78 70.65 209.99 70.72 ;
    RECT 209.78 71.01 209.99 71.08 ;
    RECT 209.78 71.37 209.99 71.44 ;
    RECT 206.92 70.65 207.13 70.72 ;
    RECT 206.92 71.01 207.13 71.08 ;
    RECT 206.92 71.37 207.13 71.44 ;
    RECT 206.46 70.65 206.67 70.72 ;
    RECT 206.46 71.01 206.67 71.08 ;
    RECT 206.46 71.37 206.67 71.44 ;
    RECT 203.6 70.65 203.81 70.72 ;
    RECT 203.6 71.01 203.81 71.08 ;
    RECT 203.6 71.37 203.81 71.44 ;
    RECT 203.14 70.65 203.35 70.72 ;
    RECT 203.14 71.01 203.35 71.08 ;
    RECT 203.14 71.37 203.35 71.44 ;
    RECT 200.28 70.65 200.49 70.72 ;
    RECT 200.28 71.01 200.49 71.08 ;
    RECT 200.28 71.37 200.49 71.44 ;
    RECT 199.82 70.65 200.03 70.72 ;
    RECT 199.82 71.01 200.03 71.08 ;
    RECT 199.82 71.37 200.03 71.44 ;
    RECT 196.96 70.65 197.17 70.72 ;
    RECT 196.96 71.01 197.17 71.08 ;
    RECT 196.96 71.37 197.17 71.44 ;
    RECT 196.5 70.65 196.71 70.72 ;
    RECT 196.5 71.01 196.71 71.08 ;
    RECT 196.5 71.37 196.71 71.44 ;
    RECT 193.64 70.65 193.85 70.72 ;
    RECT 193.64 71.01 193.85 71.08 ;
    RECT 193.64 71.37 193.85 71.44 ;
    RECT 193.18 70.65 193.39 70.72 ;
    RECT 193.18 71.01 193.39 71.08 ;
    RECT 193.18 71.37 193.39 71.44 ;
    RECT 190.32 70.65 190.53 70.72 ;
    RECT 190.32 71.01 190.53 71.08 ;
    RECT 190.32 71.37 190.53 71.44 ;
    RECT 189.86 70.65 190.07 70.72 ;
    RECT 189.86 71.01 190.07 71.08 ;
    RECT 189.86 71.37 190.07 71.44 ;
    RECT 187.0 70.65 187.21 70.72 ;
    RECT 187.0 71.01 187.21 71.08 ;
    RECT 187.0 71.37 187.21 71.44 ;
    RECT 186.54 70.65 186.75 70.72 ;
    RECT 186.54 71.01 186.75 71.08 ;
    RECT 186.54 71.37 186.75 71.44 ;
    RECT 183.68 70.65 183.89 70.72 ;
    RECT 183.68 71.01 183.89 71.08 ;
    RECT 183.68 71.37 183.89 71.44 ;
    RECT 183.22 70.65 183.43 70.72 ;
    RECT 183.22 71.01 183.43 71.08 ;
    RECT 183.22 71.37 183.43 71.44 ;
    RECT 147.485 71.01 147.555 71.08 ;
    RECT 266.68 70.65 266.89 70.72 ;
    RECT 266.68 71.01 266.89 71.08 ;
    RECT 266.68 71.37 266.89 71.44 ;
    RECT 266.22 70.65 266.43 70.72 ;
    RECT 266.22 71.01 266.43 71.08 ;
    RECT 266.22 71.37 266.43 71.44 ;
    RECT 263.36 70.65 263.57 70.72 ;
    RECT 263.36 71.01 263.57 71.08 ;
    RECT 263.36 71.37 263.57 71.44 ;
    RECT 262.9 70.65 263.11 70.72 ;
    RECT 262.9 71.01 263.11 71.08 ;
    RECT 262.9 71.37 263.11 71.44 ;
    RECT 260.04 70.65 260.25 70.72 ;
    RECT 260.04 71.01 260.25 71.08 ;
    RECT 260.04 71.37 260.25 71.44 ;
    RECT 259.58 70.65 259.79 70.72 ;
    RECT 259.58 71.01 259.79 71.08 ;
    RECT 259.58 71.37 259.79 71.44 ;
    RECT 256.72 70.65 256.93 70.72 ;
    RECT 256.72 71.01 256.93 71.08 ;
    RECT 256.72 71.37 256.93 71.44 ;
    RECT 256.26 70.65 256.47 70.72 ;
    RECT 256.26 71.01 256.47 71.08 ;
    RECT 256.26 71.37 256.47 71.44 ;
    RECT 253.4 70.65 253.61 70.72 ;
    RECT 253.4 71.01 253.61 71.08 ;
    RECT 253.4 71.37 253.61 71.44 ;
    RECT 252.94 70.65 253.15 70.72 ;
    RECT 252.94 71.01 253.15 71.08 ;
    RECT 252.94 71.37 253.15 71.44 ;
    RECT 250.08 30.31 250.29 30.38 ;
    RECT 250.08 30.67 250.29 30.74 ;
    RECT 250.08 31.03 250.29 31.1 ;
    RECT 249.62 30.31 249.83 30.38 ;
    RECT 249.62 30.67 249.83 30.74 ;
    RECT 249.62 31.03 249.83 31.1 ;
    RECT 246.76 30.31 246.97 30.38 ;
    RECT 246.76 30.67 246.97 30.74 ;
    RECT 246.76 31.03 246.97 31.1 ;
    RECT 246.3 30.31 246.51 30.38 ;
    RECT 246.3 30.67 246.51 30.74 ;
    RECT 246.3 31.03 246.51 31.1 ;
    RECT 243.44 30.31 243.65 30.38 ;
    RECT 243.44 30.67 243.65 30.74 ;
    RECT 243.44 31.03 243.65 31.1 ;
    RECT 242.98 30.31 243.19 30.38 ;
    RECT 242.98 30.67 243.19 30.74 ;
    RECT 242.98 31.03 243.19 31.1 ;
    RECT 240.12 30.31 240.33 30.38 ;
    RECT 240.12 30.67 240.33 30.74 ;
    RECT 240.12 31.03 240.33 31.1 ;
    RECT 239.66 30.31 239.87 30.38 ;
    RECT 239.66 30.67 239.87 30.74 ;
    RECT 239.66 31.03 239.87 31.1 ;
    RECT 236.8 30.31 237.01 30.38 ;
    RECT 236.8 30.67 237.01 30.74 ;
    RECT 236.8 31.03 237.01 31.1 ;
    RECT 236.34 30.31 236.55 30.38 ;
    RECT 236.34 30.67 236.55 30.74 ;
    RECT 236.34 31.03 236.55 31.1 ;
    RECT 233.48 30.31 233.69 30.38 ;
    RECT 233.48 30.67 233.69 30.74 ;
    RECT 233.48 31.03 233.69 31.1 ;
    RECT 233.02 30.31 233.23 30.38 ;
    RECT 233.02 30.67 233.23 30.74 ;
    RECT 233.02 31.03 233.23 31.1 ;
    RECT 230.16 30.31 230.37 30.38 ;
    RECT 230.16 30.67 230.37 30.74 ;
    RECT 230.16 31.03 230.37 31.1 ;
    RECT 229.7 30.31 229.91 30.38 ;
    RECT 229.7 30.67 229.91 30.74 ;
    RECT 229.7 31.03 229.91 31.1 ;
    RECT 226.84 30.31 227.05 30.38 ;
    RECT 226.84 30.67 227.05 30.74 ;
    RECT 226.84 31.03 227.05 31.1 ;
    RECT 226.38 30.31 226.59 30.38 ;
    RECT 226.38 30.67 226.59 30.74 ;
    RECT 226.38 31.03 226.59 31.1 ;
    RECT 223.52 30.31 223.73 30.38 ;
    RECT 223.52 30.67 223.73 30.74 ;
    RECT 223.52 31.03 223.73 31.1 ;
    RECT 223.06 30.31 223.27 30.38 ;
    RECT 223.06 30.67 223.27 30.74 ;
    RECT 223.06 31.03 223.27 31.1 ;
    RECT 220.2 30.31 220.41 30.38 ;
    RECT 220.2 30.67 220.41 30.74 ;
    RECT 220.2 31.03 220.41 31.1 ;
    RECT 219.74 30.31 219.95 30.38 ;
    RECT 219.74 30.67 219.95 30.74 ;
    RECT 219.74 31.03 219.95 31.1 ;
    RECT 216.88 30.31 217.09 30.38 ;
    RECT 216.88 30.67 217.09 30.74 ;
    RECT 216.88 31.03 217.09 31.1 ;
    RECT 216.42 30.31 216.63 30.38 ;
    RECT 216.42 30.67 216.63 30.74 ;
    RECT 216.42 31.03 216.63 31.1 ;
    RECT 267.91 30.67 267.98 30.74 ;
    RECT 180.36 30.31 180.57 30.38 ;
    RECT 180.36 30.67 180.57 30.74 ;
    RECT 180.36 31.03 180.57 31.1 ;
    RECT 179.9 30.31 180.11 30.38 ;
    RECT 179.9 30.67 180.11 30.74 ;
    RECT 179.9 31.03 180.11 31.1 ;
    RECT 177.04 30.31 177.25 30.38 ;
    RECT 177.04 30.67 177.25 30.74 ;
    RECT 177.04 31.03 177.25 31.1 ;
    RECT 176.58 30.31 176.79 30.38 ;
    RECT 176.58 30.67 176.79 30.74 ;
    RECT 176.58 31.03 176.79 31.1 ;
    RECT 173.72 30.31 173.93 30.38 ;
    RECT 173.72 30.67 173.93 30.74 ;
    RECT 173.72 31.03 173.93 31.1 ;
    RECT 173.26 30.31 173.47 30.38 ;
    RECT 173.26 30.67 173.47 30.74 ;
    RECT 173.26 31.03 173.47 31.1 ;
    RECT 170.4 30.31 170.61 30.38 ;
    RECT 170.4 30.67 170.61 30.74 ;
    RECT 170.4 31.03 170.61 31.1 ;
    RECT 169.94 30.31 170.15 30.38 ;
    RECT 169.94 30.67 170.15 30.74 ;
    RECT 169.94 31.03 170.15 31.1 ;
    RECT 167.08 30.31 167.29 30.38 ;
    RECT 167.08 30.67 167.29 30.74 ;
    RECT 167.08 31.03 167.29 31.1 ;
    RECT 166.62 30.31 166.83 30.38 ;
    RECT 166.62 30.67 166.83 30.74 ;
    RECT 166.62 31.03 166.83 31.1 ;
    RECT 163.76 30.31 163.97 30.38 ;
    RECT 163.76 30.67 163.97 30.74 ;
    RECT 163.76 31.03 163.97 31.1 ;
    RECT 163.3 30.31 163.51 30.38 ;
    RECT 163.3 30.67 163.51 30.74 ;
    RECT 163.3 31.03 163.51 31.1 ;
    RECT 160.44 30.31 160.65 30.38 ;
    RECT 160.44 30.67 160.65 30.74 ;
    RECT 160.44 31.03 160.65 31.1 ;
    RECT 159.98 30.31 160.19 30.38 ;
    RECT 159.98 30.67 160.19 30.74 ;
    RECT 159.98 31.03 160.19 31.1 ;
    RECT 157.12 30.31 157.33 30.38 ;
    RECT 157.12 30.67 157.33 30.74 ;
    RECT 157.12 31.03 157.33 31.1 ;
    RECT 156.66 30.31 156.87 30.38 ;
    RECT 156.66 30.67 156.87 30.74 ;
    RECT 156.66 31.03 156.87 31.1 ;
    RECT 153.8 30.31 154.01 30.38 ;
    RECT 153.8 30.67 154.01 30.74 ;
    RECT 153.8 31.03 154.01 31.1 ;
    RECT 153.34 30.31 153.55 30.38 ;
    RECT 153.34 30.67 153.55 30.74 ;
    RECT 153.34 31.03 153.55 31.1 ;
    RECT 150.48 30.31 150.69 30.38 ;
    RECT 150.48 30.67 150.69 30.74 ;
    RECT 150.48 31.03 150.69 31.1 ;
    RECT 150.02 30.31 150.23 30.38 ;
    RECT 150.02 30.67 150.23 30.74 ;
    RECT 150.02 31.03 150.23 31.1 ;
    RECT 213.56 30.31 213.77 30.38 ;
    RECT 213.56 30.67 213.77 30.74 ;
    RECT 213.56 31.03 213.77 31.1 ;
    RECT 213.1 30.31 213.31 30.38 ;
    RECT 213.1 30.67 213.31 30.74 ;
    RECT 213.1 31.03 213.31 31.1 ;
    RECT 210.24 30.31 210.45 30.38 ;
    RECT 210.24 30.67 210.45 30.74 ;
    RECT 210.24 31.03 210.45 31.1 ;
    RECT 209.78 30.31 209.99 30.38 ;
    RECT 209.78 30.67 209.99 30.74 ;
    RECT 209.78 31.03 209.99 31.1 ;
    RECT 206.92 30.31 207.13 30.38 ;
    RECT 206.92 30.67 207.13 30.74 ;
    RECT 206.92 31.03 207.13 31.1 ;
    RECT 206.46 30.31 206.67 30.38 ;
    RECT 206.46 30.67 206.67 30.74 ;
    RECT 206.46 31.03 206.67 31.1 ;
    RECT 203.6 30.31 203.81 30.38 ;
    RECT 203.6 30.67 203.81 30.74 ;
    RECT 203.6 31.03 203.81 31.1 ;
    RECT 203.14 30.31 203.35 30.38 ;
    RECT 203.14 30.67 203.35 30.74 ;
    RECT 203.14 31.03 203.35 31.1 ;
    RECT 200.28 30.31 200.49 30.38 ;
    RECT 200.28 30.67 200.49 30.74 ;
    RECT 200.28 31.03 200.49 31.1 ;
    RECT 199.82 30.31 200.03 30.38 ;
    RECT 199.82 30.67 200.03 30.74 ;
    RECT 199.82 31.03 200.03 31.1 ;
    RECT 196.96 30.31 197.17 30.38 ;
    RECT 196.96 30.67 197.17 30.74 ;
    RECT 196.96 31.03 197.17 31.1 ;
    RECT 196.5 30.31 196.71 30.38 ;
    RECT 196.5 30.67 196.71 30.74 ;
    RECT 196.5 31.03 196.71 31.1 ;
    RECT 193.64 30.31 193.85 30.38 ;
    RECT 193.64 30.67 193.85 30.74 ;
    RECT 193.64 31.03 193.85 31.1 ;
    RECT 193.18 30.31 193.39 30.38 ;
    RECT 193.18 30.67 193.39 30.74 ;
    RECT 193.18 31.03 193.39 31.1 ;
    RECT 190.32 30.31 190.53 30.38 ;
    RECT 190.32 30.67 190.53 30.74 ;
    RECT 190.32 31.03 190.53 31.1 ;
    RECT 189.86 30.31 190.07 30.38 ;
    RECT 189.86 30.67 190.07 30.74 ;
    RECT 189.86 31.03 190.07 31.1 ;
    RECT 187.0 30.31 187.21 30.38 ;
    RECT 187.0 30.67 187.21 30.74 ;
    RECT 187.0 31.03 187.21 31.1 ;
    RECT 186.54 30.31 186.75 30.38 ;
    RECT 186.54 30.67 186.75 30.74 ;
    RECT 186.54 31.03 186.75 31.1 ;
    RECT 183.68 30.31 183.89 30.38 ;
    RECT 183.68 30.67 183.89 30.74 ;
    RECT 183.68 31.03 183.89 31.1 ;
    RECT 183.22 30.31 183.43 30.38 ;
    RECT 183.22 30.67 183.43 30.74 ;
    RECT 183.22 31.03 183.43 31.1 ;
    RECT 147.485 30.67 147.555 30.74 ;
    RECT 266.68 30.31 266.89 30.38 ;
    RECT 266.68 30.67 266.89 30.74 ;
    RECT 266.68 31.03 266.89 31.1 ;
    RECT 266.22 30.31 266.43 30.38 ;
    RECT 266.22 30.67 266.43 30.74 ;
    RECT 266.22 31.03 266.43 31.1 ;
    RECT 263.36 30.31 263.57 30.38 ;
    RECT 263.36 30.67 263.57 30.74 ;
    RECT 263.36 31.03 263.57 31.1 ;
    RECT 262.9 30.31 263.11 30.38 ;
    RECT 262.9 30.67 263.11 30.74 ;
    RECT 262.9 31.03 263.11 31.1 ;
    RECT 260.04 30.31 260.25 30.38 ;
    RECT 260.04 30.67 260.25 30.74 ;
    RECT 260.04 31.03 260.25 31.1 ;
    RECT 259.58 30.31 259.79 30.38 ;
    RECT 259.58 30.67 259.79 30.74 ;
    RECT 259.58 31.03 259.79 31.1 ;
    RECT 256.72 30.31 256.93 30.38 ;
    RECT 256.72 30.67 256.93 30.74 ;
    RECT 256.72 31.03 256.93 31.1 ;
    RECT 256.26 30.31 256.47 30.38 ;
    RECT 256.26 30.67 256.47 30.74 ;
    RECT 256.26 31.03 256.47 31.1 ;
    RECT 253.4 30.31 253.61 30.38 ;
    RECT 253.4 30.67 253.61 30.74 ;
    RECT 253.4 31.03 253.61 31.1 ;
    RECT 252.94 30.31 253.15 30.38 ;
    RECT 252.94 30.67 253.15 30.74 ;
    RECT 252.94 31.03 253.15 31.1 ;
    RECT 250.08 69.93 250.29 70.0 ;
    RECT 250.08 70.29 250.29 70.36 ;
    RECT 250.08 70.65 250.29 70.72 ;
    RECT 249.62 69.93 249.83 70.0 ;
    RECT 249.62 70.29 249.83 70.36 ;
    RECT 249.62 70.65 249.83 70.72 ;
    RECT 246.76 69.93 246.97 70.0 ;
    RECT 246.76 70.29 246.97 70.36 ;
    RECT 246.76 70.65 246.97 70.72 ;
    RECT 246.3 69.93 246.51 70.0 ;
    RECT 246.3 70.29 246.51 70.36 ;
    RECT 246.3 70.65 246.51 70.72 ;
    RECT 243.44 69.93 243.65 70.0 ;
    RECT 243.44 70.29 243.65 70.36 ;
    RECT 243.44 70.65 243.65 70.72 ;
    RECT 242.98 69.93 243.19 70.0 ;
    RECT 242.98 70.29 243.19 70.36 ;
    RECT 242.98 70.65 243.19 70.72 ;
    RECT 240.12 69.93 240.33 70.0 ;
    RECT 240.12 70.29 240.33 70.36 ;
    RECT 240.12 70.65 240.33 70.72 ;
    RECT 239.66 69.93 239.87 70.0 ;
    RECT 239.66 70.29 239.87 70.36 ;
    RECT 239.66 70.65 239.87 70.72 ;
    RECT 236.8 69.93 237.01 70.0 ;
    RECT 236.8 70.29 237.01 70.36 ;
    RECT 236.8 70.65 237.01 70.72 ;
    RECT 236.34 69.93 236.55 70.0 ;
    RECT 236.34 70.29 236.55 70.36 ;
    RECT 236.34 70.65 236.55 70.72 ;
    RECT 233.48 69.93 233.69 70.0 ;
    RECT 233.48 70.29 233.69 70.36 ;
    RECT 233.48 70.65 233.69 70.72 ;
    RECT 233.02 69.93 233.23 70.0 ;
    RECT 233.02 70.29 233.23 70.36 ;
    RECT 233.02 70.65 233.23 70.72 ;
    RECT 230.16 69.93 230.37 70.0 ;
    RECT 230.16 70.29 230.37 70.36 ;
    RECT 230.16 70.65 230.37 70.72 ;
    RECT 229.7 69.93 229.91 70.0 ;
    RECT 229.7 70.29 229.91 70.36 ;
    RECT 229.7 70.65 229.91 70.72 ;
    RECT 226.84 69.93 227.05 70.0 ;
    RECT 226.84 70.29 227.05 70.36 ;
    RECT 226.84 70.65 227.05 70.72 ;
    RECT 226.38 69.93 226.59 70.0 ;
    RECT 226.38 70.29 226.59 70.36 ;
    RECT 226.38 70.65 226.59 70.72 ;
    RECT 223.52 69.93 223.73 70.0 ;
    RECT 223.52 70.29 223.73 70.36 ;
    RECT 223.52 70.65 223.73 70.72 ;
    RECT 223.06 69.93 223.27 70.0 ;
    RECT 223.06 70.29 223.27 70.36 ;
    RECT 223.06 70.65 223.27 70.72 ;
    RECT 220.2 69.93 220.41 70.0 ;
    RECT 220.2 70.29 220.41 70.36 ;
    RECT 220.2 70.65 220.41 70.72 ;
    RECT 219.74 69.93 219.95 70.0 ;
    RECT 219.74 70.29 219.95 70.36 ;
    RECT 219.74 70.65 219.95 70.72 ;
    RECT 216.88 69.93 217.09 70.0 ;
    RECT 216.88 70.29 217.09 70.36 ;
    RECT 216.88 70.65 217.09 70.72 ;
    RECT 216.42 69.93 216.63 70.0 ;
    RECT 216.42 70.29 216.63 70.36 ;
    RECT 216.42 70.65 216.63 70.72 ;
    RECT 267.91 70.29 267.98 70.36 ;
    RECT 180.36 69.93 180.57 70.0 ;
    RECT 180.36 70.29 180.57 70.36 ;
    RECT 180.36 70.65 180.57 70.72 ;
    RECT 179.9 69.93 180.11 70.0 ;
    RECT 179.9 70.29 180.11 70.36 ;
    RECT 179.9 70.65 180.11 70.72 ;
    RECT 177.04 69.93 177.25 70.0 ;
    RECT 177.04 70.29 177.25 70.36 ;
    RECT 177.04 70.65 177.25 70.72 ;
    RECT 176.58 69.93 176.79 70.0 ;
    RECT 176.58 70.29 176.79 70.36 ;
    RECT 176.58 70.65 176.79 70.72 ;
    RECT 173.72 69.93 173.93 70.0 ;
    RECT 173.72 70.29 173.93 70.36 ;
    RECT 173.72 70.65 173.93 70.72 ;
    RECT 173.26 69.93 173.47 70.0 ;
    RECT 173.26 70.29 173.47 70.36 ;
    RECT 173.26 70.65 173.47 70.72 ;
    RECT 170.4 69.93 170.61 70.0 ;
    RECT 170.4 70.29 170.61 70.36 ;
    RECT 170.4 70.65 170.61 70.72 ;
    RECT 169.94 69.93 170.15 70.0 ;
    RECT 169.94 70.29 170.15 70.36 ;
    RECT 169.94 70.65 170.15 70.72 ;
    RECT 167.08 69.93 167.29 70.0 ;
    RECT 167.08 70.29 167.29 70.36 ;
    RECT 167.08 70.65 167.29 70.72 ;
    RECT 166.62 69.93 166.83 70.0 ;
    RECT 166.62 70.29 166.83 70.36 ;
    RECT 166.62 70.65 166.83 70.72 ;
    RECT 163.76 69.93 163.97 70.0 ;
    RECT 163.76 70.29 163.97 70.36 ;
    RECT 163.76 70.65 163.97 70.72 ;
    RECT 163.3 69.93 163.51 70.0 ;
    RECT 163.3 70.29 163.51 70.36 ;
    RECT 163.3 70.65 163.51 70.72 ;
    RECT 160.44 69.93 160.65 70.0 ;
    RECT 160.44 70.29 160.65 70.36 ;
    RECT 160.44 70.65 160.65 70.72 ;
    RECT 159.98 69.93 160.19 70.0 ;
    RECT 159.98 70.29 160.19 70.36 ;
    RECT 159.98 70.65 160.19 70.72 ;
    RECT 157.12 69.93 157.33 70.0 ;
    RECT 157.12 70.29 157.33 70.36 ;
    RECT 157.12 70.65 157.33 70.72 ;
    RECT 156.66 69.93 156.87 70.0 ;
    RECT 156.66 70.29 156.87 70.36 ;
    RECT 156.66 70.65 156.87 70.72 ;
    RECT 153.8 69.93 154.01 70.0 ;
    RECT 153.8 70.29 154.01 70.36 ;
    RECT 153.8 70.65 154.01 70.72 ;
    RECT 153.34 69.93 153.55 70.0 ;
    RECT 153.34 70.29 153.55 70.36 ;
    RECT 153.34 70.65 153.55 70.72 ;
    RECT 150.48 69.93 150.69 70.0 ;
    RECT 150.48 70.29 150.69 70.36 ;
    RECT 150.48 70.65 150.69 70.72 ;
    RECT 150.02 69.93 150.23 70.0 ;
    RECT 150.02 70.29 150.23 70.36 ;
    RECT 150.02 70.65 150.23 70.72 ;
    RECT 213.56 69.93 213.77 70.0 ;
    RECT 213.56 70.29 213.77 70.36 ;
    RECT 213.56 70.65 213.77 70.72 ;
    RECT 213.1 69.93 213.31 70.0 ;
    RECT 213.1 70.29 213.31 70.36 ;
    RECT 213.1 70.65 213.31 70.72 ;
    RECT 210.24 69.93 210.45 70.0 ;
    RECT 210.24 70.29 210.45 70.36 ;
    RECT 210.24 70.65 210.45 70.72 ;
    RECT 209.78 69.93 209.99 70.0 ;
    RECT 209.78 70.29 209.99 70.36 ;
    RECT 209.78 70.65 209.99 70.72 ;
    RECT 206.92 69.93 207.13 70.0 ;
    RECT 206.92 70.29 207.13 70.36 ;
    RECT 206.92 70.65 207.13 70.72 ;
    RECT 206.46 69.93 206.67 70.0 ;
    RECT 206.46 70.29 206.67 70.36 ;
    RECT 206.46 70.65 206.67 70.72 ;
    RECT 203.6 69.93 203.81 70.0 ;
    RECT 203.6 70.29 203.81 70.36 ;
    RECT 203.6 70.65 203.81 70.72 ;
    RECT 203.14 69.93 203.35 70.0 ;
    RECT 203.14 70.29 203.35 70.36 ;
    RECT 203.14 70.65 203.35 70.72 ;
    RECT 200.28 69.93 200.49 70.0 ;
    RECT 200.28 70.29 200.49 70.36 ;
    RECT 200.28 70.65 200.49 70.72 ;
    RECT 199.82 69.93 200.03 70.0 ;
    RECT 199.82 70.29 200.03 70.36 ;
    RECT 199.82 70.65 200.03 70.72 ;
    RECT 196.96 69.93 197.17 70.0 ;
    RECT 196.96 70.29 197.17 70.36 ;
    RECT 196.96 70.65 197.17 70.72 ;
    RECT 196.5 69.93 196.71 70.0 ;
    RECT 196.5 70.29 196.71 70.36 ;
    RECT 196.5 70.65 196.71 70.72 ;
    RECT 193.64 69.93 193.85 70.0 ;
    RECT 193.64 70.29 193.85 70.36 ;
    RECT 193.64 70.65 193.85 70.72 ;
    RECT 193.18 69.93 193.39 70.0 ;
    RECT 193.18 70.29 193.39 70.36 ;
    RECT 193.18 70.65 193.39 70.72 ;
    RECT 190.32 69.93 190.53 70.0 ;
    RECT 190.32 70.29 190.53 70.36 ;
    RECT 190.32 70.65 190.53 70.72 ;
    RECT 189.86 69.93 190.07 70.0 ;
    RECT 189.86 70.29 190.07 70.36 ;
    RECT 189.86 70.65 190.07 70.72 ;
    RECT 187.0 69.93 187.21 70.0 ;
    RECT 187.0 70.29 187.21 70.36 ;
    RECT 187.0 70.65 187.21 70.72 ;
    RECT 186.54 69.93 186.75 70.0 ;
    RECT 186.54 70.29 186.75 70.36 ;
    RECT 186.54 70.65 186.75 70.72 ;
    RECT 183.68 69.93 183.89 70.0 ;
    RECT 183.68 70.29 183.89 70.36 ;
    RECT 183.68 70.65 183.89 70.72 ;
    RECT 183.22 69.93 183.43 70.0 ;
    RECT 183.22 70.29 183.43 70.36 ;
    RECT 183.22 70.65 183.43 70.72 ;
    RECT 147.485 70.29 147.555 70.36 ;
    RECT 266.68 69.93 266.89 70.0 ;
    RECT 266.68 70.29 266.89 70.36 ;
    RECT 266.68 70.65 266.89 70.72 ;
    RECT 266.22 69.93 266.43 70.0 ;
    RECT 266.22 70.29 266.43 70.36 ;
    RECT 266.22 70.65 266.43 70.72 ;
    RECT 263.36 69.93 263.57 70.0 ;
    RECT 263.36 70.29 263.57 70.36 ;
    RECT 263.36 70.65 263.57 70.72 ;
    RECT 262.9 69.93 263.11 70.0 ;
    RECT 262.9 70.29 263.11 70.36 ;
    RECT 262.9 70.65 263.11 70.72 ;
    RECT 260.04 69.93 260.25 70.0 ;
    RECT 260.04 70.29 260.25 70.36 ;
    RECT 260.04 70.65 260.25 70.72 ;
    RECT 259.58 69.93 259.79 70.0 ;
    RECT 259.58 70.29 259.79 70.36 ;
    RECT 259.58 70.65 259.79 70.72 ;
    RECT 256.72 69.93 256.93 70.0 ;
    RECT 256.72 70.29 256.93 70.36 ;
    RECT 256.72 70.65 256.93 70.72 ;
    RECT 256.26 69.93 256.47 70.0 ;
    RECT 256.26 70.29 256.47 70.36 ;
    RECT 256.26 70.65 256.47 70.72 ;
    RECT 253.4 69.93 253.61 70.0 ;
    RECT 253.4 70.29 253.61 70.36 ;
    RECT 253.4 70.65 253.61 70.72 ;
    RECT 252.94 69.93 253.15 70.0 ;
    RECT 252.94 70.29 253.15 70.36 ;
    RECT 252.94 70.65 253.15 70.72 ;
    RECT 250.08 29.59 250.29 29.66 ;
    RECT 250.08 29.95 250.29 30.02 ;
    RECT 250.08 30.31 250.29 30.38 ;
    RECT 249.62 29.59 249.83 29.66 ;
    RECT 249.62 29.95 249.83 30.02 ;
    RECT 249.62 30.31 249.83 30.38 ;
    RECT 246.76 29.59 246.97 29.66 ;
    RECT 246.76 29.95 246.97 30.02 ;
    RECT 246.76 30.31 246.97 30.38 ;
    RECT 246.3 29.59 246.51 29.66 ;
    RECT 246.3 29.95 246.51 30.02 ;
    RECT 246.3 30.31 246.51 30.38 ;
    RECT 243.44 29.59 243.65 29.66 ;
    RECT 243.44 29.95 243.65 30.02 ;
    RECT 243.44 30.31 243.65 30.38 ;
    RECT 242.98 29.59 243.19 29.66 ;
    RECT 242.98 29.95 243.19 30.02 ;
    RECT 242.98 30.31 243.19 30.38 ;
    RECT 240.12 29.59 240.33 29.66 ;
    RECT 240.12 29.95 240.33 30.02 ;
    RECT 240.12 30.31 240.33 30.38 ;
    RECT 239.66 29.59 239.87 29.66 ;
    RECT 239.66 29.95 239.87 30.02 ;
    RECT 239.66 30.31 239.87 30.38 ;
    RECT 236.8 29.59 237.01 29.66 ;
    RECT 236.8 29.95 237.01 30.02 ;
    RECT 236.8 30.31 237.01 30.38 ;
    RECT 236.34 29.59 236.55 29.66 ;
    RECT 236.34 29.95 236.55 30.02 ;
    RECT 236.34 30.31 236.55 30.38 ;
    RECT 233.48 29.59 233.69 29.66 ;
    RECT 233.48 29.95 233.69 30.02 ;
    RECT 233.48 30.31 233.69 30.38 ;
    RECT 233.02 29.59 233.23 29.66 ;
    RECT 233.02 29.95 233.23 30.02 ;
    RECT 233.02 30.31 233.23 30.38 ;
    RECT 230.16 29.59 230.37 29.66 ;
    RECT 230.16 29.95 230.37 30.02 ;
    RECT 230.16 30.31 230.37 30.38 ;
    RECT 229.7 29.59 229.91 29.66 ;
    RECT 229.7 29.95 229.91 30.02 ;
    RECT 229.7 30.31 229.91 30.38 ;
    RECT 226.84 29.59 227.05 29.66 ;
    RECT 226.84 29.95 227.05 30.02 ;
    RECT 226.84 30.31 227.05 30.38 ;
    RECT 226.38 29.59 226.59 29.66 ;
    RECT 226.38 29.95 226.59 30.02 ;
    RECT 226.38 30.31 226.59 30.38 ;
    RECT 223.52 29.59 223.73 29.66 ;
    RECT 223.52 29.95 223.73 30.02 ;
    RECT 223.52 30.31 223.73 30.38 ;
    RECT 223.06 29.59 223.27 29.66 ;
    RECT 223.06 29.95 223.27 30.02 ;
    RECT 223.06 30.31 223.27 30.38 ;
    RECT 220.2 29.59 220.41 29.66 ;
    RECT 220.2 29.95 220.41 30.02 ;
    RECT 220.2 30.31 220.41 30.38 ;
    RECT 219.74 29.59 219.95 29.66 ;
    RECT 219.74 29.95 219.95 30.02 ;
    RECT 219.74 30.31 219.95 30.38 ;
    RECT 216.88 29.59 217.09 29.66 ;
    RECT 216.88 29.95 217.09 30.02 ;
    RECT 216.88 30.31 217.09 30.38 ;
    RECT 216.42 29.59 216.63 29.66 ;
    RECT 216.42 29.95 216.63 30.02 ;
    RECT 216.42 30.31 216.63 30.38 ;
    RECT 267.91 29.95 267.98 30.02 ;
    RECT 180.36 29.59 180.57 29.66 ;
    RECT 180.36 29.95 180.57 30.02 ;
    RECT 180.36 30.31 180.57 30.38 ;
    RECT 179.9 29.59 180.11 29.66 ;
    RECT 179.9 29.95 180.11 30.02 ;
    RECT 179.9 30.31 180.11 30.38 ;
    RECT 177.04 29.59 177.25 29.66 ;
    RECT 177.04 29.95 177.25 30.02 ;
    RECT 177.04 30.31 177.25 30.38 ;
    RECT 176.58 29.59 176.79 29.66 ;
    RECT 176.58 29.95 176.79 30.02 ;
    RECT 176.58 30.31 176.79 30.38 ;
    RECT 173.72 29.59 173.93 29.66 ;
    RECT 173.72 29.95 173.93 30.02 ;
    RECT 173.72 30.31 173.93 30.38 ;
    RECT 173.26 29.59 173.47 29.66 ;
    RECT 173.26 29.95 173.47 30.02 ;
    RECT 173.26 30.31 173.47 30.38 ;
    RECT 170.4 29.59 170.61 29.66 ;
    RECT 170.4 29.95 170.61 30.02 ;
    RECT 170.4 30.31 170.61 30.38 ;
    RECT 169.94 29.59 170.15 29.66 ;
    RECT 169.94 29.95 170.15 30.02 ;
    RECT 169.94 30.31 170.15 30.38 ;
    RECT 167.08 29.59 167.29 29.66 ;
    RECT 167.08 29.95 167.29 30.02 ;
    RECT 167.08 30.31 167.29 30.38 ;
    RECT 166.62 29.59 166.83 29.66 ;
    RECT 166.62 29.95 166.83 30.02 ;
    RECT 166.62 30.31 166.83 30.38 ;
    RECT 163.76 29.59 163.97 29.66 ;
    RECT 163.76 29.95 163.97 30.02 ;
    RECT 163.76 30.31 163.97 30.38 ;
    RECT 163.3 29.59 163.51 29.66 ;
    RECT 163.3 29.95 163.51 30.02 ;
    RECT 163.3 30.31 163.51 30.38 ;
    RECT 160.44 29.59 160.65 29.66 ;
    RECT 160.44 29.95 160.65 30.02 ;
    RECT 160.44 30.31 160.65 30.38 ;
    RECT 159.98 29.59 160.19 29.66 ;
    RECT 159.98 29.95 160.19 30.02 ;
    RECT 159.98 30.31 160.19 30.38 ;
    RECT 157.12 29.59 157.33 29.66 ;
    RECT 157.12 29.95 157.33 30.02 ;
    RECT 157.12 30.31 157.33 30.38 ;
    RECT 156.66 29.59 156.87 29.66 ;
    RECT 156.66 29.95 156.87 30.02 ;
    RECT 156.66 30.31 156.87 30.38 ;
    RECT 153.8 29.59 154.01 29.66 ;
    RECT 153.8 29.95 154.01 30.02 ;
    RECT 153.8 30.31 154.01 30.38 ;
    RECT 153.34 29.59 153.55 29.66 ;
    RECT 153.34 29.95 153.55 30.02 ;
    RECT 153.34 30.31 153.55 30.38 ;
    RECT 150.48 29.59 150.69 29.66 ;
    RECT 150.48 29.95 150.69 30.02 ;
    RECT 150.48 30.31 150.69 30.38 ;
    RECT 150.02 29.59 150.23 29.66 ;
    RECT 150.02 29.95 150.23 30.02 ;
    RECT 150.02 30.31 150.23 30.38 ;
    RECT 213.56 29.59 213.77 29.66 ;
    RECT 213.56 29.95 213.77 30.02 ;
    RECT 213.56 30.31 213.77 30.38 ;
    RECT 213.1 29.59 213.31 29.66 ;
    RECT 213.1 29.95 213.31 30.02 ;
    RECT 213.1 30.31 213.31 30.38 ;
    RECT 210.24 29.59 210.45 29.66 ;
    RECT 210.24 29.95 210.45 30.02 ;
    RECT 210.24 30.31 210.45 30.38 ;
    RECT 209.78 29.59 209.99 29.66 ;
    RECT 209.78 29.95 209.99 30.02 ;
    RECT 209.78 30.31 209.99 30.38 ;
    RECT 206.92 29.59 207.13 29.66 ;
    RECT 206.92 29.95 207.13 30.02 ;
    RECT 206.92 30.31 207.13 30.38 ;
    RECT 206.46 29.59 206.67 29.66 ;
    RECT 206.46 29.95 206.67 30.02 ;
    RECT 206.46 30.31 206.67 30.38 ;
    RECT 203.6 29.59 203.81 29.66 ;
    RECT 203.6 29.95 203.81 30.02 ;
    RECT 203.6 30.31 203.81 30.38 ;
    RECT 203.14 29.59 203.35 29.66 ;
    RECT 203.14 29.95 203.35 30.02 ;
    RECT 203.14 30.31 203.35 30.38 ;
    RECT 200.28 29.59 200.49 29.66 ;
    RECT 200.28 29.95 200.49 30.02 ;
    RECT 200.28 30.31 200.49 30.38 ;
    RECT 199.82 29.59 200.03 29.66 ;
    RECT 199.82 29.95 200.03 30.02 ;
    RECT 199.82 30.31 200.03 30.38 ;
    RECT 196.96 29.59 197.17 29.66 ;
    RECT 196.96 29.95 197.17 30.02 ;
    RECT 196.96 30.31 197.17 30.38 ;
    RECT 196.5 29.59 196.71 29.66 ;
    RECT 196.5 29.95 196.71 30.02 ;
    RECT 196.5 30.31 196.71 30.38 ;
    RECT 193.64 29.59 193.85 29.66 ;
    RECT 193.64 29.95 193.85 30.02 ;
    RECT 193.64 30.31 193.85 30.38 ;
    RECT 193.18 29.59 193.39 29.66 ;
    RECT 193.18 29.95 193.39 30.02 ;
    RECT 193.18 30.31 193.39 30.38 ;
    RECT 190.32 29.59 190.53 29.66 ;
    RECT 190.32 29.95 190.53 30.02 ;
    RECT 190.32 30.31 190.53 30.38 ;
    RECT 189.86 29.59 190.07 29.66 ;
    RECT 189.86 29.95 190.07 30.02 ;
    RECT 189.86 30.31 190.07 30.38 ;
    RECT 187.0 29.59 187.21 29.66 ;
    RECT 187.0 29.95 187.21 30.02 ;
    RECT 187.0 30.31 187.21 30.38 ;
    RECT 186.54 29.59 186.75 29.66 ;
    RECT 186.54 29.95 186.75 30.02 ;
    RECT 186.54 30.31 186.75 30.38 ;
    RECT 183.68 29.59 183.89 29.66 ;
    RECT 183.68 29.95 183.89 30.02 ;
    RECT 183.68 30.31 183.89 30.38 ;
    RECT 183.22 29.59 183.43 29.66 ;
    RECT 183.22 29.95 183.43 30.02 ;
    RECT 183.22 30.31 183.43 30.38 ;
    RECT 147.485 29.95 147.555 30.02 ;
    RECT 266.68 29.59 266.89 29.66 ;
    RECT 266.68 29.95 266.89 30.02 ;
    RECT 266.68 30.31 266.89 30.38 ;
    RECT 266.22 29.59 266.43 29.66 ;
    RECT 266.22 29.95 266.43 30.02 ;
    RECT 266.22 30.31 266.43 30.38 ;
    RECT 263.36 29.59 263.57 29.66 ;
    RECT 263.36 29.95 263.57 30.02 ;
    RECT 263.36 30.31 263.57 30.38 ;
    RECT 262.9 29.59 263.11 29.66 ;
    RECT 262.9 29.95 263.11 30.02 ;
    RECT 262.9 30.31 263.11 30.38 ;
    RECT 260.04 29.59 260.25 29.66 ;
    RECT 260.04 29.95 260.25 30.02 ;
    RECT 260.04 30.31 260.25 30.38 ;
    RECT 259.58 29.59 259.79 29.66 ;
    RECT 259.58 29.95 259.79 30.02 ;
    RECT 259.58 30.31 259.79 30.38 ;
    RECT 256.72 29.59 256.93 29.66 ;
    RECT 256.72 29.95 256.93 30.02 ;
    RECT 256.72 30.31 256.93 30.38 ;
    RECT 256.26 29.59 256.47 29.66 ;
    RECT 256.26 29.95 256.47 30.02 ;
    RECT 256.26 30.31 256.47 30.38 ;
    RECT 253.4 29.59 253.61 29.66 ;
    RECT 253.4 29.95 253.61 30.02 ;
    RECT 253.4 30.31 253.61 30.38 ;
    RECT 252.94 29.59 253.15 29.66 ;
    RECT 252.94 29.95 253.15 30.02 ;
    RECT 252.94 30.31 253.15 30.38 ;
    RECT 250.08 69.21 250.29 69.28 ;
    RECT 250.08 69.57 250.29 69.64 ;
    RECT 250.08 69.93 250.29 70.0 ;
    RECT 249.62 69.21 249.83 69.28 ;
    RECT 249.62 69.57 249.83 69.64 ;
    RECT 249.62 69.93 249.83 70.0 ;
    RECT 246.76 69.21 246.97 69.28 ;
    RECT 246.76 69.57 246.97 69.64 ;
    RECT 246.76 69.93 246.97 70.0 ;
    RECT 246.3 69.21 246.51 69.28 ;
    RECT 246.3 69.57 246.51 69.64 ;
    RECT 246.3 69.93 246.51 70.0 ;
    RECT 243.44 69.21 243.65 69.28 ;
    RECT 243.44 69.57 243.65 69.64 ;
    RECT 243.44 69.93 243.65 70.0 ;
    RECT 242.98 69.21 243.19 69.28 ;
    RECT 242.98 69.57 243.19 69.64 ;
    RECT 242.98 69.93 243.19 70.0 ;
    RECT 240.12 69.21 240.33 69.28 ;
    RECT 240.12 69.57 240.33 69.64 ;
    RECT 240.12 69.93 240.33 70.0 ;
    RECT 239.66 69.21 239.87 69.28 ;
    RECT 239.66 69.57 239.87 69.64 ;
    RECT 239.66 69.93 239.87 70.0 ;
    RECT 236.8 69.21 237.01 69.28 ;
    RECT 236.8 69.57 237.01 69.64 ;
    RECT 236.8 69.93 237.01 70.0 ;
    RECT 236.34 69.21 236.55 69.28 ;
    RECT 236.34 69.57 236.55 69.64 ;
    RECT 236.34 69.93 236.55 70.0 ;
    RECT 233.48 69.21 233.69 69.28 ;
    RECT 233.48 69.57 233.69 69.64 ;
    RECT 233.48 69.93 233.69 70.0 ;
    RECT 233.02 69.21 233.23 69.28 ;
    RECT 233.02 69.57 233.23 69.64 ;
    RECT 233.02 69.93 233.23 70.0 ;
    RECT 230.16 69.21 230.37 69.28 ;
    RECT 230.16 69.57 230.37 69.64 ;
    RECT 230.16 69.93 230.37 70.0 ;
    RECT 229.7 69.21 229.91 69.28 ;
    RECT 229.7 69.57 229.91 69.64 ;
    RECT 229.7 69.93 229.91 70.0 ;
    RECT 226.84 69.21 227.05 69.28 ;
    RECT 226.84 69.57 227.05 69.64 ;
    RECT 226.84 69.93 227.05 70.0 ;
    RECT 226.38 69.21 226.59 69.28 ;
    RECT 226.38 69.57 226.59 69.64 ;
    RECT 226.38 69.93 226.59 70.0 ;
    RECT 223.52 69.21 223.73 69.28 ;
    RECT 223.52 69.57 223.73 69.64 ;
    RECT 223.52 69.93 223.73 70.0 ;
    RECT 223.06 69.21 223.27 69.28 ;
    RECT 223.06 69.57 223.27 69.64 ;
    RECT 223.06 69.93 223.27 70.0 ;
    RECT 220.2 69.21 220.41 69.28 ;
    RECT 220.2 69.57 220.41 69.64 ;
    RECT 220.2 69.93 220.41 70.0 ;
    RECT 219.74 69.21 219.95 69.28 ;
    RECT 219.74 69.57 219.95 69.64 ;
    RECT 219.74 69.93 219.95 70.0 ;
    RECT 216.88 69.21 217.09 69.28 ;
    RECT 216.88 69.57 217.09 69.64 ;
    RECT 216.88 69.93 217.09 70.0 ;
    RECT 216.42 69.21 216.63 69.28 ;
    RECT 216.42 69.57 216.63 69.64 ;
    RECT 216.42 69.93 216.63 70.0 ;
    RECT 267.91 69.57 267.98 69.64 ;
    RECT 180.36 69.21 180.57 69.28 ;
    RECT 180.36 69.57 180.57 69.64 ;
    RECT 180.36 69.93 180.57 70.0 ;
    RECT 179.9 69.21 180.11 69.28 ;
    RECT 179.9 69.57 180.11 69.64 ;
    RECT 179.9 69.93 180.11 70.0 ;
    RECT 177.04 69.21 177.25 69.28 ;
    RECT 177.04 69.57 177.25 69.64 ;
    RECT 177.04 69.93 177.25 70.0 ;
    RECT 176.58 69.21 176.79 69.28 ;
    RECT 176.58 69.57 176.79 69.64 ;
    RECT 176.58 69.93 176.79 70.0 ;
    RECT 173.72 69.21 173.93 69.28 ;
    RECT 173.72 69.57 173.93 69.64 ;
    RECT 173.72 69.93 173.93 70.0 ;
    RECT 173.26 69.21 173.47 69.28 ;
    RECT 173.26 69.57 173.47 69.64 ;
    RECT 173.26 69.93 173.47 70.0 ;
    RECT 170.4 69.21 170.61 69.28 ;
    RECT 170.4 69.57 170.61 69.64 ;
    RECT 170.4 69.93 170.61 70.0 ;
    RECT 169.94 69.21 170.15 69.28 ;
    RECT 169.94 69.57 170.15 69.64 ;
    RECT 169.94 69.93 170.15 70.0 ;
    RECT 167.08 69.21 167.29 69.28 ;
    RECT 167.08 69.57 167.29 69.64 ;
    RECT 167.08 69.93 167.29 70.0 ;
    RECT 166.62 69.21 166.83 69.28 ;
    RECT 166.62 69.57 166.83 69.64 ;
    RECT 166.62 69.93 166.83 70.0 ;
    RECT 163.76 69.21 163.97 69.28 ;
    RECT 163.76 69.57 163.97 69.64 ;
    RECT 163.76 69.93 163.97 70.0 ;
    RECT 163.3 69.21 163.51 69.28 ;
    RECT 163.3 69.57 163.51 69.64 ;
    RECT 163.3 69.93 163.51 70.0 ;
    RECT 160.44 69.21 160.65 69.28 ;
    RECT 160.44 69.57 160.65 69.64 ;
    RECT 160.44 69.93 160.65 70.0 ;
    RECT 159.98 69.21 160.19 69.28 ;
    RECT 159.98 69.57 160.19 69.64 ;
    RECT 159.98 69.93 160.19 70.0 ;
    RECT 157.12 69.21 157.33 69.28 ;
    RECT 157.12 69.57 157.33 69.64 ;
    RECT 157.12 69.93 157.33 70.0 ;
    RECT 156.66 69.21 156.87 69.28 ;
    RECT 156.66 69.57 156.87 69.64 ;
    RECT 156.66 69.93 156.87 70.0 ;
    RECT 153.8 69.21 154.01 69.28 ;
    RECT 153.8 69.57 154.01 69.64 ;
    RECT 153.8 69.93 154.01 70.0 ;
    RECT 153.34 69.21 153.55 69.28 ;
    RECT 153.34 69.57 153.55 69.64 ;
    RECT 153.34 69.93 153.55 70.0 ;
    RECT 150.48 69.21 150.69 69.28 ;
    RECT 150.48 69.57 150.69 69.64 ;
    RECT 150.48 69.93 150.69 70.0 ;
    RECT 150.02 69.21 150.23 69.28 ;
    RECT 150.02 69.57 150.23 69.64 ;
    RECT 150.02 69.93 150.23 70.0 ;
    RECT 213.56 69.21 213.77 69.28 ;
    RECT 213.56 69.57 213.77 69.64 ;
    RECT 213.56 69.93 213.77 70.0 ;
    RECT 213.1 69.21 213.31 69.28 ;
    RECT 213.1 69.57 213.31 69.64 ;
    RECT 213.1 69.93 213.31 70.0 ;
    RECT 210.24 69.21 210.45 69.28 ;
    RECT 210.24 69.57 210.45 69.64 ;
    RECT 210.24 69.93 210.45 70.0 ;
    RECT 209.78 69.21 209.99 69.28 ;
    RECT 209.78 69.57 209.99 69.64 ;
    RECT 209.78 69.93 209.99 70.0 ;
    RECT 206.92 69.21 207.13 69.28 ;
    RECT 206.92 69.57 207.13 69.64 ;
    RECT 206.92 69.93 207.13 70.0 ;
    RECT 206.46 69.21 206.67 69.28 ;
    RECT 206.46 69.57 206.67 69.64 ;
    RECT 206.46 69.93 206.67 70.0 ;
    RECT 203.6 69.21 203.81 69.28 ;
    RECT 203.6 69.57 203.81 69.64 ;
    RECT 203.6 69.93 203.81 70.0 ;
    RECT 203.14 69.21 203.35 69.28 ;
    RECT 203.14 69.57 203.35 69.64 ;
    RECT 203.14 69.93 203.35 70.0 ;
    RECT 200.28 69.21 200.49 69.28 ;
    RECT 200.28 69.57 200.49 69.64 ;
    RECT 200.28 69.93 200.49 70.0 ;
    RECT 199.82 69.21 200.03 69.28 ;
    RECT 199.82 69.57 200.03 69.64 ;
    RECT 199.82 69.93 200.03 70.0 ;
    RECT 196.96 69.21 197.17 69.28 ;
    RECT 196.96 69.57 197.17 69.64 ;
    RECT 196.96 69.93 197.17 70.0 ;
    RECT 196.5 69.21 196.71 69.28 ;
    RECT 196.5 69.57 196.71 69.64 ;
    RECT 196.5 69.93 196.71 70.0 ;
    RECT 193.64 69.21 193.85 69.28 ;
    RECT 193.64 69.57 193.85 69.64 ;
    RECT 193.64 69.93 193.85 70.0 ;
    RECT 193.18 69.21 193.39 69.28 ;
    RECT 193.18 69.57 193.39 69.64 ;
    RECT 193.18 69.93 193.39 70.0 ;
    RECT 190.32 69.21 190.53 69.28 ;
    RECT 190.32 69.57 190.53 69.64 ;
    RECT 190.32 69.93 190.53 70.0 ;
    RECT 189.86 69.21 190.07 69.28 ;
    RECT 189.86 69.57 190.07 69.64 ;
    RECT 189.86 69.93 190.07 70.0 ;
    RECT 187.0 69.21 187.21 69.28 ;
    RECT 187.0 69.57 187.21 69.64 ;
    RECT 187.0 69.93 187.21 70.0 ;
    RECT 186.54 69.21 186.75 69.28 ;
    RECT 186.54 69.57 186.75 69.64 ;
    RECT 186.54 69.93 186.75 70.0 ;
    RECT 183.68 69.21 183.89 69.28 ;
    RECT 183.68 69.57 183.89 69.64 ;
    RECT 183.68 69.93 183.89 70.0 ;
    RECT 183.22 69.21 183.43 69.28 ;
    RECT 183.22 69.57 183.43 69.64 ;
    RECT 183.22 69.93 183.43 70.0 ;
    RECT 147.485 69.57 147.555 69.64 ;
    RECT 266.68 69.21 266.89 69.28 ;
    RECT 266.68 69.57 266.89 69.64 ;
    RECT 266.68 69.93 266.89 70.0 ;
    RECT 266.22 69.21 266.43 69.28 ;
    RECT 266.22 69.57 266.43 69.64 ;
    RECT 266.22 69.93 266.43 70.0 ;
    RECT 263.36 69.21 263.57 69.28 ;
    RECT 263.36 69.57 263.57 69.64 ;
    RECT 263.36 69.93 263.57 70.0 ;
    RECT 262.9 69.21 263.11 69.28 ;
    RECT 262.9 69.57 263.11 69.64 ;
    RECT 262.9 69.93 263.11 70.0 ;
    RECT 260.04 69.21 260.25 69.28 ;
    RECT 260.04 69.57 260.25 69.64 ;
    RECT 260.04 69.93 260.25 70.0 ;
    RECT 259.58 69.21 259.79 69.28 ;
    RECT 259.58 69.57 259.79 69.64 ;
    RECT 259.58 69.93 259.79 70.0 ;
    RECT 256.72 69.21 256.93 69.28 ;
    RECT 256.72 69.57 256.93 69.64 ;
    RECT 256.72 69.93 256.93 70.0 ;
    RECT 256.26 69.21 256.47 69.28 ;
    RECT 256.26 69.57 256.47 69.64 ;
    RECT 256.26 69.93 256.47 70.0 ;
    RECT 253.4 69.21 253.61 69.28 ;
    RECT 253.4 69.57 253.61 69.64 ;
    RECT 253.4 69.93 253.61 70.0 ;
    RECT 252.94 69.21 253.15 69.28 ;
    RECT 252.94 69.57 253.15 69.64 ;
    RECT 252.94 69.93 253.15 70.0 ;
    RECT 250.08 28.87 250.29 28.94 ;
    RECT 250.08 29.23 250.29 29.3 ;
    RECT 250.08 29.59 250.29 29.66 ;
    RECT 249.62 28.87 249.83 28.94 ;
    RECT 249.62 29.23 249.83 29.3 ;
    RECT 249.62 29.59 249.83 29.66 ;
    RECT 246.76 28.87 246.97 28.94 ;
    RECT 246.76 29.23 246.97 29.3 ;
    RECT 246.76 29.59 246.97 29.66 ;
    RECT 246.3 28.87 246.51 28.94 ;
    RECT 246.3 29.23 246.51 29.3 ;
    RECT 246.3 29.59 246.51 29.66 ;
    RECT 243.44 28.87 243.65 28.94 ;
    RECT 243.44 29.23 243.65 29.3 ;
    RECT 243.44 29.59 243.65 29.66 ;
    RECT 242.98 28.87 243.19 28.94 ;
    RECT 242.98 29.23 243.19 29.3 ;
    RECT 242.98 29.59 243.19 29.66 ;
    RECT 240.12 28.87 240.33 28.94 ;
    RECT 240.12 29.23 240.33 29.3 ;
    RECT 240.12 29.59 240.33 29.66 ;
    RECT 239.66 28.87 239.87 28.94 ;
    RECT 239.66 29.23 239.87 29.3 ;
    RECT 239.66 29.59 239.87 29.66 ;
    RECT 236.8 28.87 237.01 28.94 ;
    RECT 236.8 29.23 237.01 29.3 ;
    RECT 236.8 29.59 237.01 29.66 ;
    RECT 236.34 28.87 236.55 28.94 ;
    RECT 236.34 29.23 236.55 29.3 ;
    RECT 236.34 29.59 236.55 29.66 ;
    RECT 233.48 28.87 233.69 28.94 ;
    RECT 233.48 29.23 233.69 29.3 ;
    RECT 233.48 29.59 233.69 29.66 ;
    RECT 233.02 28.87 233.23 28.94 ;
    RECT 233.02 29.23 233.23 29.3 ;
    RECT 233.02 29.59 233.23 29.66 ;
    RECT 230.16 28.87 230.37 28.94 ;
    RECT 230.16 29.23 230.37 29.3 ;
    RECT 230.16 29.59 230.37 29.66 ;
    RECT 229.7 28.87 229.91 28.94 ;
    RECT 229.7 29.23 229.91 29.3 ;
    RECT 229.7 29.59 229.91 29.66 ;
    RECT 226.84 28.87 227.05 28.94 ;
    RECT 226.84 29.23 227.05 29.3 ;
    RECT 226.84 29.59 227.05 29.66 ;
    RECT 226.38 28.87 226.59 28.94 ;
    RECT 226.38 29.23 226.59 29.3 ;
    RECT 226.38 29.59 226.59 29.66 ;
    RECT 223.52 28.87 223.73 28.94 ;
    RECT 223.52 29.23 223.73 29.3 ;
    RECT 223.52 29.59 223.73 29.66 ;
    RECT 223.06 28.87 223.27 28.94 ;
    RECT 223.06 29.23 223.27 29.3 ;
    RECT 223.06 29.59 223.27 29.66 ;
    RECT 220.2 28.87 220.41 28.94 ;
    RECT 220.2 29.23 220.41 29.3 ;
    RECT 220.2 29.59 220.41 29.66 ;
    RECT 219.74 28.87 219.95 28.94 ;
    RECT 219.74 29.23 219.95 29.3 ;
    RECT 219.74 29.59 219.95 29.66 ;
    RECT 216.88 28.87 217.09 28.94 ;
    RECT 216.88 29.23 217.09 29.3 ;
    RECT 216.88 29.59 217.09 29.66 ;
    RECT 216.42 28.87 216.63 28.94 ;
    RECT 216.42 29.23 216.63 29.3 ;
    RECT 216.42 29.59 216.63 29.66 ;
    RECT 267.91 29.23 267.98 29.3 ;
    RECT 180.36 28.87 180.57 28.94 ;
    RECT 180.36 29.23 180.57 29.3 ;
    RECT 180.36 29.59 180.57 29.66 ;
    RECT 179.9 28.87 180.11 28.94 ;
    RECT 179.9 29.23 180.11 29.3 ;
    RECT 179.9 29.59 180.11 29.66 ;
    RECT 177.04 28.87 177.25 28.94 ;
    RECT 177.04 29.23 177.25 29.3 ;
    RECT 177.04 29.59 177.25 29.66 ;
    RECT 176.58 28.87 176.79 28.94 ;
    RECT 176.58 29.23 176.79 29.3 ;
    RECT 176.58 29.59 176.79 29.66 ;
    RECT 173.72 28.87 173.93 28.94 ;
    RECT 173.72 29.23 173.93 29.3 ;
    RECT 173.72 29.59 173.93 29.66 ;
    RECT 173.26 28.87 173.47 28.94 ;
    RECT 173.26 29.23 173.47 29.3 ;
    RECT 173.26 29.59 173.47 29.66 ;
    RECT 170.4 28.87 170.61 28.94 ;
    RECT 170.4 29.23 170.61 29.3 ;
    RECT 170.4 29.59 170.61 29.66 ;
    RECT 169.94 28.87 170.15 28.94 ;
    RECT 169.94 29.23 170.15 29.3 ;
    RECT 169.94 29.59 170.15 29.66 ;
    RECT 167.08 28.87 167.29 28.94 ;
    RECT 167.08 29.23 167.29 29.3 ;
    RECT 167.08 29.59 167.29 29.66 ;
    RECT 166.62 28.87 166.83 28.94 ;
    RECT 166.62 29.23 166.83 29.3 ;
    RECT 166.62 29.59 166.83 29.66 ;
    RECT 163.76 28.87 163.97 28.94 ;
    RECT 163.76 29.23 163.97 29.3 ;
    RECT 163.76 29.59 163.97 29.66 ;
    RECT 163.3 28.87 163.51 28.94 ;
    RECT 163.3 29.23 163.51 29.3 ;
    RECT 163.3 29.59 163.51 29.66 ;
    RECT 160.44 28.87 160.65 28.94 ;
    RECT 160.44 29.23 160.65 29.3 ;
    RECT 160.44 29.59 160.65 29.66 ;
    RECT 159.98 28.87 160.19 28.94 ;
    RECT 159.98 29.23 160.19 29.3 ;
    RECT 159.98 29.59 160.19 29.66 ;
    RECT 157.12 28.87 157.33 28.94 ;
    RECT 157.12 29.23 157.33 29.3 ;
    RECT 157.12 29.59 157.33 29.66 ;
    RECT 156.66 28.87 156.87 28.94 ;
    RECT 156.66 29.23 156.87 29.3 ;
    RECT 156.66 29.59 156.87 29.66 ;
    RECT 153.8 28.87 154.01 28.94 ;
    RECT 153.8 29.23 154.01 29.3 ;
    RECT 153.8 29.59 154.01 29.66 ;
    RECT 153.34 28.87 153.55 28.94 ;
    RECT 153.34 29.23 153.55 29.3 ;
    RECT 153.34 29.59 153.55 29.66 ;
    RECT 150.48 28.87 150.69 28.94 ;
    RECT 150.48 29.23 150.69 29.3 ;
    RECT 150.48 29.59 150.69 29.66 ;
    RECT 150.02 28.87 150.23 28.94 ;
    RECT 150.02 29.23 150.23 29.3 ;
    RECT 150.02 29.59 150.23 29.66 ;
    RECT 213.56 28.87 213.77 28.94 ;
    RECT 213.56 29.23 213.77 29.3 ;
    RECT 213.56 29.59 213.77 29.66 ;
    RECT 213.1 28.87 213.31 28.94 ;
    RECT 213.1 29.23 213.31 29.3 ;
    RECT 213.1 29.59 213.31 29.66 ;
    RECT 210.24 28.87 210.45 28.94 ;
    RECT 210.24 29.23 210.45 29.3 ;
    RECT 210.24 29.59 210.45 29.66 ;
    RECT 209.78 28.87 209.99 28.94 ;
    RECT 209.78 29.23 209.99 29.3 ;
    RECT 209.78 29.59 209.99 29.66 ;
    RECT 206.92 28.87 207.13 28.94 ;
    RECT 206.92 29.23 207.13 29.3 ;
    RECT 206.92 29.59 207.13 29.66 ;
    RECT 206.46 28.87 206.67 28.94 ;
    RECT 206.46 29.23 206.67 29.3 ;
    RECT 206.46 29.59 206.67 29.66 ;
    RECT 203.6 28.87 203.81 28.94 ;
    RECT 203.6 29.23 203.81 29.3 ;
    RECT 203.6 29.59 203.81 29.66 ;
    RECT 203.14 28.87 203.35 28.94 ;
    RECT 203.14 29.23 203.35 29.3 ;
    RECT 203.14 29.59 203.35 29.66 ;
    RECT 200.28 28.87 200.49 28.94 ;
    RECT 200.28 29.23 200.49 29.3 ;
    RECT 200.28 29.59 200.49 29.66 ;
    RECT 199.82 28.87 200.03 28.94 ;
    RECT 199.82 29.23 200.03 29.3 ;
    RECT 199.82 29.59 200.03 29.66 ;
    RECT 196.96 28.87 197.17 28.94 ;
    RECT 196.96 29.23 197.17 29.3 ;
    RECT 196.96 29.59 197.17 29.66 ;
    RECT 196.5 28.87 196.71 28.94 ;
    RECT 196.5 29.23 196.71 29.3 ;
    RECT 196.5 29.59 196.71 29.66 ;
    RECT 193.64 28.87 193.85 28.94 ;
    RECT 193.64 29.23 193.85 29.3 ;
    RECT 193.64 29.59 193.85 29.66 ;
    RECT 193.18 28.87 193.39 28.94 ;
    RECT 193.18 29.23 193.39 29.3 ;
    RECT 193.18 29.59 193.39 29.66 ;
    RECT 190.32 28.87 190.53 28.94 ;
    RECT 190.32 29.23 190.53 29.3 ;
    RECT 190.32 29.59 190.53 29.66 ;
    RECT 189.86 28.87 190.07 28.94 ;
    RECT 189.86 29.23 190.07 29.3 ;
    RECT 189.86 29.59 190.07 29.66 ;
    RECT 187.0 28.87 187.21 28.94 ;
    RECT 187.0 29.23 187.21 29.3 ;
    RECT 187.0 29.59 187.21 29.66 ;
    RECT 186.54 28.87 186.75 28.94 ;
    RECT 186.54 29.23 186.75 29.3 ;
    RECT 186.54 29.59 186.75 29.66 ;
    RECT 183.68 28.87 183.89 28.94 ;
    RECT 183.68 29.23 183.89 29.3 ;
    RECT 183.68 29.59 183.89 29.66 ;
    RECT 183.22 28.87 183.43 28.94 ;
    RECT 183.22 29.23 183.43 29.3 ;
    RECT 183.22 29.59 183.43 29.66 ;
    RECT 147.485 29.23 147.555 29.3 ;
    RECT 266.68 28.87 266.89 28.94 ;
    RECT 266.68 29.23 266.89 29.3 ;
    RECT 266.68 29.59 266.89 29.66 ;
    RECT 266.22 28.87 266.43 28.94 ;
    RECT 266.22 29.23 266.43 29.3 ;
    RECT 266.22 29.59 266.43 29.66 ;
    RECT 263.36 28.87 263.57 28.94 ;
    RECT 263.36 29.23 263.57 29.3 ;
    RECT 263.36 29.59 263.57 29.66 ;
    RECT 262.9 28.87 263.11 28.94 ;
    RECT 262.9 29.23 263.11 29.3 ;
    RECT 262.9 29.59 263.11 29.66 ;
    RECT 260.04 28.87 260.25 28.94 ;
    RECT 260.04 29.23 260.25 29.3 ;
    RECT 260.04 29.59 260.25 29.66 ;
    RECT 259.58 28.87 259.79 28.94 ;
    RECT 259.58 29.23 259.79 29.3 ;
    RECT 259.58 29.59 259.79 29.66 ;
    RECT 256.72 28.87 256.93 28.94 ;
    RECT 256.72 29.23 256.93 29.3 ;
    RECT 256.72 29.59 256.93 29.66 ;
    RECT 256.26 28.87 256.47 28.94 ;
    RECT 256.26 29.23 256.47 29.3 ;
    RECT 256.26 29.59 256.47 29.66 ;
    RECT 253.4 28.87 253.61 28.94 ;
    RECT 253.4 29.23 253.61 29.3 ;
    RECT 253.4 29.59 253.61 29.66 ;
    RECT 252.94 28.87 253.15 28.94 ;
    RECT 252.94 29.23 253.15 29.3 ;
    RECT 252.94 29.59 253.15 29.66 ;
    RECT 250.08 68.49 250.29 68.56 ;
    RECT 250.08 68.85 250.29 68.92 ;
    RECT 250.08 69.21 250.29 69.28 ;
    RECT 249.62 68.49 249.83 68.56 ;
    RECT 249.62 68.85 249.83 68.92 ;
    RECT 249.62 69.21 249.83 69.28 ;
    RECT 246.76 68.49 246.97 68.56 ;
    RECT 246.76 68.85 246.97 68.92 ;
    RECT 246.76 69.21 246.97 69.28 ;
    RECT 246.3 68.49 246.51 68.56 ;
    RECT 246.3 68.85 246.51 68.92 ;
    RECT 246.3 69.21 246.51 69.28 ;
    RECT 243.44 68.49 243.65 68.56 ;
    RECT 243.44 68.85 243.65 68.92 ;
    RECT 243.44 69.21 243.65 69.28 ;
    RECT 242.98 68.49 243.19 68.56 ;
    RECT 242.98 68.85 243.19 68.92 ;
    RECT 242.98 69.21 243.19 69.28 ;
    RECT 240.12 68.49 240.33 68.56 ;
    RECT 240.12 68.85 240.33 68.92 ;
    RECT 240.12 69.21 240.33 69.28 ;
    RECT 239.66 68.49 239.87 68.56 ;
    RECT 239.66 68.85 239.87 68.92 ;
    RECT 239.66 69.21 239.87 69.28 ;
    RECT 236.8 68.49 237.01 68.56 ;
    RECT 236.8 68.85 237.01 68.92 ;
    RECT 236.8 69.21 237.01 69.28 ;
    RECT 236.34 68.49 236.55 68.56 ;
    RECT 236.34 68.85 236.55 68.92 ;
    RECT 236.34 69.21 236.55 69.28 ;
    RECT 233.48 68.49 233.69 68.56 ;
    RECT 233.48 68.85 233.69 68.92 ;
    RECT 233.48 69.21 233.69 69.28 ;
    RECT 233.02 68.49 233.23 68.56 ;
    RECT 233.02 68.85 233.23 68.92 ;
    RECT 233.02 69.21 233.23 69.28 ;
    RECT 230.16 68.49 230.37 68.56 ;
    RECT 230.16 68.85 230.37 68.92 ;
    RECT 230.16 69.21 230.37 69.28 ;
    RECT 229.7 68.49 229.91 68.56 ;
    RECT 229.7 68.85 229.91 68.92 ;
    RECT 229.7 69.21 229.91 69.28 ;
    RECT 226.84 68.49 227.05 68.56 ;
    RECT 226.84 68.85 227.05 68.92 ;
    RECT 226.84 69.21 227.05 69.28 ;
    RECT 226.38 68.49 226.59 68.56 ;
    RECT 226.38 68.85 226.59 68.92 ;
    RECT 226.38 69.21 226.59 69.28 ;
    RECT 223.52 68.49 223.73 68.56 ;
    RECT 223.52 68.85 223.73 68.92 ;
    RECT 223.52 69.21 223.73 69.28 ;
    RECT 223.06 68.49 223.27 68.56 ;
    RECT 223.06 68.85 223.27 68.92 ;
    RECT 223.06 69.21 223.27 69.28 ;
    RECT 220.2 68.49 220.41 68.56 ;
    RECT 220.2 68.85 220.41 68.92 ;
    RECT 220.2 69.21 220.41 69.28 ;
    RECT 219.74 68.49 219.95 68.56 ;
    RECT 219.74 68.85 219.95 68.92 ;
    RECT 219.74 69.21 219.95 69.28 ;
    RECT 216.88 68.49 217.09 68.56 ;
    RECT 216.88 68.85 217.09 68.92 ;
    RECT 216.88 69.21 217.09 69.28 ;
    RECT 216.42 68.49 216.63 68.56 ;
    RECT 216.42 68.85 216.63 68.92 ;
    RECT 216.42 69.21 216.63 69.28 ;
    RECT 267.91 68.85 267.98 68.92 ;
    RECT 180.36 68.49 180.57 68.56 ;
    RECT 180.36 68.85 180.57 68.92 ;
    RECT 180.36 69.21 180.57 69.28 ;
    RECT 179.9 68.49 180.11 68.56 ;
    RECT 179.9 68.85 180.11 68.92 ;
    RECT 179.9 69.21 180.11 69.28 ;
    RECT 177.04 68.49 177.25 68.56 ;
    RECT 177.04 68.85 177.25 68.92 ;
    RECT 177.04 69.21 177.25 69.28 ;
    RECT 176.58 68.49 176.79 68.56 ;
    RECT 176.58 68.85 176.79 68.92 ;
    RECT 176.58 69.21 176.79 69.28 ;
    RECT 173.72 68.49 173.93 68.56 ;
    RECT 173.72 68.85 173.93 68.92 ;
    RECT 173.72 69.21 173.93 69.28 ;
    RECT 173.26 68.49 173.47 68.56 ;
    RECT 173.26 68.85 173.47 68.92 ;
    RECT 173.26 69.21 173.47 69.28 ;
    RECT 170.4 68.49 170.61 68.56 ;
    RECT 170.4 68.85 170.61 68.92 ;
    RECT 170.4 69.21 170.61 69.28 ;
    RECT 169.94 68.49 170.15 68.56 ;
    RECT 169.94 68.85 170.15 68.92 ;
    RECT 169.94 69.21 170.15 69.28 ;
    RECT 167.08 68.49 167.29 68.56 ;
    RECT 167.08 68.85 167.29 68.92 ;
    RECT 167.08 69.21 167.29 69.28 ;
    RECT 166.62 68.49 166.83 68.56 ;
    RECT 166.62 68.85 166.83 68.92 ;
    RECT 166.62 69.21 166.83 69.28 ;
    RECT 163.76 68.49 163.97 68.56 ;
    RECT 163.76 68.85 163.97 68.92 ;
    RECT 163.76 69.21 163.97 69.28 ;
    RECT 163.3 68.49 163.51 68.56 ;
    RECT 163.3 68.85 163.51 68.92 ;
    RECT 163.3 69.21 163.51 69.28 ;
    RECT 160.44 68.49 160.65 68.56 ;
    RECT 160.44 68.85 160.65 68.92 ;
    RECT 160.44 69.21 160.65 69.28 ;
    RECT 159.98 68.49 160.19 68.56 ;
    RECT 159.98 68.85 160.19 68.92 ;
    RECT 159.98 69.21 160.19 69.28 ;
    RECT 157.12 68.49 157.33 68.56 ;
    RECT 157.12 68.85 157.33 68.92 ;
    RECT 157.12 69.21 157.33 69.28 ;
    RECT 156.66 68.49 156.87 68.56 ;
    RECT 156.66 68.85 156.87 68.92 ;
    RECT 156.66 69.21 156.87 69.28 ;
    RECT 153.8 68.49 154.01 68.56 ;
    RECT 153.8 68.85 154.01 68.92 ;
    RECT 153.8 69.21 154.01 69.28 ;
    RECT 153.34 68.49 153.55 68.56 ;
    RECT 153.34 68.85 153.55 68.92 ;
    RECT 153.34 69.21 153.55 69.28 ;
    RECT 150.48 68.49 150.69 68.56 ;
    RECT 150.48 68.85 150.69 68.92 ;
    RECT 150.48 69.21 150.69 69.28 ;
    RECT 150.02 68.49 150.23 68.56 ;
    RECT 150.02 68.85 150.23 68.92 ;
    RECT 150.02 69.21 150.23 69.28 ;
    RECT 213.56 68.49 213.77 68.56 ;
    RECT 213.56 68.85 213.77 68.92 ;
    RECT 213.56 69.21 213.77 69.28 ;
    RECT 213.1 68.49 213.31 68.56 ;
    RECT 213.1 68.85 213.31 68.92 ;
    RECT 213.1 69.21 213.31 69.28 ;
    RECT 210.24 68.49 210.45 68.56 ;
    RECT 210.24 68.85 210.45 68.92 ;
    RECT 210.24 69.21 210.45 69.28 ;
    RECT 209.78 68.49 209.99 68.56 ;
    RECT 209.78 68.85 209.99 68.92 ;
    RECT 209.78 69.21 209.99 69.28 ;
    RECT 206.92 68.49 207.13 68.56 ;
    RECT 206.92 68.85 207.13 68.92 ;
    RECT 206.92 69.21 207.13 69.28 ;
    RECT 206.46 68.49 206.67 68.56 ;
    RECT 206.46 68.85 206.67 68.92 ;
    RECT 206.46 69.21 206.67 69.28 ;
    RECT 203.6 68.49 203.81 68.56 ;
    RECT 203.6 68.85 203.81 68.92 ;
    RECT 203.6 69.21 203.81 69.28 ;
    RECT 203.14 68.49 203.35 68.56 ;
    RECT 203.14 68.85 203.35 68.92 ;
    RECT 203.14 69.21 203.35 69.28 ;
    RECT 200.28 68.49 200.49 68.56 ;
    RECT 200.28 68.85 200.49 68.92 ;
    RECT 200.28 69.21 200.49 69.28 ;
    RECT 199.82 68.49 200.03 68.56 ;
    RECT 199.82 68.85 200.03 68.92 ;
    RECT 199.82 69.21 200.03 69.28 ;
    RECT 196.96 68.49 197.17 68.56 ;
    RECT 196.96 68.85 197.17 68.92 ;
    RECT 196.96 69.21 197.17 69.28 ;
    RECT 196.5 68.49 196.71 68.56 ;
    RECT 196.5 68.85 196.71 68.92 ;
    RECT 196.5 69.21 196.71 69.28 ;
    RECT 193.64 68.49 193.85 68.56 ;
    RECT 193.64 68.85 193.85 68.92 ;
    RECT 193.64 69.21 193.85 69.28 ;
    RECT 193.18 68.49 193.39 68.56 ;
    RECT 193.18 68.85 193.39 68.92 ;
    RECT 193.18 69.21 193.39 69.28 ;
    RECT 190.32 68.49 190.53 68.56 ;
    RECT 190.32 68.85 190.53 68.92 ;
    RECT 190.32 69.21 190.53 69.28 ;
    RECT 189.86 68.49 190.07 68.56 ;
    RECT 189.86 68.85 190.07 68.92 ;
    RECT 189.86 69.21 190.07 69.28 ;
    RECT 187.0 68.49 187.21 68.56 ;
    RECT 187.0 68.85 187.21 68.92 ;
    RECT 187.0 69.21 187.21 69.28 ;
    RECT 186.54 68.49 186.75 68.56 ;
    RECT 186.54 68.85 186.75 68.92 ;
    RECT 186.54 69.21 186.75 69.28 ;
    RECT 183.68 68.49 183.89 68.56 ;
    RECT 183.68 68.85 183.89 68.92 ;
    RECT 183.68 69.21 183.89 69.28 ;
    RECT 183.22 68.49 183.43 68.56 ;
    RECT 183.22 68.85 183.43 68.92 ;
    RECT 183.22 69.21 183.43 69.28 ;
    RECT 147.485 68.85 147.555 68.92 ;
    RECT 266.68 68.49 266.89 68.56 ;
    RECT 266.68 68.85 266.89 68.92 ;
    RECT 266.68 69.21 266.89 69.28 ;
    RECT 266.22 68.49 266.43 68.56 ;
    RECT 266.22 68.85 266.43 68.92 ;
    RECT 266.22 69.21 266.43 69.28 ;
    RECT 263.36 68.49 263.57 68.56 ;
    RECT 263.36 68.85 263.57 68.92 ;
    RECT 263.36 69.21 263.57 69.28 ;
    RECT 262.9 68.49 263.11 68.56 ;
    RECT 262.9 68.85 263.11 68.92 ;
    RECT 262.9 69.21 263.11 69.28 ;
    RECT 260.04 68.49 260.25 68.56 ;
    RECT 260.04 68.85 260.25 68.92 ;
    RECT 260.04 69.21 260.25 69.28 ;
    RECT 259.58 68.49 259.79 68.56 ;
    RECT 259.58 68.85 259.79 68.92 ;
    RECT 259.58 69.21 259.79 69.28 ;
    RECT 256.72 68.49 256.93 68.56 ;
    RECT 256.72 68.85 256.93 68.92 ;
    RECT 256.72 69.21 256.93 69.28 ;
    RECT 256.26 68.49 256.47 68.56 ;
    RECT 256.26 68.85 256.47 68.92 ;
    RECT 256.26 69.21 256.47 69.28 ;
    RECT 253.4 68.49 253.61 68.56 ;
    RECT 253.4 68.85 253.61 68.92 ;
    RECT 253.4 69.21 253.61 69.28 ;
    RECT 252.94 68.49 253.15 68.56 ;
    RECT 252.94 68.85 253.15 68.92 ;
    RECT 252.94 69.21 253.15 69.28 ;
    RECT 250.08 67.77 250.29 67.84 ;
    RECT 250.08 68.13 250.29 68.2 ;
    RECT 250.08 68.49 250.29 68.56 ;
    RECT 249.62 67.77 249.83 67.84 ;
    RECT 249.62 68.13 249.83 68.2 ;
    RECT 249.62 68.49 249.83 68.56 ;
    RECT 246.76 67.77 246.97 67.84 ;
    RECT 246.76 68.13 246.97 68.2 ;
    RECT 246.76 68.49 246.97 68.56 ;
    RECT 246.3 67.77 246.51 67.84 ;
    RECT 246.3 68.13 246.51 68.2 ;
    RECT 246.3 68.49 246.51 68.56 ;
    RECT 243.44 67.77 243.65 67.84 ;
    RECT 243.44 68.13 243.65 68.2 ;
    RECT 243.44 68.49 243.65 68.56 ;
    RECT 242.98 67.77 243.19 67.84 ;
    RECT 242.98 68.13 243.19 68.2 ;
    RECT 242.98 68.49 243.19 68.56 ;
    RECT 240.12 67.77 240.33 67.84 ;
    RECT 240.12 68.13 240.33 68.2 ;
    RECT 240.12 68.49 240.33 68.56 ;
    RECT 239.66 67.77 239.87 67.84 ;
    RECT 239.66 68.13 239.87 68.2 ;
    RECT 239.66 68.49 239.87 68.56 ;
    RECT 236.8 67.77 237.01 67.84 ;
    RECT 236.8 68.13 237.01 68.2 ;
    RECT 236.8 68.49 237.01 68.56 ;
    RECT 236.34 67.77 236.55 67.84 ;
    RECT 236.34 68.13 236.55 68.2 ;
    RECT 236.34 68.49 236.55 68.56 ;
    RECT 233.48 67.77 233.69 67.84 ;
    RECT 233.48 68.13 233.69 68.2 ;
    RECT 233.48 68.49 233.69 68.56 ;
    RECT 233.02 67.77 233.23 67.84 ;
    RECT 233.02 68.13 233.23 68.2 ;
    RECT 233.02 68.49 233.23 68.56 ;
    RECT 230.16 67.77 230.37 67.84 ;
    RECT 230.16 68.13 230.37 68.2 ;
    RECT 230.16 68.49 230.37 68.56 ;
    RECT 229.7 67.77 229.91 67.84 ;
    RECT 229.7 68.13 229.91 68.2 ;
    RECT 229.7 68.49 229.91 68.56 ;
    RECT 226.84 67.77 227.05 67.84 ;
    RECT 226.84 68.13 227.05 68.2 ;
    RECT 226.84 68.49 227.05 68.56 ;
    RECT 226.38 67.77 226.59 67.84 ;
    RECT 226.38 68.13 226.59 68.2 ;
    RECT 226.38 68.49 226.59 68.56 ;
    RECT 223.52 67.77 223.73 67.84 ;
    RECT 223.52 68.13 223.73 68.2 ;
    RECT 223.52 68.49 223.73 68.56 ;
    RECT 223.06 67.77 223.27 67.84 ;
    RECT 223.06 68.13 223.27 68.2 ;
    RECT 223.06 68.49 223.27 68.56 ;
    RECT 220.2 67.77 220.41 67.84 ;
    RECT 220.2 68.13 220.41 68.2 ;
    RECT 220.2 68.49 220.41 68.56 ;
    RECT 219.74 67.77 219.95 67.84 ;
    RECT 219.74 68.13 219.95 68.2 ;
    RECT 219.74 68.49 219.95 68.56 ;
    RECT 216.88 67.77 217.09 67.84 ;
    RECT 216.88 68.13 217.09 68.2 ;
    RECT 216.88 68.49 217.09 68.56 ;
    RECT 216.42 67.77 216.63 67.84 ;
    RECT 216.42 68.13 216.63 68.2 ;
    RECT 216.42 68.49 216.63 68.56 ;
    RECT 267.91 68.13 267.98 68.2 ;
    RECT 180.36 67.77 180.57 67.84 ;
    RECT 180.36 68.13 180.57 68.2 ;
    RECT 180.36 68.49 180.57 68.56 ;
    RECT 179.9 67.77 180.11 67.84 ;
    RECT 179.9 68.13 180.11 68.2 ;
    RECT 179.9 68.49 180.11 68.56 ;
    RECT 177.04 67.77 177.25 67.84 ;
    RECT 177.04 68.13 177.25 68.2 ;
    RECT 177.04 68.49 177.25 68.56 ;
    RECT 176.58 67.77 176.79 67.84 ;
    RECT 176.58 68.13 176.79 68.2 ;
    RECT 176.58 68.49 176.79 68.56 ;
    RECT 173.72 67.77 173.93 67.84 ;
    RECT 173.72 68.13 173.93 68.2 ;
    RECT 173.72 68.49 173.93 68.56 ;
    RECT 173.26 67.77 173.47 67.84 ;
    RECT 173.26 68.13 173.47 68.2 ;
    RECT 173.26 68.49 173.47 68.56 ;
    RECT 170.4 67.77 170.61 67.84 ;
    RECT 170.4 68.13 170.61 68.2 ;
    RECT 170.4 68.49 170.61 68.56 ;
    RECT 169.94 67.77 170.15 67.84 ;
    RECT 169.94 68.13 170.15 68.2 ;
    RECT 169.94 68.49 170.15 68.56 ;
    RECT 167.08 67.77 167.29 67.84 ;
    RECT 167.08 68.13 167.29 68.2 ;
    RECT 167.08 68.49 167.29 68.56 ;
    RECT 166.62 67.77 166.83 67.84 ;
    RECT 166.62 68.13 166.83 68.2 ;
    RECT 166.62 68.49 166.83 68.56 ;
    RECT 163.76 67.77 163.97 67.84 ;
    RECT 163.76 68.13 163.97 68.2 ;
    RECT 163.76 68.49 163.97 68.56 ;
    RECT 163.3 67.77 163.51 67.84 ;
    RECT 163.3 68.13 163.51 68.2 ;
    RECT 163.3 68.49 163.51 68.56 ;
    RECT 160.44 67.77 160.65 67.84 ;
    RECT 160.44 68.13 160.65 68.2 ;
    RECT 160.44 68.49 160.65 68.56 ;
    RECT 159.98 67.77 160.19 67.84 ;
    RECT 159.98 68.13 160.19 68.2 ;
    RECT 159.98 68.49 160.19 68.56 ;
    RECT 157.12 67.77 157.33 67.84 ;
    RECT 157.12 68.13 157.33 68.2 ;
    RECT 157.12 68.49 157.33 68.56 ;
    RECT 156.66 67.77 156.87 67.84 ;
    RECT 156.66 68.13 156.87 68.2 ;
    RECT 156.66 68.49 156.87 68.56 ;
    RECT 153.8 67.77 154.01 67.84 ;
    RECT 153.8 68.13 154.01 68.2 ;
    RECT 153.8 68.49 154.01 68.56 ;
    RECT 153.34 67.77 153.55 67.84 ;
    RECT 153.34 68.13 153.55 68.2 ;
    RECT 153.34 68.49 153.55 68.56 ;
    RECT 150.48 67.77 150.69 67.84 ;
    RECT 150.48 68.13 150.69 68.2 ;
    RECT 150.48 68.49 150.69 68.56 ;
    RECT 150.02 67.77 150.23 67.84 ;
    RECT 150.02 68.13 150.23 68.2 ;
    RECT 150.02 68.49 150.23 68.56 ;
    RECT 213.56 67.77 213.77 67.84 ;
    RECT 213.56 68.13 213.77 68.2 ;
    RECT 213.56 68.49 213.77 68.56 ;
    RECT 213.1 67.77 213.31 67.84 ;
    RECT 213.1 68.13 213.31 68.2 ;
    RECT 213.1 68.49 213.31 68.56 ;
    RECT 210.24 67.77 210.45 67.84 ;
    RECT 210.24 68.13 210.45 68.2 ;
    RECT 210.24 68.49 210.45 68.56 ;
    RECT 209.78 67.77 209.99 67.84 ;
    RECT 209.78 68.13 209.99 68.2 ;
    RECT 209.78 68.49 209.99 68.56 ;
    RECT 206.92 67.77 207.13 67.84 ;
    RECT 206.92 68.13 207.13 68.2 ;
    RECT 206.92 68.49 207.13 68.56 ;
    RECT 206.46 67.77 206.67 67.84 ;
    RECT 206.46 68.13 206.67 68.2 ;
    RECT 206.46 68.49 206.67 68.56 ;
    RECT 203.6 67.77 203.81 67.84 ;
    RECT 203.6 68.13 203.81 68.2 ;
    RECT 203.6 68.49 203.81 68.56 ;
    RECT 203.14 67.77 203.35 67.84 ;
    RECT 203.14 68.13 203.35 68.2 ;
    RECT 203.14 68.49 203.35 68.56 ;
    RECT 200.28 67.77 200.49 67.84 ;
    RECT 200.28 68.13 200.49 68.2 ;
    RECT 200.28 68.49 200.49 68.56 ;
    RECT 199.82 67.77 200.03 67.84 ;
    RECT 199.82 68.13 200.03 68.2 ;
    RECT 199.82 68.49 200.03 68.56 ;
    RECT 196.96 67.77 197.17 67.84 ;
    RECT 196.96 68.13 197.17 68.2 ;
    RECT 196.96 68.49 197.17 68.56 ;
    RECT 196.5 67.77 196.71 67.84 ;
    RECT 196.5 68.13 196.71 68.2 ;
    RECT 196.5 68.49 196.71 68.56 ;
    RECT 193.64 67.77 193.85 67.84 ;
    RECT 193.64 68.13 193.85 68.2 ;
    RECT 193.64 68.49 193.85 68.56 ;
    RECT 193.18 67.77 193.39 67.84 ;
    RECT 193.18 68.13 193.39 68.2 ;
    RECT 193.18 68.49 193.39 68.56 ;
    RECT 190.32 67.77 190.53 67.84 ;
    RECT 190.32 68.13 190.53 68.2 ;
    RECT 190.32 68.49 190.53 68.56 ;
    RECT 189.86 67.77 190.07 67.84 ;
    RECT 189.86 68.13 190.07 68.2 ;
    RECT 189.86 68.49 190.07 68.56 ;
    RECT 187.0 67.77 187.21 67.84 ;
    RECT 187.0 68.13 187.21 68.2 ;
    RECT 187.0 68.49 187.21 68.56 ;
    RECT 186.54 67.77 186.75 67.84 ;
    RECT 186.54 68.13 186.75 68.2 ;
    RECT 186.54 68.49 186.75 68.56 ;
    RECT 183.68 67.77 183.89 67.84 ;
    RECT 183.68 68.13 183.89 68.2 ;
    RECT 183.68 68.49 183.89 68.56 ;
    RECT 183.22 67.77 183.43 67.84 ;
    RECT 183.22 68.13 183.43 68.2 ;
    RECT 183.22 68.49 183.43 68.56 ;
    RECT 147.485 68.13 147.555 68.2 ;
    RECT 266.68 67.77 266.89 67.84 ;
    RECT 266.68 68.13 266.89 68.2 ;
    RECT 266.68 68.49 266.89 68.56 ;
    RECT 266.22 67.77 266.43 67.84 ;
    RECT 266.22 68.13 266.43 68.2 ;
    RECT 266.22 68.49 266.43 68.56 ;
    RECT 263.36 67.77 263.57 67.84 ;
    RECT 263.36 68.13 263.57 68.2 ;
    RECT 263.36 68.49 263.57 68.56 ;
    RECT 262.9 67.77 263.11 67.84 ;
    RECT 262.9 68.13 263.11 68.2 ;
    RECT 262.9 68.49 263.11 68.56 ;
    RECT 260.04 67.77 260.25 67.84 ;
    RECT 260.04 68.13 260.25 68.2 ;
    RECT 260.04 68.49 260.25 68.56 ;
    RECT 259.58 67.77 259.79 67.84 ;
    RECT 259.58 68.13 259.79 68.2 ;
    RECT 259.58 68.49 259.79 68.56 ;
    RECT 256.72 67.77 256.93 67.84 ;
    RECT 256.72 68.13 256.93 68.2 ;
    RECT 256.72 68.49 256.93 68.56 ;
    RECT 256.26 67.77 256.47 67.84 ;
    RECT 256.26 68.13 256.47 68.2 ;
    RECT 256.26 68.49 256.47 68.56 ;
    RECT 253.4 67.77 253.61 67.84 ;
    RECT 253.4 68.13 253.61 68.2 ;
    RECT 253.4 68.49 253.61 68.56 ;
    RECT 252.94 67.77 253.15 67.84 ;
    RECT 252.94 68.13 253.15 68.2 ;
    RECT 252.94 68.49 253.15 68.56 ;
    RECT 250.08 67.05 250.29 67.12 ;
    RECT 250.08 67.41 250.29 67.48 ;
    RECT 250.08 67.77 250.29 67.84 ;
    RECT 249.62 67.05 249.83 67.12 ;
    RECT 249.62 67.41 249.83 67.48 ;
    RECT 249.62 67.77 249.83 67.84 ;
    RECT 246.76 67.05 246.97 67.12 ;
    RECT 246.76 67.41 246.97 67.48 ;
    RECT 246.76 67.77 246.97 67.84 ;
    RECT 246.3 67.05 246.51 67.12 ;
    RECT 246.3 67.41 246.51 67.48 ;
    RECT 246.3 67.77 246.51 67.84 ;
    RECT 243.44 67.05 243.65 67.12 ;
    RECT 243.44 67.41 243.65 67.48 ;
    RECT 243.44 67.77 243.65 67.84 ;
    RECT 242.98 67.05 243.19 67.12 ;
    RECT 242.98 67.41 243.19 67.48 ;
    RECT 242.98 67.77 243.19 67.84 ;
    RECT 240.12 67.05 240.33 67.12 ;
    RECT 240.12 67.41 240.33 67.48 ;
    RECT 240.12 67.77 240.33 67.84 ;
    RECT 239.66 67.05 239.87 67.12 ;
    RECT 239.66 67.41 239.87 67.48 ;
    RECT 239.66 67.77 239.87 67.84 ;
    RECT 236.8 67.05 237.01 67.12 ;
    RECT 236.8 67.41 237.01 67.48 ;
    RECT 236.8 67.77 237.01 67.84 ;
    RECT 236.34 67.05 236.55 67.12 ;
    RECT 236.34 67.41 236.55 67.48 ;
    RECT 236.34 67.77 236.55 67.84 ;
    RECT 233.48 67.05 233.69 67.12 ;
    RECT 233.48 67.41 233.69 67.48 ;
    RECT 233.48 67.77 233.69 67.84 ;
    RECT 233.02 67.05 233.23 67.12 ;
    RECT 233.02 67.41 233.23 67.48 ;
    RECT 233.02 67.77 233.23 67.84 ;
    RECT 230.16 67.05 230.37 67.12 ;
    RECT 230.16 67.41 230.37 67.48 ;
    RECT 230.16 67.77 230.37 67.84 ;
    RECT 229.7 67.05 229.91 67.12 ;
    RECT 229.7 67.41 229.91 67.48 ;
    RECT 229.7 67.77 229.91 67.84 ;
    RECT 226.84 67.05 227.05 67.12 ;
    RECT 226.84 67.41 227.05 67.48 ;
    RECT 226.84 67.77 227.05 67.84 ;
    RECT 226.38 67.05 226.59 67.12 ;
    RECT 226.38 67.41 226.59 67.48 ;
    RECT 226.38 67.77 226.59 67.84 ;
    RECT 223.52 67.05 223.73 67.12 ;
    RECT 223.52 67.41 223.73 67.48 ;
    RECT 223.52 67.77 223.73 67.84 ;
    RECT 223.06 67.05 223.27 67.12 ;
    RECT 223.06 67.41 223.27 67.48 ;
    RECT 223.06 67.77 223.27 67.84 ;
    RECT 220.2 67.05 220.41 67.12 ;
    RECT 220.2 67.41 220.41 67.48 ;
    RECT 220.2 67.77 220.41 67.84 ;
    RECT 219.74 67.05 219.95 67.12 ;
    RECT 219.74 67.41 219.95 67.48 ;
    RECT 219.74 67.77 219.95 67.84 ;
    RECT 216.88 67.05 217.09 67.12 ;
    RECT 216.88 67.41 217.09 67.48 ;
    RECT 216.88 67.77 217.09 67.84 ;
    RECT 216.42 67.05 216.63 67.12 ;
    RECT 216.42 67.41 216.63 67.48 ;
    RECT 216.42 67.77 216.63 67.84 ;
    RECT 267.91 67.41 267.98 67.48 ;
    RECT 180.36 67.05 180.57 67.12 ;
    RECT 180.36 67.41 180.57 67.48 ;
    RECT 180.36 67.77 180.57 67.84 ;
    RECT 179.9 67.05 180.11 67.12 ;
    RECT 179.9 67.41 180.11 67.48 ;
    RECT 179.9 67.77 180.11 67.84 ;
    RECT 177.04 67.05 177.25 67.12 ;
    RECT 177.04 67.41 177.25 67.48 ;
    RECT 177.04 67.77 177.25 67.84 ;
    RECT 176.58 67.05 176.79 67.12 ;
    RECT 176.58 67.41 176.79 67.48 ;
    RECT 176.58 67.77 176.79 67.84 ;
    RECT 173.72 67.05 173.93 67.12 ;
    RECT 173.72 67.41 173.93 67.48 ;
    RECT 173.72 67.77 173.93 67.84 ;
    RECT 173.26 67.05 173.47 67.12 ;
    RECT 173.26 67.41 173.47 67.48 ;
    RECT 173.26 67.77 173.47 67.84 ;
    RECT 170.4 67.05 170.61 67.12 ;
    RECT 170.4 67.41 170.61 67.48 ;
    RECT 170.4 67.77 170.61 67.84 ;
    RECT 169.94 67.05 170.15 67.12 ;
    RECT 169.94 67.41 170.15 67.48 ;
    RECT 169.94 67.77 170.15 67.84 ;
    RECT 167.08 67.05 167.29 67.12 ;
    RECT 167.08 67.41 167.29 67.48 ;
    RECT 167.08 67.77 167.29 67.84 ;
    RECT 166.62 67.05 166.83 67.12 ;
    RECT 166.62 67.41 166.83 67.48 ;
    RECT 166.62 67.77 166.83 67.84 ;
    RECT 163.76 67.05 163.97 67.12 ;
    RECT 163.76 67.41 163.97 67.48 ;
    RECT 163.76 67.77 163.97 67.84 ;
    RECT 163.3 67.05 163.51 67.12 ;
    RECT 163.3 67.41 163.51 67.48 ;
    RECT 163.3 67.77 163.51 67.84 ;
    RECT 160.44 67.05 160.65 67.12 ;
    RECT 160.44 67.41 160.65 67.48 ;
    RECT 160.44 67.77 160.65 67.84 ;
    RECT 159.98 67.05 160.19 67.12 ;
    RECT 159.98 67.41 160.19 67.48 ;
    RECT 159.98 67.77 160.19 67.84 ;
    RECT 157.12 67.05 157.33 67.12 ;
    RECT 157.12 67.41 157.33 67.48 ;
    RECT 157.12 67.77 157.33 67.84 ;
    RECT 156.66 67.05 156.87 67.12 ;
    RECT 156.66 67.41 156.87 67.48 ;
    RECT 156.66 67.77 156.87 67.84 ;
    RECT 153.8 67.05 154.01 67.12 ;
    RECT 153.8 67.41 154.01 67.48 ;
    RECT 153.8 67.77 154.01 67.84 ;
    RECT 153.34 67.05 153.55 67.12 ;
    RECT 153.34 67.41 153.55 67.48 ;
    RECT 153.34 67.77 153.55 67.84 ;
    RECT 150.48 67.05 150.69 67.12 ;
    RECT 150.48 67.41 150.69 67.48 ;
    RECT 150.48 67.77 150.69 67.84 ;
    RECT 150.02 67.05 150.23 67.12 ;
    RECT 150.02 67.41 150.23 67.48 ;
    RECT 150.02 67.77 150.23 67.84 ;
    RECT 213.56 67.05 213.77 67.12 ;
    RECT 213.56 67.41 213.77 67.48 ;
    RECT 213.56 67.77 213.77 67.84 ;
    RECT 213.1 67.05 213.31 67.12 ;
    RECT 213.1 67.41 213.31 67.48 ;
    RECT 213.1 67.77 213.31 67.84 ;
    RECT 210.24 67.05 210.45 67.12 ;
    RECT 210.24 67.41 210.45 67.48 ;
    RECT 210.24 67.77 210.45 67.84 ;
    RECT 209.78 67.05 209.99 67.12 ;
    RECT 209.78 67.41 209.99 67.48 ;
    RECT 209.78 67.77 209.99 67.84 ;
    RECT 206.92 67.05 207.13 67.12 ;
    RECT 206.92 67.41 207.13 67.48 ;
    RECT 206.92 67.77 207.13 67.84 ;
    RECT 206.46 67.05 206.67 67.12 ;
    RECT 206.46 67.41 206.67 67.48 ;
    RECT 206.46 67.77 206.67 67.84 ;
    RECT 203.6 67.05 203.81 67.12 ;
    RECT 203.6 67.41 203.81 67.48 ;
    RECT 203.6 67.77 203.81 67.84 ;
    RECT 203.14 67.05 203.35 67.12 ;
    RECT 203.14 67.41 203.35 67.48 ;
    RECT 203.14 67.77 203.35 67.84 ;
    RECT 200.28 67.05 200.49 67.12 ;
    RECT 200.28 67.41 200.49 67.48 ;
    RECT 200.28 67.77 200.49 67.84 ;
    RECT 199.82 67.05 200.03 67.12 ;
    RECT 199.82 67.41 200.03 67.48 ;
    RECT 199.82 67.77 200.03 67.84 ;
    RECT 196.96 67.05 197.17 67.12 ;
    RECT 196.96 67.41 197.17 67.48 ;
    RECT 196.96 67.77 197.17 67.84 ;
    RECT 196.5 67.05 196.71 67.12 ;
    RECT 196.5 67.41 196.71 67.48 ;
    RECT 196.5 67.77 196.71 67.84 ;
    RECT 193.64 67.05 193.85 67.12 ;
    RECT 193.64 67.41 193.85 67.48 ;
    RECT 193.64 67.77 193.85 67.84 ;
    RECT 193.18 67.05 193.39 67.12 ;
    RECT 193.18 67.41 193.39 67.48 ;
    RECT 193.18 67.77 193.39 67.84 ;
    RECT 190.32 67.05 190.53 67.12 ;
    RECT 190.32 67.41 190.53 67.48 ;
    RECT 190.32 67.77 190.53 67.84 ;
    RECT 189.86 67.05 190.07 67.12 ;
    RECT 189.86 67.41 190.07 67.48 ;
    RECT 189.86 67.77 190.07 67.84 ;
    RECT 187.0 67.05 187.21 67.12 ;
    RECT 187.0 67.41 187.21 67.48 ;
    RECT 187.0 67.77 187.21 67.84 ;
    RECT 186.54 67.05 186.75 67.12 ;
    RECT 186.54 67.41 186.75 67.48 ;
    RECT 186.54 67.77 186.75 67.84 ;
    RECT 183.68 67.05 183.89 67.12 ;
    RECT 183.68 67.41 183.89 67.48 ;
    RECT 183.68 67.77 183.89 67.84 ;
    RECT 183.22 67.05 183.43 67.12 ;
    RECT 183.22 67.41 183.43 67.48 ;
    RECT 183.22 67.77 183.43 67.84 ;
    RECT 147.485 67.41 147.555 67.48 ;
    RECT 266.68 67.05 266.89 67.12 ;
    RECT 266.68 67.41 266.89 67.48 ;
    RECT 266.68 67.77 266.89 67.84 ;
    RECT 266.22 67.05 266.43 67.12 ;
    RECT 266.22 67.41 266.43 67.48 ;
    RECT 266.22 67.77 266.43 67.84 ;
    RECT 263.36 67.05 263.57 67.12 ;
    RECT 263.36 67.41 263.57 67.48 ;
    RECT 263.36 67.77 263.57 67.84 ;
    RECT 262.9 67.05 263.11 67.12 ;
    RECT 262.9 67.41 263.11 67.48 ;
    RECT 262.9 67.77 263.11 67.84 ;
    RECT 260.04 67.05 260.25 67.12 ;
    RECT 260.04 67.41 260.25 67.48 ;
    RECT 260.04 67.77 260.25 67.84 ;
    RECT 259.58 67.05 259.79 67.12 ;
    RECT 259.58 67.41 259.79 67.48 ;
    RECT 259.58 67.77 259.79 67.84 ;
    RECT 256.72 67.05 256.93 67.12 ;
    RECT 256.72 67.41 256.93 67.48 ;
    RECT 256.72 67.77 256.93 67.84 ;
    RECT 256.26 67.05 256.47 67.12 ;
    RECT 256.26 67.41 256.47 67.48 ;
    RECT 256.26 67.77 256.47 67.84 ;
    RECT 253.4 67.05 253.61 67.12 ;
    RECT 253.4 67.41 253.61 67.48 ;
    RECT 253.4 67.77 253.61 67.84 ;
    RECT 252.94 67.05 253.15 67.12 ;
    RECT 252.94 67.41 253.15 67.48 ;
    RECT 252.94 67.77 253.15 67.84 ;
    RECT 250.08 66.33 250.29 66.4 ;
    RECT 250.08 66.69 250.29 66.76 ;
    RECT 250.08 67.05 250.29 67.12 ;
    RECT 249.62 66.33 249.83 66.4 ;
    RECT 249.62 66.69 249.83 66.76 ;
    RECT 249.62 67.05 249.83 67.12 ;
    RECT 246.76 66.33 246.97 66.4 ;
    RECT 246.76 66.69 246.97 66.76 ;
    RECT 246.76 67.05 246.97 67.12 ;
    RECT 246.3 66.33 246.51 66.4 ;
    RECT 246.3 66.69 246.51 66.76 ;
    RECT 246.3 67.05 246.51 67.12 ;
    RECT 243.44 66.33 243.65 66.4 ;
    RECT 243.44 66.69 243.65 66.76 ;
    RECT 243.44 67.05 243.65 67.12 ;
    RECT 242.98 66.33 243.19 66.4 ;
    RECT 242.98 66.69 243.19 66.76 ;
    RECT 242.98 67.05 243.19 67.12 ;
    RECT 240.12 66.33 240.33 66.4 ;
    RECT 240.12 66.69 240.33 66.76 ;
    RECT 240.12 67.05 240.33 67.12 ;
    RECT 239.66 66.33 239.87 66.4 ;
    RECT 239.66 66.69 239.87 66.76 ;
    RECT 239.66 67.05 239.87 67.12 ;
    RECT 236.8 66.33 237.01 66.4 ;
    RECT 236.8 66.69 237.01 66.76 ;
    RECT 236.8 67.05 237.01 67.12 ;
    RECT 236.34 66.33 236.55 66.4 ;
    RECT 236.34 66.69 236.55 66.76 ;
    RECT 236.34 67.05 236.55 67.12 ;
    RECT 233.48 66.33 233.69 66.4 ;
    RECT 233.48 66.69 233.69 66.76 ;
    RECT 233.48 67.05 233.69 67.12 ;
    RECT 233.02 66.33 233.23 66.4 ;
    RECT 233.02 66.69 233.23 66.76 ;
    RECT 233.02 67.05 233.23 67.12 ;
    RECT 230.16 66.33 230.37 66.4 ;
    RECT 230.16 66.69 230.37 66.76 ;
    RECT 230.16 67.05 230.37 67.12 ;
    RECT 229.7 66.33 229.91 66.4 ;
    RECT 229.7 66.69 229.91 66.76 ;
    RECT 229.7 67.05 229.91 67.12 ;
    RECT 226.84 66.33 227.05 66.4 ;
    RECT 226.84 66.69 227.05 66.76 ;
    RECT 226.84 67.05 227.05 67.12 ;
    RECT 226.38 66.33 226.59 66.4 ;
    RECT 226.38 66.69 226.59 66.76 ;
    RECT 226.38 67.05 226.59 67.12 ;
    RECT 223.52 66.33 223.73 66.4 ;
    RECT 223.52 66.69 223.73 66.76 ;
    RECT 223.52 67.05 223.73 67.12 ;
    RECT 223.06 66.33 223.27 66.4 ;
    RECT 223.06 66.69 223.27 66.76 ;
    RECT 223.06 67.05 223.27 67.12 ;
    RECT 220.2 66.33 220.41 66.4 ;
    RECT 220.2 66.69 220.41 66.76 ;
    RECT 220.2 67.05 220.41 67.12 ;
    RECT 219.74 66.33 219.95 66.4 ;
    RECT 219.74 66.69 219.95 66.76 ;
    RECT 219.74 67.05 219.95 67.12 ;
    RECT 216.88 66.33 217.09 66.4 ;
    RECT 216.88 66.69 217.09 66.76 ;
    RECT 216.88 67.05 217.09 67.12 ;
    RECT 216.42 66.33 216.63 66.4 ;
    RECT 216.42 66.69 216.63 66.76 ;
    RECT 216.42 67.05 216.63 67.12 ;
    RECT 267.91 66.69 267.98 66.76 ;
    RECT 180.36 66.33 180.57 66.4 ;
    RECT 180.36 66.69 180.57 66.76 ;
    RECT 180.36 67.05 180.57 67.12 ;
    RECT 179.9 66.33 180.11 66.4 ;
    RECT 179.9 66.69 180.11 66.76 ;
    RECT 179.9 67.05 180.11 67.12 ;
    RECT 177.04 66.33 177.25 66.4 ;
    RECT 177.04 66.69 177.25 66.76 ;
    RECT 177.04 67.05 177.25 67.12 ;
    RECT 176.58 66.33 176.79 66.4 ;
    RECT 176.58 66.69 176.79 66.76 ;
    RECT 176.58 67.05 176.79 67.12 ;
    RECT 173.72 66.33 173.93 66.4 ;
    RECT 173.72 66.69 173.93 66.76 ;
    RECT 173.72 67.05 173.93 67.12 ;
    RECT 173.26 66.33 173.47 66.4 ;
    RECT 173.26 66.69 173.47 66.76 ;
    RECT 173.26 67.05 173.47 67.12 ;
    RECT 170.4 66.33 170.61 66.4 ;
    RECT 170.4 66.69 170.61 66.76 ;
    RECT 170.4 67.05 170.61 67.12 ;
    RECT 169.94 66.33 170.15 66.4 ;
    RECT 169.94 66.69 170.15 66.76 ;
    RECT 169.94 67.05 170.15 67.12 ;
    RECT 167.08 66.33 167.29 66.4 ;
    RECT 167.08 66.69 167.29 66.76 ;
    RECT 167.08 67.05 167.29 67.12 ;
    RECT 166.62 66.33 166.83 66.4 ;
    RECT 166.62 66.69 166.83 66.76 ;
    RECT 166.62 67.05 166.83 67.12 ;
    RECT 163.76 66.33 163.97 66.4 ;
    RECT 163.76 66.69 163.97 66.76 ;
    RECT 163.76 67.05 163.97 67.12 ;
    RECT 163.3 66.33 163.51 66.4 ;
    RECT 163.3 66.69 163.51 66.76 ;
    RECT 163.3 67.05 163.51 67.12 ;
    RECT 160.44 66.33 160.65 66.4 ;
    RECT 160.44 66.69 160.65 66.76 ;
    RECT 160.44 67.05 160.65 67.12 ;
    RECT 159.98 66.33 160.19 66.4 ;
    RECT 159.98 66.69 160.19 66.76 ;
    RECT 159.98 67.05 160.19 67.12 ;
    RECT 157.12 66.33 157.33 66.4 ;
    RECT 157.12 66.69 157.33 66.76 ;
    RECT 157.12 67.05 157.33 67.12 ;
    RECT 156.66 66.33 156.87 66.4 ;
    RECT 156.66 66.69 156.87 66.76 ;
    RECT 156.66 67.05 156.87 67.12 ;
    RECT 153.8 66.33 154.01 66.4 ;
    RECT 153.8 66.69 154.01 66.76 ;
    RECT 153.8 67.05 154.01 67.12 ;
    RECT 153.34 66.33 153.55 66.4 ;
    RECT 153.34 66.69 153.55 66.76 ;
    RECT 153.34 67.05 153.55 67.12 ;
    RECT 150.48 66.33 150.69 66.4 ;
    RECT 150.48 66.69 150.69 66.76 ;
    RECT 150.48 67.05 150.69 67.12 ;
    RECT 150.02 66.33 150.23 66.4 ;
    RECT 150.02 66.69 150.23 66.76 ;
    RECT 150.02 67.05 150.23 67.12 ;
    RECT 213.56 66.33 213.77 66.4 ;
    RECT 213.56 66.69 213.77 66.76 ;
    RECT 213.56 67.05 213.77 67.12 ;
    RECT 213.1 66.33 213.31 66.4 ;
    RECT 213.1 66.69 213.31 66.76 ;
    RECT 213.1 67.05 213.31 67.12 ;
    RECT 210.24 66.33 210.45 66.4 ;
    RECT 210.24 66.69 210.45 66.76 ;
    RECT 210.24 67.05 210.45 67.12 ;
    RECT 209.78 66.33 209.99 66.4 ;
    RECT 209.78 66.69 209.99 66.76 ;
    RECT 209.78 67.05 209.99 67.12 ;
    RECT 206.92 66.33 207.13 66.4 ;
    RECT 206.92 66.69 207.13 66.76 ;
    RECT 206.92 67.05 207.13 67.12 ;
    RECT 206.46 66.33 206.67 66.4 ;
    RECT 206.46 66.69 206.67 66.76 ;
    RECT 206.46 67.05 206.67 67.12 ;
    RECT 203.6 66.33 203.81 66.4 ;
    RECT 203.6 66.69 203.81 66.76 ;
    RECT 203.6 67.05 203.81 67.12 ;
    RECT 203.14 66.33 203.35 66.4 ;
    RECT 203.14 66.69 203.35 66.76 ;
    RECT 203.14 67.05 203.35 67.12 ;
    RECT 200.28 66.33 200.49 66.4 ;
    RECT 200.28 66.69 200.49 66.76 ;
    RECT 200.28 67.05 200.49 67.12 ;
    RECT 199.82 66.33 200.03 66.4 ;
    RECT 199.82 66.69 200.03 66.76 ;
    RECT 199.82 67.05 200.03 67.12 ;
    RECT 196.96 66.33 197.17 66.4 ;
    RECT 196.96 66.69 197.17 66.76 ;
    RECT 196.96 67.05 197.17 67.12 ;
    RECT 196.5 66.33 196.71 66.4 ;
    RECT 196.5 66.69 196.71 66.76 ;
    RECT 196.5 67.05 196.71 67.12 ;
    RECT 193.64 66.33 193.85 66.4 ;
    RECT 193.64 66.69 193.85 66.76 ;
    RECT 193.64 67.05 193.85 67.12 ;
    RECT 193.18 66.33 193.39 66.4 ;
    RECT 193.18 66.69 193.39 66.76 ;
    RECT 193.18 67.05 193.39 67.12 ;
    RECT 190.32 66.33 190.53 66.4 ;
    RECT 190.32 66.69 190.53 66.76 ;
    RECT 190.32 67.05 190.53 67.12 ;
    RECT 189.86 66.33 190.07 66.4 ;
    RECT 189.86 66.69 190.07 66.76 ;
    RECT 189.86 67.05 190.07 67.12 ;
    RECT 187.0 66.33 187.21 66.4 ;
    RECT 187.0 66.69 187.21 66.76 ;
    RECT 187.0 67.05 187.21 67.12 ;
    RECT 186.54 66.33 186.75 66.4 ;
    RECT 186.54 66.69 186.75 66.76 ;
    RECT 186.54 67.05 186.75 67.12 ;
    RECT 183.68 66.33 183.89 66.4 ;
    RECT 183.68 66.69 183.89 66.76 ;
    RECT 183.68 67.05 183.89 67.12 ;
    RECT 183.22 66.33 183.43 66.4 ;
    RECT 183.22 66.69 183.43 66.76 ;
    RECT 183.22 67.05 183.43 67.12 ;
    RECT 147.485 66.69 147.555 66.76 ;
    RECT 266.68 66.33 266.89 66.4 ;
    RECT 266.68 66.69 266.89 66.76 ;
    RECT 266.68 67.05 266.89 67.12 ;
    RECT 266.22 66.33 266.43 66.4 ;
    RECT 266.22 66.69 266.43 66.76 ;
    RECT 266.22 67.05 266.43 67.12 ;
    RECT 263.36 66.33 263.57 66.4 ;
    RECT 263.36 66.69 263.57 66.76 ;
    RECT 263.36 67.05 263.57 67.12 ;
    RECT 262.9 66.33 263.11 66.4 ;
    RECT 262.9 66.69 263.11 66.76 ;
    RECT 262.9 67.05 263.11 67.12 ;
    RECT 260.04 66.33 260.25 66.4 ;
    RECT 260.04 66.69 260.25 66.76 ;
    RECT 260.04 67.05 260.25 67.12 ;
    RECT 259.58 66.33 259.79 66.4 ;
    RECT 259.58 66.69 259.79 66.76 ;
    RECT 259.58 67.05 259.79 67.12 ;
    RECT 256.72 66.33 256.93 66.4 ;
    RECT 256.72 66.69 256.93 66.76 ;
    RECT 256.72 67.05 256.93 67.12 ;
    RECT 256.26 66.33 256.47 66.4 ;
    RECT 256.26 66.69 256.47 66.76 ;
    RECT 256.26 67.05 256.47 67.12 ;
    RECT 253.4 66.33 253.61 66.4 ;
    RECT 253.4 66.69 253.61 66.76 ;
    RECT 253.4 67.05 253.61 67.12 ;
    RECT 252.94 66.33 253.15 66.4 ;
    RECT 252.94 66.69 253.15 66.76 ;
    RECT 252.94 67.05 253.15 67.12 ;
    RECT 250.08 65.61 250.29 65.68 ;
    RECT 250.08 65.97 250.29 66.04 ;
    RECT 250.08 66.33 250.29 66.4 ;
    RECT 249.62 65.61 249.83 65.68 ;
    RECT 249.62 65.97 249.83 66.04 ;
    RECT 249.62 66.33 249.83 66.4 ;
    RECT 246.76 65.61 246.97 65.68 ;
    RECT 246.76 65.97 246.97 66.04 ;
    RECT 246.76 66.33 246.97 66.4 ;
    RECT 246.3 65.61 246.51 65.68 ;
    RECT 246.3 65.97 246.51 66.04 ;
    RECT 246.3 66.33 246.51 66.4 ;
    RECT 243.44 65.61 243.65 65.68 ;
    RECT 243.44 65.97 243.65 66.04 ;
    RECT 243.44 66.33 243.65 66.4 ;
    RECT 242.98 65.61 243.19 65.68 ;
    RECT 242.98 65.97 243.19 66.04 ;
    RECT 242.98 66.33 243.19 66.4 ;
    RECT 240.12 65.61 240.33 65.68 ;
    RECT 240.12 65.97 240.33 66.04 ;
    RECT 240.12 66.33 240.33 66.4 ;
    RECT 239.66 65.61 239.87 65.68 ;
    RECT 239.66 65.97 239.87 66.04 ;
    RECT 239.66 66.33 239.87 66.4 ;
    RECT 236.8 65.61 237.01 65.68 ;
    RECT 236.8 65.97 237.01 66.04 ;
    RECT 236.8 66.33 237.01 66.4 ;
    RECT 236.34 65.61 236.55 65.68 ;
    RECT 236.34 65.97 236.55 66.04 ;
    RECT 236.34 66.33 236.55 66.4 ;
    RECT 233.48 65.61 233.69 65.68 ;
    RECT 233.48 65.97 233.69 66.04 ;
    RECT 233.48 66.33 233.69 66.4 ;
    RECT 233.02 65.61 233.23 65.68 ;
    RECT 233.02 65.97 233.23 66.04 ;
    RECT 233.02 66.33 233.23 66.4 ;
    RECT 230.16 65.61 230.37 65.68 ;
    RECT 230.16 65.97 230.37 66.04 ;
    RECT 230.16 66.33 230.37 66.4 ;
    RECT 229.7 65.61 229.91 65.68 ;
    RECT 229.7 65.97 229.91 66.04 ;
    RECT 229.7 66.33 229.91 66.4 ;
    RECT 226.84 65.61 227.05 65.68 ;
    RECT 226.84 65.97 227.05 66.04 ;
    RECT 226.84 66.33 227.05 66.4 ;
    RECT 226.38 65.61 226.59 65.68 ;
    RECT 226.38 65.97 226.59 66.04 ;
    RECT 226.38 66.33 226.59 66.4 ;
    RECT 223.52 65.61 223.73 65.68 ;
    RECT 223.52 65.97 223.73 66.04 ;
    RECT 223.52 66.33 223.73 66.4 ;
    RECT 223.06 65.61 223.27 65.68 ;
    RECT 223.06 65.97 223.27 66.04 ;
    RECT 223.06 66.33 223.27 66.4 ;
    RECT 220.2 65.61 220.41 65.68 ;
    RECT 220.2 65.97 220.41 66.04 ;
    RECT 220.2 66.33 220.41 66.4 ;
    RECT 219.74 65.61 219.95 65.68 ;
    RECT 219.74 65.97 219.95 66.04 ;
    RECT 219.74 66.33 219.95 66.4 ;
    RECT 216.88 65.61 217.09 65.68 ;
    RECT 216.88 65.97 217.09 66.04 ;
    RECT 216.88 66.33 217.09 66.4 ;
    RECT 216.42 65.61 216.63 65.68 ;
    RECT 216.42 65.97 216.63 66.04 ;
    RECT 216.42 66.33 216.63 66.4 ;
    RECT 267.91 65.97 267.98 66.04 ;
    RECT 180.36 65.61 180.57 65.68 ;
    RECT 180.36 65.97 180.57 66.04 ;
    RECT 180.36 66.33 180.57 66.4 ;
    RECT 179.9 65.61 180.11 65.68 ;
    RECT 179.9 65.97 180.11 66.04 ;
    RECT 179.9 66.33 180.11 66.4 ;
    RECT 177.04 65.61 177.25 65.68 ;
    RECT 177.04 65.97 177.25 66.04 ;
    RECT 177.04 66.33 177.25 66.4 ;
    RECT 176.58 65.61 176.79 65.68 ;
    RECT 176.58 65.97 176.79 66.04 ;
    RECT 176.58 66.33 176.79 66.4 ;
    RECT 173.72 65.61 173.93 65.68 ;
    RECT 173.72 65.97 173.93 66.04 ;
    RECT 173.72 66.33 173.93 66.4 ;
    RECT 173.26 65.61 173.47 65.68 ;
    RECT 173.26 65.97 173.47 66.04 ;
    RECT 173.26 66.33 173.47 66.4 ;
    RECT 170.4 65.61 170.61 65.68 ;
    RECT 170.4 65.97 170.61 66.04 ;
    RECT 170.4 66.33 170.61 66.4 ;
    RECT 169.94 65.61 170.15 65.68 ;
    RECT 169.94 65.97 170.15 66.04 ;
    RECT 169.94 66.33 170.15 66.4 ;
    RECT 167.08 65.61 167.29 65.68 ;
    RECT 167.08 65.97 167.29 66.04 ;
    RECT 167.08 66.33 167.29 66.4 ;
    RECT 166.62 65.61 166.83 65.68 ;
    RECT 166.62 65.97 166.83 66.04 ;
    RECT 166.62 66.33 166.83 66.4 ;
    RECT 163.76 65.61 163.97 65.68 ;
    RECT 163.76 65.97 163.97 66.04 ;
    RECT 163.76 66.33 163.97 66.4 ;
    RECT 163.3 65.61 163.51 65.68 ;
    RECT 163.3 65.97 163.51 66.04 ;
    RECT 163.3 66.33 163.51 66.4 ;
    RECT 160.44 65.61 160.65 65.68 ;
    RECT 160.44 65.97 160.65 66.04 ;
    RECT 160.44 66.33 160.65 66.4 ;
    RECT 159.98 65.61 160.19 65.68 ;
    RECT 159.98 65.97 160.19 66.04 ;
    RECT 159.98 66.33 160.19 66.4 ;
    RECT 157.12 65.61 157.33 65.68 ;
    RECT 157.12 65.97 157.33 66.04 ;
    RECT 157.12 66.33 157.33 66.4 ;
    RECT 156.66 65.61 156.87 65.68 ;
    RECT 156.66 65.97 156.87 66.04 ;
    RECT 156.66 66.33 156.87 66.4 ;
    RECT 153.8 65.61 154.01 65.68 ;
    RECT 153.8 65.97 154.01 66.04 ;
    RECT 153.8 66.33 154.01 66.4 ;
    RECT 153.34 65.61 153.55 65.68 ;
    RECT 153.34 65.97 153.55 66.04 ;
    RECT 153.34 66.33 153.55 66.4 ;
    RECT 150.48 65.61 150.69 65.68 ;
    RECT 150.48 65.97 150.69 66.04 ;
    RECT 150.48 66.33 150.69 66.4 ;
    RECT 150.02 65.61 150.23 65.68 ;
    RECT 150.02 65.97 150.23 66.04 ;
    RECT 150.02 66.33 150.23 66.4 ;
    RECT 213.56 65.61 213.77 65.68 ;
    RECT 213.56 65.97 213.77 66.04 ;
    RECT 213.56 66.33 213.77 66.4 ;
    RECT 213.1 65.61 213.31 65.68 ;
    RECT 213.1 65.97 213.31 66.04 ;
    RECT 213.1 66.33 213.31 66.4 ;
    RECT 210.24 65.61 210.45 65.68 ;
    RECT 210.24 65.97 210.45 66.04 ;
    RECT 210.24 66.33 210.45 66.4 ;
    RECT 209.78 65.61 209.99 65.68 ;
    RECT 209.78 65.97 209.99 66.04 ;
    RECT 209.78 66.33 209.99 66.4 ;
    RECT 206.92 65.61 207.13 65.68 ;
    RECT 206.92 65.97 207.13 66.04 ;
    RECT 206.92 66.33 207.13 66.4 ;
    RECT 206.46 65.61 206.67 65.68 ;
    RECT 206.46 65.97 206.67 66.04 ;
    RECT 206.46 66.33 206.67 66.4 ;
    RECT 203.6 65.61 203.81 65.68 ;
    RECT 203.6 65.97 203.81 66.04 ;
    RECT 203.6 66.33 203.81 66.4 ;
    RECT 203.14 65.61 203.35 65.68 ;
    RECT 203.14 65.97 203.35 66.04 ;
    RECT 203.14 66.33 203.35 66.4 ;
    RECT 200.28 65.61 200.49 65.68 ;
    RECT 200.28 65.97 200.49 66.04 ;
    RECT 200.28 66.33 200.49 66.4 ;
    RECT 199.82 65.61 200.03 65.68 ;
    RECT 199.82 65.97 200.03 66.04 ;
    RECT 199.82 66.33 200.03 66.4 ;
    RECT 196.96 65.61 197.17 65.68 ;
    RECT 196.96 65.97 197.17 66.04 ;
    RECT 196.96 66.33 197.17 66.4 ;
    RECT 196.5 65.61 196.71 65.68 ;
    RECT 196.5 65.97 196.71 66.04 ;
    RECT 196.5 66.33 196.71 66.4 ;
    RECT 193.64 65.61 193.85 65.68 ;
    RECT 193.64 65.97 193.85 66.04 ;
    RECT 193.64 66.33 193.85 66.4 ;
    RECT 193.18 65.61 193.39 65.68 ;
    RECT 193.18 65.97 193.39 66.04 ;
    RECT 193.18 66.33 193.39 66.4 ;
    RECT 190.32 65.61 190.53 65.68 ;
    RECT 190.32 65.97 190.53 66.04 ;
    RECT 190.32 66.33 190.53 66.4 ;
    RECT 189.86 65.61 190.07 65.68 ;
    RECT 189.86 65.97 190.07 66.04 ;
    RECT 189.86 66.33 190.07 66.4 ;
    RECT 187.0 65.61 187.21 65.68 ;
    RECT 187.0 65.97 187.21 66.04 ;
    RECT 187.0 66.33 187.21 66.4 ;
    RECT 186.54 65.61 186.75 65.68 ;
    RECT 186.54 65.97 186.75 66.04 ;
    RECT 186.54 66.33 186.75 66.4 ;
    RECT 183.68 65.61 183.89 65.68 ;
    RECT 183.68 65.97 183.89 66.04 ;
    RECT 183.68 66.33 183.89 66.4 ;
    RECT 183.22 65.61 183.43 65.68 ;
    RECT 183.22 65.97 183.43 66.04 ;
    RECT 183.22 66.33 183.43 66.4 ;
    RECT 147.485 65.97 147.555 66.04 ;
    RECT 266.68 65.61 266.89 65.68 ;
    RECT 266.68 65.97 266.89 66.04 ;
    RECT 266.68 66.33 266.89 66.4 ;
    RECT 266.22 65.61 266.43 65.68 ;
    RECT 266.22 65.97 266.43 66.04 ;
    RECT 266.22 66.33 266.43 66.4 ;
    RECT 263.36 65.61 263.57 65.68 ;
    RECT 263.36 65.97 263.57 66.04 ;
    RECT 263.36 66.33 263.57 66.4 ;
    RECT 262.9 65.61 263.11 65.68 ;
    RECT 262.9 65.97 263.11 66.04 ;
    RECT 262.9 66.33 263.11 66.4 ;
    RECT 260.04 65.61 260.25 65.68 ;
    RECT 260.04 65.97 260.25 66.04 ;
    RECT 260.04 66.33 260.25 66.4 ;
    RECT 259.58 65.61 259.79 65.68 ;
    RECT 259.58 65.97 259.79 66.04 ;
    RECT 259.58 66.33 259.79 66.4 ;
    RECT 256.72 65.61 256.93 65.68 ;
    RECT 256.72 65.97 256.93 66.04 ;
    RECT 256.72 66.33 256.93 66.4 ;
    RECT 256.26 65.61 256.47 65.68 ;
    RECT 256.26 65.97 256.47 66.04 ;
    RECT 256.26 66.33 256.47 66.4 ;
    RECT 253.4 65.61 253.61 65.68 ;
    RECT 253.4 65.97 253.61 66.04 ;
    RECT 253.4 66.33 253.61 66.4 ;
    RECT 252.94 65.61 253.15 65.68 ;
    RECT 252.94 65.97 253.15 66.04 ;
    RECT 252.94 66.33 253.15 66.4 ;
    RECT 250.08 56.23 250.29 56.3 ;
    RECT 250.08 56.59 250.29 56.66 ;
    RECT 250.08 56.95 250.29 57.02 ;
    RECT 249.62 56.23 249.83 56.3 ;
    RECT 249.62 56.59 249.83 56.66 ;
    RECT 249.62 56.95 249.83 57.02 ;
    RECT 267.91 56.59 267.98 56.66 ;
    RECT 246.76 56.23 246.97 56.3 ;
    RECT 246.76 56.59 246.97 56.66 ;
    RECT 246.76 56.95 246.97 57.02 ;
    RECT 246.3 56.23 246.51 56.3 ;
    RECT 246.3 56.59 246.51 56.66 ;
    RECT 246.3 56.95 246.51 57.02 ;
    RECT 243.44 56.23 243.65 56.3 ;
    RECT 243.44 56.59 243.65 56.66 ;
    RECT 243.44 56.95 243.65 57.02 ;
    RECT 242.98 56.23 243.19 56.3 ;
    RECT 242.98 56.59 243.19 56.66 ;
    RECT 242.98 56.95 243.19 57.02 ;
    RECT 240.12 56.23 240.33 56.3 ;
    RECT 240.12 56.59 240.33 56.66 ;
    RECT 240.12 56.95 240.33 57.02 ;
    RECT 239.66 56.23 239.87 56.3 ;
    RECT 239.66 56.59 239.87 56.66 ;
    RECT 239.66 56.95 239.87 57.02 ;
    RECT 236.8 56.23 237.01 56.3 ;
    RECT 236.8 56.59 237.01 56.66 ;
    RECT 236.8 56.95 237.01 57.02 ;
    RECT 236.34 56.23 236.55 56.3 ;
    RECT 236.34 56.59 236.55 56.66 ;
    RECT 236.34 56.95 236.55 57.02 ;
    RECT 233.48 56.23 233.69 56.3 ;
    RECT 233.48 56.59 233.69 56.66 ;
    RECT 233.48 56.95 233.69 57.02 ;
    RECT 233.02 56.23 233.23 56.3 ;
    RECT 233.02 56.59 233.23 56.66 ;
    RECT 233.02 56.95 233.23 57.02 ;
    RECT 230.16 56.23 230.37 56.3 ;
    RECT 230.16 56.59 230.37 56.66 ;
    RECT 230.16 56.95 230.37 57.02 ;
    RECT 229.7 56.23 229.91 56.3 ;
    RECT 229.7 56.59 229.91 56.66 ;
    RECT 229.7 56.95 229.91 57.02 ;
    RECT 226.84 56.23 227.05 56.3 ;
    RECT 226.84 56.59 227.05 56.66 ;
    RECT 226.84 56.95 227.05 57.02 ;
    RECT 226.38 56.23 226.59 56.3 ;
    RECT 226.38 56.59 226.59 56.66 ;
    RECT 226.38 56.95 226.59 57.02 ;
    RECT 223.52 56.23 223.73 56.3 ;
    RECT 223.52 56.59 223.73 56.66 ;
    RECT 223.52 56.95 223.73 57.02 ;
    RECT 223.06 56.23 223.27 56.3 ;
    RECT 223.06 56.59 223.27 56.66 ;
    RECT 223.06 56.95 223.27 57.02 ;
    RECT 220.2 56.23 220.41 56.3 ;
    RECT 220.2 56.59 220.41 56.66 ;
    RECT 220.2 56.95 220.41 57.02 ;
    RECT 219.74 56.23 219.95 56.3 ;
    RECT 219.74 56.59 219.95 56.66 ;
    RECT 219.74 56.95 219.95 57.02 ;
    RECT 216.88 56.23 217.09 56.3 ;
    RECT 216.88 56.59 217.09 56.66 ;
    RECT 216.88 56.95 217.09 57.02 ;
    RECT 216.42 56.23 216.63 56.3 ;
    RECT 216.42 56.59 216.63 56.66 ;
    RECT 216.42 56.95 216.63 57.02 ;
    RECT 147.485 56.59 147.555 56.66 ;
    RECT 180.36 56.23 180.57 56.3 ;
    RECT 180.36 56.59 180.57 56.66 ;
    RECT 180.36 56.95 180.57 57.02 ;
    RECT 179.9 56.23 180.11 56.3 ;
    RECT 179.9 56.59 180.11 56.66 ;
    RECT 179.9 56.95 180.11 57.02 ;
    RECT 177.04 56.23 177.25 56.3 ;
    RECT 177.04 56.59 177.25 56.66 ;
    RECT 177.04 56.95 177.25 57.02 ;
    RECT 176.58 56.23 176.79 56.3 ;
    RECT 176.58 56.59 176.79 56.66 ;
    RECT 176.58 56.95 176.79 57.02 ;
    RECT 173.72 56.23 173.93 56.3 ;
    RECT 173.72 56.59 173.93 56.66 ;
    RECT 173.72 56.95 173.93 57.02 ;
    RECT 173.26 56.23 173.47 56.3 ;
    RECT 173.26 56.59 173.47 56.66 ;
    RECT 173.26 56.95 173.47 57.02 ;
    RECT 170.4 56.23 170.61 56.3 ;
    RECT 170.4 56.59 170.61 56.66 ;
    RECT 170.4 56.95 170.61 57.02 ;
    RECT 169.94 56.23 170.15 56.3 ;
    RECT 169.94 56.59 170.15 56.66 ;
    RECT 169.94 56.95 170.15 57.02 ;
    RECT 167.08 56.23 167.29 56.3 ;
    RECT 167.08 56.59 167.29 56.66 ;
    RECT 167.08 56.95 167.29 57.02 ;
    RECT 166.62 56.23 166.83 56.3 ;
    RECT 166.62 56.59 166.83 56.66 ;
    RECT 166.62 56.95 166.83 57.02 ;
    RECT 163.76 56.23 163.97 56.3 ;
    RECT 163.76 56.59 163.97 56.66 ;
    RECT 163.76 56.95 163.97 57.02 ;
    RECT 163.3 56.23 163.51 56.3 ;
    RECT 163.3 56.59 163.51 56.66 ;
    RECT 163.3 56.95 163.51 57.02 ;
    RECT 160.44 56.23 160.65 56.3 ;
    RECT 160.44 56.59 160.65 56.66 ;
    RECT 160.44 56.95 160.65 57.02 ;
    RECT 159.98 56.23 160.19 56.3 ;
    RECT 159.98 56.59 160.19 56.66 ;
    RECT 159.98 56.95 160.19 57.02 ;
    RECT 157.12 56.23 157.33 56.3 ;
    RECT 157.12 56.59 157.33 56.66 ;
    RECT 157.12 56.95 157.33 57.02 ;
    RECT 156.66 56.23 156.87 56.3 ;
    RECT 156.66 56.59 156.87 56.66 ;
    RECT 156.66 56.95 156.87 57.02 ;
    RECT 153.8 56.23 154.01 56.3 ;
    RECT 153.8 56.59 154.01 56.66 ;
    RECT 153.8 56.95 154.01 57.02 ;
    RECT 153.34 56.23 153.55 56.3 ;
    RECT 153.34 56.59 153.55 56.66 ;
    RECT 153.34 56.95 153.55 57.02 ;
    RECT 150.48 56.23 150.69 56.3 ;
    RECT 150.48 56.59 150.69 56.66 ;
    RECT 150.48 56.95 150.69 57.02 ;
    RECT 150.02 56.23 150.23 56.3 ;
    RECT 150.02 56.59 150.23 56.66 ;
    RECT 150.02 56.95 150.23 57.02 ;
    RECT 213.56 56.23 213.77 56.3 ;
    RECT 213.56 56.59 213.77 56.66 ;
    RECT 213.56 56.95 213.77 57.02 ;
    RECT 213.1 56.23 213.31 56.3 ;
    RECT 213.1 56.59 213.31 56.66 ;
    RECT 213.1 56.95 213.31 57.02 ;
    RECT 210.24 56.23 210.45 56.3 ;
    RECT 210.24 56.59 210.45 56.66 ;
    RECT 210.24 56.95 210.45 57.02 ;
    RECT 209.78 56.23 209.99 56.3 ;
    RECT 209.78 56.59 209.99 56.66 ;
    RECT 209.78 56.95 209.99 57.02 ;
    RECT 206.92 56.23 207.13 56.3 ;
    RECT 206.92 56.59 207.13 56.66 ;
    RECT 206.92 56.95 207.13 57.02 ;
    RECT 206.46 56.23 206.67 56.3 ;
    RECT 206.46 56.59 206.67 56.66 ;
    RECT 206.46 56.95 206.67 57.02 ;
    RECT 203.6 56.23 203.81 56.3 ;
    RECT 203.6 56.59 203.81 56.66 ;
    RECT 203.6 56.95 203.81 57.02 ;
    RECT 203.14 56.23 203.35 56.3 ;
    RECT 203.14 56.59 203.35 56.66 ;
    RECT 203.14 56.95 203.35 57.02 ;
    RECT 200.28 56.23 200.49 56.3 ;
    RECT 200.28 56.59 200.49 56.66 ;
    RECT 200.28 56.95 200.49 57.02 ;
    RECT 199.82 56.23 200.03 56.3 ;
    RECT 199.82 56.59 200.03 56.66 ;
    RECT 199.82 56.95 200.03 57.02 ;
    RECT 196.96 56.23 197.17 56.3 ;
    RECT 196.96 56.59 197.17 56.66 ;
    RECT 196.96 56.95 197.17 57.02 ;
    RECT 196.5 56.23 196.71 56.3 ;
    RECT 196.5 56.59 196.71 56.66 ;
    RECT 196.5 56.95 196.71 57.02 ;
    RECT 193.64 56.23 193.85 56.3 ;
    RECT 193.64 56.59 193.85 56.66 ;
    RECT 193.64 56.95 193.85 57.02 ;
    RECT 193.18 56.23 193.39 56.3 ;
    RECT 193.18 56.59 193.39 56.66 ;
    RECT 193.18 56.95 193.39 57.02 ;
    RECT 190.32 56.23 190.53 56.3 ;
    RECT 190.32 56.59 190.53 56.66 ;
    RECT 190.32 56.95 190.53 57.02 ;
    RECT 189.86 56.23 190.07 56.3 ;
    RECT 189.86 56.59 190.07 56.66 ;
    RECT 189.86 56.95 190.07 57.02 ;
    RECT 187.0 56.23 187.21 56.3 ;
    RECT 187.0 56.59 187.21 56.66 ;
    RECT 187.0 56.95 187.21 57.02 ;
    RECT 186.54 56.23 186.75 56.3 ;
    RECT 186.54 56.59 186.75 56.66 ;
    RECT 186.54 56.95 186.75 57.02 ;
    RECT 183.68 56.23 183.89 56.3 ;
    RECT 183.68 56.59 183.89 56.66 ;
    RECT 183.68 56.95 183.89 57.02 ;
    RECT 183.22 56.23 183.43 56.3 ;
    RECT 183.22 56.59 183.43 56.66 ;
    RECT 183.22 56.95 183.43 57.02 ;
    RECT 266.68 56.23 266.89 56.3 ;
    RECT 266.68 56.59 266.89 56.66 ;
    RECT 266.68 56.95 266.89 57.02 ;
    RECT 266.22 56.23 266.43 56.3 ;
    RECT 266.22 56.59 266.43 56.66 ;
    RECT 266.22 56.95 266.43 57.02 ;
    RECT 263.36 56.23 263.57 56.3 ;
    RECT 263.36 56.59 263.57 56.66 ;
    RECT 263.36 56.95 263.57 57.02 ;
    RECT 262.9 56.23 263.11 56.3 ;
    RECT 262.9 56.59 263.11 56.66 ;
    RECT 262.9 56.95 263.11 57.02 ;
    RECT 260.04 56.23 260.25 56.3 ;
    RECT 260.04 56.59 260.25 56.66 ;
    RECT 260.04 56.95 260.25 57.02 ;
    RECT 259.58 56.23 259.79 56.3 ;
    RECT 259.58 56.59 259.79 56.66 ;
    RECT 259.58 56.95 259.79 57.02 ;
    RECT 256.72 56.23 256.93 56.3 ;
    RECT 256.72 56.59 256.93 56.66 ;
    RECT 256.72 56.95 256.93 57.02 ;
    RECT 256.26 56.23 256.47 56.3 ;
    RECT 256.26 56.59 256.47 56.66 ;
    RECT 256.26 56.95 256.47 57.02 ;
    RECT 253.4 56.23 253.61 56.3 ;
    RECT 253.4 56.59 253.61 56.66 ;
    RECT 253.4 56.95 253.61 57.02 ;
    RECT 252.94 56.23 253.15 56.3 ;
    RECT 252.94 56.59 253.15 56.66 ;
    RECT 252.94 56.95 253.15 57.02 ;
    RECT 173.26 98.97 173.47 99.04 ;
    RECT 199.33 99.23 199.54 99.3 ;
    RECT 219.25 99.23 219.46 99.3 ;
    RECT 169.45 99.23 169.66 99.3 ;
    RECT 255.77 99.49 255.98 99.56 ;
    RECT 159.49 99.49 159.7 99.56 ;
    RECT 225.89 99.49 226.1 99.56 ;
    RECT 209.78 98.97 209.99 99.04 ;
    RECT 210.24 98.97 210.45 99.04 ;
    RECT 233.02 98.97 233.23 99.04 ;
    RECT 233.48 98.97 233.69 99.04 ;
    RECT 182.73 99.49 182.94 99.56 ;
    RECT 150.02 98.97 150.23 99.04 ;
    RECT 150.48 98.97 150.69 99.04 ;
    RECT 265.73 99.23 265.94 99.3 ;
    RECT 173.72 98.97 173.93 99.04 ;
    RECT 205.97 99.49 206.18 99.56 ;
    RECT 186.54 98.97 186.75 99.04 ;
    RECT 187.0 98.97 187.21 99.04 ;
    RECT 192.69 99.23 192.9 99.3 ;
    RECT 162.81 99.23 163.02 99.3 ;
    RECT 249.13 99.49 249.34 99.56 ;
    RECT 245.81 99.23 246.02 99.3 ;
    RECT 226.38 98.97 226.59 99.04 ;
    RECT 226.84 98.97 227.05 99.04 ;
    RECT 262.9 98.97 263.11 99.04 ;
    RECT 263.36 98.97 263.57 99.04 ;
    RECT 259.09 99.23 259.3 99.3 ;
    RECT 166.62 98.97 166.83 99.04 ;
    RECT 167.08 98.97 167.29 99.04 ;
    RECT 267.135 99.75 267.355 99.82 ;
    RECT 263.815 99.75 264.035 99.82 ;
    RECT 152.85 99.49 153.06 99.56 ;
    RECT 260.495 99.75 260.715 99.82 ;
    RECT 257.175 99.75 257.395 99.82 ;
    RECT 199.33 99.49 199.54 99.56 ;
    RECT 219.25 99.49 219.46 99.56 ;
    RECT 253.855 99.75 254.075 99.82 ;
    RECT 250.535 99.75 250.755 99.82 ;
    RECT 203.14 98.97 203.35 99.04 ;
    RECT 203.6 98.97 203.81 99.04 ;
    RECT 176.09 99.49 176.3 99.56 ;
    RECT 242.49 99.49 242.7 99.56 ;
    RECT 239.17 99.23 239.38 99.3 ;
    RECT 242.98 98.97 243.19 99.04 ;
    RECT 243.44 98.97 243.65 99.04 ;
    RECT 265.73 99.49 265.94 99.56 ;
    RECT 247.215 99.75 247.435 99.82 ;
    RECT 243.895 99.75 244.115 99.82 ;
    RECT 240.575 99.75 240.795 99.82 ;
    RECT 237.255 99.75 237.475 99.82 ;
    RECT 256.26 98.97 256.47 99.04 ;
    RECT 233.935 99.75 234.155 99.82 ;
    RECT 230.615 99.75 230.835 99.82 ;
    RECT 186.05 99.23 186.26 99.3 ;
    RECT 227.295 99.75 227.515 99.82 ;
    RECT 156.17 99.23 156.38 99.3 ;
    RECT 223.975 99.75 224.195 99.82 ;
    RECT 220.655 99.75 220.875 99.82 ;
    RECT 217.335 99.75 217.555 99.82 ;
    RECT 159.98 98.97 160.19 99.04 ;
    RECT 160.44 98.97 160.65 99.04 ;
    RECT 192.69 99.49 192.9 99.56 ;
    RECT 209.29 99.23 209.5 99.3 ;
    RECT 179.41 99.23 179.62 99.3 ;
    RECT 196.5 98.97 196.71 99.04 ;
    RECT 169.45 99.49 169.66 99.56 ;
    RECT 196.96 98.97 197.17 99.04 ;
    RECT 235.85 99.49 236.06 99.56 ;
    RECT 219.74 98.97 219.95 99.04 ;
    RECT 220.2 98.97 220.41 99.04 ;
    RECT 256.72 98.97 256.93 99.04 ;
    RECT 232.53 99.23 232.74 99.3 ;
    RECT 252.45 99.23 252.66 99.3 ;
    RECT 214.015 99.75 214.235 99.82 ;
    RECT 210.695 99.75 210.915 99.82 ;
    RECT 207.375 99.75 207.595 99.82 ;
    RECT 259.09 99.49 259.3 99.56 ;
    RECT 204.055 99.75 204.275 99.82 ;
    RECT 200.735 99.75 200.955 99.82 ;
    RECT 197.415 99.75 197.635 99.82 ;
    RECT 194.095 99.75 194.315 99.82 ;
    RECT 190.775 99.75 190.995 99.82 ;
    RECT 187.455 99.75 187.675 99.82 ;
    RECT 184.135 99.75 184.355 99.82 ;
    RECT 149.53 99.23 149.74 99.3 ;
    RECT 176.58 98.97 176.79 99.04 ;
    RECT 177.04 98.97 177.25 99.04 ;
    RECT 202.65 99.23 202.86 99.3 ;
    RECT 222.57 99.23 222.78 99.3 ;
    RECT 172.77 99.23 172.98 99.3 ;
    RECT 162.81 99.49 163.02 99.56 ;
    RECT 189.86 98.97 190.07 99.04 ;
    RECT 229.21 99.49 229.42 99.56 ;
    RECT 213.1 98.97 213.31 99.04 ;
    RECT 213.56 98.97 213.77 99.04 ;
    RECT 249.62 98.97 249.83 99.04 ;
    RECT 225.89 99.23 226.1 99.3 ;
    RECT 236.34 98.97 236.55 99.04 ;
    RECT 250.08 98.97 250.29 99.04 ;
    RECT 236.8 98.97 237.01 99.04 ;
    RECT 153.34 98.97 153.55 99.04 ;
    RECT 186.05 99.49 186.26 99.56 ;
    RECT 153.8 98.97 154.01 99.04 ;
    RECT 180.815 99.75 181.035 99.82 ;
    RECT 177.495 99.75 177.715 99.82 ;
    RECT 174.175 99.75 174.395 99.82 ;
    RECT 170.855 99.75 171.075 99.82 ;
    RECT 167.535 99.75 167.755 99.82 ;
    RECT 164.215 99.75 164.435 99.82 ;
    RECT 160.895 99.75 161.115 99.82 ;
    RECT 157.575 99.75 157.795 99.82 ;
    RECT 154.255 99.75 154.475 99.82 ;
    RECT 190.32 98.97 190.53 99.04 ;
    RECT 209.29 99.49 209.5 99.56 ;
    RECT 150.935 99.75 151.155 99.82 ;
    RECT 196.01 99.23 196.22 99.3 ;
    RECT 215.93 99.23 216.14 99.3 ;
    RECT 166.13 99.23 166.34 99.3 ;
    RECT 252.45 99.49 252.66 99.56 ;
    RECT 206.46 98.97 206.67 99.04 ;
    RECT 229.7 98.97 229.91 99.04 ;
    RECT 230.16 98.97 230.37 99.04 ;
    RECT 266.22 98.97 266.43 99.04 ;
    RECT 266.68 98.97 266.89 99.04 ;
    RECT 262.41 99.23 262.62 99.3 ;
    RECT 169.94 98.97 170.15 99.04 ;
    RECT 170.4 98.97 170.61 99.04 ;
    RECT 156.17 99.49 156.38 99.56 ;
    RECT 202.65 99.49 202.86 99.56 ;
    RECT 222.57 99.49 222.78 99.56 ;
    RECT 183.22 98.97 183.43 99.04 ;
    RECT 183.68 98.97 183.89 99.04 ;
    RECT 206.92 98.97 207.13 99.04 ;
    RECT 179.41 99.49 179.62 99.56 ;
    RECT 245.81 99.49 246.02 99.56 ;
    RECT 159.49 99.23 159.7 99.3 ;
    RECT 242.49 99.23 242.7 99.3 ;
    RECT 246.3 98.97 246.51 99.04 ;
    RECT 246.76 98.97 246.97 99.04 ;
    RECT 223.06 98.97 223.27 99.04 ;
    RECT 259.58 98.97 259.79 99.04 ;
    RECT 260.04 98.97 260.25 99.04 ;
    RECT 189.37 99.23 189.58 99.3 ;
    RECT 163.3 98.97 163.51 99.04 ;
    RECT 163.76 98.97 163.97 99.04 ;
    RECT 149.53 99.49 149.74 99.56 ;
    RECT 196.01 99.49 196.22 99.56 ;
    RECT 215.93 99.49 216.14 99.56 ;
    RECT 212.61 99.23 212.82 99.3 ;
    RECT 199.82 98.97 200.03 99.04 ;
    RECT 200.28 98.97 200.49 99.04 ;
    RECT 172.77 99.49 172.98 99.56 ;
    RECT 239.17 99.49 239.38 99.56 ;
    RECT 223.52 98.97 223.73 99.04 ;
    RECT 235.85 99.23 236.06 99.3 ;
    RECT 255.77 99.23 255.98 99.3 ;
    RECT 239.66 98.97 239.87 99.04 ;
    RECT 262.41 99.49 262.62 99.56 ;
    RECT 182.73 99.23 182.94 99.3 ;
    RECT 152.85 99.23 153.06 99.3 ;
    RECT 156.66 98.97 156.87 99.04 ;
    RECT 179.9 98.97 180.11 99.04 ;
    RECT 180.36 98.97 180.57 99.04 ;
    RECT 205.97 99.23 206.18 99.3 ;
    RECT 176.09 99.23 176.3 99.3 ;
    RECT 193.18 98.97 193.39 99.04 ;
    RECT 166.13 99.49 166.34 99.56 ;
    RECT 193.64 98.97 193.85 99.04 ;
    RECT 232.53 99.49 232.74 99.56 ;
    RECT 216.42 98.97 216.63 99.04 ;
    RECT 216.88 98.97 217.09 99.04 ;
    RECT 252.94 98.97 253.15 99.04 ;
    RECT 253.4 98.97 253.61 99.04 ;
    RECT 229.21 99.23 229.42 99.3 ;
    RECT 249.13 99.23 249.34 99.3 ;
    RECT 240.12 98.97 240.33 99.04 ;
    RECT 268.12 99.23 268.19 99.3 ;
    RECT 267.91 98.97 267.98 99.04 ;
    RECT 157.12 98.97 157.33 99.04 ;
    RECT 189.37 99.49 189.58 99.56 ;
    RECT 147.275 99.23 147.345 99.3 ;
    RECT 147.485 98.97 147.555 99.04 ;
    RECT 212.61 99.49 212.82 99.56 ;
    RECT 250.08 28.15 250.29 28.22 ;
    RECT 250.08 28.51 250.29 28.58 ;
    RECT 250.08 28.87 250.29 28.94 ;
    RECT 249.62 28.15 249.83 28.22 ;
    RECT 249.62 28.51 249.83 28.58 ;
    RECT 249.62 28.87 249.83 28.94 ;
    RECT 246.76 28.15 246.97 28.22 ;
    RECT 246.76 28.51 246.97 28.58 ;
    RECT 246.76 28.87 246.97 28.94 ;
    RECT 246.3 28.15 246.51 28.22 ;
    RECT 246.3 28.51 246.51 28.58 ;
    RECT 246.3 28.87 246.51 28.94 ;
    RECT 243.44 28.15 243.65 28.22 ;
    RECT 243.44 28.51 243.65 28.58 ;
    RECT 243.44 28.87 243.65 28.94 ;
    RECT 242.98 28.15 243.19 28.22 ;
    RECT 242.98 28.51 243.19 28.58 ;
    RECT 242.98 28.87 243.19 28.94 ;
    RECT 240.12 28.15 240.33 28.22 ;
    RECT 240.12 28.51 240.33 28.58 ;
    RECT 240.12 28.87 240.33 28.94 ;
    RECT 239.66 28.15 239.87 28.22 ;
    RECT 239.66 28.51 239.87 28.58 ;
    RECT 239.66 28.87 239.87 28.94 ;
    RECT 236.8 28.15 237.01 28.22 ;
    RECT 236.8 28.51 237.01 28.58 ;
    RECT 236.8 28.87 237.01 28.94 ;
    RECT 236.34 28.15 236.55 28.22 ;
    RECT 236.34 28.51 236.55 28.58 ;
    RECT 236.34 28.87 236.55 28.94 ;
    RECT 233.48 28.15 233.69 28.22 ;
    RECT 233.48 28.51 233.69 28.58 ;
    RECT 233.48 28.87 233.69 28.94 ;
    RECT 233.02 28.15 233.23 28.22 ;
    RECT 233.02 28.51 233.23 28.58 ;
    RECT 233.02 28.87 233.23 28.94 ;
    RECT 230.16 28.15 230.37 28.22 ;
    RECT 230.16 28.51 230.37 28.58 ;
    RECT 230.16 28.87 230.37 28.94 ;
    RECT 229.7 28.15 229.91 28.22 ;
    RECT 229.7 28.51 229.91 28.58 ;
    RECT 229.7 28.87 229.91 28.94 ;
    RECT 226.84 28.15 227.05 28.22 ;
    RECT 226.84 28.51 227.05 28.58 ;
    RECT 226.84 28.87 227.05 28.94 ;
    RECT 226.38 28.15 226.59 28.22 ;
    RECT 226.38 28.51 226.59 28.58 ;
    RECT 226.38 28.87 226.59 28.94 ;
    RECT 223.52 28.15 223.73 28.22 ;
    RECT 223.52 28.51 223.73 28.58 ;
    RECT 223.52 28.87 223.73 28.94 ;
    RECT 223.06 28.15 223.27 28.22 ;
    RECT 223.06 28.51 223.27 28.58 ;
    RECT 223.06 28.87 223.27 28.94 ;
    RECT 220.2 28.15 220.41 28.22 ;
    RECT 220.2 28.51 220.41 28.58 ;
    RECT 220.2 28.87 220.41 28.94 ;
    RECT 219.74 28.15 219.95 28.22 ;
    RECT 219.74 28.51 219.95 28.58 ;
    RECT 219.74 28.87 219.95 28.94 ;
    RECT 216.88 28.15 217.09 28.22 ;
    RECT 216.88 28.51 217.09 28.58 ;
    RECT 216.88 28.87 217.09 28.94 ;
    RECT 216.42 28.15 216.63 28.22 ;
    RECT 216.42 28.51 216.63 28.58 ;
    RECT 216.42 28.87 216.63 28.94 ;
    RECT 267.91 28.51 267.98 28.58 ;
    RECT 180.36 28.15 180.57 28.22 ;
    RECT 180.36 28.51 180.57 28.58 ;
    RECT 180.36 28.87 180.57 28.94 ;
    RECT 179.9 28.15 180.11 28.22 ;
    RECT 179.9 28.51 180.11 28.58 ;
    RECT 179.9 28.87 180.11 28.94 ;
    RECT 177.04 28.15 177.25 28.22 ;
    RECT 177.04 28.51 177.25 28.58 ;
    RECT 177.04 28.87 177.25 28.94 ;
    RECT 176.58 28.15 176.79 28.22 ;
    RECT 176.58 28.51 176.79 28.58 ;
    RECT 176.58 28.87 176.79 28.94 ;
    RECT 173.72 28.15 173.93 28.22 ;
    RECT 173.72 28.51 173.93 28.58 ;
    RECT 173.72 28.87 173.93 28.94 ;
    RECT 173.26 28.15 173.47 28.22 ;
    RECT 173.26 28.51 173.47 28.58 ;
    RECT 173.26 28.87 173.47 28.94 ;
    RECT 170.4 28.15 170.61 28.22 ;
    RECT 170.4 28.51 170.61 28.58 ;
    RECT 170.4 28.87 170.61 28.94 ;
    RECT 169.94 28.15 170.15 28.22 ;
    RECT 169.94 28.51 170.15 28.58 ;
    RECT 169.94 28.87 170.15 28.94 ;
    RECT 167.08 28.15 167.29 28.22 ;
    RECT 167.08 28.51 167.29 28.58 ;
    RECT 167.08 28.87 167.29 28.94 ;
    RECT 166.62 28.15 166.83 28.22 ;
    RECT 166.62 28.51 166.83 28.58 ;
    RECT 166.62 28.87 166.83 28.94 ;
    RECT 163.76 28.15 163.97 28.22 ;
    RECT 163.76 28.51 163.97 28.58 ;
    RECT 163.76 28.87 163.97 28.94 ;
    RECT 163.3 28.15 163.51 28.22 ;
    RECT 163.3 28.51 163.51 28.58 ;
    RECT 163.3 28.87 163.51 28.94 ;
    RECT 160.44 28.15 160.65 28.22 ;
    RECT 160.44 28.51 160.65 28.58 ;
    RECT 160.44 28.87 160.65 28.94 ;
    RECT 159.98 28.15 160.19 28.22 ;
    RECT 159.98 28.51 160.19 28.58 ;
    RECT 159.98 28.87 160.19 28.94 ;
    RECT 157.12 28.15 157.33 28.22 ;
    RECT 157.12 28.51 157.33 28.58 ;
    RECT 157.12 28.87 157.33 28.94 ;
    RECT 156.66 28.15 156.87 28.22 ;
    RECT 156.66 28.51 156.87 28.58 ;
    RECT 156.66 28.87 156.87 28.94 ;
    RECT 153.8 28.15 154.01 28.22 ;
    RECT 153.8 28.51 154.01 28.58 ;
    RECT 153.8 28.87 154.01 28.94 ;
    RECT 153.34 28.15 153.55 28.22 ;
    RECT 153.34 28.51 153.55 28.58 ;
    RECT 153.34 28.87 153.55 28.94 ;
    RECT 150.48 28.15 150.69 28.22 ;
    RECT 150.48 28.51 150.69 28.58 ;
    RECT 150.48 28.87 150.69 28.94 ;
    RECT 150.02 28.15 150.23 28.22 ;
    RECT 150.02 28.51 150.23 28.58 ;
    RECT 150.02 28.87 150.23 28.94 ;
    RECT 213.56 28.15 213.77 28.22 ;
    RECT 213.56 28.51 213.77 28.58 ;
    RECT 213.56 28.87 213.77 28.94 ;
    RECT 213.1 28.15 213.31 28.22 ;
    RECT 213.1 28.51 213.31 28.58 ;
    RECT 213.1 28.87 213.31 28.94 ;
    RECT 210.24 28.15 210.45 28.22 ;
    RECT 210.24 28.51 210.45 28.58 ;
    RECT 210.24 28.87 210.45 28.94 ;
    RECT 209.78 28.15 209.99 28.22 ;
    RECT 209.78 28.51 209.99 28.58 ;
    RECT 209.78 28.87 209.99 28.94 ;
    RECT 206.92 28.15 207.13 28.22 ;
    RECT 206.92 28.51 207.13 28.58 ;
    RECT 206.92 28.87 207.13 28.94 ;
    RECT 206.46 28.15 206.67 28.22 ;
    RECT 206.46 28.51 206.67 28.58 ;
    RECT 206.46 28.87 206.67 28.94 ;
    RECT 203.6 28.15 203.81 28.22 ;
    RECT 203.6 28.51 203.81 28.58 ;
    RECT 203.6 28.87 203.81 28.94 ;
    RECT 203.14 28.15 203.35 28.22 ;
    RECT 203.14 28.51 203.35 28.58 ;
    RECT 203.14 28.87 203.35 28.94 ;
    RECT 200.28 28.15 200.49 28.22 ;
    RECT 200.28 28.51 200.49 28.58 ;
    RECT 200.28 28.87 200.49 28.94 ;
    RECT 199.82 28.15 200.03 28.22 ;
    RECT 199.82 28.51 200.03 28.58 ;
    RECT 199.82 28.87 200.03 28.94 ;
    RECT 196.96 28.15 197.17 28.22 ;
    RECT 196.96 28.51 197.17 28.58 ;
    RECT 196.96 28.87 197.17 28.94 ;
    RECT 196.5 28.15 196.71 28.22 ;
    RECT 196.5 28.51 196.71 28.58 ;
    RECT 196.5 28.87 196.71 28.94 ;
    RECT 193.64 28.15 193.85 28.22 ;
    RECT 193.64 28.51 193.85 28.58 ;
    RECT 193.64 28.87 193.85 28.94 ;
    RECT 193.18 28.15 193.39 28.22 ;
    RECT 193.18 28.51 193.39 28.58 ;
    RECT 193.18 28.87 193.39 28.94 ;
    RECT 190.32 28.15 190.53 28.22 ;
    RECT 190.32 28.51 190.53 28.58 ;
    RECT 190.32 28.87 190.53 28.94 ;
    RECT 189.86 28.15 190.07 28.22 ;
    RECT 189.86 28.51 190.07 28.58 ;
    RECT 189.86 28.87 190.07 28.94 ;
    RECT 187.0 28.15 187.21 28.22 ;
    RECT 187.0 28.51 187.21 28.58 ;
    RECT 187.0 28.87 187.21 28.94 ;
    RECT 186.54 28.15 186.75 28.22 ;
    RECT 186.54 28.51 186.75 28.58 ;
    RECT 186.54 28.87 186.75 28.94 ;
    RECT 183.68 28.15 183.89 28.22 ;
    RECT 183.68 28.51 183.89 28.58 ;
    RECT 183.68 28.87 183.89 28.94 ;
    RECT 183.22 28.15 183.43 28.22 ;
    RECT 183.22 28.51 183.43 28.58 ;
    RECT 183.22 28.87 183.43 28.94 ;
    RECT 147.485 28.51 147.555 28.58 ;
    RECT 266.68 28.15 266.89 28.22 ;
    RECT 266.68 28.51 266.89 28.58 ;
    RECT 266.68 28.87 266.89 28.94 ;
    RECT 266.22 28.15 266.43 28.22 ;
    RECT 266.22 28.51 266.43 28.58 ;
    RECT 266.22 28.87 266.43 28.94 ;
    RECT 263.36 28.15 263.57 28.22 ;
    RECT 263.36 28.51 263.57 28.58 ;
    RECT 263.36 28.87 263.57 28.94 ;
    RECT 262.9 28.15 263.11 28.22 ;
    RECT 262.9 28.51 263.11 28.58 ;
    RECT 262.9 28.87 263.11 28.94 ;
    RECT 260.04 28.15 260.25 28.22 ;
    RECT 260.04 28.51 260.25 28.58 ;
    RECT 260.04 28.87 260.25 28.94 ;
    RECT 259.58 28.15 259.79 28.22 ;
    RECT 259.58 28.51 259.79 28.58 ;
    RECT 259.58 28.87 259.79 28.94 ;
    RECT 256.72 28.15 256.93 28.22 ;
    RECT 256.72 28.51 256.93 28.58 ;
    RECT 256.72 28.87 256.93 28.94 ;
    RECT 256.26 28.15 256.47 28.22 ;
    RECT 256.26 28.51 256.47 28.58 ;
    RECT 256.26 28.87 256.47 28.94 ;
    RECT 253.4 28.15 253.61 28.22 ;
    RECT 253.4 28.51 253.61 28.58 ;
    RECT 253.4 28.87 253.61 28.94 ;
    RECT 252.94 28.15 253.15 28.22 ;
    RECT 252.94 28.51 253.15 28.58 ;
    RECT 252.94 28.87 253.15 28.94 ;
    RECT 250.08 27.43 250.29 27.5 ;
    RECT 250.08 27.79 250.29 27.86 ;
    RECT 250.08 28.15 250.29 28.22 ;
    RECT 249.62 27.43 249.83 27.5 ;
    RECT 249.62 27.79 249.83 27.86 ;
    RECT 249.62 28.15 249.83 28.22 ;
    RECT 246.76 27.43 246.97 27.5 ;
    RECT 246.76 27.79 246.97 27.86 ;
    RECT 246.76 28.15 246.97 28.22 ;
    RECT 246.3 27.43 246.51 27.5 ;
    RECT 246.3 27.79 246.51 27.86 ;
    RECT 246.3 28.15 246.51 28.22 ;
    RECT 243.44 27.43 243.65 27.5 ;
    RECT 243.44 27.79 243.65 27.86 ;
    RECT 243.44 28.15 243.65 28.22 ;
    RECT 242.98 27.43 243.19 27.5 ;
    RECT 242.98 27.79 243.19 27.86 ;
    RECT 242.98 28.15 243.19 28.22 ;
    RECT 240.12 27.43 240.33 27.5 ;
    RECT 240.12 27.79 240.33 27.86 ;
    RECT 240.12 28.15 240.33 28.22 ;
    RECT 239.66 27.43 239.87 27.5 ;
    RECT 239.66 27.79 239.87 27.86 ;
    RECT 239.66 28.15 239.87 28.22 ;
    RECT 236.8 27.43 237.01 27.5 ;
    RECT 236.8 27.79 237.01 27.86 ;
    RECT 236.8 28.15 237.01 28.22 ;
    RECT 236.34 27.43 236.55 27.5 ;
    RECT 236.34 27.79 236.55 27.86 ;
    RECT 236.34 28.15 236.55 28.22 ;
    RECT 233.48 27.43 233.69 27.5 ;
    RECT 233.48 27.79 233.69 27.86 ;
    RECT 233.48 28.15 233.69 28.22 ;
    RECT 233.02 27.43 233.23 27.5 ;
    RECT 233.02 27.79 233.23 27.86 ;
    RECT 233.02 28.15 233.23 28.22 ;
    RECT 230.16 27.43 230.37 27.5 ;
    RECT 230.16 27.79 230.37 27.86 ;
    RECT 230.16 28.15 230.37 28.22 ;
    RECT 229.7 27.43 229.91 27.5 ;
    RECT 229.7 27.79 229.91 27.86 ;
    RECT 229.7 28.15 229.91 28.22 ;
    RECT 226.84 27.43 227.05 27.5 ;
    RECT 226.84 27.79 227.05 27.86 ;
    RECT 226.84 28.15 227.05 28.22 ;
    RECT 226.38 27.43 226.59 27.5 ;
    RECT 226.38 27.79 226.59 27.86 ;
    RECT 226.38 28.15 226.59 28.22 ;
    RECT 223.52 27.43 223.73 27.5 ;
    RECT 223.52 27.79 223.73 27.86 ;
    RECT 223.52 28.15 223.73 28.22 ;
    RECT 223.06 27.43 223.27 27.5 ;
    RECT 223.06 27.79 223.27 27.86 ;
    RECT 223.06 28.15 223.27 28.22 ;
    RECT 220.2 27.43 220.41 27.5 ;
    RECT 220.2 27.79 220.41 27.86 ;
    RECT 220.2 28.15 220.41 28.22 ;
    RECT 219.74 27.43 219.95 27.5 ;
    RECT 219.74 27.79 219.95 27.86 ;
    RECT 219.74 28.15 219.95 28.22 ;
    RECT 216.88 27.43 217.09 27.5 ;
    RECT 216.88 27.79 217.09 27.86 ;
    RECT 216.88 28.15 217.09 28.22 ;
    RECT 216.42 27.43 216.63 27.5 ;
    RECT 216.42 27.79 216.63 27.86 ;
    RECT 216.42 28.15 216.63 28.22 ;
    RECT 267.91 27.79 267.98 27.86 ;
    RECT 180.36 27.43 180.57 27.5 ;
    RECT 180.36 27.79 180.57 27.86 ;
    RECT 180.36 28.15 180.57 28.22 ;
    RECT 179.9 27.43 180.11 27.5 ;
    RECT 179.9 27.79 180.11 27.86 ;
    RECT 179.9 28.15 180.11 28.22 ;
    RECT 177.04 27.43 177.25 27.5 ;
    RECT 177.04 27.79 177.25 27.86 ;
    RECT 177.04 28.15 177.25 28.22 ;
    RECT 176.58 27.43 176.79 27.5 ;
    RECT 176.58 27.79 176.79 27.86 ;
    RECT 176.58 28.15 176.79 28.22 ;
    RECT 173.72 27.43 173.93 27.5 ;
    RECT 173.72 27.79 173.93 27.86 ;
    RECT 173.72 28.15 173.93 28.22 ;
    RECT 173.26 27.43 173.47 27.5 ;
    RECT 173.26 27.79 173.47 27.86 ;
    RECT 173.26 28.15 173.47 28.22 ;
    RECT 170.4 27.43 170.61 27.5 ;
    RECT 170.4 27.79 170.61 27.86 ;
    RECT 170.4 28.15 170.61 28.22 ;
    RECT 169.94 27.43 170.15 27.5 ;
    RECT 169.94 27.79 170.15 27.86 ;
    RECT 169.94 28.15 170.15 28.22 ;
    RECT 167.08 27.43 167.29 27.5 ;
    RECT 167.08 27.79 167.29 27.86 ;
    RECT 167.08 28.15 167.29 28.22 ;
    RECT 166.62 27.43 166.83 27.5 ;
    RECT 166.62 27.79 166.83 27.86 ;
    RECT 166.62 28.15 166.83 28.22 ;
    RECT 163.76 27.43 163.97 27.5 ;
    RECT 163.76 27.79 163.97 27.86 ;
    RECT 163.76 28.15 163.97 28.22 ;
    RECT 163.3 27.43 163.51 27.5 ;
    RECT 163.3 27.79 163.51 27.86 ;
    RECT 163.3 28.15 163.51 28.22 ;
    RECT 160.44 27.43 160.65 27.5 ;
    RECT 160.44 27.79 160.65 27.86 ;
    RECT 160.44 28.15 160.65 28.22 ;
    RECT 159.98 27.43 160.19 27.5 ;
    RECT 159.98 27.79 160.19 27.86 ;
    RECT 159.98 28.15 160.19 28.22 ;
    RECT 157.12 27.43 157.33 27.5 ;
    RECT 157.12 27.79 157.33 27.86 ;
    RECT 157.12 28.15 157.33 28.22 ;
    RECT 156.66 27.43 156.87 27.5 ;
    RECT 156.66 27.79 156.87 27.86 ;
    RECT 156.66 28.15 156.87 28.22 ;
    RECT 153.8 27.43 154.01 27.5 ;
    RECT 153.8 27.79 154.01 27.86 ;
    RECT 153.8 28.15 154.01 28.22 ;
    RECT 153.34 27.43 153.55 27.5 ;
    RECT 153.34 27.79 153.55 27.86 ;
    RECT 153.34 28.15 153.55 28.22 ;
    RECT 150.48 27.43 150.69 27.5 ;
    RECT 150.48 27.79 150.69 27.86 ;
    RECT 150.48 28.15 150.69 28.22 ;
    RECT 150.02 27.43 150.23 27.5 ;
    RECT 150.02 27.79 150.23 27.86 ;
    RECT 150.02 28.15 150.23 28.22 ;
    RECT 213.56 27.43 213.77 27.5 ;
    RECT 213.56 27.79 213.77 27.86 ;
    RECT 213.56 28.15 213.77 28.22 ;
    RECT 213.1 27.43 213.31 27.5 ;
    RECT 213.1 27.79 213.31 27.86 ;
    RECT 213.1 28.15 213.31 28.22 ;
    RECT 210.24 27.43 210.45 27.5 ;
    RECT 210.24 27.79 210.45 27.86 ;
    RECT 210.24 28.15 210.45 28.22 ;
    RECT 209.78 27.43 209.99 27.5 ;
    RECT 209.78 27.79 209.99 27.86 ;
    RECT 209.78 28.15 209.99 28.22 ;
    RECT 206.92 27.43 207.13 27.5 ;
    RECT 206.92 27.79 207.13 27.86 ;
    RECT 206.92 28.15 207.13 28.22 ;
    RECT 206.46 27.43 206.67 27.5 ;
    RECT 206.46 27.79 206.67 27.86 ;
    RECT 206.46 28.15 206.67 28.22 ;
    RECT 203.6 27.43 203.81 27.5 ;
    RECT 203.6 27.79 203.81 27.86 ;
    RECT 203.6 28.15 203.81 28.22 ;
    RECT 203.14 27.43 203.35 27.5 ;
    RECT 203.14 27.79 203.35 27.86 ;
    RECT 203.14 28.15 203.35 28.22 ;
    RECT 200.28 27.43 200.49 27.5 ;
    RECT 200.28 27.79 200.49 27.86 ;
    RECT 200.28 28.15 200.49 28.22 ;
    RECT 199.82 27.43 200.03 27.5 ;
    RECT 199.82 27.79 200.03 27.86 ;
    RECT 199.82 28.15 200.03 28.22 ;
    RECT 196.96 27.43 197.17 27.5 ;
    RECT 196.96 27.79 197.17 27.86 ;
    RECT 196.96 28.15 197.17 28.22 ;
    RECT 196.5 27.43 196.71 27.5 ;
    RECT 196.5 27.79 196.71 27.86 ;
    RECT 196.5 28.15 196.71 28.22 ;
    RECT 193.64 27.43 193.85 27.5 ;
    RECT 193.64 27.79 193.85 27.86 ;
    RECT 193.64 28.15 193.85 28.22 ;
    RECT 193.18 27.43 193.39 27.5 ;
    RECT 193.18 27.79 193.39 27.86 ;
    RECT 193.18 28.15 193.39 28.22 ;
    RECT 190.32 27.43 190.53 27.5 ;
    RECT 190.32 27.79 190.53 27.86 ;
    RECT 190.32 28.15 190.53 28.22 ;
    RECT 189.86 27.43 190.07 27.5 ;
    RECT 189.86 27.79 190.07 27.86 ;
    RECT 189.86 28.15 190.07 28.22 ;
    RECT 187.0 27.43 187.21 27.5 ;
    RECT 187.0 27.79 187.21 27.86 ;
    RECT 187.0 28.15 187.21 28.22 ;
    RECT 186.54 27.43 186.75 27.5 ;
    RECT 186.54 27.79 186.75 27.86 ;
    RECT 186.54 28.15 186.75 28.22 ;
    RECT 183.68 27.43 183.89 27.5 ;
    RECT 183.68 27.79 183.89 27.86 ;
    RECT 183.68 28.15 183.89 28.22 ;
    RECT 183.22 27.43 183.43 27.5 ;
    RECT 183.22 27.79 183.43 27.86 ;
    RECT 183.22 28.15 183.43 28.22 ;
    RECT 147.485 27.79 147.555 27.86 ;
    RECT 266.68 27.43 266.89 27.5 ;
    RECT 266.68 27.79 266.89 27.86 ;
    RECT 266.68 28.15 266.89 28.22 ;
    RECT 266.22 27.43 266.43 27.5 ;
    RECT 266.22 27.79 266.43 27.86 ;
    RECT 266.22 28.15 266.43 28.22 ;
    RECT 263.36 27.43 263.57 27.5 ;
    RECT 263.36 27.79 263.57 27.86 ;
    RECT 263.36 28.15 263.57 28.22 ;
    RECT 262.9 27.43 263.11 27.5 ;
    RECT 262.9 27.79 263.11 27.86 ;
    RECT 262.9 28.15 263.11 28.22 ;
    RECT 260.04 27.43 260.25 27.5 ;
    RECT 260.04 27.79 260.25 27.86 ;
    RECT 260.04 28.15 260.25 28.22 ;
    RECT 259.58 27.43 259.79 27.5 ;
    RECT 259.58 27.79 259.79 27.86 ;
    RECT 259.58 28.15 259.79 28.22 ;
    RECT 256.72 27.43 256.93 27.5 ;
    RECT 256.72 27.79 256.93 27.86 ;
    RECT 256.72 28.15 256.93 28.22 ;
    RECT 256.26 27.43 256.47 27.5 ;
    RECT 256.26 27.79 256.47 27.86 ;
    RECT 256.26 28.15 256.47 28.22 ;
    RECT 253.4 27.43 253.61 27.5 ;
    RECT 253.4 27.79 253.61 27.86 ;
    RECT 253.4 28.15 253.61 28.22 ;
    RECT 252.94 27.43 253.15 27.5 ;
    RECT 252.94 27.79 253.15 27.86 ;
    RECT 252.94 28.15 253.15 28.22 ;
    RECT 250.08 26.71 250.29 26.78 ;
    RECT 250.08 27.07 250.29 27.14 ;
    RECT 250.08 27.43 250.29 27.5 ;
    RECT 249.62 26.71 249.83 26.78 ;
    RECT 249.62 27.07 249.83 27.14 ;
    RECT 249.62 27.43 249.83 27.5 ;
    RECT 246.76 26.71 246.97 26.78 ;
    RECT 246.76 27.07 246.97 27.14 ;
    RECT 246.76 27.43 246.97 27.5 ;
    RECT 246.3 26.71 246.51 26.78 ;
    RECT 246.3 27.07 246.51 27.14 ;
    RECT 246.3 27.43 246.51 27.5 ;
    RECT 243.44 26.71 243.65 26.78 ;
    RECT 243.44 27.07 243.65 27.14 ;
    RECT 243.44 27.43 243.65 27.5 ;
    RECT 242.98 26.71 243.19 26.78 ;
    RECT 242.98 27.07 243.19 27.14 ;
    RECT 242.98 27.43 243.19 27.5 ;
    RECT 240.12 26.71 240.33 26.78 ;
    RECT 240.12 27.07 240.33 27.14 ;
    RECT 240.12 27.43 240.33 27.5 ;
    RECT 239.66 26.71 239.87 26.78 ;
    RECT 239.66 27.07 239.87 27.14 ;
    RECT 239.66 27.43 239.87 27.5 ;
    RECT 236.8 26.71 237.01 26.78 ;
    RECT 236.8 27.07 237.01 27.14 ;
    RECT 236.8 27.43 237.01 27.5 ;
    RECT 236.34 26.71 236.55 26.78 ;
    RECT 236.34 27.07 236.55 27.14 ;
    RECT 236.34 27.43 236.55 27.5 ;
    RECT 233.48 26.71 233.69 26.78 ;
    RECT 233.48 27.07 233.69 27.14 ;
    RECT 233.48 27.43 233.69 27.5 ;
    RECT 233.02 26.71 233.23 26.78 ;
    RECT 233.02 27.07 233.23 27.14 ;
    RECT 233.02 27.43 233.23 27.5 ;
    RECT 230.16 26.71 230.37 26.78 ;
    RECT 230.16 27.07 230.37 27.14 ;
    RECT 230.16 27.43 230.37 27.5 ;
    RECT 229.7 26.71 229.91 26.78 ;
    RECT 229.7 27.07 229.91 27.14 ;
    RECT 229.7 27.43 229.91 27.5 ;
    RECT 226.84 26.71 227.05 26.78 ;
    RECT 226.84 27.07 227.05 27.14 ;
    RECT 226.84 27.43 227.05 27.5 ;
    RECT 226.38 26.71 226.59 26.78 ;
    RECT 226.38 27.07 226.59 27.14 ;
    RECT 226.38 27.43 226.59 27.5 ;
    RECT 223.52 26.71 223.73 26.78 ;
    RECT 223.52 27.07 223.73 27.14 ;
    RECT 223.52 27.43 223.73 27.5 ;
    RECT 223.06 26.71 223.27 26.78 ;
    RECT 223.06 27.07 223.27 27.14 ;
    RECT 223.06 27.43 223.27 27.5 ;
    RECT 220.2 26.71 220.41 26.78 ;
    RECT 220.2 27.07 220.41 27.14 ;
    RECT 220.2 27.43 220.41 27.5 ;
    RECT 219.74 26.71 219.95 26.78 ;
    RECT 219.74 27.07 219.95 27.14 ;
    RECT 219.74 27.43 219.95 27.5 ;
    RECT 216.88 26.71 217.09 26.78 ;
    RECT 216.88 27.07 217.09 27.14 ;
    RECT 216.88 27.43 217.09 27.5 ;
    RECT 216.42 26.71 216.63 26.78 ;
    RECT 216.42 27.07 216.63 27.14 ;
    RECT 216.42 27.43 216.63 27.5 ;
    RECT 267.91 27.07 267.98 27.14 ;
    RECT 180.36 26.71 180.57 26.78 ;
    RECT 180.36 27.07 180.57 27.14 ;
    RECT 180.36 27.43 180.57 27.5 ;
    RECT 179.9 26.71 180.11 26.78 ;
    RECT 179.9 27.07 180.11 27.14 ;
    RECT 179.9 27.43 180.11 27.5 ;
    RECT 177.04 26.71 177.25 26.78 ;
    RECT 177.04 27.07 177.25 27.14 ;
    RECT 177.04 27.43 177.25 27.5 ;
    RECT 176.58 26.71 176.79 26.78 ;
    RECT 176.58 27.07 176.79 27.14 ;
    RECT 176.58 27.43 176.79 27.5 ;
    RECT 173.72 26.71 173.93 26.78 ;
    RECT 173.72 27.07 173.93 27.14 ;
    RECT 173.72 27.43 173.93 27.5 ;
    RECT 173.26 26.71 173.47 26.78 ;
    RECT 173.26 27.07 173.47 27.14 ;
    RECT 173.26 27.43 173.47 27.5 ;
    RECT 170.4 26.71 170.61 26.78 ;
    RECT 170.4 27.07 170.61 27.14 ;
    RECT 170.4 27.43 170.61 27.5 ;
    RECT 169.94 26.71 170.15 26.78 ;
    RECT 169.94 27.07 170.15 27.14 ;
    RECT 169.94 27.43 170.15 27.5 ;
    RECT 167.08 26.71 167.29 26.78 ;
    RECT 167.08 27.07 167.29 27.14 ;
    RECT 167.08 27.43 167.29 27.5 ;
    RECT 166.62 26.71 166.83 26.78 ;
    RECT 166.62 27.07 166.83 27.14 ;
    RECT 166.62 27.43 166.83 27.5 ;
    RECT 163.76 26.71 163.97 26.78 ;
    RECT 163.76 27.07 163.97 27.14 ;
    RECT 163.76 27.43 163.97 27.5 ;
    RECT 163.3 26.71 163.51 26.78 ;
    RECT 163.3 27.07 163.51 27.14 ;
    RECT 163.3 27.43 163.51 27.5 ;
    RECT 160.44 26.71 160.65 26.78 ;
    RECT 160.44 27.07 160.65 27.14 ;
    RECT 160.44 27.43 160.65 27.5 ;
    RECT 159.98 26.71 160.19 26.78 ;
    RECT 159.98 27.07 160.19 27.14 ;
    RECT 159.98 27.43 160.19 27.5 ;
    RECT 157.12 26.71 157.33 26.78 ;
    RECT 157.12 27.07 157.33 27.14 ;
    RECT 157.12 27.43 157.33 27.5 ;
    RECT 156.66 26.71 156.87 26.78 ;
    RECT 156.66 27.07 156.87 27.14 ;
    RECT 156.66 27.43 156.87 27.5 ;
    RECT 153.8 26.71 154.01 26.78 ;
    RECT 153.8 27.07 154.01 27.14 ;
    RECT 153.8 27.43 154.01 27.5 ;
    RECT 153.34 26.71 153.55 26.78 ;
    RECT 153.34 27.07 153.55 27.14 ;
    RECT 153.34 27.43 153.55 27.5 ;
    RECT 150.48 26.71 150.69 26.78 ;
    RECT 150.48 27.07 150.69 27.14 ;
    RECT 150.48 27.43 150.69 27.5 ;
    RECT 150.02 26.71 150.23 26.78 ;
    RECT 150.02 27.07 150.23 27.14 ;
    RECT 150.02 27.43 150.23 27.5 ;
    RECT 213.56 26.71 213.77 26.78 ;
    RECT 213.56 27.07 213.77 27.14 ;
    RECT 213.56 27.43 213.77 27.5 ;
    RECT 213.1 26.71 213.31 26.78 ;
    RECT 213.1 27.07 213.31 27.14 ;
    RECT 213.1 27.43 213.31 27.5 ;
    RECT 210.24 26.71 210.45 26.78 ;
    RECT 210.24 27.07 210.45 27.14 ;
    RECT 210.24 27.43 210.45 27.5 ;
    RECT 209.78 26.71 209.99 26.78 ;
    RECT 209.78 27.07 209.99 27.14 ;
    RECT 209.78 27.43 209.99 27.5 ;
    RECT 206.92 26.71 207.13 26.78 ;
    RECT 206.92 27.07 207.13 27.14 ;
    RECT 206.92 27.43 207.13 27.5 ;
    RECT 206.46 26.71 206.67 26.78 ;
    RECT 206.46 27.07 206.67 27.14 ;
    RECT 206.46 27.43 206.67 27.5 ;
    RECT 203.6 26.71 203.81 26.78 ;
    RECT 203.6 27.07 203.81 27.14 ;
    RECT 203.6 27.43 203.81 27.5 ;
    RECT 203.14 26.71 203.35 26.78 ;
    RECT 203.14 27.07 203.35 27.14 ;
    RECT 203.14 27.43 203.35 27.5 ;
    RECT 200.28 26.71 200.49 26.78 ;
    RECT 200.28 27.07 200.49 27.14 ;
    RECT 200.28 27.43 200.49 27.5 ;
    RECT 199.82 26.71 200.03 26.78 ;
    RECT 199.82 27.07 200.03 27.14 ;
    RECT 199.82 27.43 200.03 27.5 ;
    RECT 196.96 26.71 197.17 26.78 ;
    RECT 196.96 27.07 197.17 27.14 ;
    RECT 196.96 27.43 197.17 27.5 ;
    RECT 196.5 26.71 196.71 26.78 ;
    RECT 196.5 27.07 196.71 27.14 ;
    RECT 196.5 27.43 196.71 27.5 ;
    RECT 193.64 26.71 193.85 26.78 ;
    RECT 193.64 27.07 193.85 27.14 ;
    RECT 193.64 27.43 193.85 27.5 ;
    RECT 193.18 26.71 193.39 26.78 ;
    RECT 193.18 27.07 193.39 27.14 ;
    RECT 193.18 27.43 193.39 27.5 ;
    RECT 190.32 26.71 190.53 26.78 ;
    RECT 190.32 27.07 190.53 27.14 ;
    RECT 190.32 27.43 190.53 27.5 ;
    RECT 189.86 26.71 190.07 26.78 ;
    RECT 189.86 27.07 190.07 27.14 ;
    RECT 189.86 27.43 190.07 27.5 ;
    RECT 187.0 26.71 187.21 26.78 ;
    RECT 187.0 27.07 187.21 27.14 ;
    RECT 187.0 27.43 187.21 27.5 ;
    RECT 186.54 26.71 186.75 26.78 ;
    RECT 186.54 27.07 186.75 27.14 ;
    RECT 186.54 27.43 186.75 27.5 ;
    RECT 183.68 26.71 183.89 26.78 ;
    RECT 183.68 27.07 183.89 27.14 ;
    RECT 183.68 27.43 183.89 27.5 ;
    RECT 183.22 26.71 183.43 26.78 ;
    RECT 183.22 27.07 183.43 27.14 ;
    RECT 183.22 27.43 183.43 27.5 ;
    RECT 147.485 27.07 147.555 27.14 ;
    RECT 266.68 26.71 266.89 26.78 ;
    RECT 266.68 27.07 266.89 27.14 ;
    RECT 266.68 27.43 266.89 27.5 ;
    RECT 266.22 26.71 266.43 26.78 ;
    RECT 266.22 27.07 266.43 27.14 ;
    RECT 266.22 27.43 266.43 27.5 ;
    RECT 263.36 26.71 263.57 26.78 ;
    RECT 263.36 27.07 263.57 27.14 ;
    RECT 263.36 27.43 263.57 27.5 ;
    RECT 262.9 26.71 263.11 26.78 ;
    RECT 262.9 27.07 263.11 27.14 ;
    RECT 262.9 27.43 263.11 27.5 ;
    RECT 260.04 26.71 260.25 26.78 ;
    RECT 260.04 27.07 260.25 27.14 ;
    RECT 260.04 27.43 260.25 27.5 ;
    RECT 259.58 26.71 259.79 26.78 ;
    RECT 259.58 27.07 259.79 27.14 ;
    RECT 259.58 27.43 259.79 27.5 ;
    RECT 256.72 26.71 256.93 26.78 ;
    RECT 256.72 27.07 256.93 27.14 ;
    RECT 256.72 27.43 256.93 27.5 ;
    RECT 256.26 26.71 256.47 26.78 ;
    RECT 256.26 27.07 256.47 27.14 ;
    RECT 256.26 27.43 256.47 27.5 ;
    RECT 253.4 26.71 253.61 26.78 ;
    RECT 253.4 27.07 253.61 27.14 ;
    RECT 253.4 27.43 253.61 27.5 ;
    RECT 252.94 26.71 253.15 26.78 ;
    RECT 252.94 27.07 253.15 27.14 ;
    RECT 252.94 27.43 253.15 27.5 ;
    RECT 250.08 25.99 250.29 26.06 ;
    RECT 250.08 26.35 250.29 26.42 ;
    RECT 250.08 26.71 250.29 26.78 ;
    RECT 249.62 25.99 249.83 26.06 ;
    RECT 249.62 26.35 249.83 26.42 ;
    RECT 249.62 26.71 249.83 26.78 ;
    RECT 246.76 25.99 246.97 26.06 ;
    RECT 246.76 26.35 246.97 26.42 ;
    RECT 246.76 26.71 246.97 26.78 ;
    RECT 246.3 25.99 246.51 26.06 ;
    RECT 246.3 26.35 246.51 26.42 ;
    RECT 246.3 26.71 246.51 26.78 ;
    RECT 243.44 25.99 243.65 26.06 ;
    RECT 243.44 26.35 243.65 26.42 ;
    RECT 243.44 26.71 243.65 26.78 ;
    RECT 242.98 25.99 243.19 26.06 ;
    RECT 242.98 26.35 243.19 26.42 ;
    RECT 242.98 26.71 243.19 26.78 ;
    RECT 240.12 25.99 240.33 26.06 ;
    RECT 240.12 26.35 240.33 26.42 ;
    RECT 240.12 26.71 240.33 26.78 ;
    RECT 239.66 25.99 239.87 26.06 ;
    RECT 239.66 26.35 239.87 26.42 ;
    RECT 239.66 26.71 239.87 26.78 ;
    RECT 236.8 25.99 237.01 26.06 ;
    RECT 236.8 26.35 237.01 26.42 ;
    RECT 236.8 26.71 237.01 26.78 ;
    RECT 236.34 25.99 236.55 26.06 ;
    RECT 236.34 26.35 236.55 26.42 ;
    RECT 236.34 26.71 236.55 26.78 ;
    RECT 233.48 25.99 233.69 26.06 ;
    RECT 233.48 26.35 233.69 26.42 ;
    RECT 233.48 26.71 233.69 26.78 ;
    RECT 233.02 25.99 233.23 26.06 ;
    RECT 233.02 26.35 233.23 26.42 ;
    RECT 233.02 26.71 233.23 26.78 ;
    RECT 230.16 25.99 230.37 26.06 ;
    RECT 230.16 26.35 230.37 26.42 ;
    RECT 230.16 26.71 230.37 26.78 ;
    RECT 229.7 25.99 229.91 26.06 ;
    RECT 229.7 26.35 229.91 26.42 ;
    RECT 229.7 26.71 229.91 26.78 ;
    RECT 226.84 25.99 227.05 26.06 ;
    RECT 226.84 26.35 227.05 26.42 ;
    RECT 226.84 26.71 227.05 26.78 ;
    RECT 226.38 25.99 226.59 26.06 ;
    RECT 226.38 26.35 226.59 26.42 ;
    RECT 226.38 26.71 226.59 26.78 ;
    RECT 223.52 25.99 223.73 26.06 ;
    RECT 223.52 26.35 223.73 26.42 ;
    RECT 223.52 26.71 223.73 26.78 ;
    RECT 223.06 25.99 223.27 26.06 ;
    RECT 223.06 26.35 223.27 26.42 ;
    RECT 223.06 26.71 223.27 26.78 ;
    RECT 220.2 25.99 220.41 26.06 ;
    RECT 220.2 26.35 220.41 26.42 ;
    RECT 220.2 26.71 220.41 26.78 ;
    RECT 219.74 25.99 219.95 26.06 ;
    RECT 219.74 26.35 219.95 26.42 ;
    RECT 219.74 26.71 219.95 26.78 ;
    RECT 216.88 25.99 217.09 26.06 ;
    RECT 216.88 26.35 217.09 26.42 ;
    RECT 216.88 26.71 217.09 26.78 ;
    RECT 216.42 25.99 216.63 26.06 ;
    RECT 216.42 26.35 216.63 26.42 ;
    RECT 216.42 26.71 216.63 26.78 ;
    RECT 267.91 26.35 267.98 26.42 ;
    RECT 180.36 25.99 180.57 26.06 ;
    RECT 180.36 26.35 180.57 26.42 ;
    RECT 180.36 26.71 180.57 26.78 ;
    RECT 179.9 25.99 180.11 26.06 ;
    RECT 179.9 26.35 180.11 26.42 ;
    RECT 179.9 26.71 180.11 26.78 ;
    RECT 177.04 25.99 177.25 26.06 ;
    RECT 177.04 26.35 177.25 26.42 ;
    RECT 177.04 26.71 177.25 26.78 ;
    RECT 176.58 25.99 176.79 26.06 ;
    RECT 176.58 26.35 176.79 26.42 ;
    RECT 176.58 26.71 176.79 26.78 ;
    RECT 173.72 25.99 173.93 26.06 ;
    RECT 173.72 26.35 173.93 26.42 ;
    RECT 173.72 26.71 173.93 26.78 ;
    RECT 173.26 25.99 173.47 26.06 ;
    RECT 173.26 26.35 173.47 26.42 ;
    RECT 173.26 26.71 173.47 26.78 ;
    RECT 170.4 25.99 170.61 26.06 ;
    RECT 170.4 26.35 170.61 26.42 ;
    RECT 170.4 26.71 170.61 26.78 ;
    RECT 169.94 25.99 170.15 26.06 ;
    RECT 169.94 26.35 170.15 26.42 ;
    RECT 169.94 26.71 170.15 26.78 ;
    RECT 167.08 25.99 167.29 26.06 ;
    RECT 167.08 26.35 167.29 26.42 ;
    RECT 167.08 26.71 167.29 26.78 ;
    RECT 166.62 25.99 166.83 26.06 ;
    RECT 166.62 26.35 166.83 26.42 ;
    RECT 166.62 26.71 166.83 26.78 ;
    RECT 163.76 25.99 163.97 26.06 ;
    RECT 163.76 26.35 163.97 26.42 ;
    RECT 163.76 26.71 163.97 26.78 ;
    RECT 163.3 25.99 163.51 26.06 ;
    RECT 163.3 26.35 163.51 26.42 ;
    RECT 163.3 26.71 163.51 26.78 ;
    RECT 160.44 25.99 160.65 26.06 ;
    RECT 160.44 26.35 160.65 26.42 ;
    RECT 160.44 26.71 160.65 26.78 ;
    RECT 159.98 25.99 160.19 26.06 ;
    RECT 159.98 26.35 160.19 26.42 ;
    RECT 159.98 26.71 160.19 26.78 ;
    RECT 157.12 25.99 157.33 26.06 ;
    RECT 157.12 26.35 157.33 26.42 ;
    RECT 157.12 26.71 157.33 26.78 ;
    RECT 156.66 25.99 156.87 26.06 ;
    RECT 156.66 26.35 156.87 26.42 ;
    RECT 156.66 26.71 156.87 26.78 ;
    RECT 153.8 25.99 154.01 26.06 ;
    RECT 153.8 26.35 154.01 26.42 ;
    RECT 153.8 26.71 154.01 26.78 ;
    RECT 153.34 25.99 153.55 26.06 ;
    RECT 153.34 26.35 153.55 26.42 ;
    RECT 153.34 26.71 153.55 26.78 ;
    RECT 150.48 25.99 150.69 26.06 ;
    RECT 150.48 26.35 150.69 26.42 ;
    RECT 150.48 26.71 150.69 26.78 ;
    RECT 150.02 25.99 150.23 26.06 ;
    RECT 150.02 26.35 150.23 26.42 ;
    RECT 150.02 26.71 150.23 26.78 ;
    RECT 213.56 25.99 213.77 26.06 ;
    RECT 213.56 26.35 213.77 26.42 ;
    RECT 213.56 26.71 213.77 26.78 ;
    RECT 213.1 25.99 213.31 26.06 ;
    RECT 213.1 26.35 213.31 26.42 ;
    RECT 213.1 26.71 213.31 26.78 ;
    RECT 210.24 25.99 210.45 26.06 ;
    RECT 210.24 26.35 210.45 26.42 ;
    RECT 210.24 26.71 210.45 26.78 ;
    RECT 209.78 25.99 209.99 26.06 ;
    RECT 209.78 26.35 209.99 26.42 ;
    RECT 209.78 26.71 209.99 26.78 ;
    RECT 206.92 25.99 207.13 26.06 ;
    RECT 206.92 26.35 207.13 26.42 ;
    RECT 206.92 26.71 207.13 26.78 ;
    RECT 206.46 25.99 206.67 26.06 ;
    RECT 206.46 26.35 206.67 26.42 ;
    RECT 206.46 26.71 206.67 26.78 ;
    RECT 203.6 25.99 203.81 26.06 ;
    RECT 203.6 26.35 203.81 26.42 ;
    RECT 203.6 26.71 203.81 26.78 ;
    RECT 203.14 25.99 203.35 26.06 ;
    RECT 203.14 26.35 203.35 26.42 ;
    RECT 203.14 26.71 203.35 26.78 ;
    RECT 200.28 25.99 200.49 26.06 ;
    RECT 200.28 26.35 200.49 26.42 ;
    RECT 200.28 26.71 200.49 26.78 ;
    RECT 199.82 25.99 200.03 26.06 ;
    RECT 199.82 26.35 200.03 26.42 ;
    RECT 199.82 26.71 200.03 26.78 ;
    RECT 196.96 25.99 197.17 26.06 ;
    RECT 196.96 26.35 197.17 26.42 ;
    RECT 196.96 26.71 197.17 26.78 ;
    RECT 196.5 25.99 196.71 26.06 ;
    RECT 196.5 26.35 196.71 26.42 ;
    RECT 196.5 26.71 196.71 26.78 ;
    RECT 193.64 25.99 193.85 26.06 ;
    RECT 193.64 26.35 193.85 26.42 ;
    RECT 193.64 26.71 193.85 26.78 ;
    RECT 193.18 25.99 193.39 26.06 ;
    RECT 193.18 26.35 193.39 26.42 ;
    RECT 193.18 26.71 193.39 26.78 ;
    RECT 190.32 25.99 190.53 26.06 ;
    RECT 190.32 26.35 190.53 26.42 ;
    RECT 190.32 26.71 190.53 26.78 ;
    RECT 189.86 25.99 190.07 26.06 ;
    RECT 189.86 26.35 190.07 26.42 ;
    RECT 189.86 26.71 190.07 26.78 ;
    RECT 187.0 25.99 187.21 26.06 ;
    RECT 187.0 26.35 187.21 26.42 ;
    RECT 187.0 26.71 187.21 26.78 ;
    RECT 186.54 25.99 186.75 26.06 ;
    RECT 186.54 26.35 186.75 26.42 ;
    RECT 186.54 26.71 186.75 26.78 ;
    RECT 183.68 25.99 183.89 26.06 ;
    RECT 183.68 26.35 183.89 26.42 ;
    RECT 183.68 26.71 183.89 26.78 ;
    RECT 183.22 25.99 183.43 26.06 ;
    RECT 183.22 26.35 183.43 26.42 ;
    RECT 183.22 26.71 183.43 26.78 ;
    RECT 147.485 26.35 147.555 26.42 ;
    RECT 266.68 25.99 266.89 26.06 ;
    RECT 266.68 26.35 266.89 26.42 ;
    RECT 266.68 26.71 266.89 26.78 ;
    RECT 266.22 25.99 266.43 26.06 ;
    RECT 266.22 26.35 266.43 26.42 ;
    RECT 266.22 26.71 266.43 26.78 ;
    RECT 263.36 25.99 263.57 26.06 ;
    RECT 263.36 26.35 263.57 26.42 ;
    RECT 263.36 26.71 263.57 26.78 ;
    RECT 262.9 25.99 263.11 26.06 ;
    RECT 262.9 26.35 263.11 26.42 ;
    RECT 262.9 26.71 263.11 26.78 ;
    RECT 260.04 25.99 260.25 26.06 ;
    RECT 260.04 26.35 260.25 26.42 ;
    RECT 260.04 26.71 260.25 26.78 ;
    RECT 259.58 25.99 259.79 26.06 ;
    RECT 259.58 26.35 259.79 26.42 ;
    RECT 259.58 26.71 259.79 26.78 ;
    RECT 256.72 25.99 256.93 26.06 ;
    RECT 256.72 26.35 256.93 26.42 ;
    RECT 256.72 26.71 256.93 26.78 ;
    RECT 256.26 25.99 256.47 26.06 ;
    RECT 256.26 26.35 256.47 26.42 ;
    RECT 256.26 26.71 256.47 26.78 ;
    RECT 253.4 25.99 253.61 26.06 ;
    RECT 253.4 26.35 253.61 26.42 ;
    RECT 253.4 26.71 253.61 26.78 ;
    RECT 252.94 25.99 253.15 26.06 ;
    RECT 252.94 26.35 253.15 26.42 ;
    RECT 252.94 26.71 253.15 26.78 ;
    RECT 250.08 25.27 250.29 25.34 ;
    RECT 250.08 25.63 250.29 25.7 ;
    RECT 250.08 25.99 250.29 26.06 ;
    RECT 249.62 25.27 249.83 25.34 ;
    RECT 249.62 25.63 249.83 25.7 ;
    RECT 249.62 25.99 249.83 26.06 ;
    RECT 246.76 25.27 246.97 25.34 ;
    RECT 246.76 25.63 246.97 25.7 ;
    RECT 246.76 25.99 246.97 26.06 ;
    RECT 246.3 25.27 246.51 25.34 ;
    RECT 246.3 25.63 246.51 25.7 ;
    RECT 246.3 25.99 246.51 26.06 ;
    RECT 243.44 25.27 243.65 25.34 ;
    RECT 243.44 25.63 243.65 25.7 ;
    RECT 243.44 25.99 243.65 26.06 ;
    RECT 242.98 25.27 243.19 25.34 ;
    RECT 242.98 25.63 243.19 25.7 ;
    RECT 242.98 25.99 243.19 26.06 ;
    RECT 240.12 25.27 240.33 25.34 ;
    RECT 240.12 25.63 240.33 25.7 ;
    RECT 240.12 25.99 240.33 26.06 ;
    RECT 239.66 25.27 239.87 25.34 ;
    RECT 239.66 25.63 239.87 25.7 ;
    RECT 239.66 25.99 239.87 26.06 ;
    RECT 236.8 25.27 237.01 25.34 ;
    RECT 236.8 25.63 237.01 25.7 ;
    RECT 236.8 25.99 237.01 26.06 ;
    RECT 236.34 25.27 236.55 25.34 ;
    RECT 236.34 25.63 236.55 25.7 ;
    RECT 236.34 25.99 236.55 26.06 ;
    RECT 233.48 25.27 233.69 25.34 ;
    RECT 233.48 25.63 233.69 25.7 ;
    RECT 233.48 25.99 233.69 26.06 ;
    RECT 233.02 25.27 233.23 25.34 ;
    RECT 233.02 25.63 233.23 25.7 ;
    RECT 233.02 25.99 233.23 26.06 ;
    RECT 230.16 25.27 230.37 25.34 ;
    RECT 230.16 25.63 230.37 25.7 ;
    RECT 230.16 25.99 230.37 26.06 ;
    RECT 229.7 25.27 229.91 25.34 ;
    RECT 229.7 25.63 229.91 25.7 ;
    RECT 229.7 25.99 229.91 26.06 ;
    RECT 226.84 25.27 227.05 25.34 ;
    RECT 226.84 25.63 227.05 25.7 ;
    RECT 226.84 25.99 227.05 26.06 ;
    RECT 226.38 25.27 226.59 25.34 ;
    RECT 226.38 25.63 226.59 25.7 ;
    RECT 226.38 25.99 226.59 26.06 ;
    RECT 223.52 25.27 223.73 25.34 ;
    RECT 223.52 25.63 223.73 25.7 ;
    RECT 223.52 25.99 223.73 26.06 ;
    RECT 223.06 25.27 223.27 25.34 ;
    RECT 223.06 25.63 223.27 25.7 ;
    RECT 223.06 25.99 223.27 26.06 ;
    RECT 220.2 25.27 220.41 25.34 ;
    RECT 220.2 25.63 220.41 25.7 ;
    RECT 220.2 25.99 220.41 26.06 ;
    RECT 219.74 25.27 219.95 25.34 ;
    RECT 219.74 25.63 219.95 25.7 ;
    RECT 219.74 25.99 219.95 26.06 ;
    RECT 216.88 25.27 217.09 25.34 ;
    RECT 216.88 25.63 217.09 25.7 ;
    RECT 216.88 25.99 217.09 26.06 ;
    RECT 216.42 25.27 216.63 25.34 ;
    RECT 216.42 25.63 216.63 25.7 ;
    RECT 216.42 25.99 216.63 26.06 ;
    RECT 267.91 25.63 267.98 25.7 ;
    RECT 180.36 25.27 180.57 25.34 ;
    RECT 180.36 25.63 180.57 25.7 ;
    RECT 180.36 25.99 180.57 26.06 ;
    RECT 179.9 25.27 180.11 25.34 ;
    RECT 179.9 25.63 180.11 25.7 ;
    RECT 179.9 25.99 180.11 26.06 ;
    RECT 177.04 25.27 177.25 25.34 ;
    RECT 177.04 25.63 177.25 25.7 ;
    RECT 177.04 25.99 177.25 26.06 ;
    RECT 176.58 25.27 176.79 25.34 ;
    RECT 176.58 25.63 176.79 25.7 ;
    RECT 176.58 25.99 176.79 26.06 ;
    RECT 173.72 25.27 173.93 25.34 ;
    RECT 173.72 25.63 173.93 25.7 ;
    RECT 173.72 25.99 173.93 26.06 ;
    RECT 173.26 25.27 173.47 25.34 ;
    RECT 173.26 25.63 173.47 25.7 ;
    RECT 173.26 25.99 173.47 26.06 ;
    RECT 170.4 25.27 170.61 25.34 ;
    RECT 170.4 25.63 170.61 25.7 ;
    RECT 170.4 25.99 170.61 26.06 ;
    RECT 169.94 25.27 170.15 25.34 ;
    RECT 169.94 25.63 170.15 25.7 ;
    RECT 169.94 25.99 170.15 26.06 ;
    RECT 167.08 25.27 167.29 25.34 ;
    RECT 167.08 25.63 167.29 25.7 ;
    RECT 167.08 25.99 167.29 26.06 ;
    RECT 166.62 25.27 166.83 25.34 ;
    RECT 166.62 25.63 166.83 25.7 ;
    RECT 166.62 25.99 166.83 26.06 ;
    RECT 163.76 25.27 163.97 25.34 ;
    RECT 163.76 25.63 163.97 25.7 ;
    RECT 163.76 25.99 163.97 26.06 ;
    RECT 163.3 25.27 163.51 25.34 ;
    RECT 163.3 25.63 163.51 25.7 ;
    RECT 163.3 25.99 163.51 26.06 ;
    RECT 160.44 25.27 160.65 25.34 ;
    RECT 160.44 25.63 160.65 25.7 ;
    RECT 160.44 25.99 160.65 26.06 ;
    RECT 159.98 25.27 160.19 25.34 ;
    RECT 159.98 25.63 160.19 25.7 ;
    RECT 159.98 25.99 160.19 26.06 ;
    RECT 157.12 25.27 157.33 25.34 ;
    RECT 157.12 25.63 157.33 25.7 ;
    RECT 157.12 25.99 157.33 26.06 ;
    RECT 156.66 25.27 156.87 25.34 ;
    RECT 156.66 25.63 156.87 25.7 ;
    RECT 156.66 25.99 156.87 26.06 ;
    RECT 153.8 25.27 154.01 25.34 ;
    RECT 153.8 25.63 154.01 25.7 ;
    RECT 153.8 25.99 154.01 26.06 ;
    RECT 153.34 25.27 153.55 25.34 ;
    RECT 153.34 25.63 153.55 25.7 ;
    RECT 153.34 25.99 153.55 26.06 ;
    RECT 150.48 25.27 150.69 25.34 ;
    RECT 150.48 25.63 150.69 25.7 ;
    RECT 150.48 25.99 150.69 26.06 ;
    RECT 150.02 25.27 150.23 25.34 ;
    RECT 150.02 25.63 150.23 25.7 ;
    RECT 150.02 25.99 150.23 26.06 ;
    RECT 213.56 25.27 213.77 25.34 ;
    RECT 213.56 25.63 213.77 25.7 ;
    RECT 213.56 25.99 213.77 26.06 ;
    RECT 213.1 25.27 213.31 25.34 ;
    RECT 213.1 25.63 213.31 25.7 ;
    RECT 213.1 25.99 213.31 26.06 ;
    RECT 210.24 25.27 210.45 25.34 ;
    RECT 210.24 25.63 210.45 25.7 ;
    RECT 210.24 25.99 210.45 26.06 ;
    RECT 209.78 25.27 209.99 25.34 ;
    RECT 209.78 25.63 209.99 25.7 ;
    RECT 209.78 25.99 209.99 26.06 ;
    RECT 206.92 25.27 207.13 25.34 ;
    RECT 206.92 25.63 207.13 25.7 ;
    RECT 206.92 25.99 207.13 26.06 ;
    RECT 206.46 25.27 206.67 25.34 ;
    RECT 206.46 25.63 206.67 25.7 ;
    RECT 206.46 25.99 206.67 26.06 ;
    RECT 203.6 25.27 203.81 25.34 ;
    RECT 203.6 25.63 203.81 25.7 ;
    RECT 203.6 25.99 203.81 26.06 ;
    RECT 203.14 25.27 203.35 25.34 ;
    RECT 203.14 25.63 203.35 25.7 ;
    RECT 203.14 25.99 203.35 26.06 ;
    RECT 200.28 25.27 200.49 25.34 ;
    RECT 200.28 25.63 200.49 25.7 ;
    RECT 200.28 25.99 200.49 26.06 ;
    RECT 199.82 25.27 200.03 25.34 ;
    RECT 199.82 25.63 200.03 25.7 ;
    RECT 199.82 25.99 200.03 26.06 ;
    RECT 196.96 25.27 197.17 25.34 ;
    RECT 196.96 25.63 197.17 25.7 ;
    RECT 196.96 25.99 197.17 26.06 ;
    RECT 196.5 25.27 196.71 25.34 ;
    RECT 196.5 25.63 196.71 25.7 ;
    RECT 196.5 25.99 196.71 26.06 ;
    RECT 193.64 25.27 193.85 25.34 ;
    RECT 193.64 25.63 193.85 25.7 ;
    RECT 193.64 25.99 193.85 26.06 ;
    RECT 193.18 25.27 193.39 25.34 ;
    RECT 193.18 25.63 193.39 25.7 ;
    RECT 193.18 25.99 193.39 26.06 ;
    RECT 190.32 25.27 190.53 25.34 ;
    RECT 190.32 25.63 190.53 25.7 ;
    RECT 190.32 25.99 190.53 26.06 ;
    RECT 189.86 25.27 190.07 25.34 ;
    RECT 189.86 25.63 190.07 25.7 ;
    RECT 189.86 25.99 190.07 26.06 ;
    RECT 187.0 25.27 187.21 25.34 ;
    RECT 187.0 25.63 187.21 25.7 ;
    RECT 187.0 25.99 187.21 26.06 ;
    RECT 186.54 25.27 186.75 25.34 ;
    RECT 186.54 25.63 186.75 25.7 ;
    RECT 186.54 25.99 186.75 26.06 ;
    RECT 183.68 25.27 183.89 25.34 ;
    RECT 183.68 25.63 183.89 25.7 ;
    RECT 183.68 25.99 183.89 26.06 ;
    RECT 183.22 25.27 183.43 25.34 ;
    RECT 183.22 25.63 183.43 25.7 ;
    RECT 183.22 25.99 183.43 26.06 ;
    RECT 147.485 25.63 147.555 25.7 ;
    RECT 266.68 25.27 266.89 25.34 ;
    RECT 266.68 25.63 266.89 25.7 ;
    RECT 266.68 25.99 266.89 26.06 ;
    RECT 266.22 25.27 266.43 25.34 ;
    RECT 266.22 25.63 266.43 25.7 ;
    RECT 266.22 25.99 266.43 26.06 ;
    RECT 263.36 25.27 263.57 25.34 ;
    RECT 263.36 25.63 263.57 25.7 ;
    RECT 263.36 25.99 263.57 26.06 ;
    RECT 262.9 25.27 263.11 25.34 ;
    RECT 262.9 25.63 263.11 25.7 ;
    RECT 262.9 25.99 263.11 26.06 ;
    RECT 260.04 25.27 260.25 25.34 ;
    RECT 260.04 25.63 260.25 25.7 ;
    RECT 260.04 25.99 260.25 26.06 ;
    RECT 259.58 25.27 259.79 25.34 ;
    RECT 259.58 25.63 259.79 25.7 ;
    RECT 259.58 25.99 259.79 26.06 ;
    RECT 256.72 25.27 256.93 25.34 ;
    RECT 256.72 25.63 256.93 25.7 ;
    RECT 256.72 25.99 256.93 26.06 ;
    RECT 256.26 25.27 256.47 25.34 ;
    RECT 256.26 25.63 256.47 25.7 ;
    RECT 256.26 25.99 256.47 26.06 ;
    RECT 253.4 25.27 253.61 25.34 ;
    RECT 253.4 25.63 253.61 25.7 ;
    RECT 253.4 25.99 253.61 26.06 ;
    RECT 252.94 25.27 253.15 25.34 ;
    RECT 252.94 25.63 253.15 25.7 ;
    RECT 252.94 25.99 253.15 26.06 ;
    RECT 250.08 64.89 250.29 64.96 ;
    RECT 250.08 65.25 250.29 65.32 ;
    RECT 250.08 65.61 250.29 65.68 ;
    RECT 249.62 64.89 249.83 64.96 ;
    RECT 249.62 65.25 249.83 65.32 ;
    RECT 249.62 65.61 249.83 65.68 ;
    RECT 246.76 64.89 246.97 64.96 ;
    RECT 246.76 65.25 246.97 65.32 ;
    RECT 246.76 65.61 246.97 65.68 ;
    RECT 246.3 64.89 246.51 64.96 ;
    RECT 246.3 65.25 246.51 65.32 ;
    RECT 246.3 65.61 246.51 65.68 ;
    RECT 243.44 64.89 243.65 64.96 ;
    RECT 243.44 65.25 243.65 65.32 ;
    RECT 243.44 65.61 243.65 65.68 ;
    RECT 242.98 64.89 243.19 64.96 ;
    RECT 242.98 65.25 243.19 65.32 ;
    RECT 242.98 65.61 243.19 65.68 ;
    RECT 240.12 64.89 240.33 64.96 ;
    RECT 240.12 65.25 240.33 65.32 ;
    RECT 240.12 65.61 240.33 65.68 ;
    RECT 239.66 64.89 239.87 64.96 ;
    RECT 239.66 65.25 239.87 65.32 ;
    RECT 239.66 65.61 239.87 65.68 ;
    RECT 236.8 64.89 237.01 64.96 ;
    RECT 236.8 65.25 237.01 65.32 ;
    RECT 236.8 65.61 237.01 65.68 ;
    RECT 236.34 64.89 236.55 64.96 ;
    RECT 236.34 65.25 236.55 65.32 ;
    RECT 236.34 65.61 236.55 65.68 ;
    RECT 233.48 64.89 233.69 64.96 ;
    RECT 233.48 65.25 233.69 65.32 ;
    RECT 233.48 65.61 233.69 65.68 ;
    RECT 233.02 64.89 233.23 64.96 ;
    RECT 233.02 65.25 233.23 65.32 ;
    RECT 233.02 65.61 233.23 65.68 ;
    RECT 230.16 64.89 230.37 64.96 ;
    RECT 230.16 65.25 230.37 65.32 ;
    RECT 230.16 65.61 230.37 65.68 ;
    RECT 229.7 64.89 229.91 64.96 ;
    RECT 229.7 65.25 229.91 65.32 ;
    RECT 229.7 65.61 229.91 65.68 ;
    RECT 226.84 64.89 227.05 64.96 ;
    RECT 226.84 65.25 227.05 65.32 ;
    RECT 226.84 65.61 227.05 65.68 ;
    RECT 226.38 64.89 226.59 64.96 ;
    RECT 226.38 65.25 226.59 65.32 ;
    RECT 226.38 65.61 226.59 65.68 ;
    RECT 223.52 64.89 223.73 64.96 ;
    RECT 223.52 65.25 223.73 65.32 ;
    RECT 223.52 65.61 223.73 65.68 ;
    RECT 223.06 64.89 223.27 64.96 ;
    RECT 223.06 65.25 223.27 65.32 ;
    RECT 223.06 65.61 223.27 65.68 ;
    RECT 220.2 64.89 220.41 64.96 ;
    RECT 220.2 65.25 220.41 65.32 ;
    RECT 220.2 65.61 220.41 65.68 ;
    RECT 219.74 64.89 219.95 64.96 ;
    RECT 219.74 65.25 219.95 65.32 ;
    RECT 219.74 65.61 219.95 65.68 ;
    RECT 216.88 64.89 217.09 64.96 ;
    RECT 216.88 65.25 217.09 65.32 ;
    RECT 216.88 65.61 217.09 65.68 ;
    RECT 216.42 64.89 216.63 64.96 ;
    RECT 216.42 65.25 216.63 65.32 ;
    RECT 216.42 65.61 216.63 65.68 ;
    RECT 267.91 65.25 267.98 65.32 ;
    RECT 180.36 64.89 180.57 64.96 ;
    RECT 180.36 65.25 180.57 65.32 ;
    RECT 180.36 65.61 180.57 65.68 ;
    RECT 179.9 64.89 180.11 64.96 ;
    RECT 179.9 65.25 180.11 65.32 ;
    RECT 179.9 65.61 180.11 65.68 ;
    RECT 177.04 64.89 177.25 64.96 ;
    RECT 177.04 65.25 177.25 65.32 ;
    RECT 177.04 65.61 177.25 65.68 ;
    RECT 176.58 64.89 176.79 64.96 ;
    RECT 176.58 65.25 176.79 65.32 ;
    RECT 176.58 65.61 176.79 65.68 ;
    RECT 173.72 64.89 173.93 64.96 ;
    RECT 173.72 65.25 173.93 65.32 ;
    RECT 173.72 65.61 173.93 65.68 ;
    RECT 173.26 64.89 173.47 64.96 ;
    RECT 173.26 65.25 173.47 65.32 ;
    RECT 173.26 65.61 173.47 65.68 ;
    RECT 170.4 64.89 170.61 64.96 ;
    RECT 170.4 65.25 170.61 65.32 ;
    RECT 170.4 65.61 170.61 65.68 ;
    RECT 169.94 64.89 170.15 64.96 ;
    RECT 169.94 65.25 170.15 65.32 ;
    RECT 169.94 65.61 170.15 65.68 ;
    RECT 167.08 64.89 167.29 64.96 ;
    RECT 167.08 65.25 167.29 65.32 ;
    RECT 167.08 65.61 167.29 65.68 ;
    RECT 166.62 64.89 166.83 64.96 ;
    RECT 166.62 65.25 166.83 65.32 ;
    RECT 166.62 65.61 166.83 65.68 ;
    RECT 163.76 64.89 163.97 64.96 ;
    RECT 163.76 65.25 163.97 65.32 ;
    RECT 163.76 65.61 163.97 65.68 ;
    RECT 163.3 64.89 163.51 64.96 ;
    RECT 163.3 65.25 163.51 65.32 ;
    RECT 163.3 65.61 163.51 65.68 ;
    RECT 160.44 64.89 160.65 64.96 ;
    RECT 160.44 65.25 160.65 65.32 ;
    RECT 160.44 65.61 160.65 65.68 ;
    RECT 159.98 64.89 160.19 64.96 ;
    RECT 159.98 65.25 160.19 65.32 ;
    RECT 159.98 65.61 160.19 65.68 ;
    RECT 157.12 64.89 157.33 64.96 ;
    RECT 157.12 65.25 157.33 65.32 ;
    RECT 157.12 65.61 157.33 65.68 ;
    RECT 156.66 64.89 156.87 64.96 ;
    RECT 156.66 65.25 156.87 65.32 ;
    RECT 156.66 65.61 156.87 65.68 ;
    RECT 153.8 64.89 154.01 64.96 ;
    RECT 153.8 65.25 154.01 65.32 ;
    RECT 153.8 65.61 154.01 65.68 ;
    RECT 153.34 64.89 153.55 64.96 ;
    RECT 153.34 65.25 153.55 65.32 ;
    RECT 153.34 65.61 153.55 65.68 ;
    RECT 150.48 64.89 150.69 64.96 ;
    RECT 150.48 65.25 150.69 65.32 ;
    RECT 150.48 65.61 150.69 65.68 ;
    RECT 150.02 64.89 150.23 64.96 ;
    RECT 150.02 65.25 150.23 65.32 ;
    RECT 150.02 65.61 150.23 65.68 ;
    RECT 213.56 64.89 213.77 64.96 ;
    RECT 213.56 65.25 213.77 65.32 ;
    RECT 213.56 65.61 213.77 65.68 ;
    RECT 213.1 64.89 213.31 64.96 ;
    RECT 213.1 65.25 213.31 65.32 ;
    RECT 213.1 65.61 213.31 65.68 ;
    RECT 210.24 64.89 210.45 64.96 ;
    RECT 210.24 65.25 210.45 65.32 ;
    RECT 210.24 65.61 210.45 65.68 ;
    RECT 209.78 64.89 209.99 64.96 ;
    RECT 209.78 65.25 209.99 65.32 ;
    RECT 209.78 65.61 209.99 65.68 ;
    RECT 206.92 64.89 207.13 64.96 ;
    RECT 206.92 65.25 207.13 65.32 ;
    RECT 206.92 65.61 207.13 65.68 ;
    RECT 206.46 64.89 206.67 64.96 ;
    RECT 206.46 65.25 206.67 65.32 ;
    RECT 206.46 65.61 206.67 65.68 ;
    RECT 203.6 64.89 203.81 64.96 ;
    RECT 203.6 65.25 203.81 65.32 ;
    RECT 203.6 65.61 203.81 65.68 ;
    RECT 203.14 64.89 203.35 64.96 ;
    RECT 203.14 65.25 203.35 65.32 ;
    RECT 203.14 65.61 203.35 65.68 ;
    RECT 200.28 64.89 200.49 64.96 ;
    RECT 200.28 65.25 200.49 65.32 ;
    RECT 200.28 65.61 200.49 65.68 ;
    RECT 199.82 64.89 200.03 64.96 ;
    RECT 199.82 65.25 200.03 65.32 ;
    RECT 199.82 65.61 200.03 65.68 ;
    RECT 196.96 64.89 197.17 64.96 ;
    RECT 196.96 65.25 197.17 65.32 ;
    RECT 196.96 65.61 197.17 65.68 ;
    RECT 196.5 64.89 196.71 64.96 ;
    RECT 196.5 65.25 196.71 65.32 ;
    RECT 196.5 65.61 196.71 65.68 ;
    RECT 193.64 64.89 193.85 64.96 ;
    RECT 193.64 65.25 193.85 65.32 ;
    RECT 193.64 65.61 193.85 65.68 ;
    RECT 193.18 64.89 193.39 64.96 ;
    RECT 193.18 65.25 193.39 65.32 ;
    RECT 193.18 65.61 193.39 65.68 ;
    RECT 190.32 64.89 190.53 64.96 ;
    RECT 190.32 65.25 190.53 65.32 ;
    RECT 190.32 65.61 190.53 65.68 ;
    RECT 189.86 64.89 190.07 64.96 ;
    RECT 189.86 65.25 190.07 65.32 ;
    RECT 189.86 65.61 190.07 65.68 ;
    RECT 187.0 64.89 187.21 64.96 ;
    RECT 187.0 65.25 187.21 65.32 ;
    RECT 187.0 65.61 187.21 65.68 ;
    RECT 186.54 64.89 186.75 64.96 ;
    RECT 186.54 65.25 186.75 65.32 ;
    RECT 186.54 65.61 186.75 65.68 ;
    RECT 183.68 64.89 183.89 64.96 ;
    RECT 183.68 65.25 183.89 65.32 ;
    RECT 183.68 65.61 183.89 65.68 ;
    RECT 183.22 64.89 183.43 64.96 ;
    RECT 183.22 65.25 183.43 65.32 ;
    RECT 183.22 65.61 183.43 65.68 ;
    RECT 147.485 65.25 147.555 65.32 ;
    RECT 266.68 64.89 266.89 64.96 ;
    RECT 266.68 65.25 266.89 65.32 ;
    RECT 266.68 65.61 266.89 65.68 ;
    RECT 266.22 64.89 266.43 64.96 ;
    RECT 266.22 65.25 266.43 65.32 ;
    RECT 266.22 65.61 266.43 65.68 ;
    RECT 263.36 64.89 263.57 64.96 ;
    RECT 263.36 65.25 263.57 65.32 ;
    RECT 263.36 65.61 263.57 65.68 ;
    RECT 262.9 64.89 263.11 64.96 ;
    RECT 262.9 65.25 263.11 65.32 ;
    RECT 262.9 65.61 263.11 65.68 ;
    RECT 260.04 64.89 260.25 64.96 ;
    RECT 260.04 65.25 260.25 65.32 ;
    RECT 260.04 65.61 260.25 65.68 ;
    RECT 259.58 64.89 259.79 64.96 ;
    RECT 259.58 65.25 259.79 65.32 ;
    RECT 259.58 65.61 259.79 65.68 ;
    RECT 256.72 64.89 256.93 64.96 ;
    RECT 256.72 65.25 256.93 65.32 ;
    RECT 256.72 65.61 256.93 65.68 ;
    RECT 256.26 64.89 256.47 64.96 ;
    RECT 256.26 65.25 256.47 65.32 ;
    RECT 256.26 65.61 256.47 65.68 ;
    RECT 253.4 64.89 253.61 64.96 ;
    RECT 253.4 65.25 253.61 65.32 ;
    RECT 253.4 65.61 253.61 65.68 ;
    RECT 252.94 64.89 253.15 64.96 ;
    RECT 252.94 65.25 253.15 65.32 ;
    RECT 252.94 65.61 253.15 65.68 ;
    RECT 250.08 24.55 250.29 24.62 ;
    RECT 250.08 24.91 250.29 24.98 ;
    RECT 250.08 25.27 250.29 25.34 ;
    RECT 249.62 24.55 249.83 24.62 ;
    RECT 249.62 24.91 249.83 24.98 ;
    RECT 249.62 25.27 249.83 25.34 ;
    RECT 246.76 24.55 246.97 24.62 ;
    RECT 246.76 24.91 246.97 24.98 ;
    RECT 246.76 25.27 246.97 25.34 ;
    RECT 246.3 24.55 246.51 24.62 ;
    RECT 246.3 24.91 246.51 24.98 ;
    RECT 246.3 25.27 246.51 25.34 ;
    RECT 243.44 24.55 243.65 24.62 ;
    RECT 243.44 24.91 243.65 24.98 ;
    RECT 243.44 25.27 243.65 25.34 ;
    RECT 242.98 24.55 243.19 24.62 ;
    RECT 242.98 24.91 243.19 24.98 ;
    RECT 242.98 25.27 243.19 25.34 ;
    RECT 240.12 24.55 240.33 24.62 ;
    RECT 240.12 24.91 240.33 24.98 ;
    RECT 240.12 25.27 240.33 25.34 ;
    RECT 239.66 24.55 239.87 24.62 ;
    RECT 239.66 24.91 239.87 24.98 ;
    RECT 239.66 25.27 239.87 25.34 ;
    RECT 236.8 24.55 237.01 24.62 ;
    RECT 236.8 24.91 237.01 24.98 ;
    RECT 236.8 25.27 237.01 25.34 ;
    RECT 236.34 24.55 236.55 24.62 ;
    RECT 236.34 24.91 236.55 24.98 ;
    RECT 236.34 25.27 236.55 25.34 ;
    RECT 233.48 24.55 233.69 24.62 ;
    RECT 233.48 24.91 233.69 24.98 ;
    RECT 233.48 25.27 233.69 25.34 ;
    RECT 233.02 24.55 233.23 24.62 ;
    RECT 233.02 24.91 233.23 24.98 ;
    RECT 233.02 25.27 233.23 25.34 ;
    RECT 230.16 24.55 230.37 24.62 ;
    RECT 230.16 24.91 230.37 24.98 ;
    RECT 230.16 25.27 230.37 25.34 ;
    RECT 229.7 24.55 229.91 24.62 ;
    RECT 229.7 24.91 229.91 24.98 ;
    RECT 229.7 25.27 229.91 25.34 ;
    RECT 226.84 24.55 227.05 24.62 ;
    RECT 226.84 24.91 227.05 24.98 ;
    RECT 226.84 25.27 227.05 25.34 ;
    RECT 226.38 24.55 226.59 24.62 ;
    RECT 226.38 24.91 226.59 24.98 ;
    RECT 226.38 25.27 226.59 25.34 ;
    RECT 223.52 24.55 223.73 24.62 ;
    RECT 223.52 24.91 223.73 24.98 ;
    RECT 223.52 25.27 223.73 25.34 ;
    RECT 223.06 24.55 223.27 24.62 ;
    RECT 223.06 24.91 223.27 24.98 ;
    RECT 223.06 25.27 223.27 25.34 ;
    RECT 220.2 24.55 220.41 24.62 ;
    RECT 220.2 24.91 220.41 24.98 ;
    RECT 220.2 25.27 220.41 25.34 ;
    RECT 219.74 24.55 219.95 24.62 ;
    RECT 219.74 24.91 219.95 24.98 ;
    RECT 219.74 25.27 219.95 25.34 ;
    RECT 216.88 24.55 217.09 24.62 ;
    RECT 216.88 24.91 217.09 24.98 ;
    RECT 216.88 25.27 217.09 25.34 ;
    RECT 216.42 24.55 216.63 24.62 ;
    RECT 216.42 24.91 216.63 24.98 ;
    RECT 216.42 25.27 216.63 25.34 ;
    RECT 267.91 24.91 267.98 24.98 ;
    RECT 180.36 24.55 180.57 24.62 ;
    RECT 180.36 24.91 180.57 24.98 ;
    RECT 180.36 25.27 180.57 25.34 ;
    RECT 179.9 24.55 180.11 24.62 ;
    RECT 179.9 24.91 180.11 24.98 ;
    RECT 179.9 25.27 180.11 25.34 ;
    RECT 177.04 24.55 177.25 24.62 ;
    RECT 177.04 24.91 177.25 24.98 ;
    RECT 177.04 25.27 177.25 25.34 ;
    RECT 176.58 24.55 176.79 24.62 ;
    RECT 176.58 24.91 176.79 24.98 ;
    RECT 176.58 25.27 176.79 25.34 ;
    RECT 173.72 24.55 173.93 24.62 ;
    RECT 173.72 24.91 173.93 24.98 ;
    RECT 173.72 25.27 173.93 25.34 ;
    RECT 173.26 24.55 173.47 24.62 ;
    RECT 173.26 24.91 173.47 24.98 ;
    RECT 173.26 25.27 173.47 25.34 ;
    RECT 170.4 24.55 170.61 24.62 ;
    RECT 170.4 24.91 170.61 24.98 ;
    RECT 170.4 25.27 170.61 25.34 ;
    RECT 169.94 24.55 170.15 24.62 ;
    RECT 169.94 24.91 170.15 24.98 ;
    RECT 169.94 25.27 170.15 25.34 ;
    RECT 167.08 24.55 167.29 24.62 ;
    RECT 167.08 24.91 167.29 24.98 ;
    RECT 167.08 25.27 167.29 25.34 ;
    RECT 166.62 24.55 166.83 24.62 ;
    RECT 166.62 24.91 166.83 24.98 ;
    RECT 166.62 25.27 166.83 25.34 ;
    RECT 163.76 24.55 163.97 24.62 ;
    RECT 163.76 24.91 163.97 24.98 ;
    RECT 163.76 25.27 163.97 25.34 ;
    RECT 163.3 24.55 163.51 24.62 ;
    RECT 163.3 24.91 163.51 24.98 ;
    RECT 163.3 25.27 163.51 25.34 ;
    RECT 160.44 24.55 160.65 24.62 ;
    RECT 160.44 24.91 160.65 24.98 ;
    RECT 160.44 25.27 160.65 25.34 ;
    RECT 159.98 24.55 160.19 24.62 ;
    RECT 159.98 24.91 160.19 24.98 ;
    RECT 159.98 25.27 160.19 25.34 ;
    RECT 157.12 24.55 157.33 24.62 ;
    RECT 157.12 24.91 157.33 24.98 ;
    RECT 157.12 25.27 157.33 25.34 ;
    RECT 156.66 24.55 156.87 24.62 ;
    RECT 156.66 24.91 156.87 24.98 ;
    RECT 156.66 25.27 156.87 25.34 ;
    RECT 153.8 24.55 154.01 24.62 ;
    RECT 153.8 24.91 154.01 24.98 ;
    RECT 153.8 25.27 154.01 25.34 ;
    RECT 153.34 24.55 153.55 24.62 ;
    RECT 153.34 24.91 153.55 24.98 ;
    RECT 153.34 25.27 153.55 25.34 ;
    RECT 150.48 24.55 150.69 24.62 ;
    RECT 150.48 24.91 150.69 24.98 ;
    RECT 150.48 25.27 150.69 25.34 ;
    RECT 150.02 24.55 150.23 24.62 ;
    RECT 150.02 24.91 150.23 24.98 ;
    RECT 150.02 25.27 150.23 25.34 ;
    RECT 213.56 24.55 213.77 24.62 ;
    RECT 213.56 24.91 213.77 24.98 ;
    RECT 213.56 25.27 213.77 25.34 ;
    RECT 213.1 24.55 213.31 24.62 ;
    RECT 213.1 24.91 213.31 24.98 ;
    RECT 213.1 25.27 213.31 25.34 ;
    RECT 210.24 24.55 210.45 24.62 ;
    RECT 210.24 24.91 210.45 24.98 ;
    RECT 210.24 25.27 210.45 25.34 ;
    RECT 209.78 24.55 209.99 24.62 ;
    RECT 209.78 24.91 209.99 24.98 ;
    RECT 209.78 25.27 209.99 25.34 ;
    RECT 206.92 24.55 207.13 24.62 ;
    RECT 206.92 24.91 207.13 24.98 ;
    RECT 206.92 25.27 207.13 25.34 ;
    RECT 206.46 24.55 206.67 24.62 ;
    RECT 206.46 24.91 206.67 24.98 ;
    RECT 206.46 25.27 206.67 25.34 ;
    RECT 203.6 24.55 203.81 24.62 ;
    RECT 203.6 24.91 203.81 24.98 ;
    RECT 203.6 25.27 203.81 25.34 ;
    RECT 203.14 24.55 203.35 24.62 ;
    RECT 203.14 24.91 203.35 24.98 ;
    RECT 203.14 25.27 203.35 25.34 ;
    RECT 200.28 24.55 200.49 24.62 ;
    RECT 200.28 24.91 200.49 24.98 ;
    RECT 200.28 25.27 200.49 25.34 ;
    RECT 199.82 24.55 200.03 24.62 ;
    RECT 199.82 24.91 200.03 24.98 ;
    RECT 199.82 25.27 200.03 25.34 ;
    RECT 196.96 24.55 197.17 24.62 ;
    RECT 196.96 24.91 197.17 24.98 ;
    RECT 196.96 25.27 197.17 25.34 ;
    RECT 196.5 24.55 196.71 24.62 ;
    RECT 196.5 24.91 196.71 24.98 ;
    RECT 196.5 25.27 196.71 25.34 ;
    RECT 193.64 24.55 193.85 24.62 ;
    RECT 193.64 24.91 193.85 24.98 ;
    RECT 193.64 25.27 193.85 25.34 ;
    RECT 193.18 24.55 193.39 24.62 ;
    RECT 193.18 24.91 193.39 24.98 ;
    RECT 193.18 25.27 193.39 25.34 ;
    RECT 190.32 24.55 190.53 24.62 ;
    RECT 190.32 24.91 190.53 24.98 ;
    RECT 190.32 25.27 190.53 25.34 ;
    RECT 189.86 24.55 190.07 24.62 ;
    RECT 189.86 24.91 190.07 24.98 ;
    RECT 189.86 25.27 190.07 25.34 ;
    RECT 187.0 24.55 187.21 24.62 ;
    RECT 187.0 24.91 187.21 24.98 ;
    RECT 187.0 25.27 187.21 25.34 ;
    RECT 186.54 24.55 186.75 24.62 ;
    RECT 186.54 24.91 186.75 24.98 ;
    RECT 186.54 25.27 186.75 25.34 ;
    RECT 183.68 24.55 183.89 24.62 ;
    RECT 183.68 24.91 183.89 24.98 ;
    RECT 183.68 25.27 183.89 25.34 ;
    RECT 183.22 24.55 183.43 24.62 ;
    RECT 183.22 24.91 183.43 24.98 ;
    RECT 183.22 25.27 183.43 25.34 ;
    RECT 147.485 24.91 147.555 24.98 ;
    RECT 266.68 24.55 266.89 24.62 ;
    RECT 266.68 24.91 266.89 24.98 ;
    RECT 266.68 25.27 266.89 25.34 ;
    RECT 266.22 24.55 266.43 24.62 ;
    RECT 266.22 24.91 266.43 24.98 ;
    RECT 266.22 25.27 266.43 25.34 ;
    RECT 263.36 24.55 263.57 24.62 ;
    RECT 263.36 24.91 263.57 24.98 ;
    RECT 263.36 25.27 263.57 25.34 ;
    RECT 262.9 24.55 263.11 24.62 ;
    RECT 262.9 24.91 263.11 24.98 ;
    RECT 262.9 25.27 263.11 25.34 ;
    RECT 260.04 24.55 260.25 24.62 ;
    RECT 260.04 24.91 260.25 24.98 ;
    RECT 260.04 25.27 260.25 25.34 ;
    RECT 259.58 24.55 259.79 24.62 ;
    RECT 259.58 24.91 259.79 24.98 ;
    RECT 259.58 25.27 259.79 25.34 ;
    RECT 256.72 24.55 256.93 24.62 ;
    RECT 256.72 24.91 256.93 24.98 ;
    RECT 256.72 25.27 256.93 25.34 ;
    RECT 256.26 24.55 256.47 24.62 ;
    RECT 256.26 24.91 256.47 24.98 ;
    RECT 256.26 25.27 256.47 25.34 ;
    RECT 253.4 24.55 253.61 24.62 ;
    RECT 253.4 24.91 253.61 24.98 ;
    RECT 253.4 25.27 253.61 25.34 ;
    RECT 252.94 24.55 253.15 24.62 ;
    RECT 252.94 24.91 253.15 24.98 ;
    RECT 252.94 25.27 253.15 25.34 ;
    RECT 250.08 64.17 250.29 64.24 ;
    RECT 250.08 64.53 250.29 64.6 ;
    RECT 250.08 64.89 250.29 64.96 ;
    RECT 249.62 64.17 249.83 64.24 ;
    RECT 249.62 64.53 249.83 64.6 ;
    RECT 249.62 64.89 249.83 64.96 ;
    RECT 246.76 64.17 246.97 64.24 ;
    RECT 246.76 64.53 246.97 64.6 ;
    RECT 246.76 64.89 246.97 64.96 ;
    RECT 246.3 64.17 246.51 64.24 ;
    RECT 246.3 64.53 246.51 64.6 ;
    RECT 246.3 64.89 246.51 64.96 ;
    RECT 243.44 64.17 243.65 64.24 ;
    RECT 243.44 64.53 243.65 64.6 ;
    RECT 243.44 64.89 243.65 64.96 ;
    RECT 242.98 64.17 243.19 64.24 ;
    RECT 242.98 64.53 243.19 64.6 ;
    RECT 242.98 64.89 243.19 64.96 ;
    RECT 240.12 64.17 240.33 64.24 ;
    RECT 240.12 64.53 240.33 64.6 ;
    RECT 240.12 64.89 240.33 64.96 ;
    RECT 239.66 64.17 239.87 64.24 ;
    RECT 239.66 64.53 239.87 64.6 ;
    RECT 239.66 64.89 239.87 64.96 ;
    RECT 236.8 64.17 237.01 64.24 ;
    RECT 236.8 64.53 237.01 64.6 ;
    RECT 236.8 64.89 237.01 64.96 ;
    RECT 236.34 64.17 236.55 64.24 ;
    RECT 236.34 64.53 236.55 64.6 ;
    RECT 236.34 64.89 236.55 64.96 ;
    RECT 233.48 64.17 233.69 64.24 ;
    RECT 233.48 64.53 233.69 64.6 ;
    RECT 233.48 64.89 233.69 64.96 ;
    RECT 233.02 64.17 233.23 64.24 ;
    RECT 233.02 64.53 233.23 64.6 ;
    RECT 233.02 64.89 233.23 64.96 ;
    RECT 230.16 64.17 230.37 64.24 ;
    RECT 230.16 64.53 230.37 64.6 ;
    RECT 230.16 64.89 230.37 64.96 ;
    RECT 229.7 64.17 229.91 64.24 ;
    RECT 229.7 64.53 229.91 64.6 ;
    RECT 229.7 64.89 229.91 64.96 ;
    RECT 226.84 64.17 227.05 64.24 ;
    RECT 226.84 64.53 227.05 64.6 ;
    RECT 226.84 64.89 227.05 64.96 ;
    RECT 226.38 64.17 226.59 64.24 ;
    RECT 226.38 64.53 226.59 64.6 ;
    RECT 226.38 64.89 226.59 64.96 ;
    RECT 223.52 64.17 223.73 64.24 ;
    RECT 223.52 64.53 223.73 64.6 ;
    RECT 223.52 64.89 223.73 64.96 ;
    RECT 223.06 64.17 223.27 64.24 ;
    RECT 223.06 64.53 223.27 64.6 ;
    RECT 223.06 64.89 223.27 64.96 ;
    RECT 220.2 64.17 220.41 64.24 ;
    RECT 220.2 64.53 220.41 64.6 ;
    RECT 220.2 64.89 220.41 64.96 ;
    RECT 219.74 64.17 219.95 64.24 ;
    RECT 219.74 64.53 219.95 64.6 ;
    RECT 219.74 64.89 219.95 64.96 ;
    RECT 216.88 64.17 217.09 64.24 ;
    RECT 216.88 64.53 217.09 64.6 ;
    RECT 216.88 64.89 217.09 64.96 ;
    RECT 216.42 64.17 216.63 64.24 ;
    RECT 216.42 64.53 216.63 64.6 ;
    RECT 216.42 64.89 216.63 64.96 ;
    RECT 267.91 64.53 267.98 64.6 ;
    RECT 180.36 64.17 180.57 64.24 ;
    RECT 180.36 64.53 180.57 64.6 ;
    RECT 180.36 64.89 180.57 64.96 ;
    RECT 179.9 64.17 180.11 64.24 ;
    RECT 179.9 64.53 180.11 64.6 ;
    RECT 179.9 64.89 180.11 64.96 ;
    RECT 177.04 64.17 177.25 64.24 ;
    RECT 177.04 64.53 177.25 64.6 ;
    RECT 177.04 64.89 177.25 64.96 ;
    RECT 176.58 64.17 176.79 64.24 ;
    RECT 176.58 64.53 176.79 64.6 ;
    RECT 176.58 64.89 176.79 64.96 ;
    RECT 173.72 64.17 173.93 64.24 ;
    RECT 173.72 64.53 173.93 64.6 ;
    RECT 173.72 64.89 173.93 64.96 ;
    RECT 173.26 64.17 173.47 64.24 ;
    RECT 173.26 64.53 173.47 64.6 ;
    RECT 173.26 64.89 173.47 64.96 ;
    RECT 170.4 64.17 170.61 64.24 ;
    RECT 170.4 64.53 170.61 64.6 ;
    RECT 170.4 64.89 170.61 64.96 ;
    RECT 169.94 64.17 170.15 64.24 ;
    RECT 169.94 64.53 170.15 64.6 ;
    RECT 169.94 64.89 170.15 64.96 ;
    RECT 167.08 64.17 167.29 64.24 ;
    RECT 167.08 64.53 167.29 64.6 ;
    RECT 167.08 64.89 167.29 64.96 ;
    RECT 166.62 64.17 166.83 64.24 ;
    RECT 166.62 64.53 166.83 64.6 ;
    RECT 166.62 64.89 166.83 64.96 ;
    RECT 163.76 64.17 163.97 64.24 ;
    RECT 163.76 64.53 163.97 64.6 ;
    RECT 163.76 64.89 163.97 64.96 ;
    RECT 163.3 64.17 163.51 64.24 ;
    RECT 163.3 64.53 163.51 64.6 ;
    RECT 163.3 64.89 163.51 64.96 ;
    RECT 160.44 64.17 160.65 64.24 ;
    RECT 160.44 64.53 160.65 64.6 ;
    RECT 160.44 64.89 160.65 64.96 ;
    RECT 159.98 64.17 160.19 64.24 ;
    RECT 159.98 64.53 160.19 64.6 ;
    RECT 159.98 64.89 160.19 64.96 ;
    RECT 157.12 64.17 157.33 64.24 ;
    RECT 157.12 64.53 157.33 64.6 ;
    RECT 157.12 64.89 157.33 64.96 ;
    RECT 156.66 64.17 156.87 64.24 ;
    RECT 156.66 64.53 156.87 64.6 ;
    RECT 156.66 64.89 156.87 64.96 ;
    RECT 153.8 64.17 154.01 64.24 ;
    RECT 153.8 64.53 154.01 64.6 ;
    RECT 153.8 64.89 154.01 64.96 ;
    RECT 153.34 64.17 153.55 64.24 ;
    RECT 153.34 64.53 153.55 64.6 ;
    RECT 153.34 64.89 153.55 64.96 ;
    RECT 150.48 64.17 150.69 64.24 ;
    RECT 150.48 64.53 150.69 64.6 ;
    RECT 150.48 64.89 150.69 64.96 ;
    RECT 150.02 64.17 150.23 64.24 ;
    RECT 150.02 64.53 150.23 64.6 ;
    RECT 150.02 64.89 150.23 64.96 ;
    RECT 213.56 64.17 213.77 64.24 ;
    RECT 213.56 64.53 213.77 64.6 ;
    RECT 213.56 64.89 213.77 64.96 ;
    RECT 213.1 64.17 213.31 64.24 ;
    RECT 213.1 64.53 213.31 64.6 ;
    RECT 213.1 64.89 213.31 64.96 ;
    RECT 210.24 64.17 210.45 64.24 ;
    RECT 210.24 64.53 210.45 64.6 ;
    RECT 210.24 64.89 210.45 64.96 ;
    RECT 209.78 64.17 209.99 64.24 ;
    RECT 209.78 64.53 209.99 64.6 ;
    RECT 209.78 64.89 209.99 64.96 ;
    RECT 206.92 64.17 207.13 64.24 ;
    RECT 206.92 64.53 207.13 64.6 ;
    RECT 206.92 64.89 207.13 64.96 ;
    RECT 206.46 64.17 206.67 64.24 ;
    RECT 206.46 64.53 206.67 64.6 ;
    RECT 206.46 64.89 206.67 64.96 ;
    RECT 203.6 64.17 203.81 64.24 ;
    RECT 203.6 64.53 203.81 64.6 ;
    RECT 203.6 64.89 203.81 64.96 ;
    RECT 203.14 64.17 203.35 64.24 ;
    RECT 203.14 64.53 203.35 64.6 ;
    RECT 203.14 64.89 203.35 64.96 ;
    RECT 200.28 64.17 200.49 64.24 ;
    RECT 200.28 64.53 200.49 64.6 ;
    RECT 200.28 64.89 200.49 64.96 ;
    RECT 199.82 64.17 200.03 64.24 ;
    RECT 199.82 64.53 200.03 64.6 ;
    RECT 199.82 64.89 200.03 64.96 ;
    RECT 196.96 64.17 197.17 64.24 ;
    RECT 196.96 64.53 197.17 64.6 ;
    RECT 196.96 64.89 197.17 64.96 ;
    RECT 196.5 64.17 196.71 64.24 ;
    RECT 196.5 64.53 196.71 64.6 ;
    RECT 196.5 64.89 196.71 64.96 ;
    RECT 193.64 64.17 193.85 64.24 ;
    RECT 193.64 64.53 193.85 64.6 ;
    RECT 193.64 64.89 193.85 64.96 ;
    RECT 193.18 64.17 193.39 64.24 ;
    RECT 193.18 64.53 193.39 64.6 ;
    RECT 193.18 64.89 193.39 64.96 ;
    RECT 190.32 64.17 190.53 64.24 ;
    RECT 190.32 64.53 190.53 64.6 ;
    RECT 190.32 64.89 190.53 64.96 ;
    RECT 189.86 64.17 190.07 64.24 ;
    RECT 189.86 64.53 190.07 64.6 ;
    RECT 189.86 64.89 190.07 64.96 ;
    RECT 187.0 64.17 187.21 64.24 ;
    RECT 187.0 64.53 187.21 64.6 ;
    RECT 187.0 64.89 187.21 64.96 ;
    RECT 186.54 64.17 186.75 64.24 ;
    RECT 186.54 64.53 186.75 64.6 ;
    RECT 186.54 64.89 186.75 64.96 ;
    RECT 183.68 64.17 183.89 64.24 ;
    RECT 183.68 64.53 183.89 64.6 ;
    RECT 183.68 64.89 183.89 64.96 ;
    RECT 183.22 64.17 183.43 64.24 ;
    RECT 183.22 64.53 183.43 64.6 ;
    RECT 183.22 64.89 183.43 64.96 ;
    RECT 147.485 64.53 147.555 64.6 ;
    RECT 266.68 64.17 266.89 64.24 ;
    RECT 266.68 64.53 266.89 64.6 ;
    RECT 266.68 64.89 266.89 64.96 ;
    RECT 266.22 64.17 266.43 64.24 ;
    RECT 266.22 64.53 266.43 64.6 ;
    RECT 266.22 64.89 266.43 64.96 ;
    RECT 263.36 64.17 263.57 64.24 ;
    RECT 263.36 64.53 263.57 64.6 ;
    RECT 263.36 64.89 263.57 64.96 ;
    RECT 262.9 64.17 263.11 64.24 ;
    RECT 262.9 64.53 263.11 64.6 ;
    RECT 262.9 64.89 263.11 64.96 ;
    RECT 260.04 64.17 260.25 64.24 ;
    RECT 260.04 64.53 260.25 64.6 ;
    RECT 260.04 64.89 260.25 64.96 ;
    RECT 259.58 64.17 259.79 64.24 ;
    RECT 259.58 64.53 259.79 64.6 ;
    RECT 259.58 64.89 259.79 64.96 ;
    RECT 256.72 64.17 256.93 64.24 ;
    RECT 256.72 64.53 256.93 64.6 ;
    RECT 256.72 64.89 256.93 64.96 ;
    RECT 256.26 64.17 256.47 64.24 ;
    RECT 256.26 64.53 256.47 64.6 ;
    RECT 256.26 64.89 256.47 64.96 ;
    RECT 253.4 64.17 253.61 64.24 ;
    RECT 253.4 64.53 253.61 64.6 ;
    RECT 253.4 64.89 253.61 64.96 ;
    RECT 252.94 64.17 253.15 64.24 ;
    RECT 252.94 64.53 253.15 64.6 ;
    RECT 252.94 64.89 253.15 64.96 ;
    RECT 250.08 23.83 250.29 23.9 ;
    RECT 250.08 24.19 250.29 24.26 ;
    RECT 250.08 24.55 250.29 24.62 ;
    RECT 249.62 23.83 249.83 23.9 ;
    RECT 249.62 24.19 249.83 24.26 ;
    RECT 249.62 24.55 249.83 24.62 ;
    RECT 246.76 23.83 246.97 23.9 ;
    RECT 246.76 24.19 246.97 24.26 ;
    RECT 246.76 24.55 246.97 24.62 ;
    RECT 246.3 23.83 246.51 23.9 ;
    RECT 246.3 24.19 246.51 24.26 ;
    RECT 246.3 24.55 246.51 24.62 ;
    RECT 243.44 23.83 243.65 23.9 ;
    RECT 243.44 24.19 243.65 24.26 ;
    RECT 243.44 24.55 243.65 24.62 ;
    RECT 242.98 23.83 243.19 23.9 ;
    RECT 242.98 24.19 243.19 24.26 ;
    RECT 242.98 24.55 243.19 24.62 ;
    RECT 240.12 23.83 240.33 23.9 ;
    RECT 240.12 24.19 240.33 24.26 ;
    RECT 240.12 24.55 240.33 24.62 ;
    RECT 239.66 23.83 239.87 23.9 ;
    RECT 239.66 24.19 239.87 24.26 ;
    RECT 239.66 24.55 239.87 24.62 ;
    RECT 236.8 23.83 237.01 23.9 ;
    RECT 236.8 24.19 237.01 24.26 ;
    RECT 236.8 24.55 237.01 24.62 ;
    RECT 236.34 23.83 236.55 23.9 ;
    RECT 236.34 24.19 236.55 24.26 ;
    RECT 236.34 24.55 236.55 24.62 ;
    RECT 233.48 23.83 233.69 23.9 ;
    RECT 233.48 24.19 233.69 24.26 ;
    RECT 233.48 24.55 233.69 24.62 ;
    RECT 233.02 23.83 233.23 23.9 ;
    RECT 233.02 24.19 233.23 24.26 ;
    RECT 233.02 24.55 233.23 24.62 ;
    RECT 230.16 23.83 230.37 23.9 ;
    RECT 230.16 24.19 230.37 24.26 ;
    RECT 230.16 24.55 230.37 24.62 ;
    RECT 229.7 23.83 229.91 23.9 ;
    RECT 229.7 24.19 229.91 24.26 ;
    RECT 229.7 24.55 229.91 24.62 ;
    RECT 226.84 23.83 227.05 23.9 ;
    RECT 226.84 24.19 227.05 24.26 ;
    RECT 226.84 24.55 227.05 24.62 ;
    RECT 226.38 23.83 226.59 23.9 ;
    RECT 226.38 24.19 226.59 24.26 ;
    RECT 226.38 24.55 226.59 24.62 ;
    RECT 223.52 23.83 223.73 23.9 ;
    RECT 223.52 24.19 223.73 24.26 ;
    RECT 223.52 24.55 223.73 24.62 ;
    RECT 223.06 23.83 223.27 23.9 ;
    RECT 223.06 24.19 223.27 24.26 ;
    RECT 223.06 24.55 223.27 24.62 ;
    RECT 220.2 23.83 220.41 23.9 ;
    RECT 220.2 24.19 220.41 24.26 ;
    RECT 220.2 24.55 220.41 24.62 ;
    RECT 219.74 23.83 219.95 23.9 ;
    RECT 219.74 24.19 219.95 24.26 ;
    RECT 219.74 24.55 219.95 24.62 ;
    RECT 216.88 23.83 217.09 23.9 ;
    RECT 216.88 24.19 217.09 24.26 ;
    RECT 216.88 24.55 217.09 24.62 ;
    RECT 216.42 23.83 216.63 23.9 ;
    RECT 216.42 24.19 216.63 24.26 ;
    RECT 216.42 24.55 216.63 24.62 ;
    RECT 267.91 24.19 267.98 24.26 ;
    RECT 180.36 23.83 180.57 23.9 ;
    RECT 180.36 24.19 180.57 24.26 ;
    RECT 180.36 24.55 180.57 24.62 ;
    RECT 179.9 23.83 180.11 23.9 ;
    RECT 179.9 24.19 180.11 24.26 ;
    RECT 179.9 24.55 180.11 24.62 ;
    RECT 177.04 23.83 177.25 23.9 ;
    RECT 177.04 24.19 177.25 24.26 ;
    RECT 177.04 24.55 177.25 24.62 ;
    RECT 176.58 23.83 176.79 23.9 ;
    RECT 176.58 24.19 176.79 24.26 ;
    RECT 176.58 24.55 176.79 24.62 ;
    RECT 173.72 23.83 173.93 23.9 ;
    RECT 173.72 24.19 173.93 24.26 ;
    RECT 173.72 24.55 173.93 24.62 ;
    RECT 173.26 23.83 173.47 23.9 ;
    RECT 173.26 24.19 173.47 24.26 ;
    RECT 173.26 24.55 173.47 24.62 ;
    RECT 170.4 23.83 170.61 23.9 ;
    RECT 170.4 24.19 170.61 24.26 ;
    RECT 170.4 24.55 170.61 24.62 ;
    RECT 169.94 23.83 170.15 23.9 ;
    RECT 169.94 24.19 170.15 24.26 ;
    RECT 169.94 24.55 170.15 24.62 ;
    RECT 167.08 23.83 167.29 23.9 ;
    RECT 167.08 24.19 167.29 24.26 ;
    RECT 167.08 24.55 167.29 24.62 ;
    RECT 166.62 23.83 166.83 23.9 ;
    RECT 166.62 24.19 166.83 24.26 ;
    RECT 166.62 24.55 166.83 24.62 ;
    RECT 163.76 23.83 163.97 23.9 ;
    RECT 163.76 24.19 163.97 24.26 ;
    RECT 163.76 24.55 163.97 24.62 ;
    RECT 163.3 23.83 163.51 23.9 ;
    RECT 163.3 24.19 163.51 24.26 ;
    RECT 163.3 24.55 163.51 24.62 ;
    RECT 160.44 23.83 160.65 23.9 ;
    RECT 160.44 24.19 160.65 24.26 ;
    RECT 160.44 24.55 160.65 24.62 ;
    RECT 159.98 23.83 160.19 23.9 ;
    RECT 159.98 24.19 160.19 24.26 ;
    RECT 159.98 24.55 160.19 24.62 ;
    RECT 157.12 23.83 157.33 23.9 ;
    RECT 157.12 24.19 157.33 24.26 ;
    RECT 157.12 24.55 157.33 24.62 ;
    RECT 156.66 23.83 156.87 23.9 ;
    RECT 156.66 24.19 156.87 24.26 ;
    RECT 156.66 24.55 156.87 24.62 ;
    RECT 153.8 23.83 154.01 23.9 ;
    RECT 153.8 24.19 154.01 24.26 ;
    RECT 153.8 24.55 154.01 24.62 ;
    RECT 153.34 23.83 153.55 23.9 ;
    RECT 153.34 24.19 153.55 24.26 ;
    RECT 153.34 24.55 153.55 24.62 ;
    RECT 150.48 23.83 150.69 23.9 ;
    RECT 150.48 24.19 150.69 24.26 ;
    RECT 150.48 24.55 150.69 24.62 ;
    RECT 150.02 23.83 150.23 23.9 ;
    RECT 150.02 24.19 150.23 24.26 ;
    RECT 150.02 24.55 150.23 24.62 ;
    RECT 213.56 23.83 213.77 23.9 ;
    RECT 213.56 24.19 213.77 24.26 ;
    RECT 213.56 24.55 213.77 24.62 ;
    RECT 213.1 23.83 213.31 23.9 ;
    RECT 213.1 24.19 213.31 24.26 ;
    RECT 213.1 24.55 213.31 24.62 ;
    RECT 210.24 23.83 210.45 23.9 ;
    RECT 210.24 24.19 210.45 24.26 ;
    RECT 210.24 24.55 210.45 24.62 ;
    RECT 209.78 23.83 209.99 23.9 ;
    RECT 209.78 24.19 209.99 24.26 ;
    RECT 209.78 24.55 209.99 24.62 ;
    RECT 206.92 23.83 207.13 23.9 ;
    RECT 206.92 24.19 207.13 24.26 ;
    RECT 206.92 24.55 207.13 24.62 ;
    RECT 206.46 23.83 206.67 23.9 ;
    RECT 206.46 24.19 206.67 24.26 ;
    RECT 206.46 24.55 206.67 24.62 ;
    RECT 203.6 23.83 203.81 23.9 ;
    RECT 203.6 24.19 203.81 24.26 ;
    RECT 203.6 24.55 203.81 24.62 ;
    RECT 203.14 23.83 203.35 23.9 ;
    RECT 203.14 24.19 203.35 24.26 ;
    RECT 203.14 24.55 203.35 24.62 ;
    RECT 200.28 23.83 200.49 23.9 ;
    RECT 200.28 24.19 200.49 24.26 ;
    RECT 200.28 24.55 200.49 24.62 ;
    RECT 199.82 23.83 200.03 23.9 ;
    RECT 199.82 24.19 200.03 24.26 ;
    RECT 199.82 24.55 200.03 24.62 ;
    RECT 196.96 23.83 197.17 23.9 ;
    RECT 196.96 24.19 197.17 24.26 ;
    RECT 196.96 24.55 197.17 24.62 ;
    RECT 196.5 23.83 196.71 23.9 ;
    RECT 196.5 24.19 196.71 24.26 ;
    RECT 196.5 24.55 196.71 24.62 ;
    RECT 193.64 23.83 193.85 23.9 ;
    RECT 193.64 24.19 193.85 24.26 ;
    RECT 193.64 24.55 193.85 24.62 ;
    RECT 193.18 23.83 193.39 23.9 ;
    RECT 193.18 24.19 193.39 24.26 ;
    RECT 193.18 24.55 193.39 24.62 ;
    RECT 190.32 23.83 190.53 23.9 ;
    RECT 190.32 24.19 190.53 24.26 ;
    RECT 190.32 24.55 190.53 24.62 ;
    RECT 189.86 23.83 190.07 23.9 ;
    RECT 189.86 24.19 190.07 24.26 ;
    RECT 189.86 24.55 190.07 24.62 ;
    RECT 187.0 23.83 187.21 23.9 ;
    RECT 187.0 24.19 187.21 24.26 ;
    RECT 187.0 24.55 187.21 24.62 ;
    RECT 186.54 23.83 186.75 23.9 ;
    RECT 186.54 24.19 186.75 24.26 ;
    RECT 186.54 24.55 186.75 24.62 ;
    RECT 183.68 23.83 183.89 23.9 ;
    RECT 183.68 24.19 183.89 24.26 ;
    RECT 183.68 24.55 183.89 24.62 ;
    RECT 183.22 23.83 183.43 23.9 ;
    RECT 183.22 24.19 183.43 24.26 ;
    RECT 183.22 24.55 183.43 24.62 ;
    RECT 147.485 24.19 147.555 24.26 ;
    RECT 266.68 23.83 266.89 23.9 ;
    RECT 266.68 24.19 266.89 24.26 ;
    RECT 266.68 24.55 266.89 24.62 ;
    RECT 266.22 23.83 266.43 23.9 ;
    RECT 266.22 24.19 266.43 24.26 ;
    RECT 266.22 24.55 266.43 24.62 ;
    RECT 263.36 23.83 263.57 23.9 ;
    RECT 263.36 24.19 263.57 24.26 ;
    RECT 263.36 24.55 263.57 24.62 ;
    RECT 262.9 23.83 263.11 23.9 ;
    RECT 262.9 24.19 263.11 24.26 ;
    RECT 262.9 24.55 263.11 24.62 ;
    RECT 260.04 23.83 260.25 23.9 ;
    RECT 260.04 24.19 260.25 24.26 ;
    RECT 260.04 24.55 260.25 24.62 ;
    RECT 259.58 23.83 259.79 23.9 ;
    RECT 259.58 24.19 259.79 24.26 ;
    RECT 259.58 24.55 259.79 24.62 ;
    RECT 256.72 23.83 256.93 23.9 ;
    RECT 256.72 24.19 256.93 24.26 ;
    RECT 256.72 24.55 256.93 24.62 ;
    RECT 256.26 23.83 256.47 23.9 ;
    RECT 256.26 24.19 256.47 24.26 ;
    RECT 256.26 24.55 256.47 24.62 ;
    RECT 253.4 23.83 253.61 23.9 ;
    RECT 253.4 24.19 253.61 24.26 ;
    RECT 253.4 24.55 253.61 24.62 ;
    RECT 252.94 23.83 253.15 23.9 ;
    RECT 252.94 24.19 253.15 24.26 ;
    RECT 252.94 24.55 253.15 24.62 ;
    RECT 250.08 63.45 250.29 63.52 ;
    RECT 250.08 63.81 250.29 63.88 ;
    RECT 250.08 64.17 250.29 64.24 ;
    RECT 249.62 63.45 249.83 63.52 ;
    RECT 249.62 63.81 249.83 63.88 ;
    RECT 249.62 64.17 249.83 64.24 ;
    RECT 246.76 63.45 246.97 63.52 ;
    RECT 246.76 63.81 246.97 63.88 ;
    RECT 246.76 64.17 246.97 64.24 ;
    RECT 246.3 63.45 246.51 63.52 ;
    RECT 246.3 63.81 246.51 63.88 ;
    RECT 246.3 64.17 246.51 64.24 ;
    RECT 243.44 63.45 243.65 63.52 ;
    RECT 243.44 63.81 243.65 63.88 ;
    RECT 243.44 64.17 243.65 64.24 ;
    RECT 242.98 63.45 243.19 63.52 ;
    RECT 242.98 63.81 243.19 63.88 ;
    RECT 242.98 64.17 243.19 64.24 ;
    RECT 240.12 63.45 240.33 63.52 ;
    RECT 240.12 63.81 240.33 63.88 ;
    RECT 240.12 64.17 240.33 64.24 ;
    RECT 239.66 63.45 239.87 63.52 ;
    RECT 239.66 63.81 239.87 63.88 ;
    RECT 239.66 64.17 239.87 64.24 ;
    RECT 236.8 63.45 237.01 63.52 ;
    RECT 236.8 63.81 237.01 63.88 ;
    RECT 236.8 64.17 237.01 64.24 ;
    RECT 236.34 63.45 236.55 63.52 ;
    RECT 236.34 63.81 236.55 63.88 ;
    RECT 236.34 64.17 236.55 64.24 ;
    RECT 233.48 63.45 233.69 63.52 ;
    RECT 233.48 63.81 233.69 63.88 ;
    RECT 233.48 64.17 233.69 64.24 ;
    RECT 233.02 63.45 233.23 63.52 ;
    RECT 233.02 63.81 233.23 63.88 ;
    RECT 233.02 64.17 233.23 64.24 ;
    RECT 230.16 63.45 230.37 63.52 ;
    RECT 230.16 63.81 230.37 63.88 ;
    RECT 230.16 64.17 230.37 64.24 ;
    RECT 229.7 63.45 229.91 63.52 ;
    RECT 229.7 63.81 229.91 63.88 ;
    RECT 229.7 64.17 229.91 64.24 ;
    RECT 226.84 63.45 227.05 63.52 ;
    RECT 226.84 63.81 227.05 63.88 ;
    RECT 226.84 64.17 227.05 64.24 ;
    RECT 226.38 63.45 226.59 63.52 ;
    RECT 226.38 63.81 226.59 63.88 ;
    RECT 226.38 64.17 226.59 64.24 ;
    RECT 223.52 63.45 223.73 63.52 ;
    RECT 223.52 63.81 223.73 63.88 ;
    RECT 223.52 64.17 223.73 64.24 ;
    RECT 223.06 63.45 223.27 63.52 ;
    RECT 223.06 63.81 223.27 63.88 ;
    RECT 223.06 64.17 223.27 64.24 ;
    RECT 220.2 63.45 220.41 63.52 ;
    RECT 220.2 63.81 220.41 63.88 ;
    RECT 220.2 64.17 220.41 64.24 ;
    RECT 219.74 63.45 219.95 63.52 ;
    RECT 219.74 63.81 219.95 63.88 ;
    RECT 219.74 64.17 219.95 64.24 ;
    RECT 216.88 63.45 217.09 63.52 ;
    RECT 216.88 63.81 217.09 63.88 ;
    RECT 216.88 64.17 217.09 64.24 ;
    RECT 216.42 63.45 216.63 63.52 ;
    RECT 216.42 63.81 216.63 63.88 ;
    RECT 216.42 64.17 216.63 64.24 ;
    RECT 267.91 63.81 267.98 63.88 ;
    RECT 180.36 63.45 180.57 63.52 ;
    RECT 180.36 63.81 180.57 63.88 ;
    RECT 180.36 64.17 180.57 64.24 ;
    RECT 179.9 63.45 180.11 63.52 ;
    RECT 179.9 63.81 180.11 63.88 ;
    RECT 179.9 64.17 180.11 64.24 ;
    RECT 177.04 63.45 177.25 63.52 ;
    RECT 177.04 63.81 177.25 63.88 ;
    RECT 177.04 64.17 177.25 64.24 ;
    RECT 176.58 63.45 176.79 63.52 ;
    RECT 176.58 63.81 176.79 63.88 ;
    RECT 176.58 64.17 176.79 64.24 ;
    RECT 173.72 63.45 173.93 63.52 ;
    RECT 173.72 63.81 173.93 63.88 ;
    RECT 173.72 64.17 173.93 64.24 ;
    RECT 173.26 63.45 173.47 63.52 ;
    RECT 173.26 63.81 173.47 63.88 ;
    RECT 173.26 64.17 173.47 64.24 ;
    RECT 170.4 63.45 170.61 63.52 ;
    RECT 170.4 63.81 170.61 63.88 ;
    RECT 170.4 64.17 170.61 64.24 ;
    RECT 169.94 63.45 170.15 63.52 ;
    RECT 169.94 63.81 170.15 63.88 ;
    RECT 169.94 64.17 170.15 64.24 ;
    RECT 167.08 63.45 167.29 63.52 ;
    RECT 167.08 63.81 167.29 63.88 ;
    RECT 167.08 64.17 167.29 64.24 ;
    RECT 166.62 63.45 166.83 63.52 ;
    RECT 166.62 63.81 166.83 63.88 ;
    RECT 166.62 64.17 166.83 64.24 ;
    RECT 163.76 63.45 163.97 63.52 ;
    RECT 163.76 63.81 163.97 63.88 ;
    RECT 163.76 64.17 163.97 64.24 ;
    RECT 163.3 63.45 163.51 63.52 ;
    RECT 163.3 63.81 163.51 63.88 ;
    RECT 163.3 64.17 163.51 64.24 ;
    RECT 160.44 63.45 160.65 63.52 ;
    RECT 160.44 63.81 160.65 63.88 ;
    RECT 160.44 64.17 160.65 64.24 ;
    RECT 159.98 63.45 160.19 63.52 ;
    RECT 159.98 63.81 160.19 63.88 ;
    RECT 159.98 64.17 160.19 64.24 ;
    RECT 157.12 63.45 157.33 63.52 ;
    RECT 157.12 63.81 157.33 63.88 ;
    RECT 157.12 64.17 157.33 64.24 ;
    RECT 156.66 63.45 156.87 63.52 ;
    RECT 156.66 63.81 156.87 63.88 ;
    RECT 156.66 64.17 156.87 64.24 ;
    RECT 153.8 63.45 154.01 63.52 ;
    RECT 153.8 63.81 154.01 63.88 ;
    RECT 153.8 64.17 154.01 64.24 ;
    RECT 153.34 63.45 153.55 63.52 ;
    RECT 153.34 63.81 153.55 63.88 ;
    RECT 153.34 64.17 153.55 64.24 ;
    RECT 150.48 63.45 150.69 63.52 ;
    RECT 150.48 63.81 150.69 63.88 ;
    RECT 150.48 64.17 150.69 64.24 ;
    RECT 150.02 63.45 150.23 63.52 ;
    RECT 150.02 63.81 150.23 63.88 ;
    RECT 150.02 64.17 150.23 64.24 ;
    RECT 213.56 63.45 213.77 63.52 ;
    RECT 213.56 63.81 213.77 63.88 ;
    RECT 213.56 64.17 213.77 64.24 ;
    RECT 213.1 63.45 213.31 63.52 ;
    RECT 213.1 63.81 213.31 63.88 ;
    RECT 213.1 64.17 213.31 64.24 ;
    RECT 210.24 63.45 210.45 63.52 ;
    RECT 210.24 63.81 210.45 63.88 ;
    RECT 210.24 64.17 210.45 64.24 ;
    RECT 209.78 63.45 209.99 63.52 ;
    RECT 209.78 63.81 209.99 63.88 ;
    RECT 209.78 64.17 209.99 64.24 ;
    RECT 206.92 63.45 207.13 63.52 ;
    RECT 206.92 63.81 207.13 63.88 ;
    RECT 206.92 64.17 207.13 64.24 ;
    RECT 206.46 63.45 206.67 63.52 ;
    RECT 206.46 63.81 206.67 63.88 ;
    RECT 206.46 64.17 206.67 64.24 ;
    RECT 203.6 63.45 203.81 63.52 ;
    RECT 203.6 63.81 203.81 63.88 ;
    RECT 203.6 64.17 203.81 64.24 ;
    RECT 203.14 63.45 203.35 63.52 ;
    RECT 203.14 63.81 203.35 63.88 ;
    RECT 203.14 64.17 203.35 64.24 ;
    RECT 200.28 63.45 200.49 63.52 ;
    RECT 200.28 63.81 200.49 63.88 ;
    RECT 200.28 64.17 200.49 64.24 ;
    RECT 199.82 63.45 200.03 63.52 ;
    RECT 199.82 63.81 200.03 63.88 ;
    RECT 199.82 64.17 200.03 64.24 ;
    RECT 196.96 63.45 197.17 63.52 ;
    RECT 196.96 63.81 197.17 63.88 ;
    RECT 196.96 64.17 197.17 64.24 ;
    RECT 196.5 63.45 196.71 63.52 ;
    RECT 196.5 63.81 196.71 63.88 ;
    RECT 196.5 64.17 196.71 64.24 ;
    RECT 193.64 63.45 193.85 63.52 ;
    RECT 193.64 63.81 193.85 63.88 ;
    RECT 193.64 64.17 193.85 64.24 ;
    RECT 193.18 63.45 193.39 63.52 ;
    RECT 193.18 63.81 193.39 63.88 ;
    RECT 193.18 64.17 193.39 64.24 ;
    RECT 190.32 63.45 190.53 63.52 ;
    RECT 190.32 63.81 190.53 63.88 ;
    RECT 190.32 64.17 190.53 64.24 ;
    RECT 189.86 63.45 190.07 63.52 ;
    RECT 189.86 63.81 190.07 63.88 ;
    RECT 189.86 64.17 190.07 64.24 ;
    RECT 187.0 63.45 187.21 63.52 ;
    RECT 187.0 63.81 187.21 63.88 ;
    RECT 187.0 64.17 187.21 64.24 ;
    RECT 186.54 63.45 186.75 63.52 ;
    RECT 186.54 63.81 186.75 63.88 ;
    RECT 186.54 64.17 186.75 64.24 ;
    RECT 183.68 63.45 183.89 63.52 ;
    RECT 183.68 63.81 183.89 63.88 ;
    RECT 183.68 64.17 183.89 64.24 ;
    RECT 183.22 63.45 183.43 63.52 ;
    RECT 183.22 63.81 183.43 63.88 ;
    RECT 183.22 64.17 183.43 64.24 ;
    RECT 147.485 63.81 147.555 63.88 ;
    RECT 266.68 63.45 266.89 63.52 ;
    RECT 266.68 63.81 266.89 63.88 ;
    RECT 266.68 64.17 266.89 64.24 ;
    RECT 266.22 63.45 266.43 63.52 ;
    RECT 266.22 63.81 266.43 63.88 ;
    RECT 266.22 64.17 266.43 64.24 ;
    RECT 263.36 63.45 263.57 63.52 ;
    RECT 263.36 63.81 263.57 63.88 ;
    RECT 263.36 64.17 263.57 64.24 ;
    RECT 262.9 63.45 263.11 63.52 ;
    RECT 262.9 63.81 263.11 63.88 ;
    RECT 262.9 64.17 263.11 64.24 ;
    RECT 260.04 63.45 260.25 63.52 ;
    RECT 260.04 63.81 260.25 63.88 ;
    RECT 260.04 64.17 260.25 64.24 ;
    RECT 259.58 63.45 259.79 63.52 ;
    RECT 259.58 63.81 259.79 63.88 ;
    RECT 259.58 64.17 259.79 64.24 ;
    RECT 256.72 63.45 256.93 63.52 ;
    RECT 256.72 63.81 256.93 63.88 ;
    RECT 256.72 64.17 256.93 64.24 ;
    RECT 256.26 63.45 256.47 63.52 ;
    RECT 256.26 63.81 256.47 63.88 ;
    RECT 256.26 64.17 256.47 64.24 ;
    RECT 253.4 63.45 253.61 63.52 ;
    RECT 253.4 63.81 253.61 63.88 ;
    RECT 253.4 64.17 253.61 64.24 ;
    RECT 252.94 63.45 253.15 63.52 ;
    RECT 252.94 63.81 253.15 63.88 ;
    RECT 252.94 64.17 253.15 64.24 ;
    RECT 250.08 55.51 250.29 55.58 ;
    RECT 250.08 55.87 250.29 55.94 ;
    RECT 250.08 56.23 250.29 56.3 ;
    RECT 249.62 55.51 249.83 55.58 ;
    RECT 249.62 55.87 249.83 55.94 ;
    RECT 249.62 56.23 249.83 56.3 ;
    RECT 267.91 55.87 267.98 55.94 ;
    RECT 246.76 55.51 246.97 55.58 ;
    RECT 246.76 55.87 246.97 55.94 ;
    RECT 246.76 56.23 246.97 56.3 ;
    RECT 246.3 55.51 246.51 55.58 ;
    RECT 246.3 55.87 246.51 55.94 ;
    RECT 246.3 56.23 246.51 56.3 ;
    RECT 243.44 55.51 243.65 55.58 ;
    RECT 243.44 55.87 243.65 55.94 ;
    RECT 243.44 56.23 243.65 56.3 ;
    RECT 242.98 55.51 243.19 55.58 ;
    RECT 242.98 55.87 243.19 55.94 ;
    RECT 242.98 56.23 243.19 56.3 ;
    RECT 240.12 55.51 240.33 55.58 ;
    RECT 240.12 55.87 240.33 55.94 ;
    RECT 240.12 56.23 240.33 56.3 ;
    RECT 239.66 55.51 239.87 55.58 ;
    RECT 239.66 55.87 239.87 55.94 ;
    RECT 239.66 56.23 239.87 56.3 ;
    RECT 236.8 55.51 237.01 55.58 ;
    RECT 236.8 55.87 237.01 55.94 ;
    RECT 236.8 56.23 237.01 56.3 ;
    RECT 236.34 55.51 236.55 55.58 ;
    RECT 236.34 55.87 236.55 55.94 ;
    RECT 236.34 56.23 236.55 56.3 ;
    RECT 233.48 55.51 233.69 55.58 ;
    RECT 233.48 55.87 233.69 55.94 ;
    RECT 233.48 56.23 233.69 56.3 ;
    RECT 233.02 55.51 233.23 55.58 ;
    RECT 233.02 55.87 233.23 55.94 ;
    RECT 233.02 56.23 233.23 56.3 ;
    RECT 230.16 55.51 230.37 55.58 ;
    RECT 230.16 55.87 230.37 55.94 ;
    RECT 230.16 56.23 230.37 56.3 ;
    RECT 229.7 55.51 229.91 55.58 ;
    RECT 229.7 55.87 229.91 55.94 ;
    RECT 229.7 56.23 229.91 56.3 ;
    RECT 226.84 55.51 227.05 55.58 ;
    RECT 226.84 55.87 227.05 55.94 ;
    RECT 226.84 56.23 227.05 56.3 ;
    RECT 226.38 55.51 226.59 55.58 ;
    RECT 226.38 55.87 226.59 55.94 ;
    RECT 226.38 56.23 226.59 56.3 ;
    RECT 223.52 55.51 223.73 55.58 ;
    RECT 223.52 55.87 223.73 55.94 ;
    RECT 223.52 56.23 223.73 56.3 ;
    RECT 223.06 55.51 223.27 55.58 ;
    RECT 223.06 55.87 223.27 55.94 ;
    RECT 223.06 56.23 223.27 56.3 ;
    RECT 220.2 55.51 220.41 55.58 ;
    RECT 220.2 55.87 220.41 55.94 ;
    RECT 220.2 56.23 220.41 56.3 ;
    RECT 219.74 55.51 219.95 55.58 ;
    RECT 219.74 55.87 219.95 55.94 ;
    RECT 219.74 56.23 219.95 56.3 ;
    RECT 216.88 55.51 217.09 55.58 ;
    RECT 216.88 55.87 217.09 55.94 ;
    RECT 216.88 56.23 217.09 56.3 ;
    RECT 216.42 55.51 216.63 55.58 ;
    RECT 216.42 55.87 216.63 55.94 ;
    RECT 216.42 56.23 216.63 56.3 ;
    RECT 180.36 55.51 180.57 55.58 ;
    RECT 180.36 55.87 180.57 55.94 ;
    RECT 180.36 56.23 180.57 56.3 ;
    RECT 179.9 55.51 180.11 55.58 ;
    RECT 179.9 55.87 180.11 55.94 ;
    RECT 179.9 56.23 180.11 56.3 ;
    RECT 177.04 55.51 177.25 55.58 ;
    RECT 177.04 55.87 177.25 55.94 ;
    RECT 177.04 56.23 177.25 56.3 ;
    RECT 176.58 55.51 176.79 55.58 ;
    RECT 176.58 55.87 176.79 55.94 ;
    RECT 176.58 56.23 176.79 56.3 ;
    RECT 173.72 55.51 173.93 55.58 ;
    RECT 173.72 55.87 173.93 55.94 ;
    RECT 173.72 56.23 173.93 56.3 ;
    RECT 173.26 55.51 173.47 55.58 ;
    RECT 173.26 55.87 173.47 55.94 ;
    RECT 173.26 56.23 173.47 56.3 ;
    RECT 170.4 55.51 170.61 55.58 ;
    RECT 170.4 55.87 170.61 55.94 ;
    RECT 170.4 56.23 170.61 56.3 ;
    RECT 169.94 55.51 170.15 55.58 ;
    RECT 169.94 55.87 170.15 55.94 ;
    RECT 169.94 56.23 170.15 56.3 ;
    RECT 167.08 55.51 167.29 55.58 ;
    RECT 167.08 55.87 167.29 55.94 ;
    RECT 167.08 56.23 167.29 56.3 ;
    RECT 166.62 55.51 166.83 55.58 ;
    RECT 166.62 55.87 166.83 55.94 ;
    RECT 166.62 56.23 166.83 56.3 ;
    RECT 163.76 55.51 163.97 55.58 ;
    RECT 163.76 55.87 163.97 55.94 ;
    RECT 163.76 56.23 163.97 56.3 ;
    RECT 163.3 55.51 163.51 55.58 ;
    RECT 163.3 55.87 163.51 55.94 ;
    RECT 163.3 56.23 163.51 56.3 ;
    RECT 160.44 55.51 160.65 55.58 ;
    RECT 160.44 55.87 160.65 55.94 ;
    RECT 160.44 56.23 160.65 56.3 ;
    RECT 159.98 55.51 160.19 55.58 ;
    RECT 159.98 55.87 160.19 55.94 ;
    RECT 159.98 56.23 160.19 56.3 ;
    RECT 157.12 55.51 157.33 55.58 ;
    RECT 157.12 55.87 157.33 55.94 ;
    RECT 157.12 56.23 157.33 56.3 ;
    RECT 156.66 55.51 156.87 55.58 ;
    RECT 156.66 55.87 156.87 55.94 ;
    RECT 156.66 56.23 156.87 56.3 ;
    RECT 153.8 55.51 154.01 55.58 ;
    RECT 153.8 55.87 154.01 55.94 ;
    RECT 153.8 56.23 154.01 56.3 ;
    RECT 153.34 55.51 153.55 55.58 ;
    RECT 153.34 55.87 153.55 55.94 ;
    RECT 153.34 56.23 153.55 56.3 ;
    RECT 150.48 55.51 150.69 55.58 ;
    RECT 150.48 55.87 150.69 55.94 ;
    RECT 150.48 56.23 150.69 56.3 ;
    RECT 150.02 55.51 150.23 55.58 ;
    RECT 150.02 55.87 150.23 55.94 ;
    RECT 150.02 56.23 150.23 56.3 ;
    RECT 213.56 55.51 213.77 55.58 ;
    RECT 213.56 55.87 213.77 55.94 ;
    RECT 213.56 56.23 213.77 56.3 ;
    RECT 213.1 55.51 213.31 55.58 ;
    RECT 213.1 55.87 213.31 55.94 ;
    RECT 213.1 56.23 213.31 56.3 ;
    RECT 210.24 55.51 210.45 55.58 ;
    RECT 210.24 55.87 210.45 55.94 ;
    RECT 210.24 56.23 210.45 56.3 ;
    RECT 209.78 55.51 209.99 55.58 ;
    RECT 209.78 55.87 209.99 55.94 ;
    RECT 209.78 56.23 209.99 56.3 ;
    RECT 206.92 55.51 207.13 55.58 ;
    RECT 206.92 55.87 207.13 55.94 ;
    RECT 206.92 56.23 207.13 56.3 ;
    RECT 206.46 55.51 206.67 55.58 ;
    RECT 206.46 55.87 206.67 55.94 ;
    RECT 206.46 56.23 206.67 56.3 ;
    RECT 203.6 55.51 203.81 55.58 ;
    RECT 203.6 55.87 203.81 55.94 ;
    RECT 203.6 56.23 203.81 56.3 ;
    RECT 203.14 55.51 203.35 55.58 ;
    RECT 203.14 55.87 203.35 55.94 ;
    RECT 203.14 56.23 203.35 56.3 ;
    RECT 200.28 55.51 200.49 55.58 ;
    RECT 200.28 55.87 200.49 55.94 ;
    RECT 200.28 56.23 200.49 56.3 ;
    RECT 199.82 55.51 200.03 55.58 ;
    RECT 199.82 55.87 200.03 55.94 ;
    RECT 199.82 56.23 200.03 56.3 ;
    RECT 147.485 55.87 147.555 55.94 ;
    RECT 196.96 55.51 197.17 55.58 ;
    RECT 196.96 55.87 197.17 55.94 ;
    RECT 196.96 56.23 197.17 56.3 ;
    RECT 196.5 55.51 196.71 55.58 ;
    RECT 196.5 55.87 196.71 55.94 ;
    RECT 196.5 56.23 196.71 56.3 ;
    RECT 193.64 55.51 193.85 55.58 ;
    RECT 193.64 55.87 193.85 55.94 ;
    RECT 193.64 56.23 193.85 56.3 ;
    RECT 193.18 55.51 193.39 55.58 ;
    RECT 193.18 55.87 193.39 55.94 ;
    RECT 193.18 56.23 193.39 56.3 ;
    RECT 190.32 55.51 190.53 55.58 ;
    RECT 190.32 55.87 190.53 55.94 ;
    RECT 190.32 56.23 190.53 56.3 ;
    RECT 189.86 55.51 190.07 55.58 ;
    RECT 189.86 55.87 190.07 55.94 ;
    RECT 189.86 56.23 190.07 56.3 ;
    RECT 187.0 55.51 187.21 55.58 ;
    RECT 187.0 55.87 187.21 55.94 ;
    RECT 187.0 56.23 187.21 56.3 ;
    RECT 186.54 55.51 186.75 55.58 ;
    RECT 186.54 55.87 186.75 55.94 ;
    RECT 186.54 56.23 186.75 56.3 ;
    RECT 183.68 55.51 183.89 55.58 ;
    RECT 183.68 55.87 183.89 55.94 ;
    RECT 183.68 56.23 183.89 56.3 ;
    RECT 183.22 55.51 183.43 55.58 ;
    RECT 183.22 55.87 183.43 55.94 ;
    RECT 183.22 56.23 183.43 56.3 ;
    RECT 266.68 55.51 266.89 55.58 ;
    RECT 266.68 55.87 266.89 55.94 ;
    RECT 266.68 56.23 266.89 56.3 ;
    RECT 266.22 55.51 266.43 55.58 ;
    RECT 266.22 55.87 266.43 55.94 ;
    RECT 266.22 56.23 266.43 56.3 ;
    RECT 263.36 55.51 263.57 55.58 ;
    RECT 263.36 55.87 263.57 55.94 ;
    RECT 263.36 56.23 263.57 56.3 ;
    RECT 262.9 55.51 263.11 55.58 ;
    RECT 262.9 55.87 263.11 55.94 ;
    RECT 262.9 56.23 263.11 56.3 ;
    RECT 260.04 55.51 260.25 55.58 ;
    RECT 260.04 55.87 260.25 55.94 ;
    RECT 260.04 56.23 260.25 56.3 ;
    RECT 259.58 55.51 259.79 55.58 ;
    RECT 259.58 55.87 259.79 55.94 ;
    RECT 259.58 56.23 259.79 56.3 ;
    RECT 256.72 55.51 256.93 55.58 ;
    RECT 256.72 55.87 256.93 55.94 ;
    RECT 256.72 56.23 256.93 56.3 ;
    RECT 256.26 55.51 256.47 55.58 ;
    RECT 256.26 55.87 256.47 55.94 ;
    RECT 256.26 56.23 256.47 56.3 ;
    RECT 253.4 55.51 253.61 55.58 ;
    RECT 253.4 55.87 253.61 55.94 ;
    RECT 253.4 56.23 253.61 56.3 ;
    RECT 252.94 55.51 253.15 55.58 ;
    RECT 252.94 55.87 253.15 55.94 ;
    RECT 252.94 56.23 253.15 56.3 ;
    RECT 250.08 23.11 250.29 23.18 ;
    RECT 250.08 23.47 250.29 23.54 ;
    RECT 250.08 23.83 250.29 23.9 ;
    RECT 249.62 23.11 249.83 23.18 ;
    RECT 249.62 23.47 249.83 23.54 ;
    RECT 249.62 23.83 249.83 23.9 ;
    RECT 246.76 23.11 246.97 23.18 ;
    RECT 246.76 23.47 246.97 23.54 ;
    RECT 246.76 23.83 246.97 23.9 ;
    RECT 246.3 23.11 246.51 23.18 ;
    RECT 246.3 23.47 246.51 23.54 ;
    RECT 246.3 23.83 246.51 23.9 ;
    RECT 243.44 23.11 243.65 23.18 ;
    RECT 243.44 23.47 243.65 23.54 ;
    RECT 243.44 23.83 243.65 23.9 ;
    RECT 242.98 23.11 243.19 23.18 ;
    RECT 242.98 23.47 243.19 23.54 ;
    RECT 242.98 23.83 243.19 23.9 ;
    RECT 240.12 23.11 240.33 23.18 ;
    RECT 240.12 23.47 240.33 23.54 ;
    RECT 240.12 23.83 240.33 23.9 ;
    RECT 239.66 23.11 239.87 23.18 ;
    RECT 239.66 23.47 239.87 23.54 ;
    RECT 239.66 23.83 239.87 23.9 ;
    RECT 236.8 23.11 237.01 23.18 ;
    RECT 236.8 23.47 237.01 23.54 ;
    RECT 236.8 23.83 237.01 23.9 ;
    RECT 236.34 23.11 236.55 23.18 ;
    RECT 236.34 23.47 236.55 23.54 ;
    RECT 236.34 23.83 236.55 23.9 ;
    RECT 233.48 23.11 233.69 23.18 ;
    RECT 233.48 23.47 233.69 23.54 ;
    RECT 233.48 23.83 233.69 23.9 ;
    RECT 233.02 23.11 233.23 23.18 ;
    RECT 233.02 23.47 233.23 23.54 ;
    RECT 233.02 23.83 233.23 23.9 ;
    RECT 230.16 23.11 230.37 23.18 ;
    RECT 230.16 23.47 230.37 23.54 ;
    RECT 230.16 23.83 230.37 23.9 ;
    RECT 229.7 23.11 229.91 23.18 ;
    RECT 229.7 23.47 229.91 23.54 ;
    RECT 229.7 23.83 229.91 23.9 ;
    RECT 226.84 23.11 227.05 23.18 ;
    RECT 226.84 23.47 227.05 23.54 ;
    RECT 226.84 23.83 227.05 23.9 ;
    RECT 226.38 23.11 226.59 23.18 ;
    RECT 226.38 23.47 226.59 23.54 ;
    RECT 226.38 23.83 226.59 23.9 ;
    RECT 223.52 23.11 223.73 23.18 ;
    RECT 223.52 23.47 223.73 23.54 ;
    RECT 223.52 23.83 223.73 23.9 ;
    RECT 223.06 23.11 223.27 23.18 ;
    RECT 223.06 23.47 223.27 23.54 ;
    RECT 223.06 23.83 223.27 23.9 ;
    RECT 220.2 23.11 220.41 23.18 ;
    RECT 220.2 23.47 220.41 23.54 ;
    RECT 220.2 23.83 220.41 23.9 ;
    RECT 219.74 23.11 219.95 23.18 ;
    RECT 219.74 23.47 219.95 23.54 ;
    RECT 219.74 23.83 219.95 23.9 ;
    RECT 216.88 23.11 217.09 23.18 ;
    RECT 216.88 23.47 217.09 23.54 ;
    RECT 216.88 23.83 217.09 23.9 ;
    RECT 216.42 23.11 216.63 23.18 ;
    RECT 216.42 23.47 216.63 23.54 ;
    RECT 216.42 23.83 216.63 23.9 ;
    RECT 267.91 23.47 267.98 23.54 ;
    RECT 180.36 23.11 180.57 23.18 ;
    RECT 180.36 23.47 180.57 23.54 ;
    RECT 180.36 23.83 180.57 23.9 ;
    RECT 179.9 23.11 180.11 23.18 ;
    RECT 179.9 23.47 180.11 23.54 ;
    RECT 179.9 23.83 180.11 23.9 ;
    RECT 177.04 23.11 177.25 23.18 ;
    RECT 177.04 23.47 177.25 23.54 ;
    RECT 177.04 23.83 177.25 23.9 ;
    RECT 176.58 23.11 176.79 23.18 ;
    RECT 176.58 23.47 176.79 23.54 ;
    RECT 176.58 23.83 176.79 23.9 ;
    RECT 173.72 23.11 173.93 23.18 ;
    RECT 173.72 23.47 173.93 23.54 ;
    RECT 173.72 23.83 173.93 23.9 ;
    RECT 173.26 23.11 173.47 23.18 ;
    RECT 173.26 23.47 173.47 23.54 ;
    RECT 173.26 23.83 173.47 23.9 ;
    RECT 170.4 23.11 170.61 23.18 ;
    RECT 170.4 23.47 170.61 23.54 ;
    RECT 170.4 23.83 170.61 23.9 ;
    RECT 169.94 23.11 170.15 23.18 ;
    RECT 169.94 23.47 170.15 23.54 ;
    RECT 169.94 23.83 170.15 23.9 ;
    RECT 167.08 23.11 167.29 23.18 ;
    RECT 167.08 23.47 167.29 23.54 ;
    RECT 167.08 23.83 167.29 23.9 ;
    RECT 166.62 23.11 166.83 23.18 ;
    RECT 166.62 23.47 166.83 23.54 ;
    RECT 166.62 23.83 166.83 23.9 ;
    RECT 163.76 23.11 163.97 23.18 ;
    RECT 163.76 23.47 163.97 23.54 ;
    RECT 163.76 23.83 163.97 23.9 ;
    RECT 163.3 23.11 163.51 23.18 ;
    RECT 163.3 23.47 163.51 23.54 ;
    RECT 163.3 23.83 163.51 23.9 ;
    RECT 160.44 23.11 160.65 23.18 ;
    RECT 160.44 23.47 160.65 23.54 ;
    RECT 160.44 23.83 160.65 23.9 ;
    RECT 159.98 23.11 160.19 23.18 ;
    RECT 159.98 23.47 160.19 23.54 ;
    RECT 159.98 23.83 160.19 23.9 ;
    RECT 157.12 23.11 157.33 23.18 ;
    RECT 157.12 23.47 157.33 23.54 ;
    RECT 157.12 23.83 157.33 23.9 ;
    RECT 156.66 23.11 156.87 23.18 ;
    RECT 156.66 23.47 156.87 23.54 ;
    RECT 156.66 23.83 156.87 23.9 ;
    RECT 153.8 23.11 154.01 23.18 ;
    RECT 153.8 23.47 154.01 23.54 ;
    RECT 153.8 23.83 154.01 23.9 ;
    RECT 153.34 23.11 153.55 23.18 ;
    RECT 153.34 23.47 153.55 23.54 ;
    RECT 153.34 23.83 153.55 23.9 ;
    RECT 150.48 23.11 150.69 23.18 ;
    RECT 150.48 23.47 150.69 23.54 ;
    RECT 150.48 23.83 150.69 23.9 ;
    RECT 150.02 23.11 150.23 23.18 ;
    RECT 150.02 23.47 150.23 23.54 ;
    RECT 150.02 23.83 150.23 23.9 ;
    RECT 213.56 23.11 213.77 23.18 ;
    RECT 213.56 23.47 213.77 23.54 ;
    RECT 213.56 23.83 213.77 23.9 ;
    RECT 213.1 23.11 213.31 23.18 ;
    RECT 213.1 23.47 213.31 23.54 ;
    RECT 213.1 23.83 213.31 23.9 ;
    RECT 210.24 23.11 210.45 23.18 ;
    RECT 210.24 23.47 210.45 23.54 ;
    RECT 210.24 23.83 210.45 23.9 ;
    RECT 209.78 23.11 209.99 23.18 ;
    RECT 209.78 23.47 209.99 23.54 ;
    RECT 209.78 23.83 209.99 23.9 ;
    RECT 206.92 23.11 207.13 23.18 ;
    RECT 206.92 23.47 207.13 23.54 ;
    RECT 206.92 23.83 207.13 23.9 ;
    RECT 206.46 23.11 206.67 23.18 ;
    RECT 206.46 23.47 206.67 23.54 ;
    RECT 206.46 23.83 206.67 23.9 ;
    RECT 203.6 23.11 203.81 23.18 ;
    RECT 203.6 23.47 203.81 23.54 ;
    RECT 203.6 23.83 203.81 23.9 ;
    RECT 203.14 23.11 203.35 23.18 ;
    RECT 203.14 23.47 203.35 23.54 ;
    RECT 203.14 23.83 203.35 23.9 ;
    RECT 200.28 23.11 200.49 23.18 ;
    RECT 200.28 23.47 200.49 23.54 ;
    RECT 200.28 23.83 200.49 23.9 ;
    RECT 199.82 23.11 200.03 23.18 ;
    RECT 199.82 23.47 200.03 23.54 ;
    RECT 199.82 23.83 200.03 23.9 ;
    RECT 196.96 23.11 197.17 23.18 ;
    RECT 196.96 23.47 197.17 23.54 ;
    RECT 196.96 23.83 197.17 23.9 ;
    RECT 196.5 23.11 196.71 23.18 ;
    RECT 196.5 23.47 196.71 23.54 ;
    RECT 196.5 23.83 196.71 23.9 ;
    RECT 193.64 23.11 193.85 23.18 ;
    RECT 193.64 23.47 193.85 23.54 ;
    RECT 193.64 23.83 193.85 23.9 ;
    RECT 193.18 23.11 193.39 23.18 ;
    RECT 193.18 23.47 193.39 23.54 ;
    RECT 193.18 23.83 193.39 23.9 ;
    RECT 190.32 23.11 190.53 23.18 ;
    RECT 190.32 23.47 190.53 23.54 ;
    RECT 190.32 23.83 190.53 23.9 ;
    RECT 189.86 23.11 190.07 23.18 ;
    RECT 189.86 23.47 190.07 23.54 ;
    RECT 189.86 23.83 190.07 23.9 ;
    RECT 187.0 23.11 187.21 23.18 ;
    RECT 187.0 23.47 187.21 23.54 ;
    RECT 187.0 23.83 187.21 23.9 ;
    RECT 186.54 23.11 186.75 23.18 ;
    RECT 186.54 23.47 186.75 23.54 ;
    RECT 186.54 23.83 186.75 23.9 ;
    RECT 183.68 23.11 183.89 23.18 ;
    RECT 183.68 23.47 183.89 23.54 ;
    RECT 183.68 23.83 183.89 23.9 ;
    RECT 183.22 23.11 183.43 23.18 ;
    RECT 183.22 23.47 183.43 23.54 ;
    RECT 183.22 23.83 183.43 23.9 ;
    RECT 147.485 23.47 147.555 23.54 ;
    RECT 266.68 23.11 266.89 23.18 ;
    RECT 266.68 23.47 266.89 23.54 ;
    RECT 266.68 23.83 266.89 23.9 ;
    RECT 266.22 23.11 266.43 23.18 ;
    RECT 266.22 23.47 266.43 23.54 ;
    RECT 266.22 23.83 266.43 23.9 ;
    RECT 263.36 23.11 263.57 23.18 ;
    RECT 263.36 23.47 263.57 23.54 ;
    RECT 263.36 23.83 263.57 23.9 ;
    RECT 262.9 23.11 263.11 23.18 ;
    RECT 262.9 23.47 263.11 23.54 ;
    RECT 262.9 23.83 263.11 23.9 ;
    RECT 260.04 23.11 260.25 23.18 ;
    RECT 260.04 23.47 260.25 23.54 ;
    RECT 260.04 23.83 260.25 23.9 ;
    RECT 259.58 23.11 259.79 23.18 ;
    RECT 259.58 23.47 259.79 23.54 ;
    RECT 259.58 23.83 259.79 23.9 ;
    RECT 256.72 23.11 256.93 23.18 ;
    RECT 256.72 23.47 256.93 23.54 ;
    RECT 256.72 23.83 256.93 23.9 ;
    RECT 256.26 23.11 256.47 23.18 ;
    RECT 256.26 23.47 256.47 23.54 ;
    RECT 256.26 23.83 256.47 23.9 ;
    RECT 253.4 23.11 253.61 23.18 ;
    RECT 253.4 23.47 253.61 23.54 ;
    RECT 253.4 23.83 253.61 23.9 ;
    RECT 252.94 23.11 253.15 23.18 ;
    RECT 252.94 23.47 253.15 23.54 ;
    RECT 252.94 23.83 253.15 23.9 ;
    RECT 250.08 62.73 250.29 62.8 ;
    RECT 250.08 63.09 250.29 63.16 ;
    RECT 250.08 63.45 250.29 63.52 ;
    RECT 249.62 62.73 249.83 62.8 ;
    RECT 249.62 63.09 249.83 63.16 ;
    RECT 249.62 63.45 249.83 63.52 ;
    RECT 246.76 62.73 246.97 62.8 ;
    RECT 246.76 63.09 246.97 63.16 ;
    RECT 246.76 63.45 246.97 63.52 ;
    RECT 246.3 62.73 246.51 62.8 ;
    RECT 246.3 63.09 246.51 63.16 ;
    RECT 246.3 63.45 246.51 63.52 ;
    RECT 243.44 62.73 243.65 62.8 ;
    RECT 243.44 63.09 243.65 63.16 ;
    RECT 243.44 63.45 243.65 63.52 ;
    RECT 242.98 62.73 243.19 62.8 ;
    RECT 242.98 63.09 243.19 63.16 ;
    RECT 242.98 63.45 243.19 63.52 ;
    RECT 240.12 62.73 240.33 62.8 ;
    RECT 240.12 63.09 240.33 63.16 ;
    RECT 240.12 63.45 240.33 63.52 ;
    RECT 239.66 62.73 239.87 62.8 ;
    RECT 239.66 63.09 239.87 63.16 ;
    RECT 239.66 63.45 239.87 63.52 ;
    RECT 236.8 62.73 237.01 62.8 ;
    RECT 236.8 63.09 237.01 63.16 ;
    RECT 236.8 63.45 237.01 63.52 ;
    RECT 236.34 62.73 236.55 62.8 ;
    RECT 236.34 63.09 236.55 63.16 ;
    RECT 236.34 63.45 236.55 63.52 ;
    RECT 233.48 62.73 233.69 62.8 ;
    RECT 233.48 63.09 233.69 63.16 ;
    RECT 233.48 63.45 233.69 63.52 ;
    RECT 233.02 62.73 233.23 62.8 ;
    RECT 233.02 63.09 233.23 63.16 ;
    RECT 233.02 63.45 233.23 63.52 ;
    RECT 230.16 62.73 230.37 62.8 ;
    RECT 230.16 63.09 230.37 63.16 ;
    RECT 230.16 63.45 230.37 63.52 ;
    RECT 229.7 62.73 229.91 62.8 ;
    RECT 229.7 63.09 229.91 63.16 ;
    RECT 229.7 63.45 229.91 63.52 ;
    RECT 226.84 62.73 227.05 62.8 ;
    RECT 226.84 63.09 227.05 63.16 ;
    RECT 226.84 63.45 227.05 63.52 ;
    RECT 226.38 62.73 226.59 62.8 ;
    RECT 226.38 63.09 226.59 63.16 ;
    RECT 226.38 63.45 226.59 63.52 ;
    RECT 223.52 62.73 223.73 62.8 ;
    RECT 223.52 63.09 223.73 63.16 ;
    RECT 223.52 63.45 223.73 63.52 ;
    RECT 223.06 62.73 223.27 62.8 ;
    RECT 223.06 63.09 223.27 63.16 ;
    RECT 223.06 63.45 223.27 63.52 ;
    RECT 220.2 62.73 220.41 62.8 ;
    RECT 220.2 63.09 220.41 63.16 ;
    RECT 220.2 63.45 220.41 63.52 ;
    RECT 219.74 62.73 219.95 62.8 ;
    RECT 219.74 63.09 219.95 63.16 ;
    RECT 219.74 63.45 219.95 63.52 ;
    RECT 216.88 62.73 217.09 62.8 ;
    RECT 216.88 63.09 217.09 63.16 ;
    RECT 216.88 63.45 217.09 63.52 ;
    RECT 216.42 62.73 216.63 62.8 ;
    RECT 216.42 63.09 216.63 63.16 ;
    RECT 216.42 63.45 216.63 63.52 ;
    RECT 267.91 63.09 267.98 63.16 ;
    RECT 180.36 62.73 180.57 62.8 ;
    RECT 180.36 63.09 180.57 63.16 ;
    RECT 180.36 63.45 180.57 63.52 ;
    RECT 179.9 62.73 180.11 62.8 ;
    RECT 179.9 63.09 180.11 63.16 ;
    RECT 179.9 63.45 180.11 63.52 ;
    RECT 177.04 62.73 177.25 62.8 ;
    RECT 177.04 63.09 177.25 63.16 ;
    RECT 177.04 63.45 177.25 63.52 ;
    RECT 176.58 62.73 176.79 62.8 ;
    RECT 176.58 63.09 176.79 63.16 ;
    RECT 176.58 63.45 176.79 63.52 ;
    RECT 173.72 62.73 173.93 62.8 ;
    RECT 173.72 63.09 173.93 63.16 ;
    RECT 173.72 63.45 173.93 63.52 ;
    RECT 173.26 62.73 173.47 62.8 ;
    RECT 173.26 63.09 173.47 63.16 ;
    RECT 173.26 63.45 173.47 63.52 ;
    RECT 170.4 62.73 170.61 62.8 ;
    RECT 170.4 63.09 170.61 63.16 ;
    RECT 170.4 63.45 170.61 63.52 ;
    RECT 169.94 62.73 170.15 62.8 ;
    RECT 169.94 63.09 170.15 63.16 ;
    RECT 169.94 63.45 170.15 63.52 ;
    RECT 167.08 62.73 167.29 62.8 ;
    RECT 167.08 63.09 167.29 63.16 ;
    RECT 167.08 63.45 167.29 63.52 ;
    RECT 166.62 62.73 166.83 62.8 ;
    RECT 166.62 63.09 166.83 63.16 ;
    RECT 166.62 63.45 166.83 63.52 ;
    RECT 163.76 62.73 163.97 62.8 ;
    RECT 163.76 63.09 163.97 63.16 ;
    RECT 163.76 63.45 163.97 63.52 ;
    RECT 163.3 62.73 163.51 62.8 ;
    RECT 163.3 63.09 163.51 63.16 ;
    RECT 163.3 63.45 163.51 63.52 ;
    RECT 160.44 62.73 160.65 62.8 ;
    RECT 160.44 63.09 160.65 63.16 ;
    RECT 160.44 63.45 160.65 63.52 ;
    RECT 159.98 62.73 160.19 62.8 ;
    RECT 159.98 63.09 160.19 63.16 ;
    RECT 159.98 63.45 160.19 63.52 ;
    RECT 157.12 62.73 157.33 62.8 ;
    RECT 157.12 63.09 157.33 63.16 ;
    RECT 157.12 63.45 157.33 63.52 ;
    RECT 156.66 62.73 156.87 62.8 ;
    RECT 156.66 63.09 156.87 63.16 ;
    RECT 156.66 63.45 156.87 63.52 ;
    RECT 153.8 62.73 154.01 62.8 ;
    RECT 153.8 63.09 154.01 63.16 ;
    RECT 153.8 63.45 154.01 63.52 ;
    RECT 153.34 62.73 153.55 62.8 ;
    RECT 153.34 63.09 153.55 63.16 ;
    RECT 153.34 63.45 153.55 63.52 ;
    RECT 150.48 62.73 150.69 62.8 ;
    RECT 150.48 63.09 150.69 63.16 ;
    RECT 150.48 63.45 150.69 63.52 ;
    RECT 150.02 62.73 150.23 62.8 ;
    RECT 150.02 63.09 150.23 63.16 ;
    RECT 150.02 63.45 150.23 63.52 ;
    RECT 213.56 62.73 213.77 62.8 ;
    RECT 213.56 63.09 213.77 63.16 ;
    RECT 213.56 63.45 213.77 63.52 ;
    RECT 213.1 62.73 213.31 62.8 ;
    RECT 213.1 63.09 213.31 63.16 ;
    RECT 213.1 63.45 213.31 63.52 ;
    RECT 210.24 62.73 210.45 62.8 ;
    RECT 210.24 63.09 210.45 63.16 ;
    RECT 210.24 63.45 210.45 63.52 ;
    RECT 209.78 62.73 209.99 62.8 ;
    RECT 209.78 63.09 209.99 63.16 ;
    RECT 209.78 63.45 209.99 63.52 ;
    RECT 206.92 62.73 207.13 62.8 ;
    RECT 206.92 63.09 207.13 63.16 ;
    RECT 206.92 63.45 207.13 63.52 ;
    RECT 206.46 62.73 206.67 62.8 ;
    RECT 206.46 63.09 206.67 63.16 ;
    RECT 206.46 63.45 206.67 63.52 ;
    RECT 203.6 62.73 203.81 62.8 ;
    RECT 203.6 63.09 203.81 63.16 ;
    RECT 203.6 63.45 203.81 63.52 ;
    RECT 203.14 62.73 203.35 62.8 ;
    RECT 203.14 63.09 203.35 63.16 ;
    RECT 203.14 63.45 203.35 63.52 ;
    RECT 200.28 62.73 200.49 62.8 ;
    RECT 200.28 63.09 200.49 63.16 ;
    RECT 200.28 63.45 200.49 63.52 ;
    RECT 199.82 62.73 200.03 62.8 ;
    RECT 199.82 63.09 200.03 63.16 ;
    RECT 199.82 63.45 200.03 63.52 ;
    RECT 196.96 62.73 197.17 62.8 ;
    RECT 196.96 63.09 197.17 63.16 ;
    RECT 196.96 63.45 197.17 63.52 ;
    RECT 196.5 62.73 196.71 62.8 ;
    RECT 196.5 63.09 196.71 63.16 ;
    RECT 196.5 63.45 196.71 63.52 ;
    RECT 193.64 62.73 193.85 62.8 ;
    RECT 193.64 63.09 193.85 63.16 ;
    RECT 193.64 63.45 193.85 63.52 ;
    RECT 193.18 62.73 193.39 62.8 ;
    RECT 193.18 63.09 193.39 63.16 ;
    RECT 193.18 63.45 193.39 63.52 ;
    RECT 190.32 62.73 190.53 62.8 ;
    RECT 190.32 63.09 190.53 63.16 ;
    RECT 190.32 63.45 190.53 63.52 ;
    RECT 189.86 62.73 190.07 62.8 ;
    RECT 189.86 63.09 190.07 63.16 ;
    RECT 189.86 63.45 190.07 63.52 ;
    RECT 187.0 62.73 187.21 62.8 ;
    RECT 187.0 63.09 187.21 63.16 ;
    RECT 187.0 63.45 187.21 63.52 ;
    RECT 186.54 62.73 186.75 62.8 ;
    RECT 186.54 63.09 186.75 63.16 ;
    RECT 186.54 63.45 186.75 63.52 ;
    RECT 183.68 62.73 183.89 62.8 ;
    RECT 183.68 63.09 183.89 63.16 ;
    RECT 183.68 63.45 183.89 63.52 ;
    RECT 183.22 62.73 183.43 62.8 ;
    RECT 183.22 63.09 183.43 63.16 ;
    RECT 183.22 63.45 183.43 63.52 ;
    RECT 147.485 63.09 147.555 63.16 ;
    RECT 266.68 62.73 266.89 62.8 ;
    RECT 266.68 63.09 266.89 63.16 ;
    RECT 266.68 63.45 266.89 63.52 ;
    RECT 266.22 62.73 266.43 62.8 ;
    RECT 266.22 63.09 266.43 63.16 ;
    RECT 266.22 63.45 266.43 63.52 ;
    RECT 263.36 62.73 263.57 62.8 ;
    RECT 263.36 63.09 263.57 63.16 ;
    RECT 263.36 63.45 263.57 63.52 ;
    RECT 262.9 62.73 263.11 62.8 ;
    RECT 262.9 63.09 263.11 63.16 ;
    RECT 262.9 63.45 263.11 63.52 ;
    RECT 260.04 62.73 260.25 62.8 ;
    RECT 260.04 63.09 260.25 63.16 ;
    RECT 260.04 63.45 260.25 63.52 ;
    RECT 259.58 62.73 259.79 62.8 ;
    RECT 259.58 63.09 259.79 63.16 ;
    RECT 259.58 63.45 259.79 63.52 ;
    RECT 256.72 62.73 256.93 62.8 ;
    RECT 256.72 63.09 256.93 63.16 ;
    RECT 256.72 63.45 256.93 63.52 ;
    RECT 256.26 62.73 256.47 62.8 ;
    RECT 256.26 63.09 256.47 63.16 ;
    RECT 256.26 63.45 256.47 63.52 ;
    RECT 253.4 62.73 253.61 62.8 ;
    RECT 253.4 63.09 253.61 63.16 ;
    RECT 253.4 63.45 253.61 63.52 ;
    RECT 252.94 62.73 253.15 62.8 ;
    RECT 252.94 63.09 253.15 63.16 ;
    RECT 252.94 63.45 253.15 63.52 ;
    RECT 250.08 54.79 250.29 54.86 ;
    RECT 250.08 55.15 250.29 55.22 ;
    RECT 250.08 55.51 250.29 55.58 ;
    RECT 249.62 54.79 249.83 54.86 ;
    RECT 249.62 55.15 249.83 55.22 ;
    RECT 249.62 55.51 249.83 55.58 ;
    RECT 246.76 54.79 246.97 54.86 ;
    RECT 246.76 55.15 246.97 55.22 ;
    RECT 246.76 55.51 246.97 55.58 ;
    RECT 246.3 54.79 246.51 54.86 ;
    RECT 246.3 55.15 246.51 55.22 ;
    RECT 246.3 55.51 246.51 55.58 ;
    RECT 243.44 54.79 243.65 54.86 ;
    RECT 243.44 55.15 243.65 55.22 ;
    RECT 243.44 55.51 243.65 55.58 ;
    RECT 242.98 54.79 243.19 54.86 ;
    RECT 242.98 55.15 243.19 55.22 ;
    RECT 242.98 55.51 243.19 55.58 ;
    RECT 240.12 54.79 240.33 54.86 ;
    RECT 240.12 55.15 240.33 55.22 ;
    RECT 240.12 55.51 240.33 55.58 ;
    RECT 239.66 54.79 239.87 54.86 ;
    RECT 239.66 55.15 239.87 55.22 ;
    RECT 239.66 55.51 239.87 55.58 ;
    RECT 236.8 54.79 237.01 54.86 ;
    RECT 236.8 55.15 237.01 55.22 ;
    RECT 236.8 55.51 237.01 55.58 ;
    RECT 236.34 54.79 236.55 54.86 ;
    RECT 236.34 55.15 236.55 55.22 ;
    RECT 236.34 55.51 236.55 55.58 ;
    RECT 233.48 54.79 233.69 54.86 ;
    RECT 233.48 55.15 233.69 55.22 ;
    RECT 233.48 55.51 233.69 55.58 ;
    RECT 233.02 54.79 233.23 54.86 ;
    RECT 233.02 55.15 233.23 55.22 ;
    RECT 233.02 55.51 233.23 55.58 ;
    RECT 230.16 54.79 230.37 54.86 ;
    RECT 230.16 55.15 230.37 55.22 ;
    RECT 230.16 55.51 230.37 55.58 ;
    RECT 229.7 54.79 229.91 54.86 ;
    RECT 229.7 55.15 229.91 55.22 ;
    RECT 229.7 55.51 229.91 55.58 ;
    RECT 226.84 54.79 227.05 54.86 ;
    RECT 226.84 55.15 227.05 55.22 ;
    RECT 226.84 55.51 227.05 55.58 ;
    RECT 226.38 54.79 226.59 54.86 ;
    RECT 226.38 55.15 226.59 55.22 ;
    RECT 226.38 55.51 226.59 55.58 ;
    RECT 223.52 54.79 223.73 54.86 ;
    RECT 223.52 55.15 223.73 55.22 ;
    RECT 223.52 55.51 223.73 55.58 ;
    RECT 223.06 54.79 223.27 54.86 ;
    RECT 223.06 55.15 223.27 55.22 ;
    RECT 223.06 55.51 223.27 55.58 ;
    RECT 220.2 54.79 220.41 54.86 ;
    RECT 220.2 55.15 220.41 55.22 ;
    RECT 220.2 55.51 220.41 55.58 ;
    RECT 219.74 54.79 219.95 54.86 ;
    RECT 219.74 55.15 219.95 55.22 ;
    RECT 219.74 55.51 219.95 55.58 ;
    RECT 216.88 54.79 217.09 54.86 ;
    RECT 216.88 55.15 217.09 55.22 ;
    RECT 216.88 55.51 217.09 55.58 ;
    RECT 216.42 54.79 216.63 54.86 ;
    RECT 216.42 55.15 216.63 55.22 ;
    RECT 216.42 55.51 216.63 55.58 ;
    RECT 267.91 55.15 267.98 55.22 ;
    RECT 180.36 54.79 180.57 54.86 ;
    RECT 180.36 55.15 180.57 55.22 ;
    RECT 180.36 55.51 180.57 55.58 ;
    RECT 179.9 54.79 180.11 54.86 ;
    RECT 179.9 55.15 180.11 55.22 ;
    RECT 179.9 55.51 180.11 55.58 ;
    RECT 177.04 54.79 177.25 54.86 ;
    RECT 177.04 55.15 177.25 55.22 ;
    RECT 177.04 55.51 177.25 55.58 ;
    RECT 176.58 54.79 176.79 54.86 ;
    RECT 176.58 55.15 176.79 55.22 ;
    RECT 176.58 55.51 176.79 55.58 ;
    RECT 173.72 54.79 173.93 54.86 ;
    RECT 173.72 55.15 173.93 55.22 ;
    RECT 173.72 55.51 173.93 55.58 ;
    RECT 173.26 54.79 173.47 54.86 ;
    RECT 173.26 55.15 173.47 55.22 ;
    RECT 173.26 55.51 173.47 55.58 ;
    RECT 170.4 54.79 170.61 54.86 ;
    RECT 170.4 55.15 170.61 55.22 ;
    RECT 170.4 55.51 170.61 55.58 ;
    RECT 169.94 54.79 170.15 54.86 ;
    RECT 169.94 55.15 170.15 55.22 ;
    RECT 169.94 55.51 170.15 55.58 ;
    RECT 167.08 54.79 167.29 54.86 ;
    RECT 167.08 55.15 167.29 55.22 ;
    RECT 167.08 55.51 167.29 55.58 ;
    RECT 166.62 54.79 166.83 54.86 ;
    RECT 166.62 55.15 166.83 55.22 ;
    RECT 166.62 55.51 166.83 55.58 ;
    RECT 163.76 54.79 163.97 54.86 ;
    RECT 163.76 55.15 163.97 55.22 ;
    RECT 163.76 55.51 163.97 55.58 ;
    RECT 163.3 54.79 163.51 54.86 ;
    RECT 163.3 55.15 163.51 55.22 ;
    RECT 163.3 55.51 163.51 55.58 ;
    RECT 160.44 54.79 160.65 54.86 ;
    RECT 160.44 55.15 160.65 55.22 ;
    RECT 160.44 55.51 160.65 55.58 ;
    RECT 159.98 54.79 160.19 54.86 ;
    RECT 159.98 55.15 160.19 55.22 ;
    RECT 159.98 55.51 160.19 55.58 ;
    RECT 157.12 54.79 157.33 54.86 ;
    RECT 157.12 55.15 157.33 55.22 ;
    RECT 157.12 55.51 157.33 55.58 ;
    RECT 156.66 54.79 156.87 54.86 ;
    RECT 156.66 55.15 156.87 55.22 ;
    RECT 156.66 55.51 156.87 55.58 ;
    RECT 153.8 54.79 154.01 54.86 ;
    RECT 153.8 55.15 154.01 55.22 ;
    RECT 153.8 55.51 154.01 55.58 ;
    RECT 153.34 54.79 153.55 54.86 ;
    RECT 153.34 55.15 153.55 55.22 ;
    RECT 153.34 55.51 153.55 55.58 ;
    RECT 150.48 54.79 150.69 54.86 ;
    RECT 150.48 55.15 150.69 55.22 ;
    RECT 150.48 55.51 150.69 55.58 ;
    RECT 150.02 54.79 150.23 54.86 ;
    RECT 150.02 55.15 150.23 55.22 ;
    RECT 150.02 55.51 150.23 55.58 ;
    RECT 213.56 54.79 213.77 54.86 ;
    RECT 213.56 55.15 213.77 55.22 ;
    RECT 213.56 55.51 213.77 55.58 ;
    RECT 213.1 54.79 213.31 54.86 ;
    RECT 213.1 55.15 213.31 55.22 ;
    RECT 213.1 55.51 213.31 55.58 ;
    RECT 210.24 54.79 210.45 54.86 ;
    RECT 210.24 55.15 210.45 55.22 ;
    RECT 210.24 55.51 210.45 55.58 ;
    RECT 209.78 54.79 209.99 54.86 ;
    RECT 209.78 55.15 209.99 55.22 ;
    RECT 209.78 55.51 209.99 55.58 ;
    RECT 206.92 54.79 207.13 54.86 ;
    RECT 206.92 55.15 207.13 55.22 ;
    RECT 206.92 55.51 207.13 55.58 ;
    RECT 206.46 54.79 206.67 54.86 ;
    RECT 206.46 55.15 206.67 55.22 ;
    RECT 206.46 55.51 206.67 55.58 ;
    RECT 203.6 54.79 203.81 54.86 ;
    RECT 203.6 55.15 203.81 55.22 ;
    RECT 203.6 55.51 203.81 55.58 ;
    RECT 203.14 54.79 203.35 54.86 ;
    RECT 203.14 55.15 203.35 55.22 ;
    RECT 203.14 55.51 203.35 55.58 ;
    RECT 200.28 54.79 200.49 54.86 ;
    RECT 200.28 55.15 200.49 55.22 ;
    RECT 200.28 55.51 200.49 55.58 ;
    RECT 199.82 54.79 200.03 54.86 ;
    RECT 199.82 55.15 200.03 55.22 ;
    RECT 199.82 55.51 200.03 55.58 ;
    RECT 196.96 54.79 197.17 54.86 ;
    RECT 196.96 55.15 197.17 55.22 ;
    RECT 196.96 55.51 197.17 55.58 ;
    RECT 196.5 54.79 196.71 54.86 ;
    RECT 196.5 55.15 196.71 55.22 ;
    RECT 196.5 55.51 196.71 55.58 ;
    RECT 193.64 54.79 193.85 54.86 ;
    RECT 193.64 55.15 193.85 55.22 ;
    RECT 193.64 55.51 193.85 55.58 ;
    RECT 193.18 54.79 193.39 54.86 ;
    RECT 193.18 55.15 193.39 55.22 ;
    RECT 193.18 55.51 193.39 55.58 ;
    RECT 190.32 54.79 190.53 54.86 ;
    RECT 190.32 55.15 190.53 55.22 ;
    RECT 190.32 55.51 190.53 55.58 ;
    RECT 189.86 54.79 190.07 54.86 ;
    RECT 189.86 55.15 190.07 55.22 ;
    RECT 189.86 55.51 190.07 55.58 ;
    RECT 187.0 54.79 187.21 54.86 ;
    RECT 187.0 55.15 187.21 55.22 ;
    RECT 187.0 55.51 187.21 55.58 ;
    RECT 186.54 54.79 186.75 54.86 ;
    RECT 186.54 55.15 186.75 55.22 ;
    RECT 186.54 55.51 186.75 55.58 ;
    RECT 147.485 55.15 147.555 55.22 ;
    RECT 183.68 54.79 183.89 54.86 ;
    RECT 183.68 55.15 183.89 55.22 ;
    RECT 183.68 55.51 183.89 55.58 ;
    RECT 183.22 54.79 183.43 54.86 ;
    RECT 183.22 55.15 183.43 55.22 ;
    RECT 183.22 55.51 183.43 55.58 ;
    RECT 266.68 54.79 266.89 54.86 ;
    RECT 266.68 55.15 266.89 55.22 ;
    RECT 266.68 55.51 266.89 55.58 ;
    RECT 266.22 54.79 266.43 54.86 ;
    RECT 266.22 55.15 266.43 55.22 ;
    RECT 266.22 55.51 266.43 55.58 ;
    RECT 263.36 54.79 263.57 54.86 ;
    RECT 263.36 55.15 263.57 55.22 ;
    RECT 263.36 55.51 263.57 55.58 ;
    RECT 262.9 54.79 263.11 54.86 ;
    RECT 262.9 55.15 263.11 55.22 ;
    RECT 262.9 55.51 263.11 55.58 ;
    RECT 260.04 54.79 260.25 54.86 ;
    RECT 260.04 55.15 260.25 55.22 ;
    RECT 260.04 55.51 260.25 55.58 ;
    RECT 259.58 54.79 259.79 54.86 ;
    RECT 259.58 55.15 259.79 55.22 ;
    RECT 259.58 55.51 259.79 55.58 ;
    RECT 256.72 54.79 256.93 54.86 ;
    RECT 256.72 55.15 256.93 55.22 ;
    RECT 256.72 55.51 256.93 55.58 ;
    RECT 256.26 54.79 256.47 54.86 ;
    RECT 256.26 55.15 256.47 55.22 ;
    RECT 256.26 55.51 256.47 55.58 ;
    RECT 253.4 54.79 253.61 54.86 ;
    RECT 253.4 55.15 253.61 55.22 ;
    RECT 253.4 55.51 253.61 55.58 ;
    RECT 252.94 54.79 253.15 54.86 ;
    RECT 252.94 55.15 253.15 55.22 ;
    RECT 252.94 55.51 253.15 55.58 ;
    RECT 250.08 22.39 250.29 22.46 ;
    RECT 250.08 22.75 250.29 22.82 ;
    RECT 250.08 23.11 250.29 23.18 ;
    RECT 249.62 22.39 249.83 22.46 ;
    RECT 249.62 22.75 249.83 22.82 ;
    RECT 249.62 23.11 249.83 23.18 ;
    RECT 246.76 22.39 246.97 22.46 ;
    RECT 246.76 22.75 246.97 22.82 ;
    RECT 246.76 23.11 246.97 23.18 ;
    RECT 246.3 22.39 246.51 22.46 ;
    RECT 246.3 22.75 246.51 22.82 ;
    RECT 246.3 23.11 246.51 23.18 ;
    RECT 243.44 22.39 243.65 22.46 ;
    RECT 243.44 22.75 243.65 22.82 ;
    RECT 243.44 23.11 243.65 23.18 ;
    RECT 242.98 22.39 243.19 22.46 ;
    RECT 242.98 22.75 243.19 22.82 ;
    RECT 242.98 23.11 243.19 23.18 ;
    RECT 240.12 22.39 240.33 22.46 ;
    RECT 240.12 22.75 240.33 22.82 ;
    RECT 240.12 23.11 240.33 23.18 ;
    RECT 239.66 22.39 239.87 22.46 ;
    RECT 239.66 22.75 239.87 22.82 ;
    RECT 239.66 23.11 239.87 23.18 ;
    RECT 236.8 22.39 237.01 22.46 ;
    RECT 236.8 22.75 237.01 22.82 ;
    RECT 236.8 23.11 237.01 23.18 ;
    RECT 236.34 22.39 236.55 22.46 ;
    RECT 236.34 22.75 236.55 22.82 ;
    RECT 236.34 23.11 236.55 23.18 ;
    RECT 233.48 22.39 233.69 22.46 ;
    RECT 233.48 22.75 233.69 22.82 ;
    RECT 233.48 23.11 233.69 23.18 ;
    RECT 233.02 22.39 233.23 22.46 ;
    RECT 233.02 22.75 233.23 22.82 ;
    RECT 233.02 23.11 233.23 23.18 ;
    RECT 230.16 22.39 230.37 22.46 ;
    RECT 230.16 22.75 230.37 22.82 ;
    RECT 230.16 23.11 230.37 23.18 ;
    RECT 229.7 22.39 229.91 22.46 ;
    RECT 229.7 22.75 229.91 22.82 ;
    RECT 229.7 23.11 229.91 23.18 ;
    RECT 226.84 22.39 227.05 22.46 ;
    RECT 226.84 22.75 227.05 22.82 ;
    RECT 226.84 23.11 227.05 23.18 ;
    RECT 226.38 22.39 226.59 22.46 ;
    RECT 226.38 22.75 226.59 22.82 ;
    RECT 226.38 23.11 226.59 23.18 ;
    RECT 223.52 22.39 223.73 22.46 ;
    RECT 223.52 22.75 223.73 22.82 ;
    RECT 223.52 23.11 223.73 23.18 ;
    RECT 223.06 22.39 223.27 22.46 ;
    RECT 223.06 22.75 223.27 22.82 ;
    RECT 223.06 23.11 223.27 23.18 ;
    RECT 220.2 22.39 220.41 22.46 ;
    RECT 220.2 22.75 220.41 22.82 ;
    RECT 220.2 23.11 220.41 23.18 ;
    RECT 219.74 22.39 219.95 22.46 ;
    RECT 219.74 22.75 219.95 22.82 ;
    RECT 219.74 23.11 219.95 23.18 ;
    RECT 216.88 22.39 217.09 22.46 ;
    RECT 216.88 22.75 217.09 22.82 ;
    RECT 216.88 23.11 217.09 23.18 ;
    RECT 216.42 22.39 216.63 22.46 ;
    RECT 216.42 22.75 216.63 22.82 ;
    RECT 216.42 23.11 216.63 23.18 ;
    RECT 267.91 22.75 267.98 22.82 ;
    RECT 180.36 22.39 180.57 22.46 ;
    RECT 180.36 22.75 180.57 22.82 ;
    RECT 180.36 23.11 180.57 23.18 ;
    RECT 179.9 22.39 180.11 22.46 ;
    RECT 179.9 22.75 180.11 22.82 ;
    RECT 179.9 23.11 180.11 23.18 ;
    RECT 177.04 22.39 177.25 22.46 ;
    RECT 177.04 22.75 177.25 22.82 ;
    RECT 177.04 23.11 177.25 23.18 ;
    RECT 176.58 22.39 176.79 22.46 ;
    RECT 176.58 22.75 176.79 22.82 ;
    RECT 176.58 23.11 176.79 23.18 ;
    RECT 173.72 22.39 173.93 22.46 ;
    RECT 173.72 22.75 173.93 22.82 ;
    RECT 173.72 23.11 173.93 23.18 ;
    RECT 173.26 22.39 173.47 22.46 ;
    RECT 173.26 22.75 173.47 22.82 ;
    RECT 173.26 23.11 173.47 23.18 ;
    RECT 170.4 22.39 170.61 22.46 ;
    RECT 170.4 22.75 170.61 22.82 ;
    RECT 170.4 23.11 170.61 23.18 ;
    RECT 169.94 22.39 170.15 22.46 ;
    RECT 169.94 22.75 170.15 22.82 ;
    RECT 169.94 23.11 170.15 23.18 ;
    RECT 167.08 22.39 167.29 22.46 ;
    RECT 167.08 22.75 167.29 22.82 ;
    RECT 167.08 23.11 167.29 23.18 ;
    RECT 166.62 22.39 166.83 22.46 ;
    RECT 166.62 22.75 166.83 22.82 ;
    RECT 166.62 23.11 166.83 23.18 ;
    RECT 163.76 22.39 163.97 22.46 ;
    RECT 163.76 22.75 163.97 22.82 ;
    RECT 163.76 23.11 163.97 23.18 ;
    RECT 163.3 22.39 163.51 22.46 ;
    RECT 163.3 22.75 163.51 22.82 ;
    RECT 163.3 23.11 163.51 23.18 ;
    RECT 160.44 22.39 160.65 22.46 ;
    RECT 160.44 22.75 160.65 22.82 ;
    RECT 160.44 23.11 160.65 23.18 ;
    RECT 159.98 22.39 160.19 22.46 ;
    RECT 159.98 22.75 160.19 22.82 ;
    RECT 159.98 23.11 160.19 23.18 ;
    RECT 157.12 22.39 157.33 22.46 ;
    RECT 157.12 22.75 157.33 22.82 ;
    RECT 157.12 23.11 157.33 23.18 ;
    RECT 156.66 22.39 156.87 22.46 ;
    RECT 156.66 22.75 156.87 22.82 ;
    RECT 156.66 23.11 156.87 23.18 ;
    RECT 153.8 22.39 154.01 22.46 ;
    RECT 153.8 22.75 154.01 22.82 ;
    RECT 153.8 23.11 154.01 23.18 ;
    RECT 153.34 22.39 153.55 22.46 ;
    RECT 153.34 22.75 153.55 22.82 ;
    RECT 153.34 23.11 153.55 23.18 ;
    RECT 150.48 22.39 150.69 22.46 ;
    RECT 150.48 22.75 150.69 22.82 ;
    RECT 150.48 23.11 150.69 23.18 ;
    RECT 150.02 22.39 150.23 22.46 ;
    RECT 150.02 22.75 150.23 22.82 ;
    RECT 150.02 23.11 150.23 23.18 ;
    RECT 213.56 22.39 213.77 22.46 ;
    RECT 213.56 22.75 213.77 22.82 ;
    RECT 213.56 23.11 213.77 23.18 ;
    RECT 213.1 22.39 213.31 22.46 ;
    RECT 213.1 22.75 213.31 22.82 ;
    RECT 213.1 23.11 213.31 23.18 ;
    RECT 210.24 22.39 210.45 22.46 ;
    RECT 210.24 22.75 210.45 22.82 ;
    RECT 210.24 23.11 210.45 23.18 ;
    RECT 209.78 22.39 209.99 22.46 ;
    RECT 209.78 22.75 209.99 22.82 ;
    RECT 209.78 23.11 209.99 23.18 ;
    RECT 206.92 22.39 207.13 22.46 ;
    RECT 206.92 22.75 207.13 22.82 ;
    RECT 206.92 23.11 207.13 23.18 ;
    RECT 206.46 22.39 206.67 22.46 ;
    RECT 206.46 22.75 206.67 22.82 ;
    RECT 206.46 23.11 206.67 23.18 ;
    RECT 203.6 22.39 203.81 22.46 ;
    RECT 203.6 22.75 203.81 22.82 ;
    RECT 203.6 23.11 203.81 23.18 ;
    RECT 203.14 22.39 203.35 22.46 ;
    RECT 203.14 22.75 203.35 22.82 ;
    RECT 203.14 23.11 203.35 23.18 ;
    RECT 200.28 22.39 200.49 22.46 ;
    RECT 200.28 22.75 200.49 22.82 ;
    RECT 200.28 23.11 200.49 23.18 ;
    RECT 199.82 22.39 200.03 22.46 ;
    RECT 199.82 22.75 200.03 22.82 ;
    RECT 199.82 23.11 200.03 23.18 ;
    RECT 196.96 22.39 197.17 22.46 ;
    RECT 196.96 22.75 197.17 22.82 ;
    RECT 196.96 23.11 197.17 23.18 ;
    RECT 196.5 22.39 196.71 22.46 ;
    RECT 196.5 22.75 196.71 22.82 ;
    RECT 196.5 23.11 196.71 23.18 ;
    RECT 193.64 22.39 193.85 22.46 ;
    RECT 193.64 22.75 193.85 22.82 ;
    RECT 193.64 23.11 193.85 23.18 ;
    RECT 193.18 22.39 193.39 22.46 ;
    RECT 193.18 22.75 193.39 22.82 ;
    RECT 193.18 23.11 193.39 23.18 ;
    RECT 190.32 22.39 190.53 22.46 ;
    RECT 190.32 22.75 190.53 22.82 ;
    RECT 190.32 23.11 190.53 23.18 ;
    RECT 189.86 22.39 190.07 22.46 ;
    RECT 189.86 22.75 190.07 22.82 ;
    RECT 189.86 23.11 190.07 23.18 ;
    RECT 187.0 22.39 187.21 22.46 ;
    RECT 187.0 22.75 187.21 22.82 ;
    RECT 187.0 23.11 187.21 23.18 ;
    RECT 186.54 22.39 186.75 22.46 ;
    RECT 186.54 22.75 186.75 22.82 ;
    RECT 186.54 23.11 186.75 23.18 ;
    RECT 183.68 22.39 183.89 22.46 ;
    RECT 183.68 22.75 183.89 22.82 ;
    RECT 183.68 23.11 183.89 23.18 ;
    RECT 183.22 22.39 183.43 22.46 ;
    RECT 183.22 22.75 183.43 22.82 ;
    RECT 183.22 23.11 183.43 23.18 ;
    RECT 147.485 22.75 147.555 22.82 ;
    RECT 266.68 22.39 266.89 22.46 ;
    RECT 266.68 22.75 266.89 22.82 ;
    RECT 266.68 23.11 266.89 23.18 ;
    RECT 266.22 22.39 266.43 22.46 ;
    RECT 266.22 22.75 266.43 22.82 ;
    RECT 266.22 23.11 266.43 23.18 ;
    RECT 263.36 22.39 263.57 22.46 ;
    RECT 263.36 22.75 263.57 22.82 ;
    RECT 263.36 23.11 263.57 23.18 ;
    RECT 262.9 22.39 263.11 22.46 ;
    RECT 262.9 22.75 263.11 22.82 ;
    RECT 262.9 23.11 263.11 23.18 ;
    RECT 260.04 22.39 260.25 22.46 ;
    RECT 260.04 22.75 260.25 22.82 ;
    RECT 260.04 23.11 260.25 23.18 ;
    RECT 259.58 22.39 259.79 22.46 ;
    RECT 259.58 22.75 259.79 22.82 ;
    RECT 259.58 23.11 259.79 23.18 ;
    RECT 256.72 22.39 256.93 22.46 ;
    RECT 256.72 22.75 256.93 22.82 ;
    RECT 256.72 23.11 256.93 23.18 ;
    RECT 256.26 22.39 256.47 22.46 ;
    RECT 256.26 22.75 256.47 22.82 ;
    RECT 256.26 23.11 256.47 23.18 ;
    RECT 253.4 22.39 253.61 22.46 ;
    RECT 253.4 22.75 253.61 22.82 ;
    RECT 253.4 23.11 253.61 23.18 ;
    RECT 252.94 22.39 253.15 22.46 ;
    RECT 252.94 22.75 253.15 22.82 ;
    RECT 252.94 23.11 253.15 23.18 ;
    RECT 250.08 62.01 250.29 62.08 ;
    RECT 250.08 62.37 250.29 62.44 ;
    RECT 250.08 62.73 250.29 62.8 ;
    RECT 249.62 62.01 249.83 62.08 ;
    RECT 249.62 62.37 249.83 62.44 ;
    RECT 249.62 62.73 249.83 62.8 ;
    RECT 246.76 62.01 246.97 62.08 ;
    RECT 246.76 62.37 246.97 62.44 ;
    RECT 246.76 62.73 246.97 62.8 ;
    RECT 246.3 62.01 246.51 62.08 ;
    RECT 246.3 62.37 246.51 62.44 ;
    RECT 246.3 62.73 246.51 62.8 ;
    RECT 243.44 62.01 243.65 62.08 ;
    RECT 243.44 62.37 243.65 62.44 ;
    RECT 243.44 62.73 243.65 62.8 ;
    RECT 242.98 62.01 243.19 62.08 ;
    RECT 242.98 62.37 243.19 62.44 ;
    RECT 242.98 62.73 243.19 62.8 ;
    RECT 240.12 62.01 240.33 62.08 ;
    RECT 240.12 62.37 240.33 62.44 ;
    RECT 240.12 62.73 240.33 62.8 ;
    RECT 239.66 62.01 239.87 62.08 ;
    RECT 239.66 62.37 239.87 62.44 ;
    RECT 239.66 62.73 239.87 62.8 ;
    RECT 236.8 62.01 237.01 62.08 ;
    RECT 236.8 62.37 237.01 62.44 ;
    RECT 236.8 62.73 237.01 62.8 ;
    RECT 236.34 62.01 236.55 62.08 ;
    RECT 236.34 62.37 236.55 62.44 ;
    RECT 236.34 62.73 236.55 62.8 ;
    RECT 233.48 62.01 233.69 62.08 ;
    RECT 233.48 62.37 233.69 62.44 ;
    RECT 233.48 62.73 233.69 62.8 ;
    RECT 233.02 62.01 233.23 62.08 ;
    RECT 233.02 62.37 233.23 62.44 ;
    RECT 233.02 62.73 233.23 62.8 ;
    RECT 230.16 62.01 230.37 62.08 ;
    RECT 230.16 62.37 230.37 62.44 ;
    RECT 230.16 62.73 230.37 62.8 ;
    RECT 229.7 62.01 229.91 62.08 ;
    RECT 229.7 62.37 229.91 62.44 ;
    RECT 229.7 62.73 229.91 62.8 ;
    RECT 226.84 62.01 227.05 62.08 ;
    RECT 226.84 62.37 227.05 62.44 ;
    RECT 226.84 62.73 227.05 62.8 ;
    RECT 226.38 62.01 226.59 62.08 ;
    RECT 226.38 62.37 226.59 62.44 ;
    RECT 226.38 62.73 226.59 62.8 ;
    RECT 223.52 62.01 223.73 62.08 ;
    RECT 223.52 62.37 223.73 62.44 ;
    RECT 223.52 62.73 223.73 62.8 ;
    RECT 223.06 62.01 223.27 62.08 ;
    RECT 223.06 62.37 223.27 62.44 ;
    RECT 223.06 62.73 223.27 62.8 ;
    RECT 220.2 62.01 220.41 62.08 ;
    RECT 220.2 62.37 220.41 62.44 ;
    RECT 220.2 62.73 220.41 62.8 ;
    RECT 219.74 62.01 219.95 62.08 ;
    RECT 219.74 62.37 219.95 62.44 ;
    RECT 219.74 62.73 219.95 62.8 ;
    RECT 216.88 62.01 217.09 62.08 ;
    RECT 216.88 62.37 217.09 62.44 ;
    RECT 216.88 62.73 217.09 62.8 ;
    RECT 216.42 62.01 216.63 62.08 ;
    RECT 216.42 62.37 216.63 62.44 ;
    RECT 216.42 62.73 216.63 62.8 ;
    RECT 267.91 62.37 267.98 62.44 ;
    RECT 180.36 62.01 180.57 62.08 ;
    RECT 180.36 62.37 180.57 62.44 ;
    RECT 180.36 62.73 180.57 62.8 ;
    RECT 179.9 62.01 180.11 62.08 ;
    RECT 179.9 62.37 180.11 62.44 ;
    RECT 179.9 62.73 180.11 62.8 ;
    RECT 177.04 62.01 177.25 62.08 ;
    RECT 177.04 62.37 177.25 62.44 ;
    RECT 177.04 62.73 177.25 62.8 ;
    RECT 176.58 62.01 176.79 62.08 ;
    RECT 176.58 62.37 176.79 62.44 ;
    RECT 176.58 62.73 176.79 62.8 ;
    RECT 173.72 62.01 173.93 62.08 ;
    RECT 173.72 62.37 173.93 62.44 ;
    RECT 173.72 62.73 173.93 62.8 ;
    RECT 173.26 62.01 173.47 62.08 ;
    RECT 173.26 62.37 173.47 62.44 ;
    RECT 173.26 62.73 173.47 62.8 ;
    RECT 170.4 62.01 170.61 62.08 ;
    RECT 170.4 62.37 170.61 62.44 ;
    RECT 170.4 62.73 170.61 62.8 ;
    RECT 169.94 62.01 170.15 62.08 ;
    RECT 169.94 62.37 170.15 62.44 ;
    RECT 169.94 62.73 170.15 62.8 ;
    RECT 167.08 62.01 167.29 62.08 ;
    RECT 167.08 62.37 167.29 62.44 ;
    RECT 167.08 62.73 167.29 62.8 ;
    RECT 166.62 62.01 166.83 62.08 ;
    RECT 166.62 62.37 166.83 62.44 ;
    RECT 166.62 62.73 166.83 62.8 ;
    RECT 163.76 62.01 163.97 62.08 ;
    RECT 163.76 62.37 163.97 62.44 ;
    RECT 163.76 62.73 163.97 62.8 ;
    RECT 163.3 62.01 163.51 62.08 ;
    RECT 163.3 62.37 163.51 62.44 ;
    RECT 163.3 62.73 163.51 62.8 ;
    RECT 160.44 62.01 160.65 62.08 ;
    RECT 160.44 62.37 160.65 62.44 ;
    RECT 160.44 62.73 160.65 62.8 ;
    RECT 159.98 62.01 160.19 62.08 ;
    RECT 159.98 62.37 160.19 62.44 ;
    RECT 159.98 62.73 160.19 62.8 ;
    RECT 157.12 62.01 157.33 62.08 ;
    RECT 157.12 62.37 157.33 62.44 ;
    RECT 157.12 62.73 157.33 62.8 ;
    RECT 156.66 62.01 156.87 62.08 ;
    RECT 156.66 62.37 156.87 62.44 ;
    RECT 156.66 62.73 156.87 62.8 ;
    RECT 153.8 62.01 154.01 62.08 ;
    RECT 153.8 62.37 154.01 62.44 ;
    RECT 153.8 62.73 154.01 62.8 ;
    RECT 153.34 62.01 153.55 62.08 ;
    RECT 153.34 62.37 153.55 62.44 ;
    RECT 153.34 62.73 153.55 62.8 ;
    RECT 150.48 62.01 150.69 62.08 ;
    RECT 150.48 62.37 150.69 62.44 ;
    RECT 150.48 62.73 150.69 62.8 ;
    RECT 150.02 62.01 150.23 62.08 ;
    RECT 150.02 62.37 150.23 62.44 ;
    RECT 150.02 62.73 150.23 62.8 ;
    RECT 213.56 62.01 213.77 62.08 ;
    RECT 213.56 62.37 213.77 62.44 ;
    RECT 213.56 62.73 213.77 62.8 ;
    RECT 213.1 62.01 213.31 62.08 ;
    RECT 213.1 62.37 213.31 62.44 ;
    RECT 213.1 62.73 213.31 62.8 ;
    RECT 210.24 62.01 210.45 62.08 ;
    RECT 210.24 62.37 210.45 62.44 ;
    RECT 210.24 62.73 210.45 62.8 ;
    RECT 209.78 62.01 209.99 62.08 ;
    RECT 209.78 62.37 209.99 62.44 ;
    RECT 209.78 62.73 209.99 62.8 ;
    RECT 206.92 62.01 207.13 62.08 ;
    RECT 206.92 62.37 207.13 62.44 ;
    RECT 206.92 62.73 207.13 62.8 ;
    RECT 206.46 62.01 206.67 62.08 ;
    RECT 206.46 62.37 206.67 62.44 ;
    RECT 206.46 62.73 206.67 62.8 ;
    RECT 203.6 62.01 203.81 62.08 ;
    RECT 203.6 62.37 203.81 62.44 ;
    RECT 203.6 62.73 203.81 62.8 ;
    RECT 203.14 62.01 203.35 62.08 ;
    RECT 203.14 62.37 203.35 62.44 ;
    RECT 203.14 62.73 203.35 62.8 ;
    RECT 200.28 62.01 200.49 62.08 ;
    RECT 200.28 62.37 200.49 62.44 ;
    RECT 200.28 62.73 200.49 62.8 ;
    RECT 199.82 62.01 200.03 62.08 ;
    RECT 199.82 62.37 200.03 62.44 ;
    RECT 199.82 62.73 200.03 62.8 ;
    RECT 196.96 62.01 197.17 62.08 ;
    RECT 196.96 62.37 197.17 62.44 ;
    RECT 196.96 62.73 197.17 62.8 ;
    RECT 196.5 62.01 196.71 62.08 ;
    RECT 196.5 62.37 196.71 62.44 ;
    RECT 196.5 62.73 196.71 62.8 ;
    RECT 193.64 62.01 193.85 62.08 ;
    RECT 193.64 62.37 193.85 62.44 ;
    RECT 193.64 62.73 193.85 62.8 ;
    RECT 193.18 62.01 193.39 62.08 ;
    RECT 193.18 62.37 193.39 62.44 ;
    RECT 193.18 62.73 193.39 62.8 ;
    RECT 190.32 62.01 190.53 62.08 ;
    RECT 190.32 62.37 190.53 62.44 ;
    RECT 190.32 62.73 190.53 62.8 ;
    RECT 189.86 62.01 190.07 62.08 ;
    RECT 189.86 62.37 190.07 62.44 ;
    RECT 189.86 62.73 190.07 62.8 ;
    RECT 187.0 62.01 187.21 62.08 ;
    RECT 187.0 62.37 187.21 62.44 ;
    RECT 187.0 62.73 187.21 62.8 ;
    RECT 186.54 62.01 186.75 62.08 ;
    RECT 186.54 62.37 186.75 62.44 ;
    RECT 186.54 62.73 186.75 62.8 ;
    RECT 183.68 62.01 183.89 62.08 ;
    RECT 183.68 62.37 183.89 62.44 ;
    RECT 183.68 62.73 183.89 62.8 ;
    RECT 183.22 62.01 183.43 62.08 ;
    RECT 183.22 62.37 183.43 62.44 ;
    RECT 183.22 62.73 183.43 62.8 ;
    RECT 147.485 62.37 147.555 62.44 ;
    RECT 266.68 62.01 266.89 62.08 ;
    RECT 266.68 62.37 266.89 62.44 ;
    RECT 266.68 62.73 266.89 62.8 ;
    RECT 266.22 62.01 266.43 62.08 ;
    RECT 266.22 62.37 266.43 62.44 ;
    RECT 266.22 62.73 266.43 62.8 ;
    RECT 263.36 62.01 263.57 62.08 ;
    RECT 263.36 62.37 263.57 62.44 ;
    RECT 263.36 62.73 263.57 62.8 ;
    RECT 262.9 62.01 263.11 62.08 ;
    RECT 262.9 62.37 263.11 62.44 ;
    RECT 262.9 62.73 263.11 62.8 ;
    RECT 260.04 62.01 260.25 62.08 ;
    RECT 260.04 62.37 260.25 62.44 ;
    RECT 260.04 62.73 260.25 62.8 ;
    RECT 259.58 62.01 259.79 62.08 ;
    RECT 259.58 62.37 259.79 62.44 ;
    RECT 259.58 62.73 259.79 62.8 ;
    RECT 256.72 62.01 256.93 62.08 ;
    RECT 256.72 62.37 256.93 62.44 ;
    RECT 256.72 62.73 256.93 62.8 ;
    RECT 256.26 62.01 256.47 62.08 ;
    RECT 256.26 62.37 256.47 62.44 ;
    RECT 256.26 62.73 256.47 62.8 ;
    RECT 253.4 62.01 253.61 62.08 ;
    RECT 253.4 62.37 253.61 62.44 ;
    RECT 253.4 62.73 253.61 62.8 ;
    RECT 252.94 62.01 253.15 62.08 ;
    RECT 252.94 62.37 253.15 62.44 ;
    RECT 252.94 62.73 253.15 62.8 ;
    RECT 250.08 97.29 250.29 97.36 ;
    RECT 250.08 97.65 250.29 97.72 ;
    RECT 250.08 98.01 250.29 98.08 ;
    RECT 249.62 97.29 249.83 97.36 ;
    RECT 249.62 97.65 249.83 97.72 ;
    RECT 249.62 98.01 249.83 98.08 ;
    RECT 246.76 97.29 246.97 97.36 ;
    RECT 246.76 97.65 246.97 97.72 ;
    RECT 246.76 98.01 246.97 98.08 ;
    RECT 246.3 97.29 246.51 97.36 ;
    RECT 246.3 97.65 246.51 97.72 ;
    RECT 246.3 98.01 246.51 98.08 ;
    RECT 243.44 97.29 243.65 97.36 ;
    RECT 243.44 97.65 243.65 97.72 ;
    RECT 243.44 98.01 243.65 98.08 ;
    RECT 242.98 97.29 243.19 97.36 ;
    RECT 242.98 97.65 243.19 97.72 ;
    RECT 242.98 98.01 243.19 98.08 ;
    RECT 240.12 97.29 240.33 97.36 ;
    RECT 240.12 97.65 240.33 97.72 ;
    RECT 240.12 98.01 240.33 98.08 ;
    RECT 239.66 97.29 239.87 97.36 ;
    RECT 239.66 97.65 239.87 97.72 ;
    RECT 239.66 98.01 239.87 98.08 ;
    RECT 236.8 97.29 237.01 97.36 ;
    RECT 236.8 97.65 237.01 97.72 ;
    RECT 236.8 98.01 237.01 98.08 ;
    RECT 236.34 97.29 236.55 97.36 ;
    RECT 236.34 97.65 236.55 97.72 ;
    RECT 236.34 98.01 236.55 98.08 ;
    RECT 233.48 97.29 233.69 97.36 ;
    RECT 233.48 97.65 233.69 97.72 ;
    RECT 233.48 98.01 233.69 98.08 ;
    RECT 233.02 97.29 233.23 97.36 ;
    RECT 233.02 97.65 233.23 97.72 ;
    RECT 233.02 98.01 233.23 98.08 ;
    RECT 230.16 97.29 230.37 97.36 ;
    RECT 230.16 97.65 230.37 97.72 ;
    RECT 230.16 98.01 230.37 98.08 ;
    RECT 229.7 97.29 229.91 97.36 ;
    RECT 229.7 97.65 229.91 97.72 ;
    RECT 229.7 98.01 229.91 98.08 ;
    RECT 226.84 97.29 227.05 97.36 ;
    RECT 226.84 97.65 227.05 97.72 ;
    RECT 226.84 98.01 227.05 98.08 ;
    RECT 226.38 97.29 226.59 97.36 ;
    RECT 226.38 97.65 226.59 97.72 ;
    RECT 226.38 98.01 226.59 98.08 ;
    RECT 223.52 97.29 223.73 97.36 ;
    RECT 223.52 97.65 223.73 97.72 ;
    RECT 223.52 98.01 223.73 98.08 ;
    RECT 223.06 97.29 223.27 97.36 ;
    RECT 223.06 97.65 223.27 97.72 ;
    RECT 223.06 98.01 223.27 98.08 ;
    RECT 220.2 97.29 220.41 97.36 ;
    RECT 220.2 97.65 220.41 97.72 ;
    RECT 220.2 98.01 220.41 98.08 ;
    RECT 219.74 97.29 219.95 97.36 ;
    RECT 219.74 97.65 219.95 97.72 ;
    RECT 219.74 98.01 219.95 98.08 ;
    RECT 216.88 97.29 217.09 97.36 ;
    RECT 216.88 97.65 217.09 97.72 ;
    RECT 216.88 98.01 217.09 98.08 ;
    RECT 216.42 97.29 216.63 97.36 ;
    RECT 216.42 97.65 216.63 97.72 ;
    RECT 216.42 98.01 216.63 98.08 ;
    RECT 267.91 97.65 267.98 97.72 ;
    RECT 180.36 97.29 180.57 97.36 ;
    RECT 180.36 97.65 180.57 97.72 ;
    RECT 180.36 98.01 180.57 98.08 ;
    RECT 179.9 97.29 180.11 97.36 ;
    RECT 179.9 97.65 180.11 97.72 ;
    RECT 179.9 98.01 180.11 98.08 ;
    RECT 177.04 97.29 177.25 97.36 ;
    RECT 177.04 97.65 177.25 97.72 ;
    RECT 177.04 98.01 177.25 98.08 ;
    RECT 176.58 97.29 176.79 97.36 ;
    RECT 176.58 97.65 176.79 97.72 ;
    RECT 176.58 98.01 176.79 98.08 ;
    RECT 173.72 97.29 173.93 97.36 ;
    RECT 173.72 97.65 173.93 97.72 ;
    RECT 173.72 98.01 173.93 98.08 ;
    RECT 173.26 97.29 173.47 97.36 ;
    RECT 173.26 97.65 173.47 97.72 ;
    RECT 173.26 98.01 173.47 98.08 ;
    RECT 170.4 97.29 170.61 97.36 ;
    RECT 170.4 97.65 170.61 97.72 ;
    RECT 170.4 98.01 170.61 98.08 ;
    RECT 169.94 97.29 170.15 97.36 ;
    RECT 169.94 97.65 170.15 97.72 ;
    RECT 169.94 98.01 170.15 98.08 ;
    RECT 167.08 97.29 167.29 97.36 ;
    RECT 167.08 97.65 167.29 97.72 ;
    RECT 167.08 98.01 167.29 98.08 ;
    RECT 166.62 97.29 166.83 97.36 ;
    RECT 166.62 97.65 166.83 97.72 ;
    RECT 166.62 98.01 166.83 98.08 ;
    RECT 163.76 97.29 163.97 97.36 ;
    RECT 163.76 97.65 163.97 97.72 ;
    RECT 163.76 98.01 163.97 98.08 ;
    RECT 163.3 97.29 163.51 97.36 ;
    RECT 163.3 97.65 163.51 97.72 ;
    RECT 163.3 98.01 163.51 98.08 ;
    RECT 160.44 97.29 160.65 97.36 ;
    RECT 160.44 97.65 160.65 97.72 ;
    RECT 160.44 98.01 160.65 98.08 ;
    RECT 159.98 97.29 160.19 97.36 ;
    RECT 159.98 97.65 160.19 97.72 ;
    RECT 159.98 98.01 160.19 98.08 ;
    RECT 157.12 97.29 157.33 97.36 ;
    RECT 157.12 97.65 157.33 97.72 ;
    RECT 157.12 98.01 157.33 98.08 ;
    RECT 156.66 97.29 156.87 97.36 ;
    RECT 156.66 97.65 156.87 97.72 ;
    RECT 156.66 98.01 156.87 98.08 ;
    RECT 153.8 97.29 154.01 97.36 ;
    RECT 153.8 97.65 154.01 97.72 ;
    RECT 153.8 98.01 154.01 98.08 ;
    RECT 153.34 97.29 153.55 97.36 ;
    RECT 153.34 97.65 153.55 97.72 ;
    RECT 153.34 98.01 153.55 98.08 ;
    RECT 150.48 97.29 150.69 97.36 ;
    RECT 150.48 97.65 150.69 97.72 ;
    RECT 150.48 98.01 150.69 98.08 ;
    RECT 150.02 97.29 150.23 97.36 ;
    RECT 150.02 97.65 150.23 97.72 ;
    RECT 150.02 98.01 150.23 98.08 ;
    RECT 213.56 97.29 213.77 97.36 ;
    RECT 213.56 97.65 213.77 97.72 ;
    RECT 213.56 98.01 213.77 98.08 ;
    RECT 213.1 97.29 213.31 97.36 ;
    RECT 213.1 97.65 213.31 97.72 ;
    RECT 213.1 98.01 213.31 98.08 ;
    RECT 210.24 97.29 210.45 97.36 ;
    RECT 210.24 97.65 210.45 97.72 ;
    RECT 210.24 98.01 210.45 98.08 ;
    RECT 209.78 97.29 209.99 97.36 ;
    RECT 209.78 97.65 209.99 97.72 ;
    RECT 209.78 98.01 209.99 98.08 ;
    RECT 206.92 97.29 207.13 97.36 ;
    RECT 206.92 97.65 207.13 97.72 ;
    RECT 206.92 98.01 207.13 98.08 ;
    RECT 206.46 97.29 206.67 97.36 ;
    RECT 206.46 97.65 206.67 97.72 ;
    RECT 206.46 98.01 206.67 98.08 ;
    RECT 203.6 97.29 203.81 97.36 ;
    RECT 203.6 97.65 203.81 97.72 ;
    RECT 203.6 98.01 203.81 98.08 ;
    RECT 203.14 97.29 203.35 97.36 ;
    RECT 203.14 97.65 203.35 97.72 ;
    RECT 203.14 98.01 203.35 98.08 ;
    RECT 200.28 97.29 200.49 97.36 ;
    RECT 200.28 97.65 200.49 97.72 ;
    RECT 200.28 98.01 200.49 98.08 ;
    RECT 199.82 97.29 200.03 97.36 ;
    RECT 199.82 97.65 200.03 97.72 ;
    RECT 199.82 98.01 200.03 98.08 ;
    RECT 196.96 97.29 197.17 97.36 ;
    RECT 196.96 97.65 197.17 97.72 ;
    RECT 196.96 98.01 197.17 98.08 ;
    RECT 196.5 97.29 196.71 97.36 ;
    RECT 196.5 97.65 196.71 97.72 ;
    RECT 196.5 98.01 196.71 98.08 ;
    RECT 193.64 97.29 193.85 97.36 ;
    RECT 193.64 97.65 193.85 97.72 ;
    RECT 193.64 98.01 193.85 98.08 ;
    RECT 193.18 97.29 193.39 97.36 ;
    RECT 193.18 97.65 193.39 97.72 ;
    RECT 193.18 98.01 193.39 98.08 ;
    RECT 190.32 97.29 190.53 97.36 ;
    RECT 190.32 97.65 190.53 97.72 ;
    RECT 190.32 98.01 190.53 98.08 ;
    RECT 189.86 97.29 190.07 97.36 ;
    RECT 189.86 97.65 190.07 97.72 ;
    RECT 189.86 98.01 190.07 98.08 ;
    RECT 187.0 97.29 187.21 97.36 ;
    RECT 187.0 97.65 187.21 97.72 ;
    RECT 187.0 98.01 187.21 98.08 ;
    RECT 186.54 97.29 186.75 97.36 ;
    RECT 186.54 97.65 186.75 97.72 ;
    RECT 186.54 98.01 186.75 98.08 ;
    RECT 183.68 97.29 183.89 97.36 ;
    RECT 183.68 97.65 183.89 97.72 ;
    RECT 183.68 98.01 183.89 98.08 ;
    RECT 183.22 97.29 183.43 97.36 ;
    RECT 183.22 97.65 183.43 97.72 ;
    RECT 183.22 98.01 183.43 98.08 ;
    RECT 147.485 97.65 147.555 97.72 ;
    RECT 266.68 97.29 266.89 97.36 ;
    RECT 266.68 97.65 266.89 97.72 ;
    RECT 266.68 98.01 266.89 98.08 ;
    RECT 266.22 97.29 266.43 97.36 ;
    RECT 266.22 97.65 266.43 97.72 ;
    RECT 266.22 98.01 266.43 98.08 ;
    RECT 263.36 97.29 263.57 97.36 ;
    RECT 263.36 97.65 263.57 97.72 ;
    RECT 263.36 98.01 263.57 98.08 ;
    RECT 262.9 97.29 263.11 97.36 ;
    RECT 262.9 97.65 263.11 97.72 ;
    RECT 262.9 98.01 263.11 98.08 ;
    RECT 260.04 97.29 260.25 97.36 ;
    RECT 260.04 97.65 260.25 97.72 ;
    RECT 260.04 98.01 260.25 98.08 ;
    RECT 259.58 97.29 259.79 97.36 ;
    RECT 259.58 97.65 259.79 97.72 ;
    RECT 259.58 98.01 259.79 98.08 ;
    RECT 256.72 97.29 256.93 97.36 ;
    RECT 256.72 97.65 256.93 97.72 ;
    RECT 256.72 98.01 256.93 98.08 ;
    RECT 256.26 97.29 256.47 97.36 ;
    RECT 256.26 97.65 256.47 97.72 ;
    RECT 256.26 98.01 256.47 98.08 ;
    RECT 253.4 97.29 253.61 97.36 ;
    RECT 253.4 97.65 253.61 97.72 ;
    RECT 253.4 98.01 253.61 98.08 ;
    RECT 252.94 97.29 253.15 97.36 ;
    RECT 252.94 97.65 253.15 97.72 ;
    RECT 252.94 98.01 253.15 98.08 ;
    RECT 250.08 21.67 250.29 21.74 ;
    RECT 250.08 22.03 250.29 22.1 ;
    RECT 250.08 22.39 250.29 22.46 ;
    RECT 249.62 21.67 249.83 21.74 ;
    RECT 249.62 22.03 249.83 22.1 ;
    RECT 249.62 22.39 249.83 22.46 ;
    RECT 246.76 21.67 246.97 21.74 ;
    RECT 246.76 22.03 246.97 22.1 ;
    RECT 246.76 22.39 246.97 22.46 ;
    RECT 246.3 21.67 246.51 21.74 ;
    RECT 246.3 22.03 246.51 22.1 ;
    RECT 246.3 22.39 246.51 22.46 ;
    RECT 243.44 21.67 243.65 21.74 ;
    RECT 243.44 22.03 243.65 22.1 ;
    RECT 243.44 22.39 243.65 22.46 ;
    RECT 242.98 21.67 243.19 21.74 ;
    RECT 242.98 22.03 243.19 22.1 ;
    RECT 242.98 22.39 243.19 22.46 ;
    RECT 240.12 21.67 240.33 21.74 ;
    RECT 240.12 22.03 240.33 22.1 ;
    RECT 240.12 22.39 240.33 22.46 ;
    RECT 239.66 21.67 239.87 21.74 ;
    RECT 239.66 22.03 239.87 22.1 ;
    RECT 239.66 22.39 239.87 22.46 ;
    RECT 236.8 21.67 237.01 21.74 ;
    RECT 236.8 22.03 237.01 22.1 ;
    RECT 236.8 22.39 237.01 22.46 ;
    RECT 236.34 21.67 236.55 21.74 ;
    RECT 236.34 22.03 236.55 22.1 ;
    RECT 236.34 22.39 236.55 22.46 ;
    RECT 233.48 21.67 233.69 21.74 ;
    RECT 233.48 22.03 233.69 22.1 ;
    RECT 233.48 22.39 233.69 22.46 ;
    RECT 233.02 21.67 233.23 21.74 ;
    RECT 233.02 22.03 233.23 22.1 ;
    RECT 233.02 22.39 233.23 22.46 ;
    RECT 230.16 21.67 230.37 21.74 ;
    RECT 230.16 22.03 230.37 22.1 ;
    RECT 230.16 22.39 230.37 22.46 ;
    RECT 229.7 21.67 229.91 21.74 ;
    RECT 229.7 22.03 229.91 22.1 ;
    RECT 229.7 22.39 229.91 22.46 ;
    RECT 226.84 21.67 227.05 21.74 ;
    RECT 226.84 22.03 227.05 22.1 ;
    RECT 226.84 22.39 227.05 22.46 ;
    RECT 226.38 21.67 226.59 21.74 ;
    RECT 226.38 22.03 226.59 22.1 ;
    RECT 226.38 22.39 226.59 22.46 ;
    RECT 223.52 21.67 223.73 21.74 ;
    RECT 223.52 22.03 223.73 22.1 ;
    RECT 223.52 22.39 223.73 22.46 ;
    RECT 223.06 21.67 223.27 21.74 ;
    RECT 223.06 22.03 223.27 22.1 ;
    RECT 223.06 22.39 223.27 22.46 ;
    RECT 220.2 21.67 220.41 21.74 ;
    RECT 220.2 22.03 220.41 22.1 ;
    RECT 220.2 22.39 220.41 22.46 ;
    RECT 219.74 21.67 219.95 21.74 ;
    RECT 219.74 22.03 219.95 22.1 ;
    RECT 219.74 22.39 219.95 22.46 ;
    RECT 216.88 21.67 217.09 21.74 ;
    RECT 216.88 22.03 217.09 22.1 ;
    RECT 216.88 22.39 217.09 22.46 ;
    RECT 216.42 21.67 216.63 21.74 ;
    RECT 216.42 22.03 216.63 22.1 ;
    RECT 216.42 22.39 216.63 22.46 ;
    RECT 267.91 22.03 267.98 22.1 ;
    RECT 180.36 21.67 180.57 21.74 ;
    RECT 180.36 22.03 180.57 22.1 ;
    RECT 180.36 22.39 180.57 22.46 ;
    RECT 179.9 21.67 180.11 21.74 ;
    RECT 179.9 22.03 180.11 22.1 ;
    RECT 179.9 22.39 180.11 22.46 ;
    RECT 177.04 21.67 177.25 21.74 ;
    RECT 177.04 22.03 177.25 22.1 ;
    RECT 177.04 22.39 177.25 22.46 ;
    RECT 176.58 21.67 176.79 21.74 ;
    RECT 176.58 22.03 176.79 22.1 ;
    RECT 176.58 22.39 176.79 22.46 ;
    RECT 173.72 21.67 173.93 21.74 ;
    RECT 173.72 22.03 173.93 22.1 ;
    RECT 173.72 22.39 173.93 22.46 ;
    RECT 173.26 21.67 173.47 21.74 ;
    RECT 173.26 22.03 173.47 22.1 ;
    RECT 173.26 22.39 173.47 22.46 ;
    RECT 170.4 21.67 170.61 21.74 ;
    RECT 170.4 22.03 170.61 22.1 ;
    RECT 170.4 22.39 170.61 22.46 ;
    RECT 169.94 21.67 170.15 21.74 ;
    RECT 169.94 22.03 170.15 22.1 ;
    RECT 169.94 22.39 170.15 22.46 ;
    RECT 167.08 21.67 167.29 21.74 ;
    RECT 167.08 22.03 167.29 22.1 ;
    RECT 167.08 22.39 167.29 22.46 ;
    RECT 166.62 21.67 166.83 21.74 ;
    RECT 166.62 22.03 166.83 22.1 ;
    RECT 166.62 22.39 166.83 22.46 ;
    RECT 163.76 21.67 163.97 21.74 ;
    RECT 163.76 22.03 163.97 22.1 ;
    RECT 163.76 22.39 163.97 22.46 ;
    RECT 163.3 21.67 163.51 21.74 ;
    RECT 163.3 22.03 163.51 22.1 ;
    RECT 163.3 22.39 163.51 22.46 ;
    RECT 160.44 21.67 160.65 21.74 ;
    RECT 160.44 22.03 160.65 22.1 ;
    RECT 160.44 22.39 160.65 22.46 ;
    RECT 159.98 21.67 160.19 21.74 ;
    RECT 159.98 22.03 160.19 22.1 ;
    RECT 159.98 22.39 160.19 22.46 ;
    RECT 157.12 21.67 157.33 21.74 ;
    RECT 157.12 22.03 157.33 22.1 ;
    RECT 157.12 22.39 157.33 22.46 ;
    RECT 156.66 21.67 156.87 21.74 ;
    RECT 156.66 22.03 156.87 22.1 ;
    RECT 156.66 22.39 156.87 22.46 ;
    RECT 153.8 21.67 154.01 21.74 ;
    RECT 153.8 22.03 154.01 22.1 ;
    RECT 153.8 22.39 154.01 22.46 ;
    RECT 153.34 21.67 153.55 21.74 ;
    RECT 153.34 22.03 153.55 22.1 ;
    RECT 153.34 22.39 153.55 22.46 ;
    RECT 150.48 21.67 150.69 21.74 ;
    RECT 150.48 22.03 150.69 22.1 ;
    RECT 150.48 22.39 150.69 22.46 ;
    RECT 150.02 21.67 150.23 21.74 ;
    RECT 150.02 22.03 150.23 22.1 ;
    RECT 150.02 22.39 150.23 22.46 ;
    RECT 213.56 21.67 213.77 21.74 ;
    RECT 213.56 22.03 213.77 22.1 ;
    RECT 213.56 22.39 213.77 22.46 ;
    RECT 213.1 21.67 213.31 21.74 ;
    RECT 213.1 22.03 213.31 22.1 ;
    RECT 213.1 22.39 213.31 22.46 ;
    RECT 210.24 21.67 210.45 21.74 ;
    RECT 210.24 22.03 210.45 22.1 ;
    RECT 210.24 22.39 210.45 22.46 ;
    RECT 209.78 21.67 209.99 21.74 ;
    RECT 209.78 22.03 209.99 22.1 ;
    RECT 209.78 22.39 209.99 22.46 ;
    RECT 206.92 21.67 207.13 21.74 ;
    RECT 206.92 22.03 207.13 22.1 ;
    RECT 206.92 22.39 207.13 22.46 ;
    RECT 206.46 21.67 206.67 21.74 ;
    RECT 206.46 22.03 206.67 22.1 ;
    RECT 206.46 22.39 206.67 22.46 ;
    RECT 203.6 21.67 203.81 21.74 ;
    RECT 203.6 22.03 203.81 22.1 ;
    RECT 203.6 22.39 203.81 22.46 ;
    RECT 203.14 21.67 203.35 21.74 ;
    RECT 203.14 22.03 203.35 22.1 ;
    RECT 203.14 22.39 203.35 22.46 ;
    RECT 200.28 21.67 200.49 21.74 ;
    RECT 200.28 22.03 200.49 22.1 ;
    RECT 200.28 22.39 200.49 22.46 ;
    RECT 199.82 21.67 200.03 21.74 ;
    RECT 199.82 22.03 200.03 22.1 ;
    RECT 199.82 22.39 200.03 22.46 ;
    RECT 196.96 21.67 197.17 21.74 ;
    RECT 196.96 22.03 197.17 22.1 ;
    RECT 196.96 22.39 197.17 22.46 ;
    RECT 196.5 21.67 196.71 21.74 ;
    RECT 196.5 22.03 196.71 22.1 ;
    RECT 196.5 22.39 196.71 22.46 ;
    RECT 193.64 21.67 193.85 21.74 ;
    RECT 193.64 22.03 193.85 22.1 ;
    RECT 193.64 22.39 193.85 22.46 ;
    RECT 193.18 21.67 193.39 21.74 ;
    RECT 193.18 22.03 193.39 22.1 ;
    RECT 193.18 22.39 193.39 22.46 ;
    RECT 190.32 21.67 190.53 21.74 ;
    RECT 190.32 22.03 190.53 22.1 ;
    RECT 190.32 22.39 190.53 22.46 ;
    RECT 189.86 21.67 190.07 21.74 ;
    RECT 189.86 22.03 190.07 22.1 ;
    RECT 189.86 22.39 190.07 22.46 ;
    RECT 187.0 21.67 187.21 21.74 ;
    RECT 187.0 22.03 187.21 22.1 ;
    RECT 187.0 22.39 187.21 22.46 ;
    RECT 186.54 21.67 186.75 21.74 ;
    RECT 186.54 22.03 186.75 22.1 ;
    RECT 186.54 22.39 186.75 22.46 ;
    RECT 183.68 21.67 183.89 21.74 ;
    RECT 183.68 22.03 183.89 22.1 ;
    RECT 183.68 22.39 183.89 22.46 ;
    RECT 183.22 21.67 183.43 21.74 ;
    RECT 183.22 22.03 183.43 22.1 ;
    RECT 183.22 22.39 183.43 22.46 ;
    RECT 147.485 22.03 147.555 22.1 ;
    RECT 266.68 21.67 266.89 21.74 ;
    RECT 266.68 22.03 266.89 22.1 ;
    RECT 266.68 22.39 266.89 22.46 ;
    RECT 266.22 21.67 266.43 21.74 ;
    RECT 266.22 22.03 266.43 22.1 ;
    RECT 266.22 22.39 266.43 22.46 ;
    RECT 263.36 21.67 263.57 21.74 ;
    RECT 263.36 22.03 263.57 22.1 ;
    RECT 263.36 22.39 263.57 22.46 ;
    RECT 262.9 21.67 263.11 21.74 ;
    RECT 262.9 22.03 263.11 22.1 ;
    RECT 262.9 22.39 263.11 22.46 ;
    RECT 260.04 21.67 260.25 21.74 ;
    RECT 260.04 22.03 260.25 22.1 ;
    RECT 260.04 22.39 260.25 22.46 ;
    RECT 259.58 21.67 259.79 21.74 ;
    RECT 259.58 22.03 259.79 22.1 ;
    RECT 259.58 22.39 259.79 22.46 ;
    RECT 256.72 21.67 256.93 21.74 ;
    RECT 256.72 22.03 256.93 22.1 ;
    RECT 256.72 22.39 256.93 22.46 ;
    RECT 256.26 21.67 256.47 21.74 ;
    RECT 256.26 22.03 256.47 22.1 ;
    RECT 256.26 22.39 256.47 22.46 ;
    RECT 253.4 21.67 253.61 21.74 ;
    RECT 253.4 22.03 253.61 22.1 ;
    RECT 253.4 22.39 253.61 22.46 ;
    RECT 252.94 21.67 253.15 21.74 ;
    RECT 252.94 22.03 253.15 22.1 ;
    RECT 252.94 22.39 253.15 22.46 ;
    RECT 250.08 61.29 250.29 61.36 ;
    RECT 250.08 61.65 250.29 61.72 ;
    RECT 250.08 62.01 250.29 62.08 ;
    RECT 249.62 61.29 249.83 61.36 ;
    RECT 249.62 61.65 249.83 61.72 ;
    RECT 249.62 62.01 249.83 62.08 ;
    RECT 246.76 61.29 246.97 61.36 ;
    RECT 246.76 61.65 246.97 61.72 ;
    RECT 246.76 62.01 246.97 62.08 ;
    RECT 246.3 61.29 246.51 61.36 ;
    RECT 246.3 61.65 246.51 61.72 ;
    RECT 246.3 62.01 246.51 62.08 ;
    RECT 243.44 61.29 243.65 61.36 ;
    RECT 243.44 61.65 243.65 61.72 ;
    RECT 243.44 62.01 243.65 62.08 ;
    RECT 242.98 61.29 243.19 61.36 ;
    RECT 242.98 61.65 243.19 61.72 ;
    RECT 242.98 62.01 243.19 62.08 ;
    RECT 240.12 61.29 240.33 61.36 ;
    RECT 240.12 61.65 240.33 61.72 ;
    RECT 240.12 62.01 240.33 62.08 ;
    RECT 239.66 61.29 239.87 61.36 ;
    RECT 239.66 61.65 239.87 61.72 ;
    RECT 239.66 62.01 239.87 62.08 ;
    RECT 236.8 61.29 237.01 61.36 ;
    RECT 236.8 61.65 237.01 61.72 ;
    RECT 236.8 62.01 237.01 62.08 ;
    RECT 236.34 61.29 236.55 61.36 ;
    RECT 236.34 61.65 236.55 61.72 ;
    RECT 236.34 62.01 236.55 62.08 ;
    RECT 233.48 61.29 233.69 61.36 ;
    RECT 233.48 61.65 233.69 61.72 ;
    RECT 233.48 62.01 233.69 62.08 ;
    RECT 233.02 61.29 233.23 61.36 ;
    RECT 233.02 61.65 233.23 61.72 ;
    RECT 233.02 62.01 233.23 62.08 ;
    RECT 230.16 61.29 230.37 61.36 ;
    RECT 230.16 61.65 230.37 61.72 ;
    RECT 230.16 62.01 230.37 62.08 ;
    RECT 229.7 61.29 229.91 61.36 ;
    RECT 229.7 61.65 229.91 61.72 ;
    RECT 229.7 62.01 229.91 62.08 ;
    RECT 226.84 61.29 227.05 61.36 ;
    RECT 226.84 61.65 227.05 61.72 ;
    RECT 226.84 62.01 227.05 62.08 ;
    RECT 226.38 61.29 226.59 61.36 ;
    RECT 226.38 61.65 226.59 61.72 ;
    RECT 226.38 62.01 226.59 62.08 ;
    RECT 223.52 61.29 223.73 61.36 ;
    RECT 223.52 61.65 223.73 61.72 ;
    RECT 223.52 62.01 223.73 62.08 ;
    RECT 223.06 61.29 223.27 61.36 ;
    RECT 223.06 61.65 223.27 61.72 ;
    RECT 223.06 62.01 223.27 62.08 ;
    RECT 220.2 61.29 220.41 61.36 ;
    RECT 220.2 61.65 220.41 61.72 ;
    RECT 220.2 62.01 220.41 62.08 ;
    RECT 219.74 61.29 219.95 61.36 ;
    RECT 219.74 61.65 219.95 61.72 ;
    RECT 219.74 62.01 219.95 62.08 ;
    RECT 216.88 61.29 217.09 61.36 ;
    RECT 216.88 61.65 217.09 61.72 ;
    RECT 216.88 62.01 217.09 62.08 ;
    RECT 216.42 61.29 216.63 61.36 ;
    RECT 216.42 61.65 216.63 61.72 ;
    RECT 216.42 62.01 216.63 62.08 ;
    RECT 267.91 61.65 267.98 61.72 ;
    RECT 180.36 61.29 180.57 61.36 ;
    RECT 180.36 61.65 180.57 61.72 ;
    RECT 180.36 62.01 180.57 62.08 ;
    RECT 179.9 61.29 180.11 61.36 ;
    RECT 179.9 61.65 180.11 61.72 ;
    RECT 179.9 62.01 180.11 62.08 ;
    RECT 177.04 61.29 177.25 61.36 ;
    RECT 177.04 61.65 177.25 61.72 ;
    RECT 177.04 62.01 177.25 62.08 ;
    RECT 176.58 61.29 176.79 61.36 ;
    RECT 176.58 61.65 176.79 61.72 ;
    RECT 176.58 62.01 176.79 62.08 ;
    RECT 173.72 61.29 173.93 61.36 ;
    RECT 173.72 61.65 173.93 61.72 ;
    RECT 173.72 62.01 173.93 62.08 ;
    RECT 173.26 61.29 173.47 61.36 ;
    RECT 173.26 61.65 173.47 61.72 ;
    RECT 173.26 62.01 173.47 62.08 ;
    RECT 170.4 61.29 170.61 61.36 ;
    RECT 170.4 61.65 170.61 61.72 ;
    RECT 170.4 62.01 170.61 62.08 ;
    RECT 169.94 61.29 170.15 61.36 ;
    RECT 169.94 61.65 170.15 61.72 ;
    RECT 169.94 62.01 170.15 62.08 ;
    RECT 167.08 61.29 167.29 61.36 ;
    RECT 167.08 61.65 167.29 61.72 ;
    RECT 167.08 62.01 167.29 62.08 ;
    RECT 166.62 61.29 166.83 61.36 ;
    RECT 166.62 61.65 166.83 61.72 ;
    RECT 166.62 62.01 166.83 62.08 ;
    RECT 163.76 61.29 163.97 61.36 ;
    RECT 163.76 61.65 163.97 61.72 ;
    RECT 163.76 62.01 163.97 62.08 ;
    RECT 163.3 61.29 163.51 61.36 ;
    RECT 163.3 61.65 163.51 61.72 ;
    RECT 163.3 62.01 163.51 62.08 ;
    RECT 160.44 61.29 160.65 61.36 ;
    RECT 160.44 61.65 160.65 61.72 ;
    RECT 160.44 62.01 160.65 62.08 ;
    RECT 159.98 61.29 160.19 61.36 ;
    RECT 159.98 61.65 160.19 61.72 ;
    RECT 159.98 62.01 160.19 62.08 ;
    RECT 157.12 61.29 157.33 61.36 ;
    RECT 157.12 61.65 157.33 61.72 ;
    RECT 157.12 62.01 157.33 62.08 ;
    RECT 156.66 61.29 156.87 61.36 ;
    RECT 156.66 61.65 156.87 61.72 ;
    RECT 156.66 62.01 156.87 62.08 ;
    RECT 153.8 61.29 154.01 61.36 ;
    RECT 153.8 61.65 154.01 61.72 ;
    RECT 153.8 62.01 154.01 62.08 ;
    RECT 153.34 61.29 153.55 61.36 ;
    RECT 153.34 61.65 153.55 61.72 ;
    RECT 153.34 62.01 153.55 62.08 ;
    RECT 150.48 61.29 150.69 61.36 ;
    RECT 150.48 61.65 150.69 61.72 ;
    RECT 150.48 62.01 150.69 62.08 ;
    RECT 150.02 61.29 150.23 61.36 ;
    RECT 150.02 61.65 150.23 61.72 ;
    RECT 150.02 62.01 150.23 62.08 ;
    RECT 213.56 61.29 213.77 61.36 ;
    RECT 213.56 61.65 213.77 61.72 ;
    RECT 213.56 62.01 213.77 62.08 ;
    RECT 213.1 61.29 213.31 61.36 ;
    RECT 213.1 61.65 213.31 61.72 ;
    RECT 213.1 62.01 213.31 62.08 ;
    RECT 210.24 61.29 210.45 61.36 ;
    RECT 210.24 61.65 210.45 61.72 ;
    RECT 210.24 62.01 210.45 62.08 ;
    RECT 209.78 61.29 209.99 61.36 ;
    RECT 209.78 61.65 209.99 61.72 ;
    RECT 209.78 62.01 209.99 62.08 ;
    RECT 206.92 61.29 207.13 61.36 ;
    RECT 206.92 61.65 207.13 61.72 ;
    RECT 206.92 62.01 207.13 62.08 ;
    RECT 206.46 61.29 206.67 61.36 ;
    RECT 206.46 61.65 206.67 61.72 ;
    RECT 206.46 62.01 206.67 62.08 ;
    RECT 203.6 61.29 203.81 61.36 ;
    RECT 203.6 61.65 203.81 61.72 ;
    RECT 203.6 62.01 203.81 62.08 ;
    RECT 203.14 61.29 203.35 61.36 ;
    RECT 203.14 61.65 203.35 61.72 ;
    RECT 203.14 62.01 203.35 62.08 ;
    RECT 200.28 61.29 200.49 61.36 ;
    RECT 200.28 61.65 200.49 61.72 ;
    RECT 200.28 62.01 200.49 62.08 ;
    RECT 199.82 61.29 200.03 61.36 ;
    RECT 199.82 61.65 200.03 61.72 ;
    RECT 199.82 62.01 200.03 62.08 ;
    RECT 196.96 61.29 197.17 61.36 ;
    RECT 196.96 61.65 197.17 61.72 ;
    RECT 196.96 62.01 197.17 62.08 ;
    RECT 196.5 61.29 196.71 61.36 ;
    RECT 196.5 61.65 196.71 61.72 ;
    RECT 196.5 62.01 196.71 62.08 ;
    RECT 193.64 61.29 193.85 61.36 ;
    RECT 193.64 61.65 193.85 61.72 ;
    RECT 193.64 62.01 193.85 62.08 ;
    RECT 193.18 61.29 193.39 61.36 ;
    RECT 193.18 61.65 193.39 61.72 ;
    RECT 193.18 62.01 193.39 62.08 ;
    RECT 190.32 61.29 190.53 61.36 ;
    RECT 190.32 61.65 190.53 61.72 ;
    RECT 190.32 62.01 190.53 62.08 ;
    RECT 189.86 61.29 190.07 61.36 ;
    RECT 189.86 61.65 190.07 61.72 ;
    RECT 189.86 62.01 190.07 62.08 ;
    RECT 187.0 61.29 187.21 61.36 ;
    RECT 187.0 61.65 187.21 61.72 ;
    RECT 187.0 62.01 187.21 62.08 ;
    RECT 186.54 61.29 186.75 61.36 ;
    RECT 186.54 61.65 186.75 61.72 ;
    RECT 186.54 62.01 186.75 62.08 ;
    RECT 183.68 61.29 183.89 61.36 ;
    RECT 183.68 61.65 183.89 61.72 ;
    RECT 183.68 62.01 183.89 62.08 ;
    RECT 183.22 61.29 183.43 61.36 ;
    RECT 183.22 61.65 183.43 61.72 ;
    RECT 183.22 62.01 183.43 62.08 ;
    RECT 147.485 61.65 147.555 61.72 ;
    RECT 266.68 61.29 266.89 61.36 ;
    RECT 266.68 61.65 266.89 61.72 ;
    RECT 266.68 62.01 266.89 62.08 ;
    RECT 266.22 61.29 266.43 61.36 ;
    RECT 266.22 61.65 266.43 61.72 ;
    RECT 266.22 62.01 266.43 62.08 ;
    RECT 263.36 61.29 263.57 61.36 ;
    RECT 263.36 61.65 263.57 61.72 ;
    RECT 263.36 62.01 263.57 62.08 ;
    RECT 262.9 61.29 263.11 61.36 ;
    RECT 262.9 61.65 263.11 61.72 ;
    RECT 262.9 62.01 263.11 62.08 ;
    RECT 260.04 61.29 260.25 61.36 ;
    RECT 260.04 61.65 260.25 61.72 ;
    RECT 260.04 62.01 260.25 62.08 ;
    RECT 259.58 61.29 259.79 61.36 ;
    RECT 259.58 61.65 259.79 61.72 ;
    RECT 259.58 62.01 259.79 62.08 ;
    RECT 256.72 61.29 256.93 61.36 ;
    RECT 256.72 61.65 256.93 61.72 ;
    RECT 256.72 62.01 256.93 62.08 ;
    RECT 256.26 61.29 256.47 61.36 ;
    RECT 256.26 61.65 256.47 61.72 ;
    RECT 256.26 62.01 256.47 62.08 ;
    RECT 253.4 61.29 253.61 61.36 ;
    RECT 253.4 61.65 253.61 61.72 ;
    RECT 253.4 62.01 253.61 62.08 ;
    RECT 252.94 61.29 253.15 61.36 ;
    RECT 252.94 61.65 253.15 61.72 ;
    RECT 252.94 62.01 253.15 62.08 ;
    RECT 212.61 60.79 212.82 60.86 ;
    RECT 179.9 61.05 180.11 61.12 ;
    RECT 180.36 61.05 180.57 61.12 ;
    RECT 159.49 60.79 159.7 60.86 ;
    RECT 235.85 60.79 236.06 60.86 ;
    RECT 255.77 60.79 255.98 60.86 ;
    RECT 216.42 61.05 216.63 61.12 ;
    RECT 216.88 61.05 217.09 61.12 ;
    RECT 239.66 61.05 239.87 61.12 ;
    RECT 240.12 61.05 240.33 61.12 ;
    RECT 156.66 61.05 156.87 61.12 ;
    RECT 157.12 61.05 157.33 61.12 ;
    RECT 182.73 60.79 182.94 60.86 ;
    RECT 252.94 61.05 253.15 61.12 ;
    RECT 253.4 61.05 253.61 61.12 ;
    RECT 193.18 61.05 193.39 61.12 ;
    RECT 193.64 61.05 193.85 61.12 ;
    RECT 205.97 60.79 206.18 60.86 ;
    RECT 176.09 60.79 176.3 60.86 ;
    RECT 152.85 60.79 153.06 60.86 ;
    RECT 229.21 60.79 229.42 60.86 ;
    RECT 249.13 60.79 249.34 60.86 ;
    RECT 233.02 61.05 233.23 61.12 ;
    RECT 233.48 61.05 233.69 61.12 ;
    RECT 150.02 61.05 150.23 61.12 ;
    RECT 150.48 61.05 150.69 61.12 ;
    RECT 173.26 61.05 173.47 61.12 ;
    RECT 173.72 61.05 173.93 61.12 ;
    RECT 186.54 61.05 186.75 61.12 ;
    RECT 187.0 61.05 187.21 61.12 ;
    RECT 209.78 61.05 209.99 61.12 ;
    RECT 210.24 61.05 210.45 61.12 ;
    RECT 199.33 60.79 199.54 60.86 ;
    RECT 219.25 60.79 219.46 60.86 ;
    RECT 169.45 60.79 169.66 60.86 ;
    RECT 268.12 60.79 268.19 60.86 ;
    RECT 267.91 61.05 267.98 61.12 ;
    RECT 265.73 60.79 265.94 60.86 ;
    RECT 262.9 61.05 263.11 61.12 ;
    RECT 263.36 61.05 263.57 61.12 ;
    RECT 147.275 60.79 147.345 60.86 ;
    RECT 147.485 61.05 147.555 61.12 ;
    RECT 166.62 61.05 166.83 61.12 ;
    RECT 167.08 61.05 167.29 61.12 ;
    RECT 203.14 61.05 203.35 61.12 ;
    RECT 203.6 61.05 203.81 61.12 ;
    RECT 162.81 60.79 163.02 60.86 ;
    RECT 226.38 61.05 226.59 61.12 ;
    RECT 245.81 60.79 246.02 60.86 ;
    RECT 226.84 61.05 227.05 61.12 ;
    RECT 192.69 60.79 192.9 60.86 ;
    RECT 196.5 61.05 196.71 61.12 ;
    RECT 196.96 61.05 197.17 61.12 ;
    RECT 259.09 60.79 259.3 60.86 ;
    RECT 239.17 60.79 239.38 60.86 ;
    RECT 219.74 61.05 219.95 61.12 ;
    RECT 220.2 61.05 220.41 61.12 ;
    RECT 242.98 61.05 243.19 61.12 ;
    RECT 243.44 61.05 243.65 61.12 ;
    RECT 159.98 61.05 160.19 61.12 ;
    RECT 160.44 61.05 160.65 61.12 ;
    RECT 256.26 61.05 256.47 61.12 ;
    RECT 186.05 60.79 186.26 60.86 ;
    RECT 256.72 61.05 256.93 61.12 ;
    RECT 209.29 60.79 209.5 60.86 ;
    RECT 179.41 60.79 179.62 60.86 ;
    RECT 156.17 60.79 156.38 60.86 ;
    RECT 252.45 60.79 252.66 60.86 ;
    RECT 213.1 61.05 213.31 61.12 ;
    RECT 232.53 60.79 232.74 60.86 ;
    RECT 213.56 61.05 213.77 61.12 ;
    RECT 236.34 61.05 236.55 61.12 ;
    RECT 236.8 61.05 237.01 61.12 ;
    RECT 153.34 61.05 153.55 61.12 ;
    RECT 153.8 61.05 154.01 61.12 ;
    RECT 176.58 61.05 176.79 61.12 ;
    RECT 177.04 61.05 177.25 61.12 ;
    RECT 249.62 61.05 249.83 61.12 ;
    RECT 250.08 61.05 250.29 61.12 ;
    RECT 189.86 61.05 190.07 61.12 ;
    RECT 190.32 61.05 190.53 61.12 ;
    RECT 202.65 60.79 202.86 60.86 ;
    RECT 222.57 60.79 222.78 60.86 ;
    RECT 172.77 60.79 172.98 60.86 ;
    RECT 149.53 60.79 149.74 60.86 ;
    RECT 229.7 61.05 229.91 61.12 ;
    RECT 230.16 61.05 230.37 61.12 ;
    RECT 266.22 61.05 266.43 61.12 ;
    RECT 266.68 61.05 266.89 61.12 ;
    RECT 169.94 61.05 170.15 61.12 ;
    RECT 170.4 61.05 170.61 61.12 ;
    RECT 183.22 61.05 183.43 61.12 ;
    RECT 225.89 60.79 226.1 60.86 ;
    RECT 183.68 61.05 183.89 61.12 ;
    RECT 206.46 61.05 206.67 61.12 ;
    RECT 206.92 61.05 207.13 61.12 ;
    RECT 196.01 60.79 196.22 60.86 ;
    RECT 215.93 60.79 216.14 60.86 ;
    RECT 166.13 60.79 166.34 60.86 ;
    RECT 262.41 60.79 262.62 60.86 ;
    RECT 246.3 61.05 246.51 61.12 ;
    RECT 246.76 61.05 246.97 61.12 ;
    RECT 163.3 61.05 163.51 61.12 ;
    RECT 163.76 61.05 163.97 61.12 ;
    RECT 199.82 61.05 200.03 61.12 ;
    RECT 200.28 61.05 200.49 61.12 ;
    RECT 223.06 61.05 223.27 61.12 ;
    RECT 242.49 60.79 242.7 60.86 ;
    RECT 223.52 61.05 223.73 61.12 ;
    RECT 259.58 61.05 259.79 61.12 ;
    RECT 260.04 61.05 260.25 61.12 ;
    RECT 189.37 60.79 189.58 60.86 ;
    RECT 250.08 96.57 250.29 96.64 ;
    RECT 250.08 96.93 250.29 97.0 ;
    RECT 250.08 97.29 250.29 97.36 ;
    RECT 249.62 96.57 249.83 96.64 ;
    RECT 249.62 96.93 249.83 97.0 ;
    RECT 249.62 97.29 249.83 97.36 ;
    RECT 246.76 96.57 246.97 96.64 ;
    RECT 246.76 96.93 246.97 97.0 ;
    RECT 246.76 97.29 246.97 97.36 ;
    RECT 246.3 96.57 246.51 96.64 ;
    RECT 246.3 96.93 246.51 97.0 ;
    RECT 246.3 97.29 246.51 97.36 ;
    RECT 243.44 96.57 243.65 96.64 ;
    RECT 243.44 96.93 243.65 97.0 ;
    RECT 243.44 97.29 243.65 97.36 ;
    RECT 242.98 96.57 243.19 96.64 ;
    RECT 242.98 96.93 243.19 97.0 ;
    RECT 242.98 97.29 243.19 97.36 ;
    RECT 240.12 96.57 240.33 96.64 ;
    RECT 240.12 96.93 240.33 97.0 ;
    RECT 240.12 97.29 240.33 97.36 ;
    RECT 239.66 96.57 239.87 96.64 ;
    RECT 239.66 96.93 239.87 97.0 ;
    RECT 239.66 97.29 239.87 97.36 ;
    RECT 236.8 96.57 237.01 96.64 ;
    RECT 236.8 96.93 237.01 97.0 ;
    RECT 236.8 97.29 237.01 97.36 ;
    RECT 236.34 96.57 236.55 96.64 ;
    RECT 236.34 96.93 236.55 97.0 ;
    RECT 236.34 97.29 236.55 97.36 ;
    RECT 233.48 96.57 233.69 96.64 ;
    RECT 233.48 96.93 233.69 97.0 ;
    RECT 233.48 97.29 233.69 97.36 ;
    RECT 233.02 96.57 233.23 96.64 ;
    RECT 233.02 96.93 233.23 97.0 ;
    RECT 233.02 97.29 233.23 97.36 ;
    RECT 230.16 96.57 230.37 96.64 ;
    RECT 230.16 96.93 230.37 97.0 ;
    RECT 230.16 97.29 230.37 97.36 ;
    RECT 229.7 96.57 229.91 96.64 ;
    RECT 229.7 96.93 229.91 97.0 ;
    RECT 229.7 97.29 229.91 97.36 ;
    RECT 226.84 96.57 227.05 96.64 ;
    RECT 226.84 96.93 227.05 97.0 ;
    RECT 226.84 97.29 227.05 97.36 ;
    RECT 226.38 96.57 226.59 96.64 ;
    RECT 226.38 96.93 226.59 97.0 ;
    RECT 226.38 97.29 226.59 97.36 ;
    RECT 223.52 96.57 223.73 96.64 ;
    RECT 223.52 96.93 223.73 97.0 ;
    RECT 223.52 97.29 223.73 97.36 ;
    RECT 223.06 96.57 223.27 96.64 ;
    RECT 223.06 96.93 223.27 97.0 ;
    RECT 223.06 97.29 223.27 97.36 ;
    RECT 220.2 96.57 220.41 96.64 ;
    RECT 220.2 96.93 220.41 97.0 ;
    RECT 220.2 97.29 220.41 97.36 ;
    RECT 219.74 96.57 219.95 96.64 ;
    RECT 219.74 96.93 219.95 97.0 ;
    RECT 219.74 97.29 219.95 97.36 ;
    RECT 216.88 96.57 217.09 96.64 ;
    RECT 216.88 96.93 217.09 97.0 ;
    RECT 216.88 97.29 217.09 97.36 ;
    RECT 216.42 96.57 216.63 96.64 ;
    RECT 216.42 96.93 216.63 97.0 ;
    RECT 216.42 97.29 216.63 97.36 ;
    RECT 267.91 96.93 267.98 97.0 ;
    RECT 180.36 96.57 180.57 96.64 ;
    RECT 180.36 96.93 180.57 97.0 ;
    RECT 180.36 97.29 180.57 97.36 ;
    RECT 179.9 96.57 180.11 96.64 ;
    RECT 179.9 96.93 180.11 97.0 ;
    RECT 179.9 97.29 180.11 97.36 ;
    RECT 177.04 96.57 177.25 96.64 ;
    RECT 177.04 96.93 177.25 97.0 ;
    RECT 177.04 97.29 177.25 97.36 ;
    RECT 176.58 96.57 176.79 96.64 ;
    RECT 176.58 96.93 176.79 97.0 ;
    RECT 176.58 97.29 176.79 97.36 ;
    RECT 173.72 96.57 173.93 96.64 ;
    RECT 173.72 96.93 173.93 97.0 ;
    RECT 173.72 97.29 173.93 97.36 ;
    RECT 173.26 96.57 173.47 96.64 ;
    RECT 173.26 96.93 173.47 97.0 ;
    RECT 173.26 97.29 173.47 97.36 ;
    RECT 170.4 96.57 170.61 96.64 ;
    RECT 170.4 96.93 170.61 97.0 ;
    RECT 170.4 97.29 170.61 97.36 ;
    RECT 169.94 96.57 170.15 96.64 ;
    RECT 169.94 96.93 170.15 97.0 ;
    RECT 169.94 97.29 170.15 97.36 ;
    RECT 167.08 96.57 167.29 96.64 ;
    RECT 167.08 96.93 167.29 97.0 ;
    RECT 167.08 97.29 167.29 97.36 ;
    RECT 166.62 96.57 166.83 96.64 ;
    RECT 166.62 96.93 166.83 97.0 ;
    RECT 166.62 97.29 166.83 97.36 ;
    RECT 163.76 96.57 163.97 96.64 ;
    RECT 163.76 96.93 163.97 97.0 ;
    RECT 163.76 97.29 163.97 97.36 ;
    RECT 163.3 96.57 163.51 96.64 ;
    RECT 163.3 96.93 163.51 97.0 ;
    RECT 163.3 97.29 163.51 97.36 ;
    RECT 160.44 96.57 160.65 96.64 ;
    RECT 160.44 96.93 160.65 97.0 ;
    RECT 160.44 97.29 160.65 97.36 ;
    RECT 159.98 96.57 160.19 96.64 ;
    RECT 159.98 96.93 160.19 97.0 ;
    RECT 159.98 97.29 160.19 97.36 ;
    RECT 157.12 96.57 157.33 96.64 ;
    RECT 157.12 96.93 157.33 97.0 ;
    RECT 157.12 97.29 157.33 97.36 ;
    RECT 156.66 96.57 156.87 96.64 ;
    RECT 156.66 96.93 156.87 97.0 ;
    RECT 156.66 97.29 156.87 97.36 ;
    RECT 153.8 96.57 154.01 96.64 ;
    RECT 153.8 96.93 154.01 97.0 ;
    RECT 153.8 97.29 154.01 97.36 ;
    RECT 153.34 96.57 153.55 96.64 ;
    RECT 153.34 96.93 153.55 97.0 ;
    RECT 153.34 97.29 153.55 97.36 ;
    RECT 150.48 96.57 150.69 96.64 ;
    RECT 150.48 96.93 150.69 97.0 ;
    RECT 150.48 97.29 150.69 97.36 ;
    RECT 150.02 96.57 150.23 96.64 ;
    RECT 150.02 96.93 150.23 97.0 ;
    RECT 150.02 97.29 150.23 97.36 ;
    RECT 213.56 96.57 213.77 96.64 ;
    RECT 213.56 96.93 213.77 97.0 ;
    RECT 213.56 97.29 213.77 97.36 ;
    RECT 213.1 96.57 213.31 96.64 ;
    RECT 213.1 96.93 213.31 97.0 ;
    RECT 213.1 97.29 213.31 97.36 ;
    RECT 210.24 96.57 210.45 96.64 ;
    RECT 210.24 96.93 210.45 97.0 ;
    RECT 210.24 97.29 210.45 97.36 ;
    RECT 209.78 96.57 209.99 96.64 ;
    RECT 209.78 96.93 209.99 97.0 ;
    RECT 209.78 97.29 209.99 97.36 ;
    RECT 206.92 96.57 207.13 96.64 ;
    RECT 206.92 96.93 207.13 97.0 ;
    RECT 206.92 97.29 207.13 97.36 ;
    RECT 206.46 96.57 206.67 96.64 ;
    RECT 206.46 96.93 206.67 97.0 ;
    RECT 206.46 97.29 206.67 97.36 ;
    RECT 203.6 96.57 203.81 96.64 ;
    RECT 203.6 96.93 203.81 97.0 ;
    RECT 203.6 97.29 203.81 97.36 ;
    RECT 203.14 96.57 203.35 96.64 ;
    RECT 203.14 96.93 203.35 97.0 ;
    RECT 203.14 97.29 203.35 97.36 ;
    RECT 200.28 96.57 200.49 96.64 ;
    RECT 200.28 96.93 200.49 97.0 ;
    RECT 200.28 97.29 200.49 97.36 ;
    RECT 199.82 96.57 200.03 96.64 ;
    RECT 199.82 96.93 200.03 97.0 ;
    RECT 199.82 97.29 200.03 97.36 ;
    RECT 196.96 96.57 197.17 96.64 ;
    RECT 196.96 96.93 197.17 97.0 ;
    RECT 196.96 97.29 197.17 97.36 ;
    RECT 196.5 96.57 196.71 96.64 ;
    RECT 196.5 96.93 196.71 97.0 ;
    RECT 196.5 97.29 196.71 97.36 ;
    RECT 193.64 96.57 193.85 96.64 ;
    RECT 193.64 96.93 193.85 97.0 ;
    RECT 193.64 97.29 193.85 97.36 ;
    RECT 193.18 96.57 193.39 96.64 ;
    RECT 193.18 96.93 193.39 97.0 ;
    RECT 193.18 97.29 193.39 97.36 ;
    RECT 190.32 96.57 190.53 96.64 ;
    RECT 190.32 96.93 190.53 97.0 ;
    RECT 190.32 97.29 190.53 97.36 ;
    RECT 189.86 96.57 190.07 96.64 ;
    RECT 189.86 96.93 190.07 97.0 ;
    RECT 189.86 97.29 190.07 97.36 ;
    RECT 187.0 96.57 187.21 96.64 ;
    RECT 187.0 96.93 187.21 97.0 ;
    RECT 187.0 97.29 187.21 97.36 ;
    RECT 186.54 96.57 186.75 96.64 ;
    RECT 186.54 96.93 186.75 97.0 ;
    RECT 186.54 97.29 186.75 97.36 ;
    RECT 183.68 96.57 183.89 96.64 ;
    RECT 183.68 96.93 183.89 97.0 ;
    RECT 183.68 97.29 183.89 97.36 ;
    RECT 183.22 96.57 183.43 96.64 ;
    RECT 183.22 96.93 183.43 97.0 ;
    RECT 183.22 97.29 183.43 97.36 ;
    RECT 147.485 96.93 147.555 97.0 ;
    RECT 266.68 96.57 266.89 96.64 ;
    RECT 266.68 96.93 266.89 97.0 ;
    RECT 266.68 97.29 266.89 97.36 ;
    RECT 266.22 96.57 266.43 96.64 ;
    RECT 266.22 96.93 266.43 97.0 ;
    RECT 266.22 97.29 266.43 97.36 ;
    RECT 263.36 96.57 263.57 96.64 ;
    RECT 263.36 96.93 263.57 97.0 ;
    RECT 263.36 97.29 263.57 97.36 ;
    RECT 262.9 96.57 263.11 96.64 ;
    RECT 262.9 96.93 263.11 97.0 ;
    RECT 262.9 97.29 263.11 97.36 ;
    RECT 260.04 96.57 260.25 96.64 ;
    RECT 260.04 96.93 260.25 97.0 ;
    RECT 260.04 97.29 260.25 97.36 ;
    RECT 259.58 96.57 259.79 96.64 ;
    RECT 259.58 96.93 259.79 97.0 ;
    RECT 259.58 97.29 259.79 97.36 ;
    RECT 256.72 96.57 256.93 96.64 ;
    RECT 256.72 96.93 256.93 97.0 ;
    RECT 256.72 97.29 256.93 97.36 ;
    RECT 256.26 96.57 256.47 96.64 ;
    RECT 256.26 96.93 256.47 97.0 ;
    RECT 256.26 97.29 256.47 97.36 ;
    RECT 253.4 96.57 253.61 96.64 ;
    RECT 253.4 96.93 253.61 97.0 ;
    RECT 253.4 97.29 253.61 97.36 ;
    RECT 252.94 96.57 253.15 96.64 ;
    RECT 252.94 96.93 253.15 97.0 ;
    RECT 252.94 97.29 253.15 97.36 ;
    RECT 250.08 59.83 250.29 59.9 ;
    RECT 250.08 60.19 250.29 60.26 ;
    RECT 250.08 60.55 250.29 60.62 ;
    RECT 249.62 59.83 249.83 59.9 ;
    RECT 249.62 60.19 249.83 60.26 ;
    RECT 249.62 60.55 249.83 60.62 ;
    RECT 246.76 59.83 246.97 59.9 ;
    RECT 246.76 60.19 246.97 60.26 ;
    RECT 246.76 60.55 246.97 60.62 ;
    RECT 246.3 59.83 246.51 59.9 ;
    RECT 246.3 60.19 246.51 60.26 ;
    RECT 246.3 60.55 246.51 60.62 ;
    RECT 243.44 59.83 243.65 59.9 ;
    RECT 243.44 60.19 243.65 60.26 ;
    RECT 243.44 60.55 243.65 60.62 ;
    RECT 242.98 59.83 243.19 59.9 ;
    RECT 242.98 60.19 243.19 60.26 ;
    RECT 242.98 60.55 243.19 60.62 ;
    RECT 240.12 59.83 240.33 59.9 ;
    RECT 240.12 60.19 240.33 60.26 ;
    RECT 240.12 60.55 240.33 60.62 ;
    RECT 239.66 59.83 239.87 59.9 ;
    RECT 239.66 60.19 239.87 60.26 ;
    RECT 239.66 60.55 239.87 60.62 ;
    RECT 236.8 59.83 237.01 59.9 ;
    RECT 236.8 60.19 237.01 60.26 ;
    RECT 236.8 60.55 237.01 60.62 ;
    RECT 236.34 59.83 236.55 59.9 ;
    RECT 236.34 60.19 236.55 60.26 ;
    RECT 236.34 60.55 236.55 60.62 ;
    RECT 233.48 59.83 233.69 59.9 ;
    RECT 233.48 60.19 233.69 60.26 ;
    RECT 233.48 60.55 233.69 60.62 ;
    RECT 233.02 59.83 233.23 59.9 ;
    RECT 233.02 60.19 233.23 60.26 ;
    RECT 233.02 60.55 233.23 60.62 ;
    RECT 230.16 59.83 230.37 59.9 ;
    RECT 230.16 60.19 230.37 60.26 ;
    RECT 230.16 60.55 230.37 60.62 ;
    RECT 229.7 59.83 229.91 59.9 ;
    RECT 229.7 60.19 229.91 60.26 ;
    RECT 229.7 60.55 229.91 60.62 ;
    RECT 226.84 59.83 227.05 59.9 ;
    RECT 226.84 60.19 227.05 60.26 ;
    RECT 226.84 60.55 227.05 60.62 ;
    RECT 226.38 59.83 226.59 59.9 ;
    RECT 226.38 60.19 226.59 60.26 ;
    RECT 226.38 60.55 226.59 60.62 ;
    RECT 223.52 59.83 223.73 59.9 ;
    RECT 223.52 60.19 223.73 60.26 ;
    RECT 223.52 60.55 223.73 60.62 ;
    RECT 223.06 59.83 223.27 59.9 ;
    RECT 223.06 60.19 223.27 60.26 ;
    RECT 223.06 60.55 223.27 60.62 ;
    RECT 220.2 59.83 220.41 59.9 ;
    RECT 220.2 60.19 220.41 60.26 ;
    RECT 220.2 60.55 220.41 60.62 ;
    RECT 219.74 59.83 219.95 59.9 ;
    RECT 219.74 60.19 219.95 60.26 ;
    RECT 219.74 60.55 219.95 60.62 ;
    RECT 216.88 59.83 217.09 59.9 ;
    RECT 216.88 60.19 217.09 60.26 ;
    RECT 216.88 60.55 217.09 60.62 ;
    RECT 216.42 59.83 216.63 59.9 ;
    RECT 216.42 60.19 216.63 60.26 ;
    RECT 216.42 60.55 216.63 60.62 ;
    RECT 267.91 60.19 267.98 60.26 ;
    RECT 180.36 59.83 180.57 59.9 ;
    RECT 180.36 60.19 180.57 60.26 ;
    RECT 180.36 60.55 180.57 60.62 ;
    RECT 179.9 59.83 180.11 59.9 ;
    RECT 179.9 60.19 180.11 60.26 ;
    RECT 179.9 60.55 180.11 60.62 ;
    RECT 177.04 59.83 177.25 59.9 ;
    RECT 177.04 60.19 177.25 60.26 ;
    RECT 177.04 60.55 177.25 60.62 ;
    RECT 176.58 59.83 176.79 59.9 ;
    RECT 176.58 60.19 176.79 60.26 ;
    RECT 176.58 60.55 176.79 60.62 ;
    RECT 173.72 59.83 173.93 59.9 ;
    RECT 173.72 60.19 173.93 60.26 ;
    RECT 173.72 60.55 173.93 60.62 ;
    RECT 173.26 59.83 173.47 59.9 ;
    RECT 173.26 60.19 173.47 60.26 ;
    RECT 173.26 60.55 173.47 60.62 ;
    RECT 170.4 59.83 170.61 59.9 ;
    RECT 170.4 60.19 170.61 60.26 ;
    RECT 170.4 60.55 170.61 60.62 ;
    RECT 169.94 59.83 170.15 59.9 ;
    RECT 169.94 60.19 170.15 60.26 ;
    RECT 169.94 60.55 170.15 60.62 ;
    RECT 167.08 59.83 167.29 59.9 ;
    RECT 167.08 60.19 167.29 60.26 ;
    RECT 167.08 60.55 167.29 60.62 ;
    RECT 166.62 59.83 166.83 59.9 ;
    RECT 166.62 60.19 166.83 60.26 ;
    RECT 166.62 60.55 166.83 60.62 ;
    RECT 163.76 59.83 163.97 59.9 ;
    RECT 163.76 60.19 163.97 60.26 ;
    RECT 163.76 60.55 163.97 60.62 ;
    RECT 163.3 59.83 163.51 59.9 ;
    RECT 163.3 60.19 163.51 60.26 ;
    RECT 163.3 60.55 163.51 60.62 ;
    RECT 160.44 59.83 160.65 59.9 ;
    RECT 160.44 60.19 160.65 60.26 ;
    RECT 160.44 60.55 160.65 60.62 ;
    RECT 159.98 59.83 160.19 59.9 ;
    RECT 159.98 60.19 160.19 60.26 ;
    RECT 159.98 60.55 160.19 60.62 ;
    RECT 157.12 59.83 157.33 59.9 ;
    RECT 157.12 60.19 157.33 60.26 ;
    RECT 157.12 60.55 157.33 60.62 ;
    RECT 156.66 59.83 156.87 59.9 ;
    RECT 156.66 60.19 156.87 60.26 ;
    RECT 156.66 60.55 156.87 60.62 ;
    RECT 153.8 59.83 154.01 59.9 ;
    RECT 153.8 60.19 154.01 60.26 ;
    RECT 153.8 60.55 154.01 60.62 ;
    RECT 153.34 59.83 153.55 59.9 ;
    RECT 153.34 60.19 153.55 60.26 ;
    RECT 153.34 60.55 153.55 60.62 ;
    RECT 150.48 59.83 150.69 59.9 ;
    RECT 150.48 60.19 150.69 60.26 ;
    RECT 150.48 60.55 150.69 60.62 ;
    RECT 150.02 59.83 150.23 59.9 ;
    RECT 150.02 60.19 150.23 60.26 ;
    RECT 150.02 60.55 150.23 60.62 ;
    RECT 213.56 59.83 213.77 59.9 ;
    RECT 213.56 60.19 213.77 60.26 ;
    RECT 213.56 60.55 213.77 60.62 ;
    RECT 213.1 59.83 213.31 59.9 ;
    RECT 213.1 60.19 213.31 60.26 ;
    RECT 213.1 60.55 213.31 60.62 ;
    RECT 210.24 59.83 210.45 59.9 ;
    RECT 210.24 60.19 210.45 60.26 ;
    RECT 210.24 60.55 210.45 60.62 ;
    RECT 209.78 59.83 209.99 59.9 ;
    RECT 209.78 60.19 209.99 60.26 ;
    RECT 209.78 60.55 209.99 60.62 ;
    RECT 206.92 59.83 207.13 59.9 ;
    RECT 206.92 60.19 207.13 60.26 ;
    RECT 206.92 60.55 207.13 60.62 ;
    RECT 206.46 59.83 206.67 59.9 ;
    RECT 206.46 60.19 206.67 60.26 ;
    RECT 206.46 60.55 206.67 60.62 ;
    RECT 203.6 59.83 203.81 59.9 ;
    RECT 203.6 60.19 203.81 60.26 ;
    RECT 203.6 60.55 203.81 60.62 ;
    RECT 203.14 59.83 203.35 59.9 ;
    RECT 203.14 60.19 203.35 60.26 ;
    RECT 203.14 60.55 203.35 60.62 ;
    RECT 200.28 59.83 200.49 59.9 ;
    RECT 200.28 60.19 200.49 60.26 ;
    RECT 200.28 60.55 200.49 60.62 ;
    RECT 199.82 59.83 200.03 59.9 ;
    RECT 199.82 60.19 200.03 60.26 ;
    RECT 199.82 60.55 200.03 60.62 ;
    RECT 196.96 59.83 197.17 59.9 ;
    RECT 196.96 60.19 197.17 60.26 ;
    RECT 196.96 60.55 197.17 60.62 ;
    RECT 196.5 59.83 196.71 59.9 ;
    RECT 196.5 60.19 196.71 60.26 ;
    RECT 196.5 60.55 196.71 60.62 ;
    RECT 193.64 59.83 193.85 59.9 ;
    RECT 193.64 60.19 193.85 60.26 ;
    RECT 193.64 60.55 193.85 60.62 ;
    RECT 193.18 59.83 193.39 59.9 ;
    RECT 193.18 60.19 193.39 60.26 ;
    RECT 193.18 60.55 193.39 60.62 ;
    RECT 190.32 59.83 190.53 59.9 ;
    RECT 190.32 60.19 190.53 60.26 ;
    RECT 190.32 60.55 190.53 60.62 ;
    RECT 189.86 59.83 190.07 59.9 ;
    RECT 189.86 60.19 190.07 60.26 ;
    RECT 189.86 60.55 190.07 60.62 ;
    RECT 187.0 59.83 187.21 59.9 ;
    RECT 187.0 60.19 187.21 60.26 ;
    RECT 187.0 60.55 187.21 60.62 ;
    RECT 186.54 59.83 186.75 59.9 ;
    RECT 186.54 60.19 186.75 60.26 ;
    RECT 186.54 60.55 186.75 60.62 ;
    RECT 183.68 59.83 183.89 59.9 ;
    RECT 183.68 60.19 183.89 60.26 ;
    RECT 183.68 60.55 183.89 60.62 ;
    RECT 183.22 59.83 183.43 59.9 ;
    RECT 183.22 60.19 183.43 60.26 ;
    RECT 183.22 60.55 183.43 60.62 ;
    RECT 147.485 60.19 147.555 60.26 ;
    RECT 266.68 59.83 266.89 59.9 ;
    RECT 266.68 60.19 266.89 60.26 ;
    RECT 266.68 60.55 266.89 60.62 ;
    RECT 266.22 59.83 266.43 59.9 ;
    RECT 266.22 60.19 266.43 60.26 ;
    RECT 266.22 60.55 266.43 60.62 ;
    RECT 263.36 59.83 263.57 59.9 ;
    RECT 263.36 60.19 263.57 60.26 ;
    RECT 263.36 60.55 263.57 60.62 ;
    RECT 262.9 59.83 263.11 59.9 ;
    RECT 262.9 60.19 263.11 60.26 ;
    RECT 262.9 60.55 263.11 60.62 ;
    RECT 260.04 59.83 260.25 59.9 ;
    RECT 260.04 60.19 260.25 60.26 ;
    RECT 260.04 60.55 260.25 60.62 ;
    RECT 259.58 59.83 259.79 59.9 ;
    RECT 259.58 60.19 259.79 60.26 ;
    RECT 259.58 60.55 259.79 60.62 ;
    RECT 256.72 59.83 256.93 59.9 ;
    RECT 256.72 60.19 256.93 60.26 ;
    RECT 256.72 60.55 256.93 60.62 ;
    RECT 256.26 59.83 256.47 59.9 ;
    RECT 256.26 60.19 256.47 60.26 ;
    RECT 256.26 60.55 256.47 60.62 ;
    RECT 253.4 59.83 253.61 59.9 ;
    RECT 253.4 60.19 253.61 60.26 ;
    RECT 253.4 60.55 253.61 60.62 ;
    RECT 252.94 59.83 253.15 59.9 ;
    RECT 252.94 60.19 253.15 60.26 ;
    RECT 252.94 60.55 253.15 60.62 ;
    RECT 250.08 95.85 250.29 95.92 ;
    RECT 250.08 96.21 250.29 96.28 ;
    RECT 250.08 96.57 250.29 96.64 ;
    RECT 249.62 95.85 249.83 95.92 ;
    RECT 249.62 96.21 249.83 96.28 ;
    RECT 249.62 96.57 249.83 96.64 ;
    RECT 246.76 95.85 246.97 95.92 ;
    RECT 246.76 96.21 246.97 96.28 ;
    RECT 246.76 96.57 246.97 96.64 ;
    RECT 246.3 95.85 246.51 95.92 ;
    RECT 246.3 96.21 246.51 96.28 ;
    RECT 246.3 96.57 246.51 96.64 ;
    RECT 243.44 95.85 243.65 95.92 ;
    RECT 243.44 96.21 243.65 96.28 ;
    RECT 243.44 96.57 243.65 96.64 ;
    RECT 242.98 95.85 243.19 95.92 ;
    RECT 242.98 96.21 243.19 96.28 ;
    RECT 242.98 96.57 243.19 96.64 ;
    RECT 240.12 95.85 240.33 95.92 ;
    RECT 240.12 96.21 240.33 96.28 ;
    RECT 240.12 96.57 240.33 96.64 ;
    RECT 239.66 95.85 239.87 95.92 ;
    RECT 239.66 96.21 239.87 96.28 ;
    RECT 239.66 96.57 239.87 96.64 ;
    RECT 236.8 95.85 237.01 95.92 ;
    RECT 236.8 96.21 237.01 96.28 ;
    RECT 236.8 96.57 237.01 96.64 ;
    RECT 236.34 95.85 236.55 95.92 ;
    RECT 236.34 96.21 236.55 96.28 ;
    RECT 236.34 96.57 236.55 96.64 ;
    RECT 233.48 95.85 233.69 95.92 ;
    RECT 233.48 96.21 233.69 96.28 ;
    RECT 233.48 96.57 233.69 96.64 ;
    RECT 233.02 95.85 233.23 95.92 ;
    RECT 233.02 96.21 233.23 96.28 ;
    RECT 233.02 96.57 233.23 96.64 ;
    RECT 230.16 95.85 230.37 95.92 ;
    RECT 230.16 96.21 230.37 96.28 ;
    RECT 230.16 96.57 230.37 96.64 ;
    RECT 229.7 95.85 229.91 95.92 ;
    RECT 229.7 96.21 229.91 96.28 ;
    RECT 229.7 96.57 229.91 96.64 ;
    RECT 226.84 95.85 227.05 95.92 ;
    RECT 226.84 96.21 227.05 96.28 ;
    RECT 226.84 96.57 227.05 96.64 ;
    RECT 226.38 95.85 226.59 95.92 ;
    RECT 226.38 96.21 226.59 96.28 ;
    RECT 226.38 96.57 226.59 96.64 ;
    RECT 223.52 95.85 223.73 95.92 ;
    RECT 223.52 96.21 223.73 96.28 ;
    RECT 223.52 96.57 223.73 96.64 ;
    RECT 223.06 95.85 223.27 95.92 ;
    RECT 223.06 96.21 223.27 96.28 ;
    RECT 223.06 96.57 223.27 96.64 ;
    RECT 220.2 95.85 220.41 95.92 ;
    RECT 220.2 96.21 220.41 96.28 ;
    RECT 220.2 96.57 220.41 96.64 ;
    RECT 219.74 95.85 219.95 95.92 ;
    RECT 219.74 96.21 219.95 96.28 ;
    RECT 219.74 96.57 219.95 96.64 ;
    RECT 216.88 95.85 217.09 95.92 ;
    RECT 216.88 96.21 217.09 96.28 ;
    RECT 216.88 96.57 217.09 96.64 ;
    RECT 216.42 95.85 216.63 95.92 ;
    RECT 216.42 96.21 216.63 96.28 ;
    RECT 216.42 96.57 216.63 96.64 ;
    RECT 267.91 96.21 267.98 96.28 ;
    RECT 180.36 95.85 180.57 95.92 ;
    RECT 180.36 96.21 180.57 96.28 ;
    RECT 180.36 96.57 180.57 96.64 ;
    RECT 179.9 95.85 180.11 95.92 ;
    RECT 179.9 96.21 180.11 96.28 ;
    RECT 179.9 96.57 180.11 96.64 ;
    RECT 177.04 95.85 177.25 95.92 ;
    RECT 177.04 96.21 177.25 96.28 ;
    RECT 177.04 96.57 177.25 96.64 ;
    RECT 176.58 95.85 176.79 95.92 ;
    RECT 176.58 96.21 176.79 96.28 ;
    RECT 176.58 96.57 176.79 96.64 ;
    RECT 173.72 95.85 173.93 95.92 ;
    RECT 173.72 96.21 173.93 96.28 ;
    RECT 173.72 96.57 173.93 96.64 ;
    RECT 173.26 95.85 173.47 95.92 ;
    RECT 173.26 96.21 173.47 96.28 ;
    RECT 173.26 96.57 173.47 96.64 ;
    RECT 170.4 95.85 170.61 95.92 ;
    RECT 170.4 96.21 170.61 96.28 ;
    RECT 170.4 96.57 170.61 96.64 ;
    RECT 169.94 95.85 170.15 95.92 ;
    RECT 169.94 96.21 170.15 96.28 ;
    RECT 169.94 96.57 170.15 96.64 ;
    RECT 167.08 95.85 167.29 95.92 ;
    RECT 167.08 96.21 167.29 96.28 ;
    RECT 167.08 96.57 167.29 96.64 ;
    RECT 166.62 95.85 166.83 95.92 ;
    RECT 166.62 96.21 166.83 96.28 ;
    RECT 166.62 96.57 166.83 96.64 ;
    RECT 163.76 95.85 163.97 95.92 ;
    RECT 163.76 96.21 163.97 96.28 ;
    RECT 163.76 96.57 163.97 96.64 ;
    RECT 163.3 95.85 163.51 95.92 ;
    RECT 163.3 96.21 163.51 96.28 ;
    RECT 163.3 96.57 163.51 96.64 ;
    RECT 160.44 95.85 160.65 95.92 ;
    RECT 160.44 96.21 160.65 96.28 ;
    RECT 160.44 96.57 160.65 96.64 ;
    RECT 159.98 95.85 160.19 95.92 ;
    RECT 159.98 96.21 160.19 96.28 ;
    RECT 159.98 96.57 160.19 96.64 ;
    RECT 157.12 95.85 157.33 95.92 ;
    RECT 157.12 96.21 157.33 96.28 ;
    RECT 157.12 96.57 157.33 96.64 ;
    RECT 156.66 95.85 156.87 95.92 ;
    RECT 156.66 96.21 156.87 96.28 ;
    RECT 156.66 96.57 156.87 96.64 ;
    RECT 153.8 95.85 154.01 95.92 ;
    RECT 153.8 96.21 154.01 96.28 ;
    RECT 153.8 96.57 154.01 96.64 ;
    RECT 153.34 95.85 153.55 95.92 ;
    RECT 153.34 96.21 153.55 96.28 ;
    RECT 153.34 96.57 153.55 96.64 ;
    RECT 150.48 95.85 150.69 95.92 ;
    RECT 150.48 96.21 150.69 96.28 ;
    RECT 150.48 96.57 150.69 96.64 ;
    RECT 150.02 95.85 150.23 95.92 ;
    RECT 150.02 96.21 150.23 96.28 ;
    RECT 150.02 96.57 150.23 96.64 ;
    RECT 213.56 95.85 213.77 95.92 ;
    RECT 213.56 96.21 213.77 96.28 ;
    RECT 213.56 96.57 213.77 96.64 ;
    RECT 213.1 95.85 213.31 95.92 ;
    RECT 213.1 96.21 213.31 96.28 ;
    RECT 213.1 96.57 213.31 96.64 ;
    RECT 210.24 95.85 210.45 95.92 ;
    RECT 210.24 96.21 210.45 96.28 ;
    RECT 210.24 96.57 210.45 96.64 ;
    RECT 209.78 95.85 209.99 95.92 ;
    RECT 209.78 96.21 209.99 96.28 ;
    RECT 209.78 96.57 209.99 96.64 ;
    RECT 206.92 95.85 207.13 95.92 ;
    RECT 206.92 96.21 207.13 96.28 ;
    RECT 206.92 96.57 207.13 96.64 ;
    RECT 206.46 95.85 206.67 95.92 ;
    RECT 206.46 96.21 206.67 96.28 ;
    RECT 206.46 96.57 206.67 96.64 ;
    RECT 203.6 95.85 203.81 95.92 ;
    RECT 203.6 96.21 203.81 96.28 ;
    RECT 203.6 96.57 203.81 96.64 ;
    RECT 203.14 95.85 203.35 95.92 ;
    RECT 203.14 96.21 203.35 96.28 ;
    RECT 203.14 96.57 203.35 96.64 ;
    RECT 200.28 95.85 200.49 95.92 ;
    RECT 200.28 96.21 200.49 96.28 ;
    RECT 200.28 96.57 200.49 96.64 ;
    RECT 199.82 95.85 200.03 95.92 ;
    RECT 199.82 96.21 200.03 96.28 ;
    RECT 199.82 96.57 200.03 96.64 ;
    RECT 196.96 95.85 197.17 95.92 ;
    RECT 196.96 96.21 197.17 96.28 ;
    RECT 196.96 96.57 197.17 96.64 ;
    RECT 196.5 95.85 196.71 95.92 ;
    RECT 196.5 96.21 196.71 96.28 ;
    RECT 196.5 96.57 196.71 96.64 ;
    RECT 193.64 95.85 193.85 95.92 ;
    RECT 193.64 96.21 193.85 96.28 ;
    RECT 193.64 96.57 193.85 96.64 ;
    RECT 193.18 95.85 193.39 95.92 ;
    RECT 193.18 96.21 193.39 96.28 ;
    RECT 193.18 96.57 193.39 96.64 ;
    RECT 190.32 95.85 190.53 95.92 ;
    RECT 190.32 96.21 190.53 96.28 ;
    RECT 190.32 96.57 190.53 96.64 ;
    RECT 189.86 95.85 190.07 95.92 ;
    RECT 189.86 96.21 190.07 96.28 ;
    RECT 189.86 96.57 190.07 96.64 ;
    RECT 187.0 95.85 187.21 95.92 ;
    RECT 187.0 96.21 187.21 96.28 ;
    RECT 187.0 96.57 187.21 96.64 ;
    RECT 186.54 95.85 186.75 95.92 ;
    RECT 186.54 96.21 186.75 96.28 ;
    RECT 186.54 96.57 186.75 96.64 ;
    RECT 183.68 95.85 183.89 95.92 ;
    RECT 183.68 96.21 183.89 96.28 ;
    RECT 183.68 96.57 183.89 96.64 ;
    RECT 183.22 95.85 183.43 95.92 ;
    RECT 183.22 96.21 183.43 96.28 ;
    RECT 183.22 96.57 183.43 96.64 ;
    RECT 147.485 96.21 147.555 96.28 ;
    RECT 266.68 95.85 266.89 95.92 ;
    RECT 266.68 96.21 266.89 96.28 ;
    RECT 266.68 96.57 266.89 96.64 ;
    RECT 266.22 95.85 266.43 95.92 ;
    RECT 266.22 96.21 266.43 96.28 ;
    RECT 266.22 96.57 266.43 96.64 ;
    RECT 263.36 95.85 263.57 95.92 ;
    RECT 263.36 96.21 263.57 96.28 ;
    RECT 263.36 96.57 263.57 96.64 ;
    RECT 262.9 95.85 263.11 95.92 ;
    RECT 262.9 96.21 263.11 96.28 ;
    RECT 262.9 96.57 263.11 96.64 ;
    RECT 260.04 95.85 260.25 95.92 ;
    RECT 260.04 96.21 260.25 96.28 ;
    RECT 260.04 96.57 260.25 96.64 ;
    RECT 259.58 95.85 259.79 95.92 ;
    RECT 259.58 96.21 259.79 96.28 ;
    RECT 259.58 96.57 259.79 96.64 ;
    RECT 256.72 95.85 256.93 95.92 ;
    RECT 256.72 96.21 256.93 96.28 ;
    RECT 256.72 96.57 256.93 96.64 ;
    RECT 256.26 95.85 256.47 95.92 ;
    RECT 256.26 96.21 256.47 96.28 ;
    RECT 256.26 96.57 256.47 96.64 ;
    RECT 253.4 95.85 253.61 95.92 ;
    RECT 253.4 96.21 253.61 96.28 ;
    RECT 253.4 96.57 253.61 96.64 ;
    RECT 252.94 95.85 253.15 95.92 ;
    RECT 252.94 96.21 253.15 96.28 ;
    RECT 252.94 96.57 253.15 96.64 ;
    RECT 250.08 59.11 250.29 59.18 ;
    RECT 250.08 59.47 250.29 59.54 ;
    RECT 250.08 59.83 250.29 59.9 ;
    RECT 249.62 59.11 249.83 59.18 ;
    RECT 249.62 59.47 249.83 59.54 ;
    RECT 249.62 59.83 249.83 59.9 ;
    RECT 246.76 59.11 246.97 59.18 ;
    RECT 246.76 59.47 246.97 59.54 ;
    RECT 246.76 59.83 246.97 59.9 ;
    RECT 246.3 59.11 246.51 59.18 ;
    RECT 246.3 59.47 246.51 59.54 ;
    RECT 246.3 59.83 246.51 59.9 ;
    RECT 243.44 59.11 243.65 59.18 ;
    RECT 243.44 59.47 243.65 59.54 ;
    RECT 243.44 59.83 243.65 59.9 ;
    RECT 242.98 59.11 243.19 59.18 ;
    RECT 242.98 59.47 243.19 59.54 ;
    RECT 242.98 59.83 243.19 59.9 ;
    RECT 240.12 59.11 240.33 59.18 ;
    RECT 240.12 59.47 240.33 59.54 ;
    RECT 240.12 59.83 240.33 59.9 ;
    RECT 239.66 59.11 239.87 59.18 ;
    RECT 239.66 59.47 239.87 59.54 ;
    RECT 239.66 59.83 239.87 59.9 ;
    RECT 236.8 59.11 237.01 59.18 ;
    RECT 236.8 59.47 237.01 59.54 ;
    RECT 236.8 59.83 237.01 59.9 ;
    RECT 236.34 59.11 236.55 59.18 ;
    RECT 236.34 59.47 236.55 59.54 ;
    RECT 236.34 59.83 236.55 59.9 ;
    RECT 233.48 59.11 233.69 59.18 ;
    RECT 233.48 59.47 233.69 59.54 ;
    RECT 233.48 59.83 233.69 59.9 ;
    RECT 233.02 59.11 233.23 59.18 ;
    RECT 233.02 59.47 233.23 59.54 ;
    RECT 233.02 59.83 233.23 59.9 ;
    RECT 230.16 59.11 230.37 59.18 ;
    RECT 230.16 59.47 230.37 59.54 ;
    RECT 230.16 59.83 230.37 59.9 ;
    RECT 229.7 59.11 229.91 59.18 ;
    RECT 229.7 59.47 229.91 59.54 ;
    RECT 229.7 59.83 229.91 59.9 ;
    RECT 226.84 59.11 227.05 59.18 ;
    RECT 226.84 59.47 227.05 59.54 ;
    RECT 226.84 59.83 227.05 59.9 ;
    RECT 226.38 59.11 226.59 59.18 ;
    RECT 226.38 59.47 226.59 59.54 ;
    RECT 226.38 59.83 226.59 59.9 ;
    RECT 223.52 59.11 223.73 59.18 ;
    RECT 223.52 59.47 223.73 59.54 ;
    RECT 223.52 59.83 223.73 59.9 ;
    RECT 223.06 59.11 223.27 59.18 ;
    RECT 223.06 59.47 223.27 59.54 ;
    RECT 223.06 59.83 223.27 59.9 ;
    RECT 220.2 59.11 220.41 59.18 ;
    RECT 220.2 59.47 220.41 59.54 ;
    RECT 220.2 59.83 220.41 59.9 ;
    RECT 219.74 59.11 219.95 59.18 ;
    RECT 219.74 59.47 219.95 59.54 ;
    RECT 219.74 59.83 219.95 59.9 ;
    RECT 216.88 59.11 217.09 59.18 ;
    RECT 216.88 59.47 217.09 59.54 ;
    RECT 216.88 59.83 217.09 59.9 ;
    RECT 216.42 59.11 216.63 59.18 ;
    RECT 216.42 59.47 216.63 59.54 ;
    RECT 216.42 59.83 216.63 59.9 ;
    RECT 267.91 59.47 267.98 59.54 ;
    RECT 180.36 59.11 180.57 59.18 ;
    RECT 180.36 59.47 180.57 59.54 ;
    RECT 180.36 59.83 180.57 59.9 ;
    RECT 179.9 59.11 180.11 59.18 ;
    RECT 179.9 59.47 180.11 59.54 ;
    RECT 179.9 59.83 180.11 59.9 ;
    RECT 177.04 59.11 177.25 59.18 ;
    RECT 177.04 59.47 177.25 59.54 ;
    RECT 177.04 59.83 177.25 59.9 ;
    RECT 176.58 59.11 176.79 59.18 ;
    RECT 176.58 59.47 176.79 59.54 ;
    RECT 176.58 59.83 176.79 59.9 ;
    RECT 173.72 59.11 173.93 59.18 ;
    RECT 173.72 59.47 173.93 59.54 ;
    RECT 173.72 59.83 173.93 59.9 ;
    RECT 173.26 59.11 173.47 59.18 ;
    RECT 173.26 59.47 173.47 59.54 ;
    RECT 173.26 59.83 173.47 59.9 ;
    RECT 170.4 59.11 170.61 59.18 ;
    RECT 170.4 59.47 170.61 59.54 ;
    RECT 170.4 59.83 170.61 59.9 ;
    RECT 169.94 59.11 170.15 59.18 ;
    RECT 169.94 59.47 170.15 59.54 ;
    RECT 169.94 59.83 170.15 59.9 ;
    RECT 167.08 59.11 167.29 59.18 ;
    RECT 167.08 59.47 167.29 59.54 ;
    RECT 167.08 59.83 167.29 59.9 ;
    RECT 166.62 59.11 166.83 59.18 ;
    RECT 166.62 59.47 166.83 59.54 ;
    RECT 166.62 59.83 166.83 59.9 ;
    RECT 163.76 59.11 163.97 59.18 ;
    RECT 163.76 59.47 163.97 59.54 ;
    RECT 163.76 59.83 163.97 59.9 ;
    RECT 163.3 59.11 163.51 59.18 ;
    RECT 163.3 59.47 163.51 59.54 ;
    RECT 163.3 59.83 163.51 59.9 ;
    RECT 160.44 59.11 160.65 59.18 ;
    RECT 160.44 59.47 160.65 59.54 ;
    RECT 160.44 59.83 160.65 59.9 ;
    RECT 159.98 59.11 160.19 59.18 ;
    RECT 159.98 59.47 160.19 59.54 ;
    RECT 159.98 59.83 160.19 59.9 ;
    RECT 157.12 59.11 157.33 59.18 ;
    RECT 157.12 59.47 157.33 59.54 ;
    RECT 157.12 59.83 157.33 59.9 ;
    RECT 156.66 59.11 156.87 59.18 ;
    RECT 156.66 59.47 156.87 59.54 ;
    RECT 156.66 59.83 156.87 59.9 ;
    RECT 153.8 59.11 154.01 59.18 ;
    RECT 153.8 59.47 154.01 59.54 ;
    RECT 153.8 59.83 154.01 59.9 ;
    RECT 153.34 59.11 153.55 59.18 ;
    RECT 153.34 59.47 153.55 59.54 ;
    RECT 153.34 59.83 153.55 59.9 ;
    RECT 150.48 59.11 150.69 59.18 ;
    RECT 150.48 59.47 150.69 59.54 ;
    RECT 150.48 59.83 150.69 59.9 ;
    RECT 150.02 59.11 150.23 59.18 ;
    RECT 150.02 59.47 150.23 59.54 ;
    RECT 150.02 59.83 150.23 59.9 ;
    RECT 213.56 59.11 213.77 59.18 ;
    RECT 213.56 59.47 213.77 59.54 ;
    RECT 213.56 59.83 213.77 59.9 ;
    RECT 213.1 59.11 213.31 59.18 ;
    RECT 213.1 59.47 213.31 59.54 ;
    RECT 213.1 59.83 213.31 59.9 ;
    RECT 210.24 59.11 210.45 59.18 ;
    RECT 210.24 59.47 210.45 59.54 ;
    RECT 210.24 59.83 210.45 59.9 ;
    RECT 209.78 59.11 209.99 59.18 ;
    RECT 209.78 59.47 209.99 59.54 ;
    RECT 209.78 59.83 209.99 59.9 ;
    RECT 206.92 59.11 207.13 59.18 ;
    RECT 206.92 59.47 207.13 59.54 ;
    RECT 206.92 59.83 207.13 59.9 ;
    RECT 206.46 59.11 206.67 59.18 ;
    RECT 206.46 59.47 206.67 59.54 ;
    RECT 206.46 59.83 206.67 59.9 ;
    RECT 203.6 59.11 203.81 59.18 ;
    RECT 203.6 59.47 203.81 59.54 ;
    RECT 203.6 59.83 203.81 59.9 ;
    RECT 203.14 59.11 203.35 59.18 ;
    RECT 203.14 59.47 203.35 59.54 ;
    RECT 203.14 59.83 203.35 59.9 ;
    RECT 200.28 59.11 200.49 59.18 ;
    RECT 200.28 59.47 200.49 59.54 ;
    RECT 200.28 59.83 200.49 59.9 ;
    RECT 199.82 59.11 200.03 59.18 ;
    RECT 199.82 59.47 200.03 59.54 ;
    RECT 199.82 59.83 200.03 59.9 ;
    RECT 196.96 59.11 197.17 59.18 ;
    RECT 196.96 59.47 197.17 59.54 ;
    RECT 196.96 59.83 197.17 59.9 ;
    RECT 196.5 59.11 196.71 59.18 ;
    RECT 196.5 59.47 196.71 59.54 ;
    RECT 196.5 59.83 196.71 59.9 ;
    RECT 193.64 59.11 193.85 59.18 ;
    RECT 193.64 59.47 193.85 59.54 ;
    RECT 193.64 59.83 193.85 59.9 ;
    RECT 193.18 59.11 193.39 59.18 ;
    RECT 193.18 59.47 193.39 59.54 ;
    RECT 193.18 59.83 193.39 59.9 ;
    RECT 190.32 59.11 190.53 59.18 ;
    RECT 190.32 59.47 190.53 59.54 ;
    RECT 190.32 59.83 190.53 59.9 ;
    RECT 189.86 59.11 190.07 59.18 ;
    RECT 189.86 59.47 190.07 59.54 ;
    RECT 189.86 59.83 190.07 59.9 ;
    RECT 187.0 59.11 187.21 59.18 ;
    RECT 187.0 59.47 187.21 59.54 ;
    RECT 187.0 59.83 187.21 59.9 ;
    RECT 186.54 59.11 186.75 59.18 ;
    RECT 186.54 59.47 186.75 59.54 ;
    RECT 186.54 59.83 186.75 59.9 ;
    RECT 183.68 59.11 183.89 59.18 ;
    RECT 183.68 59.47 183.89 59.54 ;
    RECT 183.68 59.83 183.89 59.9 ;
    RECT 183.22 59.11 183.43 59.18 ;
    RECT 183.22 59.47 183.43 59.54 ;
    RECT 183.22 59.83 183.43 59.9 ;
    RECT 147.485 59.47 147.555 59.54 ;
    RECT 266.68 59.11 266.89 59.18 ;
    RECT 266.68 59.47 266.89 59.54 ;
    RECT 266.68 59.83 266.89 59.9 ;
    RECT 266.22 59.11 266.43 59.18 ;
    RECT 266.22 59.47 266.43 59.54 ;
    RECT 266.22 59.83 266.43 59.9 ;
    RECT 263.36 59.11 263.57 59.18 ;
    RECT 263.36 59.47 263.57 59.54 ;
    RECT 263.36 59.83 263.57 59.9 ;
    RECT 262.9 59.11 263.11 59.18 ;
    RECT 262.9 59.47 263.11 59.54 ;
    RECT 262.9 59.83 263.11 59.9 ;
    RECT 260.04 59.11 260.25 59.18 ;
    RECT 260.04 59.47 260.25 59.54 ;
    RECT 260.04 59.83 260.25 59.9 ;
    RECT 259.58 59.11 259.79 59.18 ;
    RECT 259.58 59.47 259.79 59.54 ;
    RECT 259.58 59.83 259.79 59.9 ;
    RECT 256.72 59.11 256.93 59.18 ;
    RECT 256.72 59.47 256.93 59.54 ;
    RECT 256.72 59.83 256.93 59.9 ;
    RECT 256.26 59.11 256.47 59.18 ;
    RECT 256.26 59.47 256.47 59.54 ;
    RECT 256.26 59.83 256.47 59.9 ;
    RECT 253.4 59.11 253.61 59.18 ;
    RECT 253.4 59.47 253.61 59.54 ;
    RECT 253.4 59.83 253.61 59.9 ;
    RECT 252.94 59.11 253.15 59.18 ;
    RECT 252.94 59.47 253.15 59.54 ;
    RECT 252.94 59.83 253.15 59.9 ;
    RECT 250.08 95.13 250.29 95.2 ;
    RECT 250.08 95.49 250.29 95.56 ;
    RECT 250.08 95.85 250.29 95.92 ;
    RECT 249.62 95.13 249.83 95.2 ;
    RECT 249.62 95.49 249.83 95.56 ;
    RECT 249.62 95.85 249.83 95.92 ;
    RECT 246.76 95.13 246.97 95.2 ;
    RECT 246.76 95.49 246.97 95.56 ;
    RECT 246.76 95.85 246.97 95.92 ;
    RECT 246.3 95.13 246.51 95.2 ;
    RECT 246.3 95.49 246.51 95.56 ;
    RECT 246.3 95.85 246.51 95.92 ;
    RECT 243.44 95.13 243.65 95.2 ;
    RECT 243.44 95.49 243.65 95.56 ;
    RECT 243.44 95.85 243.65 95.92 ;
    RECT 242.98 95.13 243.19 95.2 ;
    RECT 242.98 95.49 243.19 95.56 ;
    RECT 242.98 95.85 243.19 95.92 ;
    RECT 240.12 95.13 240.33 95.2 ;
    RECT 240.12 95.49 240.33 95.56 ;
    RECT 240.12 95.85 240.33 95.92 ;
    RECT 239.66 95.13 239.87 95.2 ;
    RECT 239.66 95.49 239.87 95.56 ;
    RECT 239.66 95.85 239.87 95.92 ;
    RECT 236.8 95.13 237.01 95.2 ;
    RECT 236.8 95.49 237.01 95.56 ;
    RECT 236.8 95.85 237.01 95.92 ;
    RECT 236.34 95.13 236.55 95.2 ;
    RECT 236.34 95.49 236.55 95.56 ;
    RECT 236.34 95.85 236.55 95.92 ;
    RECT 233.48 95.13 233.69 95.2 ;
    RECT 233.48 95.49 233.69 95.56 ;
    RECT 233.48 95.85 233.69 95.92 ;
    RECT 233.02 95.13 233.23 95.2 ;
    RECT 233.02 95.49 233.23 95.56 ;
    RECT 233.02 95.85 233.23 95.92 ;
    RECT 230.16 95.13 230.37 95.2 ;
    RECT 230.16 95.49 230.37 95.56 ;
    RECT 230.16 95.85 230.37 95.92 ;
    RECT 229.7 95.13 229.91 95.2 ;
    RECT 229.7 95.49 229.91 95.56 ;
    RECT 229.7 95.85 229.91 95.92 ;
    RECT 226.84 95.13 227.05 95.2 ;
    RECT 226.84 95.49 227.05 95.56 ;
    RECT 226.84 95.85 227.05 95.92 ;
    RECT 226.38 95.13 226.59 95.2 ;
    RECT 226.38 95.49 226.59 95.56 ;
    RECT 226.38 95.85 226.59 95.92 ;
    RECT 223.52 95.13 223.73 95.2 ;
    RECT 223.52 95.49 223.73 95.56 ;
    RECT 223.52 95.85 223.73 95.92 ;
    RECT 223.06 95.13 223.27 95.2 ;
    RECT 223.06 95.49 223.27 95.56 ;
    RECT 223.06 95.85 223.27 95.92 ;
    RECT 220.2 95.13 220.41 95.2 ;
    RECT 220.2 95.49 220.41 95.56 ;
    RECT 220.2 95.85 220.41 95.92 ;
    RECT 219.74 95.13 219.95 95.2 ;
    RECT 219.74 95.49 219.95 95.56 ;
    RECT 219.74 95.85 219.95 95.92 ;
    RECT 216.88 95.13 217.09 95.2 ;
    RECT 216.88 95.49 217.09 95.56 ;
    RECT 216.88 95.85 217.09 95.92 ;
    RECT 216.42 95.13 216.63 95.2 ;
    RECT 216.42 95.49 216.63 95.56 ;
    RECT 216.42 95.85 216.63 95.92 ;
    RECT 267.91 95.49 267.98 95.56 ;
    RECT 180.36 95.13 180.57 95.2 ;
    RECT 180.36 95.49 180.57 95.56 ;
    RECT 180.36 95.85 180.57 95.92 ;
    RECT 179.9 95.13 180.11 95.2 ;
    RECT 179.9 95.49 180.11 95.56 ;
    RECT 179.9 95.85 180.11 95.92 ;
    RECT 177.04 95.13 177.25 95.2 ;
    RECT 177.04 95.49 177.25 95.56 ;
    RECT 177.04 95.85 177.25 95.92 ;
    RECT 176.58 95.13 176.79 95.2 ;
    RECT 176.58 95.49 176.79 95.56 ;
    RECT 176.58 95.85 176.79 95.92 ;
    RECT 173.72 95.13 173.93 95.2 ;
    RECT 173.72 95.49 173.93 95.56 ;
    RECT 173.72 95.85 173.93 95.92 ;
    RECT 173.26 95.13 173.47 95.2 ;
    RECT 173.26 95.49 173.47 95.56 ;
    RECT 173.26 95.85 173.47 95.92 ;
    RECT 170.4 95.13 170.61 95.2 ;
    RECT 170.4 95.49 170.61 95.56 ;
    RECT 170.4 95.85 170.61 95.92 ;
    RECT 169.94 95.13 170.15 95.2 ;
    RECT 169.94 95.49 170.15 95.56 ;
    RECT 169.94 95.85 170.15 95.92 ;
    RECT 167.08 95.13 167.29 95.2 ;
    RECT 167.08 95.49 167.29 95.56 ;
    RECT 167.08 95.85 167.29 95.92 ;
    RECT 166.62 95.13 166.83 95.2 ;
    RECT 166.62 95.49 166.83 95.56 ;
    RECT 166.62 95.85 166.83 95.92 ;
    RECT 163.76 95.13 163.97 95.2 ;
    RECT 163.76 95.49 163.97 95.56 ;
    RECT 163.76 95.85 163.97 95.92 ;
    RECT 163.3 95.13 163.51 95.2 ;
    RECT 163.3 95.49 163.51 95.56 ;
    RECT 163.3 95.85 163.51 95.92 ;
    RECT 160.44 95.13 160.65 95.2 ;
    RECT 160.44 95.49 160.65 95.56 ;
    RECT 160.44 95.85 160.65 95.92 ;
    RECT 159.98 95.13 160.19 95.2 ;
    RECT 159.98 95.49 160.19 95.56 ;
    RECT 159.98 95.85 160.19 95.92 ;
    RECT 157.12 95.13 157.33 95.2 ;
    RECT 157.12 95.49 157.33 95.56 ;
    RECT 157.12 95.85 157.33 95.92 ;
    RECT 156.66 95.13 156.87 95.2 ;
    RECT 156.66 95.49 156.87 95.56 ;
    RECT 156.66 95.85 156.87 95.92 ;
    RECT 153.8 95.13 154.01 95.2 ;
    RECT 153.8 95.49 154.01 95.56 ;
    RECT 153.8 95.85 154.01 95.92 ;
    RECT 153.34 95.13 153.55 95.2 ;
    RECT 153.34 95.49 153.55 95.56 ;
    RECT 153.34 95.85 153.55 95.92 ;
    RECT 150.48 95.13 150.69 95.2 ;
    RECT 150.48 95.49 150.69 95.56 ;
    RECT 150.48 95.85 150.69 95.92 ;
    RECT 150.02 95.13 150.23 95.2 ;
    RECT 150.02 95.49 150.23 95.56 ;
    RECT 150.02 95.85 150.23 95.92 ;
    RECT 213.56 95.13 213.77 95.2 ;
    RECT 213.56 95.49 213.77 95.56 ;
    RECT 213.56 95.85 213.77 95.92 ;
    RECT 213.1 95.13 213.31 95.2 ;
    RECT 213.1 95.49 213.31 95.56 ;
    RECT 213.1 95.85 213.31 95.92 ;
    RECT 210.24 95.13 210.45 95.2 ;
    RECT 210.24 95.49 210.45 95.56 ;
    RECT 210.24 95.85 210.45 95.92 ;
    RECT 209.78 95.13 209.99 95.2 ;
    RECT 209.78 95.49 209.99 95.56 ;
    RECT 209.78 95.85 209.99 95.92 ;
    RECT 206.92 95.13 207.13 95.2 ;
    RECT 206.92 95.49 207.13 95.56 ;
    RECT 206.92 95.85 207.13 95.92 ;
    RECT 206.46 95.13 206.67 95.2 ;
    RECT 206.46 95.49 206.67 95.56 ;
    RECT 206.46 95.85 206.67 95.92 ;
    RECT 203.6 95.13 203.81 95.2 ;
    RECT 203.6 95.49 203.81 95.56 ;
    RECT 203.6 95.85 203.81 95.92 ;
    RECT 203.14 95.13 203.35 95.2 ;
    RECT 203.14 95.49 203.35 95.56 ;
    RECT 203.14 95.85 203.35 95.92 ;
    RECT 200.28 95.13 200.49 95.2 ;
    RECT 200.28 95.49 200.49 95.56 ;
    RECT 200.28 95.85 200.49 95.92 ;
    RECT 199.82 95.13 200.03 95.2 ;
    RECT 199.82 95.49 200.03 95.56 ;
    RECT 199.82 95.85 200.03 95.92 ;
    RECT 196.96 95.13 197.17 95.2 ;
    RECT 196.96 95.49 197.17 95.56 ;
    RECT 196.96 95.85 197.17 95.92 ;
    RECT 196.5 95.13 196.71 95.2 ;
    RECT 196.5 95.49 196.71 95.56 ;
    RECT 196.5 95.85 196.71 95.92 ;
    RECT 193.64 95.13 193.85 95.2 ;
    RECT 193.64 95.49 193.85 95.56 ;
    RECT 193.64 95.85 193.85 95.92 ;
    RECT 193.18 95.13 193.39 95.2 ;
    RECT 193.18 95.49 193.39 95.56 ;
    RECT 193.18 95.85 193.39 95.92 ;
    RECT 190.32 95.13 190.53 95.2 ;
    RECT 190.32 95.49 190.53 95.56 ;
    RECT 190.32 95.85 190.53 95.92 ;
    RECT 189.86 95.13 190.07 95.2 ;
    RECT 189.86 95.49 190.07 95.56 ;
    RECT 189.86 95.85 190.07 95.92 ;
    RECT 187.0 95.13 187.21 95.2 ;
    RECT 187.0 95.49 187.21 95.56 ;
    RECT 187.0 95.85 187.21 95.92 ;
    RECT 186.54 95.13 186.75 95.2 ;
    RECT 186.54 95.49 186.75 95.56 ;
    RECT 186.54 95.85 186.75 95.92 ;
    RECT 183.68 95.13 183.89 95.2 ;
    RECT 183.68 95.49 183.89 95.56 ;
    RECT 183.68 95.85 183.89 95.92 ;
    RECT 183.22 95.13 183.43 95.2 ;
    RECT 183.22 95.49 183.43 95.56 ;
    RECT 183.22 95.85 183.43 95.92 ;
    RECT 147.485 95.49 147.555 95.56 ;
    RECT 266.68 95.13 266.89 95.2 ;
    RECT 266.68 95.49 266.89 95.56 ;
    RECT 266.68 95.85 266.89 95.92 ;
    RECT 266.22 95.13 266.43 95.2 ;
    RECT 266.22 95.49 266.43 95.56 ;
    RECT 266.22 95.85 266.43 95.92 ;
    RECT 263.36 95.13 263.57 95.2 ;
    RECT 263.36 95.49 263.57 95.56 ;
    RECT 263.36 95.85 263.57 95.92 ;
    RECT 262.9 95.13 263.11 95.2 ;
    RECT 262.9 95.49 263.11 95.56 ;
    RECT 262.9 95.85 263.11 95.92 ;
    RECT 260.04 95.13 260.25 95.2 ;
    RECT 260.04 95.49 260.25 95.56 ;
    RECT 260.04 95.85 260.25 95.92 ;
    RECT 259.58 95.13 259.79 95.2 ;
    RECT 259.58 95.49 259.79 95.56 ;
    RECT 259.58 95.85 259.79 95.92 ;
    RECT 256.72 95.13 256.93 95.2 ;
    RECT 256.72 95.49 256.93 95.56 ;
    RECT 256.72 95.85 256.93 95.92 ;
    RECT 256.26 95.13 256.47 95.2 ;
    RECT 256.26 95.49 256.47 95.56 ;
    RECT 256.26 95.85 256.47 95.92 ;
    RECT 253.4 95.13 253.61 95.2 ;
    RECT 253.4 95.49 253.61 95.56 ;
    RECT 253.4 95.85 253.61 95.92 ;
    RECT 252.94 95.13 253.15 95.2 ;
    RECT 252.94 95.49 253.15 95.56 ;
    RECT 252.94 95.85 253.15 95.92 ;
    RECT 250.08 58.39 250.29 58.46 ;
    RECT 250.08 58.75 250.29 58.82 ;
    RECT 250.08 59.11 250.29 59.18 ;
    RECT 249.62 58.39 249.83 58.46 ;
    RECT 249.62 58.75 249.83 58.82 ;
    RECT 249.62 59.11 249.83 59.18 ;
    RECT 246.76 58.39 246.97 58.46 ;
    RECT 246.76 58.75 246.97 58.82 ;
    RECT 246.76 59.11 246.97 59.18 ;
    RECT 246.3 58.39 246.51 58.46 ;
    RECT 246.3 58.75 246.51 58.82 ;
    RECT 246.3 59.11 246.51 59.18 ;
    RECT 243.44 58.39 243.65 58.46 ;
    RECT 243.44 58.75 243.65 58.82 ;
    RECT 243.44 59.11 243.65 59.18 ;
    RECT 242.98 58.39 243.19 58.46 ;
    RECT 242.98 58.75 243.19 58.82 ;
    RECT 242.98 59.11 243.19 59.18 ;
    RECT 240.12 58.39 240.33 58.46 ;
    RECT 240.12 58.75 240.33 58.82 ;
    RECT 240.12 59.11 240.33 59.18 ;
    RECT 239.66 58.39 239.87 58.46 ;
    RECT 239.66 58.75 239.87 58.82 ;
    RECT 239.66 59.11 239.87 59.18 ;
    RECT 236.8 58.39 237.01 58.46 ;
    RECT 236.8 58.75 237.01 58.82 ;
    RECT 236.8 59.11 237.01 59.18 ;
    RECT 236.34 58.39 236.55 58.46 ;
    RECT 236.34 58.75 236.55 58.82 ;
    RECT 236.34 59.11 236.55 59.18 ;
    RECT 233.48 58.39 233.69 58.46 ;
    RECT 233.48 58.75 233.69 58.82 ;
    RECT 233.48 59.11 233.69 59.18 ;
    RECT 233.02 58.39 233.23 58.46 ;
    RECT 233.02 58.75 233.23 58.82 ;
    RECT 233.02 59.11 233.23 59.18 ;
    RECT 230.16 58.39 230.37 58.46 ;
    RECT 230.16 58.75 230.37 58.82 ;
    RECT 230.16 59.11 230.37 59.18 ;
    RECT 229.7 58.39 229.91 58.46 ;
    RECT 229.7 58.75 229.91 58.82 ;
    RECT 229.7 59.11 229.91 59.18 ;
    RECT 226.84 58.39 227.05 58.46 ;
    RECT 226.84 58.75 227.05 58.82 ;
    RECT 226.84 59.11 227.05 59.18 ;
    RECT 226.38 58.39 226.59 58.46 ;
    RECT 226.38 58.75 226.59 58.82 ;
    RECT 226.38 59.11 226.59 59.18 ;
    RECT 223.52 58.39 223.73 58.46 ;
    RECT 223.52 58.75 223.73 58.82 ;
    RECT 223.52 59.11 223.73 59.18 ;
    RECT 223.06 58.39 223.27 58.46 ;
    RECT 223.06 58.75 223.27 58.82 ;
    RECT 223.06 59.11 223.27 59.18 ;
    RECT 220.2 58.39 220.41 58.46 ;
    RECT 220.2 58.75 220.41 58.82 ;
    RECT 220.2 59.11 220.41 59.18 ;
    RECT 219.74 58.39 219.95 58.46 ;
    RECT 219.74 58.75 219.95 58.82 ;
    RECT 219.74 59.11 219.95 59.18 ;
    RECT 216.88 58.39 217.09 58.46 ;
    RECT 216.88 58.75 217.09 58.82 ;
    RECT 216.88 59.11 217.09 59.18 ;
    RECT 216.42 58.39 216.63 58.46 ;
    RECT 216.42 58.75 216.63 58.82 ;
    RECT 216.42 59.11 216.63 59.18 ;
    RECT 267.91 58.75 267.98 58.82 ;
    RECT 180.36 58.39 180.57 58.46 ;
    RECT 180.36 58.75 180.57 58.82 ;
    RECT 180.36 59.11 180.57 59.18 ;
    RECT 179.9 58.39 180.11 58.46 ;
    RECT 179.9 58.75 180.11 58.82 ;
    RECT 179.9 59.11 180.11 59.18 ;
    RECT 177.04 58.39 177.25 58.46 ;
    RECT 177.04 58.75 177.25 58.82 ;
    RECT 177.04 59.11 177.25 59.18 ;
    RECT 176.58 58.39 176.79 58.46 ;
    RECT 176.58 58.75 176.79 58.82 ;
    RECT 176.58 59.11 176.79 59.18 ;
    RECT 173.72 58.39 173.93 58.46 ;
    RECT 173.72 58.75 173.93 58.82 ;
    RECT 173.72 59.11 173.93 59.18 ;
    RECT 173.26 58.39 173.47 58.46 ;
    RECT 173.26 58.75 173.47 58.82 ;
    RECT 173.26 59.11 173.47 59.18 ;
    RECT 170.4 58.39 170.61 58.46 ;
    RECT 170.4 58.75 170.61 58.82 ;
    RECT 170.4 59.11 170.61 59.18 ;
    RECT 169.94 58.39 170.15 58.46 ;
    RECT 169.94 58.75 170.15 58.82 ;
    RECT 169.94 59.11 170.15 59.18 ;
    RECT 167.08 58.39 167.29 58.46 ;
    RECT 167.08 58.75 167.29 58.82 ;
    RECT 167.08 59.11 167.29 59.18 ;
    RECT 166.62 58.39 166.83 58.46 ;
    RECT 166.62 58.75 166.83 58.82 ;
    RECT 166.62 59.11 166.83 59.18 ;
    RECT 163.76 58.39 163.97 58.46 ;
    RECT 163.76 58.75 163.97 58.82 ;
    RECT 163.76 59.11 163.97 59.18 ;
    RECT 163.3 58.39 163.51 58.46 ;
    RECT 163.3 58.75 163.51 58.82 ;
    RECT 163.3 59.11 163.51 59.18 ;
    RECT 160.44 58.39 160.65 58.46 ;
    RECT 160.44 58.75 160.65 58.82 ;
    RECT 160.44 59.11 160.65 59.18 ;
    RECT 159.98 58.39 160.19 58.46 ;
    RECT 159.98 58.75 160.19 58.82 ;
    RECT 159.98 59.11 160.19 59.18 ;
    RECT 157.12 58.39 157.33 58.46 ;
    RECT 157.12 58.75 157.33 58.82 ;
    RECT 157.12 59.11 157.33 59.18 ;
    RECT 156.66 58.39 156.87 58.46 ;
    RECT 156.66 58.75 156.87 58.82 ;
    RECT 156.66 59.11 156.87 59.18 ;
    RECT 153.8 58.39 154.01 58.46 ;
    RECT 153.8 58.75 154.01 58.82 ;
    RECT 153.8 59.11 154.01 59.18 ;
    RECT 153.34 58.39 153.55 58.46 ;
    RECT 153.34 58.75 153.55 58.82 ;
    RECT 153.34 59.11 153.55 59.18 ;
    RECT 150.48 58.39 150.69 58.46 ;
    RECT 150.48 58.75 150.69 58.82 ;
    RECT 150.48 59.11 150.69 59.18 ;
    RECT 150.02 58.39 150.23 58.46 ;
    RECT 150.02 58.75 150.23 58.82 ;
    RECT 150.02 59.11 150.23 59.18 ;
    RECT 213.56 58.39 213.77 58.46 ;
    RECT 213.56 58.75 213.77 58.82 ;
    RECT 213.56 59.11 213.77 59.18 ;
    RECT 213.1 58.39 213.31 58.46 ;
    RECT 213.1 58.75 213.31 58.82 ;
    RECT 213.1 59.11 213.31 59.18 ;
    RECT 210.24 58.39 210.45 58.46 ;
    RECT 210.24 58.75 210.45 58.82 ;
    RECT 210.24 59.11 210.45 59.18 ;
    RECT 209.78 58.39 209.99 58.46 ;
    RECT 209.78 58.75 209.99 58.82 ;
    RECT 209.78 59.11 209.99 59.18 ;
    RECT 206.92 58.39 207.13 58.46 ;
    RECT 206.92 58.75 207.13 58.82 ;
    RECT 206.92 59.11 207.13 59.18 ;
    RECT 206.46 58.39 206.67 58.46 ;
    RECT 206.46 58.75 206.67 58.82 ;
    RECT 206.46 59.11 206.67 59.18 ;
    RECT 203.6 58.39 203.81 58.46 ;
    RECT 203.6 58.75 203.81 58.82 ;
    RECT 203.6 59.11 203.81 59.18 ;
    RECT 203.14 58.39 203.35 58.46 ;
    RECT 203.14 58.75 203.35 58.82 ;
    RECT 203.14 59.11 203.35 59.18 ;
    RECT 200.28 58.39 200.49 58.46 ;
    RECT 200.28 58.75 200.49 58.82 ;
    RECT 200.28 59.11 200.49 59.18 ;
    RECT 199.82 58.39 200.03 58.46 ;
    RECT 199.82 58.75 200.03 58.82 ;
    RECT 199.82 59.11 200.03 59.18 ;
    RECT 196.96 58.39 197.17 58.46 ;
    RECT 196.96 58.75 197.17 58.82 ;
    RECT 196.96 59.11 197.17 59.18 ;
    RECT 196.5 58.39 196.71 58.46 ;
    RECT 196.5 58.75 196.71 58.82 ;
    RECT 196.5 59.11 196.71 59.18 ;
    RECT 193.64 58.39 193.85 58.46 ;
    RECT 193.64 58.75 193.85 58.82 ;
    RECT 193.64 59.11 193.85 59.18 ;
    RECT 193.18 58.39 193.39 58.46 ;
    RECT 193.18 58.75 193.39 58.82 ;
    RECT 193.18 59.11 193.39 59.18 ;
    RECT 190.32 58.39 190.53 58.46 ;
    RECT 190.32 58.75 190.53 58.82 ;
    RECT 190.32 59.11 190.53 59.18 ;
    RECT 189.86 58.39 190.07 58.46 ;
    RECT 189.86 58.75 190.07 58.82 ;
    RECT 189.86 59.11 190.07 59.18 ;
    RECT 187.0 58.39 187.21 58.46 ;
    RECT 187.0 58.75 187.21 58.82 ;
    RECT 187.0 59.11 187.21 59.18 ;
    RECT 186.54 58.39 186.75 58.46 ;
    RECT 186.54 58.75 186.75 58.82 ;
    RECT 186.54 59.11 186.75 59.18 ;
    RECT 183.68 58.39 183.89 58.46 ;
    RECT 183.68 58.75 183.89 58.82 ;
    RECT 183.68 59.11 183.89 59.18 ;
    RECT 183.22 58.39 183.43 58.46 ;
    RECT 183.22 58.75 183.43 58.82 ;
    RECT 183.22 59.11 183.43 59.18 ;
    RECT 147.485 58.75 147.555 58.82 ;
    RECT 266.68 58.39 266.89 58.46 ;
    RECT 266.68 58.75 266.89 58.82 ;
    RECT 266.68 59.11 266.89 59.18 ;
    RECT 266.22 58.39 266.43 58.46 ;
    RECT 266.22 58.75 266.43 58.82 ;
    RECT 266.22 59.11 266.43 59.18 ;
    RECT 263.36 58.39 263.57 58.46 ;
    RECT 263.36 58.75 263.57 58.82 ;
    RECT 263.36 59.11 263.57 59.18 ;
    RECT 262.9 58.39 263.11 58.46 ;
    RECT 262.9 58.75 263.11 58.82 ;
    RECT 262.9 59.11 263.11 59.18 ;
    RECT 260.04 58.39 260.25 58.46 ;
    RECT 260.04 58.75 260.25 58.82 ;
    RECT 260.04 59.11 260.25 59.18 ;
    RECT 259.58 58.39 259.79 58.46 ;
    RECT 259.58 58.75 259.79 58.82 ;
    RECT 259.58 59.11 259.79 59.18 ;
    RECT 256.72 58.39 256.93 58.46 ;
    RECT 256.72 58.75 256.93 58.82 ;
    RECT 256.72 59.11 256.93 59.18 ;
    RECT 256.26 58.39 256.47 58.46 ;
    RECT 256.26 58.75 256.47 58.82 ;
    RECT 256.26 59.11 256.47 59.18 ;
    RECT 253.4 58.39 253.61 58.46 ;
    RECT 253.4 58.75 253.61 58.82 ;
    RECT 253.4 59.11 253.61 59.18 ;
    RECT 252.94 58.39 253.15 58.46 ;
    RECT 252.94 58.75 253.15 58.82 ;
    RECT 252.94 59.11 253.15 59.18 ;
    RECT 250.08 94.41 250.29 94.48 ;
    RECT 250.08 94.77 250.29 94.84 ;
    RECT 250.08 95.13 250.29 95.2 ;
    RECT 249.62 94.41 249.83 94.48 ;
    RECT 249.62 94.77 249.83 94.84 ;
    RECT 249.62 95.13 249.83 95.2 ;
    RECT 246.76 94.41 246.97 94.48 ;
    RECT 246.76 94.77 246.97 94.84 ;
    RECT 246.76 95.13 246.97 95.2 ;
    RECT 246.3 94.41 246.51 94.48 ;
    RECT 246.3 94.77 246.51 94.84 ;
    RECT 246.3 95.13 246.51 95.2 ;
    RECT 243.44 94.41 243.65 94.48 ;
    RECT 243.44 94.77 243.65 94.84 ;
    RECT 243.44 95.13 243.65 95.2 ;
    RECT 242.98 94.41 243.19 94.48 ;
    RECT 242.98 94.77 243.19 94.84 ;
    RECT 242.98 95.13 243.19 95.2 ;
    RECT 240.12 94.41 240.33 94.48 ;
    RECT 240.12 94.77 240.33 94.84 ;
    RECT 240.12 95.13 240.33 95.2 ;
    RECT 239.66 94.41 239.87 94.48 ;
    RECT 239.66 94.77 239.87 94.84 ;
    RECT 239.66 95.13 239.87 95.2 ;
    RECT 236.8 94.41 237.01 94.48 ;
    RECT 236.8 94.77 237.01 94.84 ;
    RECT 236.8 95.13 237.01 95.2 ;
    RECT 236.34 94.41 236.55 94.48 ;
    RECT 236.34 94.77 236.55 94.84 ;
    RECT 236.34 95.13 236.55 95.2 ;
    RECT 233.48 94.41 233.69 94.48 ;
    RECT 233.48 94.77 233.69 94.84 ;
    RECT 233.48 95.13 233.69 95.2 ;
    RECT 233.02 94.41 233.23 94.48 ;
    RECT 233.02 94.77 233.23 94.84 ;
    RECT 233.02 95.13 233.23 95.2 ;
    RECT 230.16 94.41 230.37 94.48 ;
    RECT 230.16 94.77 230.37 94.84 ;
    RECT 230.16 95.13 230.37 95.2 ;
    RECT 229.7 94.41 229.91 94.48 ;
    RECT 229.7 94.77 229.91 94.84 ;
    RECT 229.7 95.13 229.91 95.2 ;
    RECT 226.84 94.41 227.05 94.48 ;
    RECT 226.84 94.77 227.05 94.84 ;
    RECT 226.84 95.13 227.05 95.2 ;
    RECT 226.38 94.41 226.59 94.48 ;
    RECT 226.38 94.77 226.59 94.84 ;
    RECT 226.38 95.13 226.59 95.2 ;
    RECT 223.52 94.41 223.73 94.48 ;
    RECT 223.52 94.77 223.73 94.84 ;
    RECT 223.52 95.13 223.73 95.2 ;
    RECT 223.06 94.41 223.27 94.48 ;
    RECT 223.06 94.77 223.27 94.84 ;
    RECT 223.06 95.13 223.27 95.2 ;
    RECT 220.2 94.41 220.41 94.48 ;
    RECT 220.2 94.77 220.41 94.84 ;
    RECT 220.2 95.13 220.41 95.2 ;
    RECT 219.74 94.41 219.95 94.48 ;
    RECT 219.74 94.77 219.95 94.84 ;
    RECT 219.74 95.13 219.95 95.2 ;
    RECT 216.88 94.41 217.09 94.48 ;
    RECT 216.88 94.77 217.09 94.84 ;
    RECT 216.88 95.13 217.09 95.2 ;
    RECT 216.42 94.41 216.63 94.48 ;
    RECT 216.42 94.77 216.63 94.84 ;
    RECT 216.42 95.13 216.63 95.2 ;
    RECT 267.91 94.77 267.98 94.84 ;
    RECT 180.36 94.41 180.57 94.48 ;
    RECT 180.36 94.77 180.57 94.84 ;
    RECT 180.36 95.13 180.57 95.2 ;
    RECT 179.9 94.41 180.11 94.48 ;
    RECT 179.9 94.77 180.11 94.84 ;
    RECT 179.9 95.13 180.11 95.2 ;
    RECT 177.04 94.41 177.25 94.48 ;
    RECT 177.04 94.77 177.25 94.84 ;
    RECT 177.04 95.13 177.25 95.2 ;
    RECT 176.58 94.41 176.79 94.48 ;
    RECT 176.58 94.77 176.79 94.84 ;
    RECT 176.58 95.13 176.79 95.2 ;
    RECT 173.72 94.41 173.93 94.48 ;
    RECT 173.72 94.77 173.93 94.84 ;
    RECT 173.72 95.13 173.93 95.2 ;
    RECT 173.26 94.41 173.47 94.48 ;
    RECT 173.26 94.77 173.47 94.84 ;
    RECT 173.26 95.13 173.47 95.2 ;
    RECT 170.4 94.41 170.61 94.48 ;
    RECT 170.4 94.77 170.61 94.84 ;
    RECT 170.4 95.13 170.61 95.2 ;
    RECT 169.94 94.41 170.15 94.48 ;
    RECT 169.94 94.77 170.15 94.84 ;
    RECT 169.94 95.13 170.15 95.2 ;
    RECT 167.08 94.41 167.29 94.48 ;
    RECT 167.08 94.77 167.29 94.84 ;
    RECT 167.08 95.13 167.29 95.2 ;
    RECT 166.62 94.41 166.83 94.48 ;
    RECT 166.62 94.77 166.83 94.84 ;
    RECT 166.62 95.13 166.83 95.2 ;
    RECT 163.76 94.41 163.97 94.48 ;
    RECT 163.76 94.77 163.97 94.84 ;
    RECT 163.76 95.13 163.97 95.2 ;
    RECT 163.3 94.41 163.51 94.48 ;
    RECT 163.3 94.77 163.51 94.84 ;
    RECT 163.3 95.13 163.51 95.2 ;
    RECT 160.44 94.41 160.65 94.48 ;
    RECT 160.44 94.77 160.65 94.84 ;
    RECT 160.44 95.13 160.65 95.2 ;
    RECT 159.98 94.41 160.19 94.48 ;
    RECT 159.98 94.77 160.19 94.84 ;
    RECT 159.98 95.13 160.19 95.2 ;
    RECT 157.12 94.41 157.33 94.48 ;
    RECT 157.12 94.77 157.33 94.84 ;
    RECT 157.12 95.13 157.33 95.2 ;
    RECT 156.66 94.41 156.87 94.48 ;
    RECT 156.66 94.77 156.87 94.84 ;
    RECT 156.66 95.13 156.87 95.2 ;
    RECT 153.8 94.41 154.01 94.48 ;
    RECT 153.8 94.77 154.01 94.84 ;
    RECT 153.8 95.13 154.01 95.2 ;
    RECT 153.34 94.41 153.55 94.48 ;
    RECT 153.34 94.77 153.55 94.84 ;
    RECT 153.34 95.13 153.55 95.2 ;
    RECT 150.48 94.41 150.69 94.48 ;
    RECT 150.48 94.77 150.69 94.84 ;
    RECT 150.48 95.13 150.69 95.2 ;
    RECT 150.02 94.41 150.23 94.48 ;
    RECT 150.02 94.77 150.23 94.84 ;
    RECT 150.02 95.13 150.23 95.2 ;
    RECT 213.56 94.41 213.77 94.48 ;
    RECT 213.56 94.77 213.77 94.84 ;
    RECT 213.56 95.13 213.77 95.2 ;
    RECT 213.1 94.41 213.31 94.48 ;
    RECT 213.1 94.77 213.31 94.84 ;
    RECT 213.1 95.13 213.31 95.2 ;
    RECT 210.24 94.41 210.45 94.48 ;
    RECT 210.24 94.77 210.45 94.84 ;
    RECT 210.24 95.13 210.45 95.2 ;
    RECT 209.78 94.41 209.99 94.48 ;
    RECT 209.78 94.77 209.99 94.84 ;
    RECT 209.78 95.13 209.99 95.2 ;
    RECT 206.92 94.41 207.13 94.48 ;
    RECT 206.92 94.77 207.13 94.84 ;
    RECT 206.92 95.13 207.13 95.2 ;
    RECT 206.46 94.41 206.67 94.48 ;
    RECT 206.46 94.77 206.67 94.84 ;
    RECT 206.46 95.13 206.67 95.2 ;
    RECT 203.6 94.41 203.81 94.48 ;
    RECT 203.6 94.77 203.81 94.84 ;
    RECT 203.6 95.13 203.81 95.2 ;
    RECT 203.14 94.41 203.35 94.48 ;
    RECT 203.14 94.77 203.35 94.84 ;
    RECT 203.14 95.13 203.35 95.2 ;
    RECT 200.28 94.41 200.49 94.48 ;
    RECT 200.28 94.77 200.49 94.84 ;
    RECT 200.28 95.13 200.49 95.2 ;
    RECT 199.82 94.41 200.03 94.48 ;
    RECT 199.82 94.77 200.03 94.84 ;
    RECT 199.82 95.13 200.03 95.2 ;
    RECT 196.96 94.41 197.17 94.48 ;
    RECT 196.96 94.77 197.17 94.84 ;
    RECT 196.96 95.13 197.17 95.2 ;
    RECT 196.5 94.41 196.71 94.48 ;
    RECT 196.5 94.77 196.71 94.84 ;
    RECT 196.5 95.13 196.71 95.2 ;
    RECT 193.64 94.41 193.85 94.48 ;
    RECT 193.64 94.77 193.85 94.84 ;
    RECT 193.64 95.13 193.85 95.2 ;
    RECT 193.18 94.41 193.39 94.48 ;
    RECT 193.18 94.77 193.39 94.84 ;
    RECT 193.18 95.13 193.39 95.2 ;
    RECT 190.32 94.41 190.53 94.48 ;
    RECT 190.32 94.77 190.53 94.84 ;
    RECT 190.32 95.13 190.53 95.2 ;
    RECT 189.86 94.41 190.07 94.48 ;
    RECT 189.86 94.77 190.07 94.84 ;
    RECT 189.86 95.13 190.07 95.2 ;
    RECT 187.0 94.41 187.21 94.48 ;
    RECT 187.0 94.77 187.21 94.84 ;
    RECT 187.0 95.13 187.21 95.2 ;
    RECT 186.54 94.41 186.75 94.48 ;
    RECT 186.54 94.77 186.75 94.84 ;
    RECT 186.54 95.13 186.75 95.2 ;
    RECT 183.68 94.41 183.89 94.48 ;
    RECT 183.68 94.77 183.89 94.84 ;
    RECT 183.68 95.13 183.89 95.2 ;
    RECT 183.22 94.41 183.43 94.48 ;
    RECT 183.22 94.77 183.43 94.84 ;
    RECT 183.22 95.13 183.43 95.2 ;
    RECT 147.485 94.77 147.555 94.84 ;
    RECT 266.68 94.41 266.89 94.48 ;
    RECT 266.68 94.77 266.89 94.84 ;
    RECT 266.68 95.13 266.89 95.2 ;
    RECT 266.22 94.41 266.43 94.48 ;
    RECT 266.22 94.77 266.43 94.84 ;
    RECT 266.22 95.13 266.43 95.2 ;
    RECT 263.36 94.41 263.57 94.48 ;
    RECT 263.36 94.77 263.57 94.84 ;
    RECT 263.36 95.13 263.57 95.2 ;
    RECT 262.9 94.41 263.11 94.48 ;
    RECT 262.9 94.77 263.11 94.84 ;
    RECT 262.9 95.13 263.11 95.2 ;
    RECT 260.04 94.41 260.25 94.48 ;
    RECT 260.04 94.77 260.25 94.84 ;
    RECT 260.04 95.13 260.25 95.2 ;
    RECT 259.58 94.41 259.79 94.48 ;
    RECT 259.58 94.77 259.79 94.84 ;
    RECT 259.58 95.13 259.79 95.2 ;
    RECT 256.72 94.41 256.93 94.48 ;
    RECT 256.72 94.77 256.93 94.84 ;
    RECT 256.72 95.13 256.93 95.2 ;
    RECT 256.26 94.41 256.47 94.48 ;
    RECT 256.26 94.77 256.47 94.84 ;
    RECT 256.26 95.13 256.47 95.2 ;
    RECT 253.4 94.41 253.61 94.48 ;
    RECT 253.4 94.77 253.61 94.84 ;
    RECT 253.4 95.13 253.61 95.2 ;
    RECT 252.94 94.41 253.15 94.48 ;
    RECT 252.94 94.77 253.15 94.84 ;
    RECT 252.94 95.13 253.15 95.2 ;
    RECT 250.08 57.67 250.29 57.74 ;
    RECT 250.08 58.03 250.29 58.1 ;
    RECT 250.08 58.39 250.29 58.46 ;
    RECT 249.62 57.67 249.83 57.74 ;
    RECT 249.62 58.03 249.83 58.1 ;
    RECT 249.62 58.39 249.83 58.46 ;
    RECT 246.76 57.67 246.97 57.74 ;
    RECT 246.76 58.03 246.97 58.1 ;
    RECT 246.76 58.39 246.97 58.46 ;
    RECT 246.3 57.67 246.51 57.74 ;
    RECT 246.3 58.03 246.51 58.1 ;
    RECT 246.3 58.39 246.51 58.46 ;
    RECT 243.44 57.67 243.65 57.74 ;
    RECT 243.44 58.03 243.65 58.1 ;
    RECT 243.44 58.39 243.65 58.46 ;
    RECT 242.98 57.67 243.19 57.74 ;
    RECT 242.98 58.03 243.19 58.1 ;
    RECT 242.98 58.39 243.19 58.46 ;
    RECT 240.12 57.67 240.33 57.74 ;
    RECT 240.12 58.03 240.33 58.1 ;
    RECT 240.12 58.39 240.33 58.46 ;
    RECT 239.66 57.67 239.87 57.74 ;
    RECT 239.66 58.03 239.87 58.1 ;
    RECT 239.66 58.39 239.87 58.46 ;
    RECT 236.8 57.67 237.01 57.74 ;
    RECT 236.8 58.03 237.01 58.1 ;
    RECT 236.8 58.39 237.01 58.46 ;
    RECT 236.34 57.67 236.55 57.74 ;
    RECT 236.34 58.03 236.55 58.1 ;
    RECT 236.34 58.39 236.55 58.46 ;
    RECT 233.48 57.67 233.69 57.74 ;
    RECT 233.48 58.03 233.69 58.1 ;
    RECT 233.48 58.39 233.69 58.46 ;
    RECT 233.02 57.67 233.23 57.74 ;
    RECT 233.02 58.03 233.23 58.1 ;
    RECT 233.02 58.39 233.23 58.46 ;
    RECT 230.16 57.67 230.37 57.74 ;
    RECT 230.16 58.03 230.37 58.1 ;
    RECT 230.16 58.39 230.37 58.46 ;
    RECT 229.7 57.67 229.91 57.74 ;
    RECT 229.7 58.03 229.91 58.1 ;
    RECT 229.7 58.39 229.91 58.46 ;
    RECT 226.84 57.67 227.05 57.74 ;
    RECT 226.84 58.03 227.05 58.1 ;
    RECT 226.84 58.39 227.05 58.46 ;
    RECT 226.38 57.67 226.59 57.74 ;
    RECT 226.38 58.03 226.59 58.1 ;
    RECT 226.38 58.39 226.59 58.46 ;
    RECT 223.52 57.67 223.73 57.74 ;
    RECT 223.52 58.03 223.73 58.1 ;
    RECT 223.52 58.39 223.73 58.46 ;
    RECT 223.06 57.67 223.27 57.74 ;
    RECT 223.06 58.03 223.27 58.1 ;
    RECT 223.06 58.39 223.27 58.46 ;
    RECT 220.2 57.67 220.41 57.74 ;
    RECT 220.2 58.03 220.41 58.1 ;
    RECT 220.2 58.39 220.41 58.46 ;
    RECT 219.74 57.67 219.95 57.74 ;
    RECT 219.74 58.03 219.95 58.1 ;
    RECT 219.74 58.39 219.95 58.46 ;
    RECT 216.88 57.67 217.09 57.74 ;
    RECT 216.88 58.03 217.09 58.1 ;
    RECT 216.88 58.39 217.09 58.46 ;
    RECT 216.42 57.67 216.63 57.74 ;
    RECT 216.42 58.03 216.63 58.1 ;
    RECT 216.42 58.39 216.63 58.46 ;
    RECT 267.91 58.03 267.98 58.1 ;
    RECT 180.36 57.67 180.57 57.74 ;
    RECT 180.36 58.03 180.57 58.1 ;
    RECT 180.36 58.39 180.57 58.46 ;
    RECT 179.9 57.67 180.11 57.74 ;
    RECT 179.9 58.03 180.11 58.1 ;
    RECT 179.9 58.39 180.11 58.46 ;
    RECT 177.04 57.67 177.25 57.74 ;
    RECT 177.04 58.03 177.25 58.1 ;
    RECT 177.04 58.39 177.25 58.46 ;
    RECT 176.58 57.67 176.79 57.74 ;
    RECT 176.58 58.03 176.79 58.1 ;
    RECT 176.58 58.39 176.79 58.46 ;
    RECT 173.72 57.67 173.93 57.74 ;
    RECT 173.72 58.03 173.93 58.1 ;
    RECT 173.72 58.39 173.93 58.46 ;
    RECT 173.26 57.67 173.47 57.74 ;
    RECT 173.26 58.03 173.47 58.1 ;
    RECT 173.26 58.39 173.47 58.46 ;
    RECT 170.4 57.67 170.61 57.74 ;
    RECT 170.4 58.03 170.61 58.1 ;
    RECT 170.4 58.39 170.61 58.46 ;
    RECT 169.94 57.67 170.15 57.74 ;
    RECT 169.94 58.03 170.15 58.1 ;
    RECT 169.94 58.39 170.15 58.46 ;
    RECT 167.08 57.67 167.29 57.74 ;
    RECT 167.08 58.03 167.29 58.1 ;
    RECT 167.08 58.39 167.29 58.46 ;
    RECT 166.62 57.67 166.83 57.74 ;
    RECT 166.62 58.03 166.83 58.1 ;
    RECT 166.62 58.39 166.83 58.46 ;
    RECT 163.76 57.67 163.97 57.74 ;
    RECT 163.76 58.03 163.97 58.1 ;
    RECT 163.76 58.39 163.97 58.46 ;
    RECT 163.3 57.67 163.51 57.74 ;
    RECT 163.3 58.03 163.51 58.1 ;
    RECT 163.3 58.39 163.51 58.46 ;
    RECT 160.44 57.67 160.65 57.74 ;
    RECT 160.44 58.03 160.65 58.1 ;
    RECT 160.44 58.39 160.65 58.46 ;
    RECT 159.98 57.67 160.19 57.74 ;
    RECT 159.98 58.03 160.19 58.1 ;
    RECT 159.98 58.39 160.19 58.46 ;
    RECT 157.12 57.67 157.33 57.74 ;
    RECT 157.12 58.03 157.33 58.1 ;
    RECT 157.12 58.39 157.33 58.46 ;
    RECT 156.66 57.67 156.87 57.74 ;
    RECT 156.66 58.03 156.87 58.1 ;
    RECT 156.66 58.39 156.87 58.46 ;
    RECT 153.8 57.67 154.01 57.74 ;
    RECT 153.8 58.03 154.01 58.1 ;
    RECT 153.8 58.39 154.01 58.46 ;
    RECT 153.34 57.67 153.55 57.74 ;
    RECT 153.34 58.03 153.55 58.1 ;
    RECT 153.34 58.39 153.55 58.46 ;
    RECT 150.48 57.67 150.69 57.74 ;
    RECT 150.48 58.03 150.69 58.1 ;
    RECT 150.48 58.39 150.69 58.46 ;
    RECT 150.02 57.67 150.23 57.74 ;
    RECT 150.02 58.03 150.23 58.1 ;
    RECT 150.02 58.39 150.23 58.46 ;
    RECT 213.56 57.67 213.77 57.74 ;
    RECT 213.56 58.03 213.77 58.1 ;
    RECT 213.56 58.39 213.77 58.46 ;
    RECT 213.1 57.67 213.31 57.74 ;
    RECT 213.1 58.03 213.31 58.1 ;
    RECT 213.1 58.39 213.31 58.46 ;
    RECT 210.24 57.67 210.45 57.74 ;
    RECT 210.24 58.03 210.45 58.1 ;
    RECT 210.24 58.39 210.45 58.46 ;
    RECT 209.78 57.67 209.99 57.74 ;
    RECT 209.78 58.03 209.99 58.1 ;
    RECT 209.78 58.39 209.99 58.46 ;
    RECT 206.92 57.67 207.13 57.74 ;
    RECT 206.92 58.03 207.13 58.1 ;
    RECT 206.92 58.39 207.13 58.46 ;
    RECT 206.46 57.67 206.67 57.74 ;
    RECT 206.46 58.03 206.67 58.1 ;
    RECT 206.46 58.39 206.67 58.46 ;
    RECT 203.6 57.67 203.81 57.74 ;
    RECT 203.6 58.03 203.81 58.1 ;
    RECT 203.6 58.39 203.81 58.46 ;
    RECT 203.14 57.67 203.35 57.74 ;
    RECT 203.14 58.03 203.35 58.1 ;
    RECT 203.14 58.39 203.35 58.46 ;
    RECT 200.28 57.67 200.49 57.74 ;
    RECT 200.28 58.03 200.49 58.1 ;
    RECT 200.28 58.39 200.49 58.46 ;
    RECT 199.82 57.67 200.03 57.74 ;
    RECT 199.82 58.03 200.03 58.1 ;
    RECT 199.82 58.39 200.03 58.46 ;
    RECT 196.96 57.67 197.17 57.74 ;
    RECT 196.96 58.03 197.17 58.1 ;
    RECT 196.96 58.39 197.17 58.46 ;
    RECT 196.5 57.67 196.71 57.74 ;
    RECT 196.5 58.03 196.71 58.1 ;
    RECT 196.5 58.39 196.71 58.46 ;
    RECT 193.64 57.67 193.85 57.74 ;
    RECT 193.64 58.03 193.85 58.1 ;
    RECT 193.64 58.39 193.85 58.46 ;
    RECT 193.18 57.67 193.39 57.74 ;
    RECT 193.18 58.03 193.39 58.1 ;
    RECT 193.18 58.39 193.39 58.46 ;
    RECT 190.32 57.67 190.53 57.74 ;
    RECT 190.32 58.03 190.53 58.1 ;
    RECT 190.32 58.39 190.53 58.46 ;
    RECT 189.86 57.67 190.07 57.74 ;
    RECT 189.86 58.03 190.07 58.1 ;
    RECT 189.86 58.39 190.07 58.46 ;
    RECT 187.0 57.67 187.21 57.74 ;
    RECT 187.0 58.03 187.21 58.1 ;
    RECT 187.0 58.39 187.21 58.46 ;
    RECT 186.54 57.67 186.75 57.74 ;
    RECT 186.54 58.03 186.75 58.1 ;
    RECT 186.54 58.39 186.75 58.46 ;
    RECT 183.68 57.67 183.89 57.74 ;
    RECT 183.68 58.03 183.89 58.1 ;
    RECT 183.68 58.39 183.89 58.46 ;
    RECT 183.22 57.67 183.43 57.74 ;
    RECT 183.22 58.03 183.43 58.1 ;
    RECT 183.22 58.39 183.43 58.46 ;
    RECT 147.485 58.03 147.555 58.1 ;
    RECT 266.68 57.67 266.89 57.74 ;
    RECT 266.68 58.03 266.89 58.1 ;
    RECT 266.68 58.39 266.89 58.46 ;
    RECT 266.22 57.67 266.43 57.74 ;
    RECT 266.22 58.03 266.43 58.1 ;
    RECT 266.22 58.39 266.43 58.46 ;
    RECT 263.36 57.67 263.57 57.74 ;
    RECT 263.36 58.03 263.57 58.1 ;
    RECT 263.36 58.39 263.57 58.46 ;
    RECT 262.9 57.67 263.11 57.74 ;
    RECT 262.9 58.03 263.11 58.1 ;
    RECT 262.9 58.39 263.11 58.46 ;
    RECT 260.04 57.67 260.25 57.74 ;
    RECT 260.04 58.03 260.25 58.1 ;
    RECT 260.04 58.39 260.25 58.46 ;
    RECT 259.58 57.67 259.79 57.74 ;
    RECT 259.58 58.03 259.79 58.1 ;
    RECT 259.58 58.39 259.79 58.46 ;
    RECT 256.72 57.67 256.93 57.74 ;
    RECT 256.72 58.03 256.93 58.1 ;
    RECT 256.72 58.39 256.93 58.46 ;
    RECT 256.26 57.67 256.47 57.74 ;
    RECT 256.26 58.03 256.47 58.1 ;
    RECT 256.26 58.39 256.47 58.46 ;
    RECT 253.4 57.67 253.61 57.74 ;
    RECT 253.4 58.03 253.61 58.1 ;
    RECT 253.4 58.39 253.61 58.46 ;
    RECT 252.94 57.67 253.15 57.74 ;
    RECT 252.94 58.03 253.15 58.1 ;
    RECT 252.94 58.39 253.15 58.46 ;
    RECT 250.08 93.69 250.29 93.76 ;
    RECT 250.08 94.05 250.29 94.12 ;
    RECT 250.08 94.41 250.29 94.48 ;
    RECT 249.62 93.69 249.83 93.76 ;
    RECT 249.62 94.05 249.83 94.12 ;
    RECT 249.62 94.41 249.83 94.48 ;
    RECT 246.76 93.69 246.97 93.76 ;
    RECT 246.76 94.05 246.97 94.12 ;
    RECT 246.76 94.41 246.97 94.48 ;
    RECT 246.3 93.69 246.51 93.76 ;
    RECT 246.3 94.05 246.51 94.12 ;
    RECT 246.3 94.41 246.51 94.48 ;
    RECT 243.44 93.69 243.65 93.76 ;
    RECT 243.44 94.05 243.65 94.12 ;
    RECT 243.44 94.41 243.65 94.48 ;
    RECT 242.98 93.69 243.19 93.76 ;
    RECT 242.98 94.05 243.19 94.12 ;
    RECT 242.98 94.41 243.19 94.48 ;
    RECT 240.12 93.69 240.33 93.76 ;
    RECT 240.12 94.05 240.33 94.12 ;
    RECT 240.12 94.41 240.33 94.48 ;
    RECT 239.66 93.69 239.87 93.76 ;
    RECT 239.66 94.05 239.87 94.12 ;
    RECT 239.66 94.41 239.87 94.48 ;
    RECT 236.8 93.69 237.01 93.76 ;
    RECT 236.8 94.05 237.01 94.12 ;
    RECT 236.8 94.41 237.01 94.48 ;
    RECT 236.34 93.69 236.55 93.76 ;
    RECT 236.34 94.05 236.55 94.12 ;
    RECT 236.34 94.41 236.55 94.48 ;
    RECT 233.48 93.69 233.69 93.76 ;
    RECT 233.48 94.05 233.69 94.12 ;
    RECT 233.48 94.41 233.69 94.48 ;
    RECT 233.02 93.69 233.23 93.76 ;
    RECT 233.02 94.05 233.23 94.12 ;
    RECT 233.02 94.41 233.23 94.48 ;
    RECT 230.16 93.69 230.37 93.76 ;
    RECT 230.16 94.05 230.37 94.12 ;
    RECT 230.16 94.41 230.37 94.48 ;
    RECT 229.7 93.69 229.91 93.76 ;
    RECT 229.7 94.05 229.91 94.12 ;
    RECT 229.7 94.41 229.91 94.48 ;
    RECT 226.84 93.69 227.05 93.76 ;
    RECT 226.84 94.05 227.05 94.12 ;
    RECT 226.84 94.41 227.05 94.48 ;
    RECT 226.38 93.69 226.59 93.76 ;
    RECT 226.38 94.05 226.59 94.12 ;
    RECT 226.38 94.41 226.59 94.48 ;
    RECT 223.52 93.69 223.73 93.76 ;
    RECT 223.52 94.05 223.73 94.12 ;
    RECT 223.52 94.41 223.73 94.48 ;
    RECT 223.06 93.69 223.27 93.76 ;
    RECT 223.06 94.05 223.27 94.12 ;
    RECT 223.06 94.41 223.27 94.48 ;
    RECT 220.2 93.69 220.41 93.76 ;
    RECT 220.2 94.05 220.41 94.12 ;
    RECT 220.2 94.41 220.41 94.48 ;
    RECT 219.74 93.69 219.95 93.76 ;
    RECT 219.74 94.05 219.95 94.12 ;
    RECT 219.74 94.41 219.95 94.48 ;
    RECT 216.88 93.69 217.09 93.76 ;
    RECT 216.88 94.05 217.09 94.12 ;
    RECT 216.88 94.41 217.09 94.48 ;
    RECT 216.42 93.69 216.63 93.76 ;
    RECT 216.42 94.05 216.63 94.12 ;
    RECT 216.42 94.41 216.63 94.48 ;
    RECT 267.91 94.05 267.98 94.12 ;
    RECT 180.36 93.69 180.57 93.76 ;
    RECT 180.36 94.05 180.57 94.12 ;
    RECT 180.36 94.41 180.57 94.48 ;
    RECT 179.9 93.69 180.11 93.76 ;
    RECT 179.9 94.05 180.11 94.12 ;
    RECT 179.9 94.41 180.11 94.48 ;
    RECT 177.04 93.69 177.25 93.76 ;
    RECT 177.04 94.05 177.25 94.12 ;
    RECT 177.04 94.41 177.25 94.48 ;
    RECT 176.58 93.69 176.79 93.76 ;
    RECT 176.58 94.05 176.79 94.12 ;
    RECT 176.58 94.41 176.79 94.48 ;
    RECT 173.72 93.69 173.93 93.76 ;
    RECT 173.72 94.05 173.93 94.12 ;
    RECT 173.72 94.41 173.93 94.48 ;
    RECT 173.26 93.69 173.47 93.76 ;
    RECT 173.26 94.05 173.47 94.12 ;
    RECT 173.26 94.41 173.47 94.48 ;
    RECT 170.4 93.69 170.61 93.76 ;
    RECT 170.4 94.05 170.61 94.12 ;
    RECT 170.4 94.41 170.61 94.48 ;
    RECT 169.94 93.69 170.15 93.76 ;
    RECT 169.94 94.05 170.15 94.12 ;
    RECT 169.94 94.41 170.15 94.48 ;
    RECT 167.08 93.69 167.29 93.76 ;
    RECT 167.08 94.05 167.29 94.12 ;
    RECT 167.08 94.41 167.29 94.48 ;
    RECT 166.62 93.69 166.83 93.76 ;
    RECT 166.62 94.05 166.83 94.12 ;
    RECT 166.62 94.41 166.83 94.48 ;
    RECT 163.76 93.69 163.97 93.76 ;
    RECT 163.76 94.05 163.97 94.12 ;
    RECT 163.76 94.41 163.97 94.48 ;
    RECT 163.3 93.69 163.51 93.76 ;
    RECT 163.3 94.05 163.51 94.12 ;
    RECT 163.3 94.41 163.51 94.48 ;
    RECT 160.44 93.69 160.65 93.76 ;
    RECT 160.44 94.05 160.65 94.12 ;
    RECT 160.44 94.41 160.65 94.48 ;
    RECT 159.98 93.69 160.19 93.76 ;
    RECT 159.98 94.05 160.19 94.12 ;
    RECT 159.98 94.41 160.19 94.48 ;
    RECT 157.12 93.69 157.33 93.76 ;
    RECT 157.12 94.05 157.33 94.12 ;
    RECT 157.12 94.41 157.33 94.48 ;
    RECT 156.66 93.69 156.87 93.76 ;
    RECT 156.66 94.05 156.87 94.12 ;
    RECT 156.66 94.41 156.87 94.48 ;
    RECT 153.8 93.69 154.01 93.76 ;
    RECT 153.8 94.05 154.01 94.12 ;
    RECT 153.8 94.41 154.01 94.48 ;
    RECT 153.34 93.69 153.55 93.76 ;
    RECT 153.34 94.05 153.55 94.12 ;
    RECT 153.34 94.41 153.55 94.48 ;
    RECT 150.48 93.69 150.69 93.76 ;
    RECT 150.48 94.05 150.69 94.12 ;
    RECT 150.48 94.41 150.69 94.48 ;
    RECT 150.02 93.69 150.23 93.76 ;
    RECT 150.02 94.05 150.23 94.12 ;
    RECT 150.02 94.41 150.23 94.48 ;
    RECT 213.56 93.69 213.77 93.76 ;
    RECT 213.56 94.05 213.77 94.12 ;
    RECT 213.56 94.41 213.77 94.48 ;
    RECT 213.1 93.69 213.31 93.76 ;
    RECT 213.1 94.05 213.31 94.12 ;
    RECT 213.1 94.41 213.31 94.48 ;
    RECT 210.24 93.69 210.45 93.76 ;
    RECT 210.24 94.05 210.45 94.12 ;
    RECT 210.24 94.41 210.45 94.48 ;
    RECT 209.78 93.69 209.99 93.76 ;
    RECT 209.78 94.05 209.99 94.12 ;
    RECT 209.78 94.41 209.99 94.48 ;
    RECT 206.92 93.69 207.13 93.76 ;
    RECT 206.92 94.05 207.13 94.12 ;
    RECT 206.92 94.41 207.13 94.48 ;
    RECT 206.46 93.69 206.67 93.76 ;
    RECT 206.46 94.05 206.67 94.12 ;
    RECT 206.46 94.41 206.67 94.48 ;
    RECT 203.6 93.69 203.81 93.76 ;
    RECT 203.6 94.05 203.81 94.12 ;
    RECT 203.6 94.41 203.81 94.48 ;
    RECT 203.14 93.69 203.35 93.76 ;
    RECT 203.14 94.05 203.35 94.12 ;
    RECT 203.14 94.41 203.35 94.48 ;
    RECT 200.28 93.69 200.49 93.76 ;
    RECT 200.28 94.05 200.49 94.12 ;
    RECT 200.28 94.41 200.49 94.48 ;
    RECT 199.82 93.69 200.03 93.76 ;
    RECT 199.82 94.05 200.03 94.12 ;
    RECT 199.82 94.41 200.03 94.48 ;
    RECT 196.96 93.69 197.17 93.76 ;
    RECT 196.96 94.05 197.17 94.12 ;
    RECT 196.96 94.41 197.17 94.48 ;
    RECT 196.5 93.69 196.71 93.76 ;
    RECT 196.5 94.05 196.71 94.12 ;
    RECT 196.5 94.41 196.71 94.48 ;
    RECT 193.64 93.69 193.85 93.76 ;
    RECT 193.64 94.05 193.85 94.12 ;
    RECT 193.64 94.41 193.85 94.48 ;
    RECT 193.18 93.69 193.39 93.76 ;
    RECT 193.18 94.05 193.39 94.12 ;
    RECT 193.18 94.41 193.39 94.48 ;
    RECT 190.32 93.69 190.53 93.76 ;
    RECT 190.32 94.05 190.53 94.12 ;
    RECT 190.32 94.41 190.53 94.48 ;
    RECT 189.86 93.69 190.07 93.76 ;
    RECT 189.86 94.05 190.07 94.12 ;
    RECT 189.86 94.41 190.07 94.48 ;
    RECT 187.0 93.69 187.21 93.76 ;
    RECT 187.0 94.05 187.21 94.12 ;
    RECT 187.0 94.41 187.21 94.48 ;
    RECT 186.54 93.69 186.75 93.76 ;
    RECT 186.54 94.05 186.75 94.12 ;
    RECT 186.54 94.41 186.75 94.48 ;
    RECT 183.68 93.69 183.89 93.76 ;
    RECT 183.68 94.05 183.89 94.12 ;
    RECT 183.68 94.41 183.89 94.48 ;
    RECT 183.22 93.69 183.43 93.76 ;
    RECT 183.22 94.05 183.43 94.12 ;
    RECT 183.22 94.41 183.43 94.48 ;
    RECT 147.485 94.05 147.555 94.12 ;
    RECT 266.68 93.69 266.89 93.76 ;
    RECT 266.68 94.05 266.89 94.12 ;
    RECT 266.68 94.41 266.89 94.48 ;
    RECT 266.22 93.69 266.43 93.76 ;
    RECT 266.22 94.05 266.43 94.12 ;
    RECT 266.22 94.41 266.43 94.48 ;
    RECT 263.36 93.69 263.57 93.76 ;
    RECT 263.36 94.05 263.57 94.12 ;
    RECT 263.36 94.41 263.57 94.48 ;
    RECT 262.9 93.69 263.11 93.76 ;
    RECT 262.9 94.05 263.11 94.12 ;
    RECT 262.9 94.41 263.11 94.48 ;
    RECT 260.04 93.69 260.25 93.76 ;
    RECT 260.04 94.05 260.25 94.12 ;
    RECT 260.04 94.41 260.25 94.48 ;
    RECT 259.58 93.69 259.79 93.76 ;
    RECT 259.58 94.05 259.79 94.12 ;
    RECT 259.58 94.41 259.79 94.48 ;
    RECT 256.72 93.69 256.93 93.76 ;
    RECT 256.72 94.05 256.93 94.12 ;
    RECT 256.72 94.41 256.93 94.48 ;
    RECT 256.26 93.69 256.47 93.76 ;
    RECT 256.26 94.05 256.47 94.12 ;
    RECT 256.26 94.41 256.47 94.48 ;
    RECT 253.4 93.69 253.61 93.76 ;
    RECT 253.4 94.05 253.61 94.12 ;
    RECT 253.4 94.41 253.61 94.48 ;
    RECT 252.94 93.69 253.15 93.76 ;
    RECT 252.94 94.05 253.15 94.12 ;
    RECT 252.94 94.41 253.15 94.48 ;
    RECT 250.08 56.95 250.29 57.02 ;
    RECT 250.08 57.31 250.29 57.38 ;
    RECT 250.08 57.67 250.29 57.74 ;
    RECT 249.62 56.95 249.83 57.02 ;
    RECT 249.62 57.31 249.83 57.38 ;
    RECT 249.62 57.67 249.83 57.74 ;
    RECT 246.76 56.95 246.97 57.02 ;
    RECT 246.76 57.31 246.97 57.38 ;
    RECT 246.76 57.67 246.97 57.74 ;
    RECT 246.3 56.95 246.51 57.02 ;
    RECT 246.3 57.31 246.51 57.38 ;
    RECT 246.3 57.67 246.51 57.74 ;
    RECT 243.44 56.95 243.65 57.02 ;
    RECT 243.44 57.31 243.65 57.38 ;
    RECT 243.44 57.67 243.65 57.74 ;
    RECT 242.98 56.95 243.19 57.02 ;
    RECT 242.98 57.31 243.19 57.38 ;
    RECT 242.98 57.67 243.19 57.74 ;
    RECT 240.12 56.95 240.33 57.02 ;
    RECT 240.12 57.31 240.33 57.38 ;
    RECT 240.12 57.67 240.33 57.74 ;
    RECT 239.66 56.95 239.87 57.02 ;
    RECT 239.66 57.31 239.87 57.38 ;
    RECT 239.66 57.67 239.87 57.74 ;
    RECT 236.8 56.95 237.01 57.02 ;
    RECT 236.8 57.31 237.01 57.38 ;
    RECT 236.8 57.67 237.01 57.74 ;
    RECT 236.34 56.95 236.55 57.02 ;
    RECT 236.34 57.31 236.55 57.38 ;
    RECT 236.34 57.67 236.55 57.74 ;
    RECT 233.48 56.95 233.69 57.02 ;
    RECT 233.48 57.31 233.69 57.38 ;
    RECT 233.48 57.67 233.69 57.74 ;
    RECT 233.02 56.95 233.23 57.02 ;
    RECT 233.02 57.31 233.23 57.38 ;
    RECT 233.02 57.67 233.23 57.74 ;
    RECT 230.16 56.95 230.37 57.02 ;
    RECT 230.16 57.31 230.37 57.38 ;
    RECT 230.16 57.67 230.37 57.74 ;
    RECT 229.7 56.95 229.91 57.02 ;
    RECT 229.7 57.31 229.91 57.38 ;
    RECT 229.7 57.67 229.91 57.74 ;
    RECT 226.84 56.95 227.05 57.02 ;
    RECT 226.84 57.31 227.05 57.38 ;
    RECT 226.84 57.67 227.05 57.74 ;
    RECT 226.38 56.95 226.59 57.02 ;
    RECT 226.38 57.31 226.59 57.38 ;
    RECT 226.38 57.67 226.59 57.74 ;
    RECT 223.52 56.95 223.73 57.02 ;
    RECT 223.52 57.31 223.73 57.38 ;
    RECT 223.52 57.67 223.73 57.74 ;
    RECT 223.06 56.95 223.27 57.02 ;
    RECT 223.06 57.31 223.27 57.38 ;
    RECT 223.06 57.67 223.27 57.74 ;
    RECT 220.2 56.95 220.41 57.02 ;
    RECT 220.2 57.31 220.41 57.38 ;
    RECT 220.2 57.67 220.41 57.74 ;
    RECT 219.74 56.95 219.95 57.02 ;
    RECT 219.74 57.31 219.95 57.38 ;
    RECT 219.74 57.67 219.95 57.74 ;
    RECT 216.88 56.95 217.09 57.02 ;
    RECT 216.88 57.31 217.09 57.38 ;
    RECT 216.88 57.67 217.09 57.74 ;
    RECT 216.42 56.95 216.63 57.02 ;
    RECT 216.42 57.31 216.63 57.38 ;
    RECT 216.42 57.67 216.63 57.74 ;
    RECT 267.91 57.31 267.98 57.38 ;
    RECT 180.36 56.95 180.57 57.02 ;
    RECT 180.36 57.31 180.57 57.38 ;
    RECT 180.36 57.67 180.57 57.74 ;
    RECT 179.9 56.95 180.11 57.02 ;
    RECT 179.9 57.31 180.11 57.38 ;
    RECT 179.9 57.67 180.11 57.74 ;
    RECT 177.04 56.95 177.25 57.02 ;
    RECT 177.04 57.31 177.25 57.38 ;
    RECT 177.04 57.67 177.25 57.74 ;
    RECT 176.58 56.95 176.79 57.02 ;
    RECT 176.58 57.31 176.79 57.38 ;
    RECT 176.58 57.67 176.79 57.74 ;
    RECT 173.72 56.95 173.93 57.02 ;
    RECT 173.72 57.31 173.93 57.38 ;
    RECT 173.72 57.67 173.93 57.74 ;
    RECT 173.26 56.95 173.47 57.02 ;
    RECT 173.26 57.31 173.47 57.38 ;
    RECT 173.26 57.67 173.47 57.74 ;
    RECT 170.4 56.95 170.61 57.02 ;
    RECT 170.4 57.31 170.61 57.38 ;
    RECT 170.4 57.67 170.61 57.74 ;
    RECT 169.94 56.95 170.15 57.02 ;
    RECT 169.94 57.31 170.15 57.38 ;
    RECT 169.94 57.67 170.15 57.74 ;
    RECT 167.08 56.95 167.29 57.02 ;
    RECT 167.08 57.31 167.29 57.38 ;
    RECT 167.08 57.67 167.29 57.74 ;
    RECT 166.62 56.95 166.83 57.02 ;
    RECT 166.62 57.31 166.83 57.38 ;
    RECT 166.62 57.67 166.83 57.74 ;
    RECT 163.76 56.95 163.97 57.02 ;
    RECT 163.76 57.31 163.97 57.38 ;
    RECT 163.76 57.67 163.97 57.74 ;
    RECT 163.3 56.95 163.51 57.02 ;
    RECT 163.3 57.31 163.51 57.38 ;
    RECT 163.3 57.67 163.51 57.74 ;
    RECT 160.44 56.95 160.65 57.02 ;
    RECT 160.44 57.31 160.65 57.38 ;
    RECT 160.44 57.67 160.65 57.74 ;
    RECT 159.98 56.95 160.19 57.02 ;
    RECT 159.98 57.31 160.19 57.38 ;
    RECT 159.98 57.67 160.19 57.74 ;
    RECT 157.12 56.95 157.33 57.02 ;
    RECT 157.12 57.31 157.33 57.38 ;
    RECT 157.12 57.67 157.33 57.74 ;
    RECT 156.66 56.95 156.87 57.02 ;
    RECT 156.66 57.31 156.87 57.38 ;
    RECT 156.66 57.67 156.87 57.74 ;
    RECT 153.8 56.95 154.01 57.02 ;
    RECT 153.8 57.31 154.01 57.38 ;
    RECT 153.8 57.67 154.01 57.74 ;
    RECT 153.34 56.95 153.55 57.02 ;
    RECT 153.34 57.31 153.55 57.38 ;
    RECT 153.34 57.67 153.55 57.74 ;
    RECT 150.48 56.95 150.69 57.02 ;
    RECT 150.48 57.31 150.69 57.38 ;
    RECT 150.48 57.67 150.69 57.74 ;
    RECT 150.02 56.95 150.23 57.02 ;
    RECT 150.02 57.31 150.23 57.38 ;
    RECT 150.02 57.67 150.23 57.74 ;
    RECT 213.56 56.95 213.77 57.02 ;
    RECT 213.56 57.31 213.77 57.38 ;
    RECT 213.56 57.67 213.77 57.74 ;
    RECT 213.1 56.95 213.31 57.02 ;
    RECT 213.1 57.31 213.31 57.38 ;
    RECT 213.1 57.67 213.31 57.74 ;
    RECT 210.24 56.95 210.45 57.02 ;
    RECT 210.24 57.31 210.45 57.38 ;
    RECT 210.24 57.67 210.45 57.74 ;
    RECT 209.78 56.95 209.99 57.02 ;
    RECT 209.78 57.31 209.99 57.38 ;
    RECT 209.78 57.67 209.99 57.74 ;
    RECT 206.92 56.95 207.13 57.02 ;
    RECT 206.92 57.31 207.13 57.38 ;
    RECT 206.92 57.67 207.13 57.74 ;
    RECT 206.46 56.95 206.67 57.02 ;
    RECT 206.46 57.31 206.67 57.38 ;
    RECT 206.46 57.67 206.67 57.74 ;
    RECT 203.6 56.95 203.81 57.02 ;
    RECT 203.6 57.31 203.81 57.38 ;
    RECT 203.6 57.67 203.81 57.74 ;
    RECT 203.14 56.95 203.35 57.02 ;
    RECT 203.14 57.31 203.35 57.38 ;
    RECT 203.14 57.67 203.35 57.74 ;
    RECT 200.28 56.95 200.49 57.02 ;
    RECT 200.28 57.31 200.49 57.38 ;
    RECT 200.28 57.67 200.49 57.74 ;
    RECT 199.82 56.95 200.03 57.02 ;
    RECT 199.82 57.31 200.03 57.38 ;
    RECT 199.82 57.67 200.03 57.74 ;
    RECT 196.96 56.95 197.17 57.02 ;
    RECT 196.96 57.31 197.17 57.38 ;
    RECT 196.96 57.67 197.17 57.74 ;
    RECT 196.5 56.95 196.71 57.02 ;
    RECT 196.5 57.31 196.71 57.38 ;
    RECT 196.5 57.67 196.71 57.74 ;
    RECT 193.64 56.95 193.85 57.02 ;
    RECT 193.64 57.31 193.85 57.38 ;
    RECT 193.64 57.67 193.85 57.74 ;
    RECT 193.18 56.95 193.39 57.02 ;
    RECT 193.18 57.31 193.39 57.38 ;
    RECT 193.18 57.67 193.39 57.74 ;
    RECT 190.32 56.95 190.53 57.02 ;
    RECT 190.32 57.31 190.53 57.38 ;
    RECT 190.32 57.67 190.53 57.74 ;
    RECT 189.86 56.95 190.07 57.02 ;
    RECT 189.86 57.31 190.07 57.38 ;
    RECT 189.86 57.67 190.07 57.74 ;
    RECT 187.0 56.95 187.21 57.02 ;
    RECT 187.0 57.31 187.21 57.38 ;
    RECT 187.0 57.67 187.21 57.74 ;
    RECT 186.54 56.95 186.75 57.02 ;
    RECT 186.54 57.31 186.75 57.38 ;
    RECT 186.54 57.67 186.75 57.74 ;
    RECT 183.68 56.95 183.89 57.02 ;
    RECT 183.68 57.31 183.89 57.38 ;
    RECT 183.68 57.67 183.89 57.74 ;
    RECT 183.22 56.95 183.43 57.02 ;
    RECT 183.22 57.31 183.43 57.38 ;
    RECT 183.22 57.67 183.43 57.74 ;
    RECT 147.485 57.31 147.555 57.38 ;
    RECT 266.68 56.95 266.89 57.02 ;
    RECT 266.68 57.31 266.89 57.38 ;
    RECT 266.68 57.67 266.89 57.74 ;
    RECT 266.22 56.95 266.43 57.02 ;
    RECT 266.22 57.31 266.43 57.38 ;
    RECT 266.22 57.67 266.43 57.74 ;
    RECT 263.36 56.95 263.57 57.02 ;
    RECT 263.36 57.31 263.57 57.38 ;
    RECT 263.36 57.67 263.57 57.74 ;
    RECT 262.9 56.95 263.11 57.02 ;
    RECT 262.9 57.31 263.11 57.38 ;
    RECT 262.9 57.67 263.11 57.74 ;
    RECT 260.04 56.95 260.25 57.02 ;
    RECT 260.04 57.31 260.25 57.38 ;
    RECT 260.04 57.67 260.25 57.74 ;
    RECT 259.58 56.95 259.79 57.02 ;
    RECT 259.58 57.31 259.79 57.38 ;
    RECT 259.58 57.67 259.79 57.74 ;
    RECT 256.72 56.95 256.93 57.02 ;
    RECT 256.72 57.31 256.93 57.38 ;
    RECT 256.72 57.67 256.93 57.74 ;
    RECT 256.26 56.95 256.47 57.02 ;
    RECT 256.26 57.31 256.47 57.38 ;
    RECT 256.26 57.67 256.47 57.74 ;
    RECT 253.4 56.95 253.61 57.02 ;
    RECT 253.4 57.31 253.61 57.38 ;
    RECT 253.4 57.67 253.61 57.74 ;
    RECT 252.94 56.95 253.15 57.02 ;
    RECT 252.94 57.31 253.15 57.38 ;
    RECT 252.94 57.67 253.15 57.74 ;
    RECT 250.08 92.97 250.29 93.04 ;
    RECT 250.08 93.33 250.29 93.4 ;
    RECT 250.08 93.69 250.29 93.76 ;
    RECT 249.62 92.97 249.83 93.04 ;
    RECT 249.62 93.33 249.83 93.4 ;
    RECT 249.62 93.69 249.83 93.76 ;
    RECT 246.76 92.97 246.97 93.04 ;
    RECT 246.76 93.33 246.97 93.4 ;
    RECT 246.76 93.69 246.97 93.76 ;
    RECT 246.3 92.97 246.51 93.04 ;
    RECT 246.3 93.33 246.51 93.4 ;
    RECT 246.3 93.69 246.51 93.76 ;
    RECT 243.44 92.97 243.65 93.04 ;
    RECT 243.44 93.33 243.65 93.4 ;
    RECT 243.44 93.69 243.65 93.76 ;
    RECT 242.98 92.97 243.19 93.04 ;
    RECT 242.98 93.33 243.19 93.4 ;
    RECT 242.98 93.69 243.19 93.76 ;
    RECT 240.12 92.97 240.33 93.04 ;
    RECT 240.12 93.33 240.33 93.4 ;
    RECT 240.12 93.69 240.33 93.76 ;
    RECT 239.66 92.97 239.87 93.04 ;
    RECT 239.66 93.33 239.87 93.4 ;
    RECT 239.66 93.69 239.87 93.76 ;
    RECT 236.8 92.97 237.01 93.04 ;
    RECT 236.8 93.33 237.01 93.4 ;
    RECT 236.8 93.69 237.01 93.76 ;
    RECT 236.34 92.97 236.55 93.04 ;
    RECT 236.34 93.33 236.55 93.4 ;
    RECT 236.34 93.69 236.55 93.76 ;
    RECT 233.48 92.97 233.69 93.04 ;
    RECT 233.48 93.33 233.69 93.4 ;
    RECT 233.48 93.69 233.69 93.76 ;
    RECT 233.02 92.97 233.23 93.04 ;
    RECT 233.02 93.33 233.23 93.4 ;
    RECT 233.02 93.69 233.23 93.76 ;
    RECT 230.16 92.97 230.37 93.04 ;
    RECT 230.16 93.33 230.37 93.4 ;
    RECT 230.16 93.69 230.37 93.76 ;
    RECT 229.7 92.97 229.91 93.04 ;
    RECT 229.7 93.33 229.91 93.4 ;
    RECT 229.7 93.69 229.91 93.76 ;
    RECT 226.84 92.97 227.05 93.04 ;
    RECT 226.84 93.33 227.05 93.4 ;
    RECT 226.84 93.69 227.05 93.76 ;
    RECT 226.38 92.97 226.59 93.04 ;
    RECT 226.38 93.33 226.59 93.4 ;
    RECT 226.38 93.69 226.59 93.76 ;
    RECT 223.52 92.97 223.73 93.04 ;
    RECT 223.52 93.33 223.73 93.4 ;
    RECT 223.52 93.69 223.73 93.76 ;
    RECT 223.06 92.97 223.27 93.04 ;
    RECT 223.06 93.33 223.27 93.4 ;
    RECT 223.06 93.69 223.27 93.76 ;
    RECT 220.2 92.97 220.41 93.04 ;
    RECT 220.2 93.33 220.41 93.4 ;
    RECT 220.2 93.69 220.41 93.76 ;
    RECT 219.74 92.97 219.95 93.04 ;
    RECT 219.74 93.33 219.95 93.4 ;
    RECT 219.74 93.69 219.95 93.76 ;
    RECT 216.88 92.97 217.09 93.04 ;
    RECT 216.88 93.33 217.09 93.4 ;
    RECT 216.88 93.69 217.09 93.76 ;
    RECT 216.42 92.97 216.63 93.04 ;
    RECT 216.42 93.33 216.63 93.4 ;
    RECT 216.42 93.69 216.63 93.76 ;
    RECT 267.91 93.33 267.98 93.4 ;
    RECT 180.36 92.97 180.57 93.04 ;
    RECT 180.36 93.33 180.57 93.4 ;
    RECT 180.36 93.69 180.57 93.76 ;
    RECT 179.9 92.97 180.11 93.04 ;
    RECT 179.9 93.33 180.11 93.4 ;
    RECT 179.9 93.69 180.11 93.76 ;
    RECT 177.04 92.97 177.25 93.04 ;
    RECT 177.04 93.33 177.25 93.4 ;
    RECT 177.04 93.69 177.25 93.76 ;
    RECT 176.58 92.97 176.79 93.04 ;
    RECT 176.58 93.33 176.79 93.4 ;
    RECT 176.58 93.69 176.79 93.76 ;
    RECT 173.72 92.97 173.93 93.04 ;
    RECT 173.72 93.33 173.93 93.4 ;
    RECT 173.72 93.69 173.93 93.76 ;
    RECT 173.26 92.97 173.47 93.04 ;
    RECT 173.26 93.33 173.47 93.4 ;
    RECT 173.26 93.69 173.47 93.76 ;
    RECT 170.4 92.97 170.61 93.04 ;
    RECT 170.4 93.33 170.61 93.4 ;
    RECT 170.4 93.69 170.61 93.76 ;
    RECT 169.94 92.97 170.15 93.04 ;
    RECT 169.94 93.33 170.15 93.4 ;
    RECT 169.94 93.69 170.15 93.76 ;
    RECT 167.08 92.97 167.29 93.04 ;
    RECT 167.08 93.33 167.29 93.4 ;
    RECT 167.08 93.69 167.29 93.76 ;
    RECT 166.62 92.97 166.83 93.04 ;
    RECT 166.62 93.33 166.83 93.4 ;
    RECT 166.62 93.69 166.83 93.76 ;
    RECT 163.76 92.97 163.97 93.04 ;
    RECT 163.76 93.33 163.97 93.4 ;
    RECT 163.76 93.69 163.97 93.76 ;
    RECT 163.3 92.97 163.51 93.04 ;
    RECT 163.3 93.33 163.51 93.4 ;
    RECT 163.3 93.69 163.51 93.76 ;
    RECT 160.44 92.97 160.65 93.04 ;
    RECT 160.44 93.33 160.65 93.4 ;
    RECT 160.44 93.69 160.65 93.76 ;
    RECT 159.98 92.97 160.19 93.04 ;
    RECT 159.98 93.33 160.19 93.4 ;
    RECT 159.98 93.69 160.19 93.76 ;
    RECT 157.12 92.97 157.33 93.04 ;
    RECT 157.12 93.33 157.33 93.4 ;
    RECT 157.12 93.69 157.33 93.76 ;
    RECT 156.66 92.97 156.87 93.04 ;
    RECT 156.66 93.33 156.87 93.4 ;
    RECT 156.66 93.69 156.87 93.76 ;
    RECT 153.8 92.97 154.01 93.04 ;
    RECT 153.8 93.33 154.01 93.4 ;
    RECT 153.8 93.69 154.01 93.76 ;
    RECT 153.34 92.97 153.55 93.04 ;
    RECT 153.34 93.33 153.55 93.4 ;
    RECT 153.34 93.69 153.55 93.76 ;
    RECT 150.48 92.97 150.69 93.04 ;
    RECT 150.48 93.33 150.69 93.4 ;
    RECT 150.48 93.69 150.69 93.76 ;
    RECT 150.02 92.97 150.23 93.04 ;
    RECT 150.02 93.33 150.23 93.4 ;
    RECT 150.02 93.69 150.23 93.76 ;
    RECT 213.56 92.97 213.77 93.04 ;
    RECT 213.56 93.33 213.77 93.4 ;
    RECT 213.56 93.69 213.77 93.76 ;
    RECT 213.1 92.97 213.31 93.04 ;
    RECT 213.1 93.33 213.31 93.4 ;
    RECT 213.1 93.69 213.31 93.76 ;
    RECT 210.24 92.97 210.45 93.04 ;
    RECT 210.24 93.33 210.45 93.4 ;
    RECT 210.24 93.69 210.45 93.76 ;
    RECT 209.78 92.97 209.99 93.04 ;
    RECT 209.78 93.33 209.99 93.4 ;
    RECT 209.78 93.69 209.99 93.76 ;
    RECT 206.92 92.97 207.13 93.04 ;
    RECT 206.92 93.33 207.13 93.4 ;
    RECT 206.92 93.69 207.13 93.76 ;
    RECT 206.46 92.97 206.67 93.04 ;
    RECT 206.46 93.33 206.67 93.4 ;
    RECT 206.46 93.69 206.67 93.76 ;
    RECT 203.6 92.97 203.81 93.04 ;
    RECT 203.6 93.33 203.81 93.4 ;
    RECT 203.6 93.69 203.81 93.76 ;
    RECT 203.14 92.97 203.35 93.04 ;
    RECT 203.14 93.33 203.35 93.4 ;
    RECT 203.14 93.69 203.35 93.76 ;
    RECT 200.28 92.97 200.49 93.04 ;
    RECT 200.28 93.33 200.49 93.4 ;
    RECT 200.28 93.69 200.49 93.76 ;
    RECT 199.82 92.97 200.03 93.04 ;
    RECT 199.82 93.33 200.03 93.4 ;
    RECT 199.82 93.69 200.03 93.76 ;
    RECT 196.96 92.97 197.17 93.04 ;
    RECT 196.96 93.33 197.17 93.4 ;
    RECT 196.96 93.69 197.17 93.76 ;
    RECT 196.5 92.97 196.71 93.04 ;
    RECT 196.5 93.33 196.71 93.4 ;
    RECT 196.5 93.69 196.71 93.76 ;
    RECT 193.64 92.97 193.85 93.04 ;
    RECT 193.64 93.33 193.85 93.4 ;
    RECT 193.64 93.69 193.85 93.76 ;
    RECT 193.18 92.97 193.39 93.04 ;
    RECT 193.18 93.33 193.39 93.4 ;
    RECT 193.18 93.69 193.39 93.76 ;
    RECT 190.32 92.97 190.53 93.04 ;
    RECT 190.32 93.33 190.53 93.4 ;
    RECT 190.32 93.69 190.53 93.76 ;
    RECT 189.86 92.97 190.07 93.04 ;
    RECT 189.86 93.33 190.07 93.4 ;
    RECT 189.86 93.69 190.07 93.76 ;
    RECT 187.0 92.97 187.21 93.04 ;
    RECT 187.0 93.33 187.21 93.4 ;
    RECT 187.0 93.69 187.21 93.76 ;
    RECT 186.54 92.97 186.75 93.04 ;
    RECT 186.54 93.33 186.75 93.4 ;
    RECT 186.54 93.69 186.75 93.76 ;
    RECT 183.68 92.97 183.89 93.04 ;
    RECT 183.68 93.33 183.89 93.4 ;
    RECT 183.68 93.69 183.89 93.76 ;
    RECT 183.22 92.97 183.43 93.04 ;
    RECT 183.22 93.33 183.43 93.4 ;
    RECT 183.22 93.69 183.43 93.76 ;
    RECT 147.485 93.33 147.555 93.4 ;
    RECT 266.68 92.97 266.89 93.04 ;
    RECT 266.68 93.33 266.89 93.4 ;
    RECT 266.68 93.69 266.89 93.76 ;
    RECT 266.22 92.97 266.43 93.04 ;
    RECT 266.22 93.33 266.43 93.4 ;
    RECT 266.22 93.69 266.43 93.76 ;
    RECT 263.36 92.97 263.57 93.04 ;
    RECT 263.36 93.33 263.57 93.4 ;
    RECT 263.36 93.69 263.57 93.76 ;
    RECT 262.9 92.97 263.11 93.04 ;
    RECT 262.9 93.33 263.11 93.4 ;
    RECT 262.9 93.69 263.11 93.76 ;
    RECT 260.04 92.97 260.25 93.04 ;
    RECT 260.04 93.33 260.25 93.4 ;
    RECT 260.04 93.69 260.25 93.76 ;
    RECT 259.58 92.97 259.79 93.04 ;
    RECT 259.58 93.33 259.79 93.4 ;
    RECT 259.58 93.69 259.79 93.76 ;
    RECT 256.72 92.97 256.93 93.04 ;
    RECT 256.72 93.33 256.93 93.4 ;
    RECT 256.72 93.69 256.93 93.76 ;
    RECT 256.26 92.97 256.47 93.04 ;
    RECT 256.26 93.33 256.47 93.4 ;
    RECT 256.26 93.69 256.47 93.76 ;
    RECT 253.4 92.97 253.61 93.04 ;
    RECT 253.4 93.33 253.61 93.4 ;
    RECT 253.4 93.69 253.61 93.76 ;
    RECT 252.94 92.97 253.15 93.04 ;
    RECT 252.94 93.33 253.15 93.4 ;
    RECT 252.94 93.69 253.15 93.76 ;
    RECT 250.08 92.25 250.29 92.32 ;
    RECT 250.08 92.61 250.29 92.68 ;
    RECT 250.08 92.97 250.29 93.04 ;
    RECT 249.62 92.25 249.83 92.32 ;
    RECT 249.62 92.61 249.83 92.68 ;
    RECT 249.62 92.97 249.83 93.04 ;
    RECT 246.76 92.25 246.97 92.32 ;
    RECT 246.76 92.61 246.97 92.68 ;
    RECT 246.76 92.97 246.97 93.04 ;
    RECT 246.3 92.25 246.51 92.32 ;
    RECT 246.3 92.61 246.51 92.68 ;
    RECT 246.3 92.97 246.51 93.04 ;
    RECT 243.44 92.25 243.65 92.32 ;
    RECT 243.44 92.61 243.65 92.68 ;
    RECT 243.44 92.97 243.65 93.04 ;
    RECT 242.98 92.25 243.19 92.32 ;
    RECT 242.98 92.61 243.19 92.68 ;
    RECT 242.98 92.97 243.19 93.04 ;
    RECT 240.12 92.25 240.33 92.32 ;
    RECT 240.12 92.61 240.33 92.68 ;
    RECT 240.12 92.97 240.33 93.04 ;
    RECT 239.66 92.25 239.87 92.32 ;
    RECT 239.66 92.61 239.87 92.68 ;
    RECT 239.66 92.97 239.87 93.04 ;
    RECT 236.8 92.25 237.01 92.32 ;
    RECT 236.8 92.61 237.01 92.68 ;
    RECT 236.8 92.97 237.01 93.04 ;
    RECT 236.34 92.25 236.55 92.32 ;
    RECT 236.34 92.61 236.55 92.68 ;
    RECT 236.34 92.97 236.55 93.04 ;
    RECT 233.48 92.25 233.69 92.32 ;
    RECT 233.48 92.61 233.69 92.68 ;
    RECT 233.48 92.97 233.69 93.04 ;
    RECT 233.02 92.25 233.23 92.32 ;
    RECT 233.02 92.61 233.23 92.68 ;
    RECT 233.02 92.97 233.23 93.04 ;
    RECT 230.16 92.25 230.37 92.32 ;
    RECT 230.16 92.61 230.37 92.68 ;
    RECT 230.16 92.97 230.37 93.04 ;
    RECT 229.7 92.25 229.91 92.32 ;
    RECT 229.7 92.61 229.91 92.68 ;
    RECT 229.7 92.97 229.91 93.04 ;
    RECT 226.84 92.25 227.05 92.32 ;
    RECT 226.84 92.61 227.05 92.68 ;
    RECT 226.84 92.97 227.05 93.04 ;
    RECT 226.38 92.25 226.59 92.32 ;
    RECT 226.38 92.61 226.59 92.68 ;
    RECT 226.38 92.97 226.59 93.04 ;
    RECT 223.52 92.25 223.73 92.32 ;
    RECT 223.52 92.61 223.73 92.68 ;
    RECT 223.52 92.97 223.73 93.04 ;
    RECT 223.06 92.25 223.27 92.32 ;
    RECT 223.06 92.61 223.27 92.68 ;
    RECT 223.06 92.97 223.27 93.04 ;
    RECT 220.2 92.25 220.41 92.32 ;
    RECT 220.2 92.61 220.41 92.68 ;
    RECT 220.2 92.97 220.41 93.04 ;
    RECT 219.74 92.25 219.95 92.32 ;
    RECT 219.74 92.61 219.95 92.68 ;
    RECT 219.74 92.97 219.95 93.04 ;
    RECT 216.88 92.25 217.09 92.32 ;
    RECT 216.88 92.61 217.09 92.68 ;
    RECT 216.88 92.97 217.09 93.04 ;
    RECT 216.42 92.25 216.63 92.32 ;
    RECT 216.42 92.61 216.63 92.68 ;
    RECT 216.42 92.97 216.63 93.04 ;
    RECT 267.91 92.61 267.98 92.68 ;
    RECT 180.36 92.25 180.57 92.32 ;
    RECT 180.36 92.61 180.57 92.68 ;
    RECT 180.36 92.97 180.57 93.04 ;
    RECT 179.9 92.25 180.11 92.32 ;
    RECT 179.9 92.61 180.11 92.68 ;
    RECT 179.9 92.97 180.11 93.04 ;
    RECT 177.04 92.25 177.25 92.32 ;
    RECT 177.04 92.61 177.25 92.68 ;
    RECT 177.04 92.97 177.25 93.04 ;
    RECT 176.58 92.25 176.79 92.32 ;
    RECT 176.58 92.61 176.79 92.68 ;
    RECT 176.58 92.97 176.79 93.04 ;
    RECT 173.72 92.25 173.93 92.32 ;
    RECT 173.72 92.61 173.93 92.68 ;
    RECT 173.72 92.97 173.93 93.04 ;
    RECT 173.26 92.25 173.47 92.32 ;
    RECT 173.26 92.61 173.47 92.68 ;
    RECT 173.26 92.97 173.47 93.04 ;
    RECT 170.4 92.25 170.61 92.32 ;
    RECT 170.4 92.61 170.61 92.68 ;
    RECT 170.4 92.97 170.61 93.04 ;
    RECT 169.94 92.25 170.15 92.32 ;
    RECT 169.94 92.61 170.15 92.68 ;
    RECT 169.94 92.97 170.15 93.04 ;
    RECT 167.08 92.25 167.29 92.32 ;
    RECT 167.08 92.61 167.29 92.68 ;
    RECT 167.08 92.97 167.29 93.04 ;
    RECT 166.62 92.25 166.83 92.32 ;
    RECT 166.62 92.61 166.83 92.68 ;
    RECT 166.62 92.97 166.83 93.04 ;
    RECT 163.76 92.25 163.97 92.32 ;
    RECT 163.76 92.61 163.97 92.68 ;
    RECT 163.76 92.97 163.97 93.04 ;
    RECT 163.3 92.25 163.51 92.32 ;
    RECT 163.3 92.61 163.51 92.68 ;
    RECT 163.3 92.97 163.51 93.04 ;
    RECT 160.44 92.25 160.65 92.32 ;
    RECT 160.44 92.61 160.65 92.68 ;
    RECT 160.44 92.97 160.65 93.04 ;
    RECT 159.98 92.25 160.19 92.32 ;
    RECT 159.98 92.61 160.19 92.68 ;
    RECT 159.98 92.97 160.19 93.04 ;
    RECT 157.12 92.25 157.33 92.32 ;
    RECT 157.12 92.61 157.33 92.68 ;
    RECT 157.12 92.97 157.33 93.04 ;
    RECT 156.66 92.25 156.87 92.32 ;
    RECT 156.66 92.61 156.87 92.68 ;
    RECT 156.66 92.97 156.87 93.04 ;
    RECT 153.8 92.25 154.01 92.32 ;
    RECT 153.8 92.61 154.01 92.68 ;
    RECT 153.8 92.97 154.01 93.04 ;
    RECT 153.34 92.25 153.55 92.32 ;
    RECT 153.34 92.61 153.55 92.68 ;
    RECT 153.34 92.97 153.55 93.04 ;
    RECT 150.48 92.25 150.69 92.32 ;
    RECT 150.48 92.61 150.69 92.68 ;
    RECT 150.48 92.97 150.69 93.04 ;
    RECT 150.02 92.25 150.23 92.32 ;
    RECT 150.02 92.61 150.23 92.68 ;
    RECT 150.02 92.97 150.23 93.04 ;
    RECT 213.56 92.25 213.77 92.32 ;
    RECT 213.56 92.61 213.77 92.68 ;
    RECT 213.56 92.97 213.77 93.04 ;
    RECT 213.1 92.25 213.31 92.32 ;
    RECT 213.1 92.61 213.31 92.68 ;
    RECT 213.1 92.97 213.31 93.04 ;
    RECT 210.24 92.25 210.45 92.32 ;
    RECT 210.24 92.61 210.45 92.68 ;
    RECT 210.24 92.97 210.45 93.04 ;
    RECT 209.78 92.25 209.99 92.32 ;
    RECT 209.78 92.61 209.99 92.68 ;
    RECT 209.78 92.97 209.99 93.04 ;
    RECT 206.92 92.25 207.13 92.32 ;
    RECT 206.92 92.61 207.13 92.68 ;
    RECT 206.92 92.97 207.13 93.04 ;
    RECT 206.46 92.25 206.67 92.32 ;
    RECT 206.46 92.61 206.67 92.68 ;
    RECT 206.46 92.97 206.67 93.04 ;
    RECT 203.6 92.25 203.81 92.32 ;
    RECT 203.6 92.61 203.81 92.68 ;
    RECT 203.6 92.97 203.81 93.04 ;
    RECT 203.14 92.25 203.35 92.32 ;
    RECT 203.14 92.61 203.35 92.68 ;
    RECT 203.14 92.97 203.35 93.04 ;
    RECT 200.28 92.25 200.49 92.32 ;
    RECT 200.28 92.61 200.49 92.68 ;
    RECT 200.28 92.97 200.49 93.04 ;
    RECT 199.82 92.25 200.03 92.32 ;
    RECT 199.82 92.61 200.03 92.68 ;
    RECT 199.82 92.97 200.03 93.04 ;
    RECT 196.96 92.25 197.17 92.32 ;
    RECT 196.96 92.61 197.17 92.68 ;
    RECT 196.96 92.97 197.17 93.04 ;
    RECT 196.5 92.25 196.71 92.32 ;
    RECT 196.5 92.61 196.71 92.68 ;
    RECT 196.5 92.97 196.71 93.04 ;
    RECT 193.64 92.25 193.85 92.32 ;
    RECT 193.64 92.61 193.85 92.68 ;
    RECT 193.64 92.97 193.85 93.04 ;
    RECT 193.18 92.25 193.39 92.32 ;
    RECT 193.18 92.61 193.39 92.68 ;
    RECT 193.18 92.97 193.39 93.04 ;
    RECT 190.32 92.25 190.53 92.32 ;
    RECT 190.32 92.61 190.53 92.68 ;
    RECT 190.32 92.97 190.53 93.04 ;
    RECT 189.86 92.25 190.07 92.32 ;
    RECT 189.86 92.61 190.07 92.68 ;
    RECT 189.86 92.97 190.07 93.04 ;
    RECT 187.0 92.25 187.21 92.32 ;
    RECT 187.0 92.61 187.21 92.68 ;
    RECT 187.0 92.97 187.21 93.04 ;
    RECT 186.54 92.25 186.75 92.32 ;
    RECT 186.54 92.61 186.75 92.68 ;
    RECT 186.54 92.97 186.75 93.04 ;
    RECT 183.68 92.25 183.89 92.32 ;
    RECT 183.68 92.61 183.89 92.68 ;
    RECT 183.68 92.97 183.89 93.04 ;
    RECT 183.22 92.25 183.43 92.32 ;
    RECT 183.22 92.61 183.43 92.68 ;
    RECT 183.22 92.97 183.43 93.04 ;
    RECT 147.485 92.61 147.555 92.68 ;
    RECT 266.68 92.25 266.89 92.32 ;
    RECT 266.68 92.61 266.89 92.68 ;
    RECT 266.68 92.97 266.89 93.04 ;
    RECT 266.22 92.25 266.43 92.32 ;
    RECT 266.22 92.61 266.43 92.68 ;
    RECT 266.22 92.97 266.43 93.04 ;
    RECT 263.36 92.25 263.57 92.32 ;
    RECT 263.36 92.61 263.57 92.68 ;
    RECT 263.36 92.97 263.57 93.04 ;
    RECT 262.9 92.25 263.11 92.32 ;
    RECT 262.9 92.61 263.11 92.68 ;
    RECT 262.9 92.97 263.11 93.04 ;
    RECT 260.04 92.25 260.25 92.32 ;
    RECT 260.04 92.61 260.25 92.68 ;
    RECT 260.04 92.97 260.25 93.04 ;
    RECT 259.58 92.25 259.79 92.32 ;
    RECT 259.58 92.61 259.79 92.68 ;
    RECT 259.58 92.97 259.79 93.04 ;
    RECT 256.72 92.25 256.93 92.32 ;
    RECT 256.72 92.61 256.93 92.68 ;
    RECT 256.72 92.97 256.93 93.04 ;
    RECT 256.26 92.25 256.47 92.32 ;
    RECT 256.26 92.61 256.47 92.68 ;
    RECT 256.26 92.97 256.47 93.04 ;
    RECT 253.4 92.25 253.61 92.32 ;
    RECT 253.4 92.61 253.61 92.68 ;
    RECT 253.4 92.97 253.61 93.04 ;
    RECT 252.94 92.25 253.15 92.32 ;
    RECT 252.94 92.61 253.15 92.68 ;
    RECT 252.94 92.97 253.15 93.04 ;
    RECT 250.08 91.53 250.29 91.6 ;
    RECT 250.08 91.89 250.29 91.96 ;
    RECT 250.08 92.25 250.29 92.32 ;
    RECT 249.62 91.53 249.83 91.6 ;
    RECT 249.62 91.89 249.83 91.96 ;
    RECT 249.62 92.25 249.83 92.32 ;
    RECT 246.76 91.53 246.97 91.6 ;
    RECT 246.76 91.89 246.97 91.96 ;
    RECT 246.76 92.25 246.97 92.32 ;
    RECT 246.3 91.53 246.51 91.6 ;
    RECT 246.3 91.89 246.51 91.96 ;
    RECT 246.3 92.25 246.51 92.32 ;
    RECT 243.44 91.53 243.65 91.6 ;
    RECT 243.44 91.89 243.65 91.96 ;
    RECT 243.44 92.25 243.65 92.32 ;
    RECT 242.98 91.53 243.19 91.6 ;
    RECT 242.98 91.89 243.19 91.96 ;
    RECT 242.98 92.25 243.19 92.32 ;
    RECT 240.12 91.53 240.33 91.6 ;
    RECT 240.12 91.89 240.33 91.96 ;
    RECT 240.12 92.25 240.33 92.32 ;
    RECT 239.66 91.53 239.87 91.6 ;
    RECT 239.66 91.89 239.87 91.96 ;
    RECT 239.66 92.25 239.87 92.32 ;
    RECT 236.8 91.53 237.01 91.6 ;
    RECT 236.8 91.89 237.01 91.96 ;
    RECT 236.8 92.25 237.01 92.32 ;
    RECT 236.34 91.53 236.55 91.6 ;
    RECT 236.34 91.89 236.55 91.96 ;
    RECT 236.34 92.25 236.55 92.32 ;
    RECT 233.48 91.53 233.69 91.6 ;
    RECT 233.48 91.89 233.69 91.96 ;
    RECT 233.48 92.25 233.69 92.32 ;
    RECT 233.02 91.53 233.23 91.6 ;
    RECT 233.02 91.89 233.23 91.96 ;
    RECT 233.02 92.25 233.23 92.32 ;
    RECT 230.16 91.53 230.37 91.6 ;
    RECT 230.16 91.89 230.37 91.96 ;
    RECT 230.16 92.25 230.37 92.32 ;
    RECT 229.7 91.53 229.91 91.6 ;
    RECT 229.7 91.89 229.91 91.96 ;
    RECT 229.7 92.25 229.91 92.32 ;
    RECT 226.84 91.53 227.05 91.6 ;
    RECT 226.84 91.89 227.05 91.96 ;
    RECT 226.84 92.25 227.05 92.32 ;
    RECT 226.38 91.53 226.59 91.6 ;
    RECT 226.38 91.89 226.59 91.96 ;
    RECT 226.38 92.25 226.59 92.32 ;
    RECT 223.52 91.53 223.73 91.6 ;
    RECT 223.52 91.89 223.73 91.96 ;
    RECT 223.52 92.25 223.73 92.32 ;
    RECT 223.06 91.53 223.27 91.6 ;
    RECT 223.06 91.89 223.27 91.96 ;
    RECT 223.06 92.25 223.27 92.32 ;
    RECT 220.2 91.53 220.41 91.6 ;
    RECT 220.2 91.89 220.41 91.96 ;
    RECT 220.2 92.25 220.41 92.32 ;
    RECT 219.74 91.53 219.95 91.6 ;
    RECT 219.74 91.89 219.95 91.96 ;
    RECT 219.74 92.25 219.95 92.32 ;
    RECT 216.88 91.53 217.09 91.6 ;
    RECT 216.88 91.89 217.09 91.96 ;
    RECT 216.88 92.25 217.09 92.32 ;
    RECT 216.42 91.53 216.63 91.6 ;
    RECT 216.42 91.89 216.63 91.96 ;
    RECT 216.42 92.25 216.63 92.32 ;
    RECT 267.91 91.89 267.98 91.96 ;
    RECT 180.36 91.53 180.57 91.6 ;
    RECT 180.36 91.89 180.57 91.96 ;
    RECT 180.36 92.25 180.57 92.32 ;
    RECT 179.9 91.53 180.11 91.6 ;
    RECT 179.9 91.89 180.11 91.96 ;
    RECT 179.9 92.25 180.11 92.32 ;
    RECT 177.04 91.53 177.25 91.6 ;
    RECT 177.04 91.89 177.25 91.96 ;
    RECT 177.04 92.25 177.25 92.32 ;
    RECT 176.58 91.53 176.79 91.6 ;
    RECT 176.58 91.89 176.79 91.96 ;
    RECT 176.58 92.25 176.79 92.32 ;
    RECT 173.72 91.53 173.93 91.6 ;
    RECT 173.72 91.89 173.93 91.96 ;
    RECT 173.72 92.25 173.93 92.32 ;
    RECT 173.26 91.53 173.47 91.6 ;
    RECT 173.26 91.89 173.47 91.96 ;
    RECT 173.26 92.25 173.47 92.32 ;
    RECT 170.4 91.53 170.61 91.6 ;
    RECT 170.4 91.89 170.61 91.96 ;
    RECT 170.4 92.25 170.61 92.32 ;
    RECT 169.94 91.53 170.15 91.6 ;
    RECT 169.94 91.89 170.15 91.96 ;
    RECT 169.94 92.25 170.15 92.32 ;
    RECT 167.08 91.53 167.29 91.6 ;
    RECT 167.08 91.89 167.29 91.96 ;
    RECT 167.08 92.25 167.29 92.32 ;
    RECT 166.62 91.53 166.83 91.6 ;
    RECT 166.62 91.89 166.83 91.96 ;
    RECT 166.62 92.25 166.83 92.32 ;
    RECT 163.76 91.53 163.97 91.6 ;
    RECT 163.76 91.89 163.97 91.96 ;
    RECT 163.76 92.25 163.97 92.32 ;
    RECT 163.3 91.53 163.51 91.6 ;
    RECT 163.3 91.89 163.51 91.96 ;
    RECT 163.3 92.25 163.51 92.32 ;
    RECT 160.44 91.53 160.65 91.6 ;
    RECT 160.44 91.89 160.65 91.96 ;
    RECT 160.44 92.25 160.65 92.32 ;
    RECT 159.98 91.53 160.19 91.6 ;
    RECT 159.98 91.89 160.19 91.96 ;
    RECT 159.98 92.25 160.19 92.32 ;
    RECT 157.12 91.53 157.33 91.6 ;
    RECT 157.12 91.89 157.33 91.96 ;
    RECT 157.12 92.25 157.33 92.32 ;
    RECT 156.66 91.53 156.87 91.6 ;
    RECT 156.66 91.89 156.87 91.96 ;
    RECT 156.66 92.25 156.87 92.32 ;
    RECT 153.8 91.53 154.01 91.6 ;
    RECT 153.8 91.89 154.01 91.96 ;
    RECT 153.8 92.25 154.01 92.32 ;
    RECT 153.34 91.53 153.55 91.6 ;
    RECT 153.34 91.89 153.55 91.96 ;
    RECT 153.34 92.25 153.55 92.32 ;
    RECT 150.48 91.53 150.69 91.6 ;
    RECT 150.48 91.89 150.69 91.96 ;
    RECT 150.48 92.25 150.69 92.32 ;
    RECT 150.02 91.53 150.23 91.6 ;
    RECT 150.02 91.89 150.23 91.96 ;
    RECT 150.02 92.25 150.23 92.32 ;
    RECT 213.56 91.53 213.77 91.6 ;
    RECT 213.56 91.89 213.77 91.96 ;
    RECT 213.56 92.25 213.77 92.32 ;
    RECT 213.1 91.53 213.31 91.6 ;
    RECT 213.1 91.89 213.31 91.96 ;
    RECT 213.1 92.25 213.31 92.32 ;
    RECT 210.24 91.53 210.45 91.6 ;
    RECT 210.24 91.89 210.45 91.96 ;
    RECT 210.24 92.25 210.45 92.32 ;
    RECT 209.78 91.53 209.99 91.6 ;
    RECT 209.78 91.89 209.99 91.96 ;
    RECT 209.78 92.25 209.99 92.32 ;
    RECT 206.92 91.53 207.13 91.6 ;
    RECT 206.92 91.89 207.13 91.96 ;
    RECT 206.92 92.25 207.13 92.32 ;
    RECT 206.46 91.53 206.67 91.6 ;
    RECT 206.46 91.89 206.67 91.96 ;
    RECT 206.46 92.25 206.67 92.32 ;
    RECT 203.6 91.53 203.81 91.6 ;
    RECT 203.6 91.89 203.81 91.96 ;
    RECT 203.6 92.25 203.81 92.32 ;
    RECT 203.14 91.53 203.35 91.6 ;
    RECT 203.14 91.89 203.35 91.96 ;
    RECT 203.14 92.25 203.35 92.32 ;
    RECT 200.28 91.53 200.49 91.6 ;
    RECT 200.28 91.89 200.49 91.96 ;
    RECT 200.28 92.25 200.49 92.32 ;
    RECT 199.82 91.53 200.03 91.6 ;
    RECT 199.82 91.89 200.03 91.96 ;
    RECT 199.82 92.25 200.03 92.32 ;
    RECT 196.96 91.53 197.17 91.6 ;
    RECT 196.96 91.89 197.17 91.96 ;
    RECT 196.96 92.25 197.17 92.32 ;
    RECT 196.5 91.53 196.71 91.6 ;
    RECT 196.5 91.89 196.71 91.96 ;
    RECT 196.5 92.25 196.71 92.32 ;
    RECT 193.64 91.53 193.85 91.6 ;
    RECT 193.64 91.89 193.85 91.96 ;
    RECT 193.64 92.25 193.85 92.32 ;
    RECT 193.18 91.53 193.39 91.6 ;
    RECT 193.18 91.89 193.39 91.96 ;
    RECT 193.18 92.25 193.39 92.32 ;
    RECT 190.32 91.53 190.53 91.6 ;
    RECT 190.32 91.89 190.53 91.96 ;
    RECT 190.32 92.25 190.53 92.32 ;
    RECT 189.86 91.53 190.07 91.6 ;
    RECT 189.86 91.89 190.07 91.96 ;
    RECT 189.86 92.25 190.07 92.32 ;
    RECT 187.0 91.53 187.21 91.6 ;
    RECT 187.0 91.89 187.21 91.96 ;
    RECT 187.0 92.25 187.21 92.32 ;
    RECT 186.54 91.53 186.75 91.6 ;
    RECT 186.54 91.89 186.75 91.96 ;
    RECT 186.54 92.25 186.75 92.32 ;
    RECT 183.68 91.53 183.89 91.6 ;
    RECT 183.68 91.89 183.89 91.96 ;
    RECT 183.68 92.25 183.89 92.32 ;
    RECT 183.22 91.53 183.43 91.6 ;
    RECT 183.22 91.89 183.43 91.96 ;
    RECT 183.22 92.25 183.43 92.32 ;
    RECT 147.485 91.89 147.555 91.96 ;
    RECT 266.68 91.53 266.89 91.6 ;
    RECT 266.68 91.89 266.89 91.96 ;
    RECT 266.68 92.25 266.89 92.32 ;
    RECT 266.22 91.53 266.43 91.6 ;
    RECT 266.22 91.89 266.43 91.96 ;
    RECT 266.22 92.25 266.43 92.32 ;
    RECT 263.36 91.53 263.57 91.6 ;
    RECT 263.36 91.89 263.57 91.96 ;
    RECT 263.36 92.25 263.57 92.32 ;
    RECT 262.9 91.53 263.11 91.6 ;
    RECT 262.9 91.89 263.11 91.96 ;
    RECT 262.9 92.25 263.11 92.32 ;
    RECT 260.04 91.53 260.25 91.6 ;
    RECT 260.04 91.89 260.25 91.96 ;
    RECT 260.04 92.25 260.25 92.32 ;
    RECT 259.58 91.53 259.79 91.6 ;
    RECT 259.58 91.89 259.79 91.96 ;
    RECT 259.58 92.25 259.79 92.32 ;
    RECT 256.72 91.53 256.93 91.6 ;
    RECT 256.72 91.89 256.93 91.96 ;
    RECT 256.72 92.25 256.93 92.32 ;
    RECT 256.26 91.53 256.47 91.6 ;
    RECT 256.26 91.89 256.47 91.96 ;
    RECT 256.26 92.25 256.47 92.32 ;
    RECT 253.4 91.53 253.61 91.6 ;
    RECT 253.4 91.89 253.61 91.96 ;
    RECT 253.4 92.25 253.61 92.32 ;
    RECT 252.94 91.53 253.15 91.6 ;
    RECT 252.94 91.89 253.15 91.96 ;
    RECT 252.94 92.25 253.15 92.32 ;
    RECT 250.08 90.81 250.29 90.88 ;
    RECT 250.08 91.17 250.29 91.24 ;
    RECT 250.08 91.53 250.29 91.6 ;
    RECT 249.62 90.81 249.83 90.88 ;
    RECT 249.62 91.17 249.83 91.24 ;
    RECT 249.62 91.53 249.83 91.6 ;
    RECT 246.76 90.81 246.97 90.88 ;
    RECT 246.76 91.17 246.97 91.24 ;
    RECT 246.76 91.53 246.97 91.6 ;
    RECT 246.3 90.81 246.51 90.88 ;
    RECT 246.3 91.17 246.51 91.24 ;
    RECT 246.3 91.53 246.51 91.6 ;
    RECT 243.44 90.81 243.65 90.88 ;
    RECT 243.44 91.17 243.65 91.24 ;
    RECT 243.44 91.53 243.65 91.6 ;
    RECT 242.98 90.81 243.19 90.88 ;
    RECT 242.98 91.17 243.19 91.24 ;
    RECT 242.98 91.53 243.19 91.6 ;
    RECT 240.12 90.81 240.33 90.88 ;
    RECT 240.12 91.17 240.33 91.24 ;
    RECT 240.12 91.53 240.33 91.6 ;
    RECT 239.66 90.81 239.87 90.88 ;
    RECT 239.66 91.17 239.87 91.24 ;
    RECT 239.66 91.53 239.87 91.6 ;
    RECT 236.8 90.81 237.01 90.88 ;
    RECT 236.8 91.17 237.01 91.24 ;
    RECT 236.8 91.53 237.01 91.6 ;
    RECT 236.34 90.81 236.55 90.88 ;
    RECT 236.34 91.17 236.55 91.24 ;
    RECT 236.34 91.53 236.55 91.6 ;
    RECT 233.48 90.81 233.69 90.88 ;
    RECT 233.48 91.17 233.69 91.24 ;
    RECT 233.48 91.53 233.69 91.6 ;
    RECT 233.02 90.81 233.23 90.88 ;
    RECT 233.02 91.17 233.23 91.24 ;
    RECT 233.02 91.53 233.23 91.6 ;
    RECT 230.16 90.81 230.37 90.88 ;
    RECT 230.16 91.17 230.37 91.24 ;
    RECT 230.16 91.53 230.37 91.6 ;
    RECT 229.7 90.81 229.91 90.88 ;
    RECT 229.7 91.17 229.91 91.24 ;
    RECT 229.7 91.53 229.91 91.6 ;
    RECT 226.84 90.81 227.05 90.88 ;
    RECT 226.84 91.17 227.05 91.24 ;
    RECT 226.84 91.53 227.05 91.6 ;
    RECT 226.38 90.81 226.59 90.88 ;
    RECT 226.38 91.17 226.59 91.24 ;
    RECT 226.38 91.53 226.59 91.6 ;
    RECT 223.52 90.81 223.73 90.88 ;
    RECT 223.52 91.17 223.73 91.24 ;
    RECT 223.52 91.53 223.73 91.6 ;
    RECT 223.06 90.81 223.27 90.88 ;
    RECT 223.06 91.17 223.27 91.24 ;
    RECT 223.06 91.53 223.27 91.6 ;
    RECT 220.2 90.81 220.41 90.88 ;
    RECT 220.2 91.17 220.41 91.24 ;
    RECT 220.2 91.53 220.41 91.6 ;
    RECT 219.74 90.81 219.95 90.88 ;
    RECT 219.74 91.17 219.95 91.24 ;
    RECT 219.74 91.53 219.95 91.6 ;
    RECT 216.88 90.81 217.09 90.88 ;
    RECT 216.88 91.17 217.09 91.24 ;
    RECT 216.88 91.53 217.09 91.6 ;
    RECT 216.42 90.81 216.63 90.88 ;
    RECT 216.42 91.17 216.63 91.24 ;
    RECT 216.42 91.53 216.63 91.6 ;
    RECT 267.91 91.17 267.98 91.24 ;
    RECT 180.36 90.81 180.57 90.88 ;
    RECT 180.36 91.17 180.57 91.24 ;
    RECT 180.36 91.53 180.57 91.6 ;
    RECT 179.9 90.81 180.11 90.88 ;
    RECT 179.9 91.17 180.11 91.24 ;
    RECT 179.9 91.53 180.11 91.6 ;
    RECT 177.04 90.81 177.25 90.88 ;
    RECT 177.04 91.17 177.25 91.24 ;
    RECT 177.04 91.53 177.25 91.6 ;
    RECT 176.58 90.81 176.79 90.88 ;
    RECT 176.58 91.17 176.79 91.24 ;
    RECT 176.58 91.53 176.79 91.6 ;
    RECT 173.72 90.81 173.93 90.88 ;
    RECT 173.72 91.17 173.93 91.24 ;
    RECT 173.72 91.53 173.93 91.6 ;
    RECT 173.26 90.81 173.47 90.88 ;
    RECT 173.26 91.17 173.47 91.24 ;
    RECT 173.26 91.53 173.47 91.6 ;
    RECT 170.4 90.81 170.61 90.88 ;
    RECT 170.4 91.17 170.61 91.24 ;
    RECT 170.4 91.53 170.61 91.6 ;
    RECT 169.94 90.81 170.15 90.88 ;
    RECT 169.94 91.17 170.15 91.24 ;
    RECT 169.94 91.53 170.15 91.6 ;
    RECT 167.08 90.81 167.29 90.88 ;
    RECT 167.08 91.17 167.29 91.24 ;
    RECT 167.08 91.53 167.29 91.6 ;
    RECT 166.62 90.81 166.83 90.88 ;
    RECT 166.62 91.17 166.83 91.24 ;
    RECT 166.62 91.53 166.83 91.6 ;
    RECT 163.76 90.81 163.97 90.88 ;
    RECT 163.76 91.17 163.97 91.24 ;
    RECT 163.76 91.53 163.97 91.6 ;
    RECT 163.3 90.81 163.51 90.88 ;
    RECT 163.3 91.17 163.51 91.24 ;
    RECT 163.3 91.53 163.51 91.6 ;
    RECT 160.44 90.81 160.65 90.88 ;
    RECT 160.44 91.17 160.65 91.24 ;
    RECT 160.44 91.53 160.65 91.6 ;
    RECT 159.98 90.81 160.19 90.88 ;
    RECT 159.98 91.17 160.19 91.24 ;
    RECT 159.98 91.53 160.19 91.6 ;
    RECT 157.12 90.81 157.33 90.88 ;
    RECT 157.12 91.17 157.33 91.24 ;
    RECT 157.12 91.53 157.33 91.6 ;
    RECT 156.66 90.81 156.87 90.88 ;
    RECT 156.66 91.17 156.87 91.24 ;
    RECT 156.66 91.53 156.87 91.6 ;
    RECT 153.8 90.81 154.01 90.88 ;
    RECT 153.8 91.17 154.01 91.24 ;
    RECT 153.8 91.53 154.01 91.6 ;
    RECT 153.34 90.81 153.55 90.88 ;
    RECT 153.34 91.17 153.55 91.24 ;
    RECT 153.34 91.53 153.55 91.6 ;
    RECT 150.48 90.81 150.69 90.88 ;
    RECT 150.48 91.17 150.69 91.24 ;
    RECT 150.48 91.53 150.69 91.6 ;
    RECT 150.02 90.81 150.23 90.88 ;
    RECT 150.02 91.17 150.23 91.24 ;
    RECT 150.02 91.53 150.23 91.6 ;
    RECT 213.56 90.81 213.77 90.88 ;
    RECT 213.56 91.17 213.77 91.24 ;
    RECT 213.56 91.53 213.77 91.6 ;
    RECT 213.1 90.81 213.31 90.88 ;
    RECT 213.1 91.17 213.31 91.24 ;
    RECT 213.1 91.53 213.31 91.6 ;
    RECT 210.24 90.81 210.45 90.88 ;
    RECT 210.24 91.17 210.45 91.24 ;
    RECT 210.24 91.53 210.45 91.6 ;
    RECT 209.78 90.81 209.99 90.88 ;
    RECT 209.78 91.17 209.99 91.24 ;
    RECT 209.78 91.53 209.99 91.6 ;
    RECT 206.92 90.81 207.13 90.88 ;
    RECT 206.92 91.17 207.13 91.24 ;
    RECT 206.92 91.53 207.13 91.6 ;
    RECT 206.46 90.81 206.67 90.88 ;
    RECT 206.46 91.17 206.67 91.24 ;
    RECT 206.46 91.53 206.67 91.6 ;
    RECT 203.6 90.81 203.81 90.88 ;
    RECT 203.6 91.17 203.81 91.24 ;
    RECT 203.6 91.53 203.81 91.6 ;
    RECT 203.14 90.81 203.35 90.88 ;
    RECT 203.14 91.17 203.35 91.24 ;
    RECT 203.14 91.53 203.35 91.6 ;
    RECT 200.28 90.81 200.49 90.88 ;
    RECT 200.28 91.17 200.49 91.24 ;
    RECT 200.28 91.53 200.49 91.6 ;
    RECT 199.82 90.81 200.03 90.88 ;
    RECT 199.82 91.17 200.03 91.24 ;
    RECT 199.82 91.53 200.03 91.6 ;
    RECT 196.96 90.81 197.17 90.88 ;
    RECT 196.96 91.17 197.17 91.24 ;
    RECT 196.96 91.53 197.17 91.6 ;
    RECT 196.5 90.81 196.71 90.88 ;
    RECT 196.5 91.17 196.71 91.24 ;
    RECT 196.5 91.53 196.71 91.6 ;
    RECT 193.64 90.81 193.85 90.88 ;
    RECT 193.64 91.17 193.85 91.24 ;
    RECT 193.64 91.53 193.85 91.6 ;
    RECT 193.18 90.81 193.39 90.88 ;
    RECT 193.18 91.17 193.39 91.24 ;
    RECT 193.18 91.53 193.39 91.6 ;
    RECT 190.32 90.81 190.53 90.88 ;
    RECT 190.32 91.17 190.53 91.24 ;
    RECT 190.32 91.53 190.53 91.6 ;
    RECT 189.86 90.81 190.07 90.88 ;
    RECT 189.86 91.17 190.07 91.24 ;
    RECT 189.86 91.53 190.07 91.6 ;
    RECT 187.0 90.81 187.21 90.88 ;
    RECT 187.0 91.17 187.21 91.24 ;
    RECT 187.0 91.53 187.21 91.6 ;
    RECT 186.54 90.81 186.75 90.88 ;
    RECT 186.54 91.17 186.75 91.24 ;
    RECT 186.54 91.53 186.75 91.6 ;
    RECT 183.68 90.81 183.89 90.88 ;
    RECT 183.68 91.17 183.89 91.24 ;
    RECT 183.68 91.53 183.89 91.6 ;
    RECT 183.22 90.81 183.43 90.88 ;
    RECT 183.22 91.17 183.43 91.24 ;
    RECT 183.22 91.53 183.43 91.6 ;
    RECT 147.485 91.17 147.555 91.24 ;
    RECT 266.68 90.81 266.89 90.88 ;
    RECT 266.68 91.17 266.89 91.24 ;
    RECT 266.68 91.53 266.89 91.6 ;
    RECT 266.22 90.81 266.43 90.88 ;
    RECT 266.22 91.17 266.43 91.24 ;
    RECT 266.22 91.53 266.43 91.6 ;
    RECT 263.36 90.81 263.57 90.88 ;
    RECT 263.36 91.17 263.57 91.24 ;
    RECT 263.36 91.53 263.57 91.6 ;
    RECT 262.9 90.81 263.11 90.88 ;
    RECT 262.9 91.17 263.11 91.24 ;
    RECT 262.9 91.53 263.11 91.6 ;
    RECT 260.04 90.81 260.25 90.88 ;
    RECT 260.04 91.17 260.25 91.24 ;
    RECT 260.04 91.53 260.25 91.6 ;
    RECT 259.58 90.81 259.79 90.88 ;
    RECT 259.58 91.17 259.79 91.24 ;
    RECT 259.58 91.53 259.79 91.6 ;
    RECT 256.72 90.81 256.93 90.88 ;
    RECT 256.72 91.17 256.93 91.24 ;
    RECT 256.72 91.53 256.93 91.6 ;
    RECT 256.26 90.81 256.47 90.88 ;
    RECT 256.26 91.17 256.47 91.24 ;
    RECT 256.26 91.53 256.47 91.6 ;
    RECT 253.4 90.81 253.61 90.88 ;
    RECT 253.4 91.17 253.61 91.24 ;
    RECT 253.4 91.53 253.61 91.6 ;
    RECT 252.94 90.81 253.15 90.88 ;
    RECT 252.94 91.17 253.15 91.24 ;
    RECT 252.94 91.53 253.15 91.6 ;
    RECT 250.08 54.07 250.29 54.14 ;
    RECT 250.08 54.43 250.29 54.5 ;
    RECT 250.08 54.79 250.29 54.86 ;
    RECT 249.62 54.07 249.83 54.14 ;
    RECT 249.62 54.43 249.83 54.5 ;
    RECT 249.62 54.79 249.83 54.86 ;
    RECT 246.76 54.07 246.97 54.14 ;
    RECT 246.76 54.43 246.97 54.5 ;
    RECT 246.76 54.79 246.97 54.86 ;
    RECT 246.3 54.07 246.51 54.14 ;
    RECT 246.3 54.43 246.51 54.5 ;
    RECT 246.3 54.79 246.51 54.86 ;
    RECT 243.44 54.07 243.65 54.14 ;
    RECT 243.44 54.43 243.65 54.5 ;
    RECT 243.44 54.79 243.65 54.86 ;
    RECT 242.98 54.07 243.19 54.14 ;
    RECT 242.98 54.43 243.19 54.5 ;
    RECT 242.98 54.79 243.19 54.86 ;
    RECT 240.12 54.07 240.33 54.14 ;
    RECT 240.12 54.43 240.33 54.5 ;
    RECT 240.12 54.79 240.33 54.86 ;
    RECT 239.66 54.07 239.87 54.14 ;
    RECT 239.66 54.43 239.87 54.5 ;
    RECT 239.66 54.79 239.87 54.86 ;
    RECT 236.8 54.07 237.01 54.14 ;
    RECT 236.8 54.43 237.01 54.5 ;
    RECT 236.8 54.79 237.01 54.86 ;
    RECT 236.34 54.07 236.55 54.14 ;
    RECT 236.34 54.43 236.55 54.5 ;
    RECT 236.34 54.79 236.55 54.86 ;
    RECT 233.48 54.07 233.69 54.14 ;
    RECT 233.48 54.43 233.69 54.5 ;
    RECT 233.48 54.79 233.69 54.86 ;
    RECT 233.02 54.07 233.23 54.14 ;
    RECT 233.02 54.43 233.23 54.5 ;
    RECT 233.02 54.79 233.23 54.86 ;
    RECT 230.16 54.07 230.37 54.14 ;
    RECT 230.16 54.43 230.37 54.5 ;
    RECT 230.16 54.79 230.37 54.86 ;
    RECT 229.7 54.07 229.91 54.14 ;
    RECT 229.7 54.43 229.91 54.5 ;
    RECT 229.7 54.79 229.91 54.86 ;
    RECT 226.84 54.07 227.05 54.14 ;
    RECT 226.84 54.43 227.05 54.5 ;
    RECT 226.84 54.79 227.05 54.86 ;
    RECT 226.38 54.07 226.59 54.14 ;
    RECT 226.38 54.43 226.59 54.5 ;
    RECT 226.38 54.79 226.59 54.86 ;
    RECT 223.52 54.07 223.73 54.14 ;
    RECT 223.52 54.43 223.73 54.5 ;
    RECT 223.52 54.79 223.73 54.86 ;
    RECT 223.06 54.07 223.27 54.14 ;
    RECT 223.06 54.43 223.27 54.5 ;
    RECT 223.06 54.79 223.27 54.86 ;
    RECT 220.2 54.07 220.41 54.14 ;
    RECT 220.2 54.43 220.41 54.5 ;
    RECT 220.2 54.79 220.41 54.86 ;
    RECT 219.74 54.07 219.95 54.14 ;
    RECT 219.74 54.43 219.95 54.5 ;
    RECT 219.74 54.79 219.95 54.86 ;
    RECT 216.88 54.07 217.09 54.14 ;
    RECT 216.88 54.43 217.09 54.5 ;
    RECT 216.88 54.79 217.09 54.86 ;
    RECT 216.42 54.07 216.63 54.14 ;
    RECT 216.42 54.43 216.63 54.5 ;
    RECT 216.42 54.79 216.63 54.86 ;
    RECT 267.91 54.43 267.98 54.5 ;
    RECT 180.36 54.07 180.57 54.14 ;
    RECT 180.36 54.43 180.57 54.5 ;
    RECT 180.36 54.79 180.57 54.86 ;
    RECT 179.9 54.07 180.11 54.14 ;
    RECT 179.9 54.43 180.11 54.5 ;
    RECT 179.9 54.79 180.11 54.86 ;
    RECT 177.04 54.07 177.25 54.14 ;
    RECT 177.04 54.43 177.25 54.5 ;
    RECT 177.04 54.79 177.25 54.86 ;
    RECT 176.58 54.07 176.79 54.14 ;
    RECT 176.58 54.43 176.79 54.5 ;
    RECT 176.58 54.79 176.79 54.86 ;
    RECT 173.72 54.07 173.93 54.14 ;
    RECT 173.72 54.43 173.93 54.5 ;
    RECT 173.72 54.79 173.93 54.86 ;
    RECT 173.26 54.07 173.47 54.14 ;
    RECT 173.26 54.43 173.47 54.5 ;
    RECT 173.26 54.79 173.47 54.86 ;
    RECT 170.4 54.07 170.61 54.14 ;
    RECT 170.4 54.43 170.61 54.5 ;
    RECT 170.4 54.79 170.61 54.86 ;
    RECT 169.94 54.07 170.15 54.14 ;
    RECT 169.94 54.43 170.15 54.5 ;
    RECT 169.94 54.79 170.15 54.86 ;
    RECT 167.08 54.07 167.29 54.14 ;
    RECT 167.08 54.43 167.29 54.5 ;
    RECT 167.08 54.79 167.29 54.86 ;
    RECT 166.62 54.07 166.83 54.14 ;
    RECT 166.62 54.43 166.83 54.5 ;
    RECT 166.62 54.79 166.83 54.86 ;
    RECT 163.76 54.07 163.97 54.14 ;
    RECT 163.76 54.43 163.97 54.5 ;
    RECT 163.76 54.79 163.97 54.86 ;
    RECT 163.3 54.07 163.51 54.14 ;
    RECT 163.3 54.43 163.51 54.5 ;
    RECT 163.3 54.79 163.51 54.86 ;
    RECT 160.44 54.07 160.65 54.14 ;
    RECT 160.44 54.43 160.65 54.5 ;
    RECT 160.44 54.79 160.65 54.86 ;
    RECT 159.98 54.07 160.19 54.14 ;
    RECT 159.98 54.43 160.19 54.5 ;
    RECT 159.98 54.79 160.19 54.86 ;
    RECT 157.12 54.07 157.33 54.14 ;
    RECT 157.12 54.43 157.33 54.5 ;
    RECT 157.12 54.79 157.33 54.86 ;
    RECT 156.66 54.07 156.87 54.14 ;
    RECT 156.66 54.43 156.87 54.5 ;
    RECT 156.66 54.79 156.87 54.86 ;
    RECT 153.8 54.07 154.01 54.14 ;
    RECT 153.8 54.43 154.01 54.5 ;
    RECT 153.8 54.79 154.01 54.86 ;
    RECT 153.34 54.07 153.55 54.14 ;
    RECT 153.34 54.43 153.55 54.5 ;
    RECT 153.34 54.79 153.55 54.86 ;
    RECT 150.48 54.07 150.69 54.14 ;
    RECT 150.48 54.43 150.69 54.5 ;
    RECT 150.48 54.79 150.69 54.86 ;
    RECT 150.02 54.07 150.23 54.14 ;
    RECT 150.02 54.43 150.23 54.5 ;
    RECT 150.02 54.79 150.23 54.86 ;
    RECT 213.56 54.07 213.77 54.14 ;
    RECT 213.56 54.43 213.77 54.5 ;
    RECT 213.56 54.79 213.77 54.86 ;
    RECT 213.1 54.07 213.31 54.14 ;
    RECT 213.1 54.43 213.31 54.5 ;
    RECT 213.1 54.79 213.31 54.86 ;
    RECT 210.24 54.07 210.45 54.14 ;
    RECT 210.24 54.43 210.45 54.5 ;
    RECT 210.24 54.79 210.45 54.86 ;
    RECT 209.78 54.07 209.99 54.14 ;
    RECT 209.78 54.43 209.99 54.5 ;
    RECT 209.78 54.79 209.99 54.86 ;
    RECT 206.92 54.07 207.13 54.14 ;
    RECT 206.92 54.43 207.13 54.5 ;
    RECT 206.92 54.79 207.13 54.86 ;
    RECT 206.46 54.07 206.67 54.14 ;
    RECT 206.46 54.43 206.67 54.5 ;
    RECT 206.46 54.79 206.67 54.86 ;
    RECT 203.6 54.07 203.81 54.14 ;
    RECT 203.6 54.43 203.81 54.5 ;
    RECT 203.6 54.79 203.81 54.86 ;
    RECT 203.14 54.07 203.35 54.14 ;
    RECT 203.14 54.43 203.35 54.5 ;
    RECT 203.14 54.79 203.35 54.86 ;
    RECT 200.28 54.07 200.49 54.14 ;
    RECT 200.28 54.43 200.49 54.5 ;
    RECT 200.28 54.79 200.49 54.86 ;
    RECT 199.82 54.07 200.03 54.14 ;
    RECT 199.82 54.43 200.03 54.5 ;
    RECT 199.82 54.79 200.03 54.86 ;
    RECT 196.96 54.07 197.17 54.14 ;
    RECT 196.96 54.43 197.17 54.5 ;
    RECT 196.96 54.79 197.17 54.86 ;
    RECT 196.5 54.07 196.71 54.14 ;
    RECT 196.5 54.43 196.71 54.5 ;
    RECT 196.5 54.79 196.71 54.86 ;
    RECT 193.64 54.07 193.85 54.14 ;
    RECT 193.64 54.43 193.85 54.5 ;
    RECT 193.64 54.79 193.85 54.86 ;
    RECT 193.18 54.07 193.39 54.14 ;
    RECT 193.18 54.43 193.39 54.5 ;
    RECT 193.18 54.79 193.39 54.86 ;
    RECT 190.32 54.07 190.53 54.14 ;
    RECT 190.32 54.43 190.53 54.5 ;
    RECT 190.32 54.79 190.53 54.86 ;
    RECT 189.86 54.07 190.07 54.14 ;
    RECT 189.86 54.43 190.07 54.5 ;
    RECT 189.86 54.79 190.07 54.86 ;
    RECT 187.0 54.07 187.21 54.14 ;
    RECT 187.0 54.43 187.21 54.5 ;
    RECT 187.0 54.79 187.21 54.86 ;
    RECT 186.54 54.07 186.75 54.14 ;
    RECT 186.54 54.43 186.75 54.5 ;
    RECT 186.54 54.79 186.75 54.86 ;
    RECT 183.68 54.07 183.89 54.14 ;
    RECT 183.68 54.43 183.89 54.5 ;
    RECT 183.68 54.79 183.89 54.86 ;
    RECT 183.22 54.07 183.43 54.14 ;
    RECT 183.22 54.43 183.43 54.5 ;
    RECT 183.22 54.79 183.43 54.86 ;
    RECT 147.485 54.43 147.555 54.5 ;
    RECT 266.68 54.07 266.89 54.14 ;
    RECT 266.68 54.43 266.89 54.5 ;
    RECT 266.68 54.79 266.89 54.86 ;
    RECT 266.22 54.07 266.43 54.14 ;
    RECT 266.22 54.43 266.43 54.5 ;
    RECT 266.22 54.79 266.43 54.86 ;
    RECT 263.36 54.07 263.57 54.14 ;
    RECT 263.36 54.43 263.57 54.5 ;
    RECT 263.36 54.79 263.57 54.86 ;
    RECT 262.9 54.07 263.11 54.14 ;
    RECT 262.9 54.43 263.11 54.5 ;
    RECT 262.9 54.79 263.11 54.86 ;
    RECT 260.04 54.07 260.25 54.14 ;
    RECT 260.04 54.43 260.25 54.5 ;
    RECT 260.04 54.79 260.25 54.86 ;
    RECT 259.58 54.07 259.79 54.14 ;
    RECT 259.58 54.43 259.79 54.5 ;
    RECT 259.58 54.79 259.79 54.86 ;
    RECT 256.72 54.07 256.93 54.14 ;
    RECT 256.72 54.43 256.93 54.5 ;
    RECT 256.72 54.79 256.93 54.86 ;
    RECT 256.26 54.07 256.47 54.14 ;
    RECT 256.26 54.43 256.47 54.5 ;
    RECT 256.26 54.79 256.47 54.86 ;
    RECT 253.4 54.07 253.61 54.14 ;
    RECT 253.4 54.43 253.61 54.5 ;
    RECT 253.4 54.79 253.61 54.86 ;
    RECT 252.94 54.07 253.15 54.14 ;
    RECT 252.94 54.43 253.15 54.5 ;
    RECT 252.94 54.79 253.15 54.86 ;
    RECT 250.08 90.09 250.29 90.16 ;
    RECT 250.08 90.45 250.29 90.52 ;
    RECT 250.08 90.81 250.29 90.88 ;
    RECT 249.62 90.09 249.83 90.16 ;
    RECT 249.62 90.45 249.83 90.52 ;
    RECT 249.62 90.81 249.83 90.88 ;
    RECT 246.76 90.09 246.97 90.16 ;
    RECT 246.76 90.45 246.97 90.52 ;
    RECT 246.76 90.81 246.97 90.88 ;
    RECT 246.3 90.09 246.51 90.16 ;
    RECT 246.3 90.45 246.51 90.52 ;
    RECT 246.3 90.81 246.51 90.88 ;
    RECT 243.44 90.09 243.65 90.16 ;
    RECT 243.44 90.45 243.65 90.52 ;
    RECT 243.44 90.81 243.65 90.88 ;
    RECT 242.98 90.09 243.19 90.16 ;
    RECT 242.98 90.45 243.19 90.52 ;
    RECT 242.98 90.81 243.19 90.88 ;
    RECT 240.12 90.09 240.33 90.16 ;
    RECT 240.12 90.45 240.33 90.52 ;
    RECT 240.12 90.81 240.33 90.88 ;
    RECT 239.66 90.09 239.87 90.16 ;
    RECT 239.66 90.45 239.87 90.52 ;
    RECT 239.66 90.81 239.87 90.88 ;
    RECT 236.8 90.09 237.01 90.16 ;
    RECT 236.8 90.45 237.01 90.52 ;
    RECT 236.8 90.81 237.01 90.88 ;
    RECT 236.34 90.09 236.55 90.16 ;
    RECT 236.34 90.45 236.55 90.52 ;
    RECT 236.34 90.81 236.55 90.88 ;
    RECT 233.48 90.09 233.69 90.16 ;
    RECT 233.48 90.45 233.69 90.52 ;
    RECT 233.48 90.81 233.69 90.88 ;
    RECT 233.02 90.09 233.23 90.16 ;
    RECT 233.02 90.45 233.23 90.52 ;
    RECT 233.02 90.81 233.23 90.88 ;
    RECT 230.16 90.09 230.37 90.16 ;
    RECT 230.16 90.45 230.37 90.52 ;
    RECT 230.16 90.81 230.37 90.88 ;
    RECT 229.7 90.09 229.91 90.16 ;
    RECT 229.7 90.45 229.91 90.52 ;
    RECT 229.7 90.81 229.91 90.88 ;
    RECT 226.84 90.09 227.05 90.16 ;
    RECT 226.84 90.45 227.05 90.52 ;
    RECT 226.84 90.81 227.05 90.88 ;
    RECT 226.38 90.09 226.59 90.16 ;
    RECT 226.38 90.45 226.59 90.52 ;
    RECT 226.38 90.81 226.59 90.88 ;
    RECT 223.52 90.09 223.73 90.16 ;
    RECT 223.52 90.45 223.73 90.52 ;
    RECT 223.52 90.81 223.73 90.88 ;
    RECT 223.06 90.09 223.27 90.16 ;
    RECT 223.06 90.45 223.27 90.52 ;
    RECT 223.06 90.81 223.27 90.88 ;
    RECT 220.2 90.09 220.41 90.16 ;
    RECT 220.2 90.45 220.41 90.52 ;
    RECT 220.2 90.81 220.41 90.88 ;
    RECT 219.74 90.09 219.95 90.16 ;
    RECT 219.74 90.45 219.95 90.52 ;
    RECT 219.74 90.81 219.95 90.88 ;
    RECT 216.88 90.09 217.09 90.16 ;
    RECT 216.88 90.45 217.09 90.52 ;
    RECT 216.88 90.81 217.09 90.88 ;
    RECT 216.42 90.09 216.63 90.16 ;
    RECT 216.42 90.45 216.63 90.52 ;
    RECT 216.42 90.81 216.63 90.88 ;
    RECT 267.91 90.45 267.98 90.52 ;
    RECT 180.36 90.09 180.57 90.16 ;
    RECT 180.36 90.45 180.57 90.52 ;
    RECT 180.36 90.81 180.57 90.88 ;
    RECT 179.9 90.09 180.11 90.16 ;
    RECT 179.9 90.45 180.11 90.52 ;
    RECT 179.9 90.81 180.11 90.88 ;
    RECT 177.04 90.09 177.25 90.16 ;
    RECT 177.04 90.45 177.25 90.52 ;
    RECT 177.04 90.81 177.25 90.88 ;
    RECT 176.58 90.09 176.79 90.16 ;
    RECT 176.58 90.45 176.79 90.52 ;
    RECT 176.58 90.81 176.79 90.88 ;
    RECT 173.72 90.09 173.93 90.16 ;
    RECT 173.72 90.45 173.93 90.52 ;
    RECT 173.72 90.81 173.93 90.88 ;
    RECT 173.26 90.09 173.47 90.16 ;
    RECT 173.26 90.45 173.47 90.52 ;
    RECT 173.26 90.81 173.47 90.88 ;
    RECT 170.4 90.09 170.61 90.16 ;
    RECT 170.4 90.45 170.61 90.52 ;
    RECT 170.4 90.81 170.61 90.88 ;
    RECT 169.94 90.09 170.15 90.16 ;
    RECT 169.94 90.45 170.15 90.52 ;
    RECT 169.94 90.81 170.15 90.88 ;
    RECT 167.08 90.09 167.29 90.16 ;
    RECT 167.08 90.45 167.29 90.52 ;
    RECT 167.08 90.81 167.29 90.88 ;
    RECT 166.62 90.09 166.83 90.16 ;
    RECT 166.62 90.45 166.83 90.52 ;
    RECT 166.62 90.81 166.83 90.88 ;
    RECT 163.76 90.09 163.97 90.16 ;
    RECT 163.76 90.45 163.97 90.52 ;
    RECT 163.76 90.81 163.97 90.88 ;
    RECT 163.3 90.09 163.51 90.16 ;
    RECT 163.3 90.45 163.51 90.52 ;
    RECT 163.3 90.81 163.51 90.88 ;
    RECT 160.44 90.09 160.65 90.16 ;
    RECT 160.44 90.45 160.65 90.52 ;
    RECT 160.44 90.81 160.65 90.88 ;
    RECT 159.98 90.09 160.19 90.16 ;
    RECT 159.98 90.45 160.19 90.52 ;
    RECT 159.98 90.81 160.19 90.88 ;
    RECT 157.12 90.09 157.33 90.16 ;
    RECT 157.12 90.45 157.33 90.52 ;
    RECT 157.12 90.81 157.33 90.88 ;
    RECT 156.66 90.09 156.87 90.16 ;
    RECT 156.66 90.45 156.87 90.52 ;
    RECT 156.66 90.81 156.87 90.88 ;
    RECT 153.8 90.09 154.01 90.16 ;
    RECT 153.8 90.45 154.01 90.52 ;
    RECT 153.8 90.81 154.01 90.88 ;
    RECT 153.34 90.09 153.55 90.16 ;
    RECT 153.34 90.45 153.55 90.52 ;
    RECT 153.34 90.81 153.55 90.88 ;
    RECT 150.48 90.09 150.69 90.16 ;
    RECT 150.48 90.45 150.69 90.52 ;
    RECT 150.48 90.81 150.69 90.88 ;
    RECT 150.02 90.09 150.23 90.16 ;
    RECT 150.02 90.45 150.23 90.52 ;
    RECT 150.02 90.81 150.23 90.88 ;
    RECT 213.56 90.09 213.77 90.16 ;
    RECT 213.56 90.45 213.77 90.52 ;
    RECT 213.56 90.81 213.77 90.88 ;
    RECT 213.1 90.09 213.31 90.16 ;
    RECT 213.1 90.45 213.31 90.52 ;
    RECT 213.1 90.81 213.31 90.88 ;
    RECT 210.24 90.09 210.45 90.16 ;
    RECT 210.24 90.45 210.45 90.52 ;
    RECT 210.24 90.81 210.45 90.88 ;
    RECT 209.78 90.09 209.99 90.16 ;
    RECT 209.78 90.45 209.99 90.52 ;
    RECT 209.78 90.81 209.99 90.88 ;
    RECT 206.92 90.09 207.13 90.16 ;
    RECT 206.92 90.45 207.13 90.52 ;
    RECT 206.92 90.81 207.13 90.88 ;
    RECT 206.46 90.09 206.67 90.16 ;
    RECT 206.46 90.45 206.67 90.52 ;
    RECT 206.46 90.81 206.67 90.88 ;
    RECT 203.6 90.09 203.81 90.16 ;
    RECT 203.6 90.45 203.81 90.52 ;
    RECT 203.6 90.81 203.81 90.88 ;
    RECT 203.14 90.09 203.35 90.16 ;
    RECT 203.14 90.45 203.35 90.52 ;
    RECT 203.14 90.81 203.35 90.88 ;
    RECT 200.28 90.09 200.49 90.16 ;
    RECT 200.28 90.45 200.49 90.52 ;
    RECT 200.28 90.81 200.49 90.88 ;
    RECT 199.82 90.09 200.03 90.16 ;
    RECT 199.82 90.45 200.03 90.52 ;
    RECT 199.82 90.81 200.03 90.88 ;
    RECT 196.96 90.09 197.17 90.16 ;
    RECT 196.96 90.45 197.17 90.52 ;
    RECT 196.96 90.81 197.17 90.88 ;
    RECT 196.5 90.09 196.71 90.16 ;
    RECT 196.5 90.45 196.71 90.52 ;
    RECT 196.5 90.81 196.71 90.88 ;
    RECT 193.64 90.09 193.85 90.16 ;
    RECT 193.64 90.45 193.85 90.52 ;
    RECT 193.64 90.81 193.85 90.88 ;
    RECT 193.18 90.09 193.39 90.16 ;
    RECT 193.18 90.45 193.39 90.52 ;
    RECT 193.18 90.81 193.39 90.88 ;
    RECT 190.32 90.09 190.53 90.16 ;
    RECT 190.32 90.45 190.53 90.52 ;
    RECT 190.32 90.81 190.53 90.88 ;
    RECT 189.86 90.09 190.07 90.16 ;
    RECT 189.86 90.45 190.07 90.52 ;
    RECT 189.86 90.81 190.07 90.88 ;
    RECT 187.0 90.09 187.21 90.16 ;
    RECT 187.0 90.45 187.21 90.52 ;
    RECT 187.0 90.81 187.21 90.88 ;
    RECT 186.54 90.09 186.75 90.16 ;
    RECT 186.54 90.45 186.75 90.52 ;
    RECT 186.54 90.81 186.75 90.88 ;
    RECT 183.68 90.09 183.89 90.16 ;
    RECT 183.68 90.45 183.89 90.52 ;
    RECT 183.68 90.81 183.89 90.88 ;
    RECT 183.22 90.09 183.43 90.16 ;
    RECT 183.22 90.45 183.43 90.52 ;
    RECT 183.22 90.81 183.43 90.88 ;
    RECT 147.485 90.45 147.555 90.52 ;
    RECT 266.68 90.09 266.89 90.16 ;
    RECT 266.68 90.45 266.89 90.52 ;
    RECT 266.68 90.81 266.89 90.88 ;
    RECT 266.22 90.09 266.43 90.16 ;
    RECT 266.22 90.45 266.43 90.52 ;
    RECT 266.22 90.81 266.43 90.88 ;
    RECT 263.36 90.09 263.57 90.16 ;
    RECT 263.36 90.45 263.57 90.52 ;
    RECT 263.36 90.81 263.57 90.88 ;
    RECT 262.9 90.09 263.11 90.16 ;
    RECT 262.9 90.45 263.11 90.52 ;
    RECT 262.9 90.81 263.11 90.88 ;
    RECT 260.04 90.09 260.25 90.16 ;
    RECT 260.04 90.45 260.25 90.52 ;
    RECT 260.04 90.81 260.25 90.88 ;
    RECT 259.58 90.09 259.79 90.16 ;
    RECT 259.58 90.45 259.79 90.52 ;
    RECT 259.58 90.81 259.79 90.88 ;
    RECT 256.72 90.09 256.93 90.16 ;
    RECT 256.72 90.45 256.93 90.52 ;
    RECT 256.72 90.81 256.93 90.88 ;
    RECT 256.26 90.09 256.47 90.16 ;
    RECT 256.26 90.45 256.47 90.52 ;
    RECT 256.26 90.81 256.47 90.88 ;
    RECT 253.4 90.09 253.61 90.16 ;
    RECT 253.4 90.45 253.61 90.52 ;
    RECT 253.4 90.81 253.61 90.88 ;
    RECT 252.94 90.09 253.15 90.16 ;
    RECT 252.94 90.45 253.15 90.52 ;
    RECT 252.94 90.81 253.15 90.88 ;
    RECT 250.08 53.35 250.29 53.42 ;
    RECT 250.08 53.71 250.29 53.78 ;
    RECT 250.08 54.07 250.29 54.14 ;
    RECT 249.62 53.35 249.83 53.42 ;
    RECT 249.62 53.71 249.83 53.78 ;
    RECT 249.62 54.07 249.83 54.14 ;
    RECT 246.76 53.35 246.97 53.42 ;
    RECT 246.76 53.71 246.97 53.78 ;
    RECT 246.76 54.07 246.97 54.14 ;
    RECT 246.3 53.35 246.51 53.42 ;
    RECT 246.3 53.71 246.51 53.78 ;
    RECT 246.3 54.07 246.51 54.14 ;
    RECT 243.44 53.35 243.65 53.42 ;
    RECT 243.44 53.71 243.65 53.78 ;
    RECT 243.44 54.07 243.65 54.14 ;
    RECT 242.98 53.35 243.19 53.42 ;
    RECT 242.98 53.71 243.19 53.78 ;
    RECT 242.98 54.07 243.19 54.14 ;
    RECT 240.12 53.35 240.33 53.42 ;
    RECT 240.12 53.71 240.33 53.78 ;
    RECT 240.12 54.07 240.33 54.14 ;
    RECT 239.66 53.35 239.87 53.42 ;
    RECT 239.66 53.71 239.87 53.78 ;
    RECT 239.66 54.07 239.87 54.14 ;
    RECT 236.8 53.35 237.01 53.42 ;
    RECT 236.8 53.71 237.01 53.78 ;
    RECT 236.8 54.07 237.01 54.14 ;
    RECT 236.34 53.35 236.55 53.42 ;
    RECT 236.34 53.71 236.55 53.78 ;
    RECT 236.34 54.07 236.55 54.14 ;
    RECT 233.48 53.35 233.69 53.42 ;
    RECT 233.48 53.71 233.69 53.78 ;
    RECT 233.48 54.07 233.69 54.14 ;
    RECT 233.02 53.35 233.23 53.42 ;
    RECT 233.02 53.71 233.23 53.78 ;
    RECT 233.02 54.07 233.23 54.14 ;
    RECT 230.16 53.35 230.37 53.42 ;
    RECT 230.16 53.71 230.37 53.78 ;
    RECT 230.16 54.07 230.37 54.14 ;
    RECT 229.7 53.35 229.91 53.42 ;
    RECT 229.7 53.71 229.91 53.78 ;
    RECT 229.7 54.07 229.91 54.14 ;
    RECT 226.84 53.35 227.05 53.42 ;
    RECT 226.84 53.71 227.05 53.78 ;
    RECT 226.84 54.07 227.05 54.14 ;
    RECT 226.38 53.35 226.59 53.42 ;
    RECT 226.38 53.71 226.59 53.78 ;
    RECT 226.38 54.07 226.59 54.14 ;
    RECT 223.52 53.35 223.73 53.42 ;
    RECT 223.52 53.71 223.73 53.78 ;
    RECT 223.52 54.07 223.73 54.14 ;
    RECT 223.06 53.35 223.27 53.42 ;
    RECT 223.06 53.71 223.27 53.78 ;
    RECT 223.06 54.07 223.27 54.14 ;
    RECT 220.2 53.35 220.41 53.42 ;
    RECT 220.2 53.71 220.41 53.78 ;
    RECT 220.2 54.07 220.41 54.14 ;
    RECT 219.74 53.35 219.95 53.42 ;
    RECT 219.74 53.71 219.95 53.78 ;
    RECT 219.74 54.07 219.95 54.14 ;
    RECT 216.88 53.35 217.09 53.42 ;
    RECT 216.88 53.71 217.09 53.78 ;
    RECT 216.88 54.07 217.09 54.14 ;
    RECT 216.42 53.35 216.63 53.42 ;
    RECT 216.42 53.71 216.63 53.78 ;
    RECT 216.42 54.07 216.63 54.14 ;
    RECT 267.91 53.71 267.98 53.78 ;
    RECT 180.36 53.35 180.57 53.42 ;
    RECT 180.36 53.71 180.57 53.78 ;
    RECT 180.36 54.07 180.57 54.14 ;
    RECT 179.9 53.35 180.11 53.42 ;
    RECT 179.9 53.71 180.11 53.78 ;
    RECT 179.9 54.07 180.11 54.14 ;
    RECT 177.04 53.35 177.25 53.42 ;
    RECT 177.04 53.71 177.25 53.78 ;
    RECT 177.04 54.07 177.25 54.14 ;
    RECT 176.58 53.35 176.79 53.42 ;
    RECT 176.58 53.71 176.79 53.78 ;
    RECT 176.58 54.07 176.79 54.14 ;
    RECT 173.72 53.35 173.93 53.42 ;
    RECT 173.72 53.71 173.93 53.78 ;
    RECT 173.72 54.07 173.93 54.14 ;
    RECT 173.26 53.35 173.47 53.42 ;
    RECT 173.26 53.71 173.47 53.78 ;
    RECT 173.26 54.07 173.47 54.14 ;
    RECT 170.4 53.35 170.61 53.42 ;
    RECT 170.4 53.71 170.61 53.78 ;
    RECT 170.4 54.07 170.61 54.14 ;
    RECT 169.94 53.35 170.15 53.42 ;
    RECT 169.94 53.71 170.15 53.78 ;
    RECT 169.94 54.07 170.15 54.14 ;
    RECT 167.08 53.35 167.29 53.42 ;
    RECT 167.08 53.71 167.29 53.78 ;
    RECT 167.08 54.07 167.29 54.14 ;
    RECT 166.62 53.35 166.83 53.42 ;
    RECT 166.62 53.71 166.83 53.78 ;
    RECT 166.62 54.07 166.83 54.14 ;
    RECT 163.76 53.35 163.97 53.42 ;
    RECT 163.76 53.71 163.97 53.78 ;
    RECT 163.76 54.07 163.97 54.14 ;
    RECT 163.3 53.35 163.51 53.42 ;
    RECT 163.3 53.71 163.51 53.78 ;
    RECT 163.3 54.07 163.51 54.14 ;
    RECT 160.44 53.35 160.65 53.42 ;
    RECT 160.44 53.71 160.65 53.78 ;
    RECT 160.44 54.07 160.65 54.14 ;
    RECT 159.98 53.35 160.19 53.42 ;
    RECT 159.98 53.71 160.19 53.78 ;
    RECT 159.98 54.07 160.19 54.14 ;
    RECT 157.12 53.35 157.33 53.42 ;
    RECT 157.12 53.71 157.33 53.78 ;
    RECT 157.12 54.07 157.33 54.14 ;
    RECT 156.66 53.35 156.87 53.42 ;
    RECT 156.66 53.71 156.87 53.78 ;
    RECT 156.66 54.07 156.87 54.14 ;
    RECT 153.8 53.35 154.01 53.42 ;
    RECT 153.8 53.71 154.01 53.78 ;
    RECT 153.8 54.07 154.01 54.14 ;
    RECT 153.34 53.35 153.55 53.42 ;
    RECT 153.34 53.71 153.55 53.78 ;
    RECT 153.34 54.07 153.55 54.14 ;
    RECT 150.48 53.35 150.69 53.42 ;
    RECT 150.48 53.71 150.69 53.78 ;
    RECT 150.48 54.07 150.69 54.14 ;
    RECT 150.02 53.35 150.23 53.42 ;
    RECT 150.02 53.71 150.23 53.78 ;
    RECT 150.02 54.07 150.23 54.14 ;
    RECT 213.56 53.35 213.77 53.42 ;
    RECT 213.56 53.71 213.77 53.78 ;
    RECT 213.56 54.07 213.77 54.14 ;
    RECT 213.1 53.35 213.31 53.42 ;
    RECT 213.1 53.71 213.31 53.78 ;
    RECT 213.1 54.07 213.31 54.14 ;
    RECT 210.24 53.35 210.45 53.42 ;
    RECT 210.24 53.71 210.45 53.78 ;
    RECT 210.24 54.07 210.45 54.14 ;
    RECT 209.78 53.35 209.99 53.42 ;
    RECT 209.78 53.71 209.99 53.78 ;
    RECT 209.78 54.07 209.99 54.14 ;
    RECT 206.92 53.35 207.13 53.42 ;
    RECT 206.92 53.71 207.13 53.78 ;
    RECT 206.92 54.07 207.13 54.14 ;
    RECT 206.46 53.35 206.67 53.42 ;
    RECT 206.46 53.71 206.67 53.78 ;
    RECT 206.46 54.07 206.67 54.14 ;
    RECT 203.6 53.35 203.81 53.42 ;
    RECT 203.6 53.71 203.81 53.78 ;
    RECT 203.6 54.07 203.81 54.14 ;
    RECT 203.14 53.35 203.35 53.42 ;
    RECT 203.14 53.71 203.35 53.78 ;
    RECT 203.14 54.07 203.35 54.14 ;
    RECT 200.28 53.35 200.49 53.42 ;
    RECT 200.28 53.71 200.49 53.78 ;
    RECT 200.28 54.07 200.49 54.14 ;
    RECT 199.82 53.35 200.03 53.42 ;
    RECT 199.82 53.71 200.03 53.78 ;
    RECT 199.82 54.07 200.03 54.14 ;
    RECT 196.96 53.35 197.17 53.42 ;
    RECT 196.96 53.71 197.17 53.78 ;
    RECT 196.96 54.07 197.17 54.14 ;
    RECT 196.5 53.35 196.71 53.42 ;
    RECT 196.5 53.71 196.71 53.78 ;
    RECT 196.5 54.07 196.71 54.14 ;
    RECT 193.64 53.35 193.85 53.42 ;
    RECT 193.64 53.71 193.85 53.78 ;
    RECT 193.64 54.07 193.85 54.14 ;
    RECT 193.18 53.35 193.39 53.42 ;
    RECT 193.18 53.71 193.39 53.78 ;
    RECT 193.18 54.07 193.39 54.14 ;
    RECT 190.32 53.35 190.53 53.42 ;
    RECT 190.32 53.71 190.53 53.78 ;
    RECT 190.32 54.07 190.53 54.14 ;
    RECT 189.86 53.35 190.07 53.42 ;
    RECT 189.86 53.71 190.07 53.78 ;
    RECT 189.86 54.07 190.07 54.14 ;
    RECT 187.0 53.35 187.21 53.42 ;
    RECT 187.0 53.71 187.21 53.78 ;
    RECT 187.0 54.07 187.21 54.14 ;
    RECT 186.54 53.35 186.75 53.42 ;
    RECT 186.54 53.71 186.75 53.78 ;
    RECT 186.54 54.07 186.75 54.14 ;
    RECT 183.68 53.35 183.89 53.42 ;
    RECT 183.68 53.71 183.89 53.78 ;
    RECT 183.68 54.07 183.89 54.14 ;
    RECT 183.22 53.35 183.43 53.42 ;
    RECT 183.22 53.71 183.43 53.78 ;
    RECT 183.22 54.07 183.43 54.14 ;
    RECT 147.485 53.71 147.555 53.78 ;
    RECT 266.68 53.35 266.89 53.42 ;
    RECT 266.68 53.71 266.89 53.78 ;
    RECT 266.68 54.07 266.89 54.14 ;
    RECT 266.22 53.35 266.43 53.42 ;
    RECT 266.22 53.71 266.43 53.78 ;
    RECT 266.22 54.07 266.43 54.14 ;
    RECT 263.36 53.35 263.57 53.42 ;
    RECT 263.36 53.71 263.57 53.78 ;
    RECT 263.36 54.07 263.57 54.14 ;
    RECT 262.9 53.35 263.11 53.42 ;
    RECT 262.9 53.71 263.11 53.78 ;
    RECT 262.9 54.07 263.11 54.14 ;
    RECT 260.04 53.35 260.25 53.42 ;
    RECT 260.04 53.71 260.25 53.78 ;
    RECT 260.04 54.07 260.25 54.14 ;
    RECT 259.58 53.35 259.79 53.42 ;
    RECT 259.58 53.71 259.79 53.78 ;
    RECT 259.58 54.07 259.79 54.14 ;
    RECT 256.72 53.35 256.93 53.42 ;
    RECT 256.72 53.71 256.93 53.78 ;
    RECT 256.72 54.07 256.93 54.14 ;
    RECT 256.26 53.35 256.47 53.42 ;
    RECT 256.26 53.71 256.47 53.78 ;
    RECT 256.26 54.07 256.47 54.14 ;
    RECT 253.4 53.35 253.61 53.42 ;
    RECT 253.4 53.71 253.61 53.78 ;
    RECT 253.4 54.07 253.61 54.14 ;
    RECT 252.94 53.35 253.15 53.42 ;
    RECT 252.94 53.71 253.15 53.78 ;
    RECT 252.94 54.07 253.15 54.14 ;
    RECT 250.08 14.47 250.29 14.54 ;
    RECT 250.08 14.83 250.29 14.9 ;
    RECT 250.08 15.19 250.29 15.26 ;
    RECT 249.62 14.47 249.83 14.54 ;
    RECT 249.62 14.83 249.83 14.9 ;
    RECT 249.62 15.19 249.83 15.26 ;
    RECT 147.485 14.83 147.555 14.9 ;
    RECT 246.76 14.47 246.97 14.54 ;
    RECT 246.76 14.83 246.97 14.9 ;
    RECT 246.76 15.19 246.97 15.26 ;
    RECT 246.3 14.47 246.51 14.54 ;
    RECT 246.3 14.83 246.51 14.9 ;
    RECT 246.3 15.19 246.51 15.26 ;
    RECT 243.44 14.47 243.65 14.54 ;
    RECT 243.44 14.83 243.65 14.9 ;
    RECT 243.44 15.19 243.65 15.26 ;
    RECT 242.98 14.47 243.19 14.54 ;
    RECT 242.98 14.83 243.19 14.9 ;
    RECT 242.98 15.19 243.19 15.26 ;
    RECT 240.12 14.47 240.33 14.54 ;
    RECT 240.12 14.83 240.33 14.9 ;
    RECT 240.12 15.19 240.33 15.26 ;
    RECT 239.66 14.47 239.87 14.54 ;
    RECT 239.66 14.83 239.87 14.9 ;
    RECT 239.66 15.19 239.87 15.26 ;
    RECT 236.8 14.47 237.01 14.54 ;
    RECT 236.8 14.83 237.01 14.9 ;
    RECT 236.8 15.19 237.01 15.26 ;
    RECT 236.34 14.47 236.55 14.54 ;
    RECT 236.34 14.83 236.55 14.9 ;
    RECT 236.34 15.19 236.55 15.26 ;
    RECT 233.48 14.47 233.69 14.54 ;
    RECT 233.48 14.83 233.69 14.9 ;
    RECT 233.48 15.19 233.69 15.26 ;
    RECT 233.02 14.47 233.23 14.54 ;
    RECT 233.02 14.83 233.23 14.9 ;
    RECT 233.02 15.19 233.23 15.26 ;
    RECT 230.16 14.47 230.37 14.54 ;
    RECT 230.16 14.83 230.37 14.9 ;
    RECT 230.16 15.19 230.37 15.26 ;
    RECT 229.7 14.47 229.91 14.54 ;
    RECT 229.7 14.83 229.91 14.9 ;
    RECT 229.7 15.19 229.91 15.26 ;
    RECT 226.84 14.47 227.05 14.54 ;
    RECT 226.84 14.83 227.05 14.9 ;
    RECT 226.84 15.19 227.05 15.26 ;
    RECT 226.38 14.47 226.59 14.54 ;
    RECT 226.38 14.83 226.59 14.9 ;
    RECT 226.38 15.19 226.59 15.26 ;
    RECT 223.52 14.47 223.73 14.54 ;
    RECT 223.52 14.83 223.73 14.9 ;
    RECT 223.52 15.19 223.73 15.26 ;
    RECT 223.06 14.47 223.27 14.54 ;
    RECT 223.06 14.83 223.27 14.9 ;
    RECT 223.06 15.19 223.27 15.26 ;
    RECT 220.2 14.47 220.41 14.54 ;
    RECT 220.2 14.83 220.41 14.9 ;
    RECT 220.2 15.19 220.41 15.26 ;
    RECT 219.74 14.47 219.95 14.54 ;
    RECT 219.74 14.83 219.95 14.9 ;
    RECT 219.74 15.19 219.95 15.26 ;
    RECT 216.88 14.47 217.09 14.54 ;
    RECT 216.88 14.83 217.09 14.9 ;
    RECT 216.88 15.19 217.09 15.26 ;
    RECT 216.42 14.47 216.63 14.54 ;
    RECT 216.42 14.83 216.63 14.9 ;
    RECT 216.42 15.19 216.63 15.26 ;
    RECT 180.36 14.47 180.57 14.54 ;
    RECT 180.36 14.83 180.57 14.9 ;
    RECT 180.36 15.19 180.57 15.26 ;
    RECT 179.9 14.47 180.11 14.54 ;
    RECT 179.9 14.83 180.11 14.9 ;
    RECT 179.9 15.19 180.11 15.26 ;
    RECT 177.04 14.47 177.25 14.54 ;
    RECT 177.04 14.83 177.25 14.9 ;
    RECT 177.04 15.19 177.25 15.26 ;
    RECT 176.58 14.47 176.79 14.54 ;
    RECT 176.58 14.83 176.79 14.9 ;
    RECT 176.58 15.19 176.79 15.26 ;
    RECT 173.72 14.47 173.93 14.54 ;
    RECT 173.72 14.83 173.93 14.9 ;
    RECT 173.72 15.19 173.93 15.26 ;
    RECT 173.26 14.47 173.47 14.54 ;
    RECT 173.26 14.83 173.47 14.9 ;
    RECT 173.26 15.19 173.47 15.26 ;
    RECT 267.91 14.83 267.98 14.9 ;
    RECT 170.4 14.47 170.61 14.54 ;
    RECT 170.4 14.83 170.61 14.9 ;
    RECT 170.4 15.19 170.61 15.26 ;
    RECT 169.94 14.47 170.15 14.54 ;
    RECT 169.94 14.83 170.15 14.9 ;
    RECT 169.94 15.19 170.15 15.26 ;
    RECT 167.08 14.47 167.29 14.54 ;
    RECT 167.08 14.83 167.29 14.9 ;
    RECT 167.08 15.19 167.29 15.26 ;
    RECT 166.62 14.47 166.83 14.54 ;
    RECT 166.62 14.83 166.83 14.9 ;
    RECT 166.62 15.19 166.83 15.26 ;
    RECT 163.76 14.47 163.97 14.54 ;
    RECT 163.76 14.83 163.97 14.9 ;
    RECT 163.76 15.19 163.97 15.26 ;
    RECT 163.3 14.47 163.51 14.54 ;
    RECT 163.3 14.83 163.51 14.9 ;
    RECT 163.3 15.19 163.51 15.26 ;
    RECT 160.44 14.47 160.65 14.54 ;
    RECT 160.44 14.83 160.65 14.9 ;
    RECT 160.44 15.19 160.65 15.26 ;
    RECT 159.98 14.47 160.19 14.54 ;
    RECT 159.98 14.83 160.19 14.9 ;
    RECT 159.98 15.19 160.19 15.26 ;
    RECT 157.12 14.47 157.33 14.54 ;
    RECT 157.12 14.83 157.33 14.9 ;
    RECT 157.12 15.19 157.33 15.26 ;
    RECT 156.66 14.47 156.87 14.54 ;
    RECT 156.66 14.83 156.87 14.9 ;
    RECT 156.66 15.19 156.87 15.26 ;
    RECT 153.8 14.47 154.01 14.54 ;
    RECT 153.8 14.83 154.01 14.9 ;
    RECT 153.8 15.19 154.01 15.26 ;
    RECT 153.34 14.47 153.55 14.54 ;
    RECT 153.34 14.83 153.55 14.9 ;
    RECT 153.34 15.19 153.55 15.26 ;
    RECT 213.56 14.47 213.77 14.54 ;
    RECT 213.56 14.83 213.77 14.9 ;
    RECT 213.56 15.19 213.77 15.26 ;
    RECT 213.1 14.47 213.31 14.54 ;
    RECT 213.1 14.83 213.31 14.9 ;
    RECT 213.1 15.19 213.31 15.26 ;
    RECT 210.24 14.47 210.45 14.54 ;
    RECT 210.24 14.83 210.45 14.9 ;
    RECT 210.24 15.19 210.45 15.26 ;
    RECT 209.78 14.47 209.99 14.54 ;
    RECT 209.78 14.83 209.99 14.9 ;
    RECT 209.78 15.19 209.99 15.26 ;
    RECT 266.68 14.47 266.89 14.54 ;
    RECT 266.68 14.83 266.89 14.9 ;
    RECT 266.68 15.19 266.89 15.26 ;
    RECT 266.22 14.47 266.43 14.54 ;
    RECT 266.22 14.83 266.43 14.9 ;
    RECT 266.22 15.19 266.43 15.26 ;
    RECT 206.92 14.47 207.13 14.54 ;
    RECT 206.92 14.83 207.13 14.9 ;
    RECT 206.92 15.19 207.13 15.26 ;
    RECT 206.46 14.47 206.67 14.54 ;
    RECT 206.46 14.83 206.67 14.9 ;
    RECT 206.46 15.19 206.67 15.26 ;
    RECT 203.6 14.47 203.81 14.54 ;
    RECT 203.6 14.83 203.81 14.9 ;
    RECT 203.6 15.19 203.81 15.26 ;
    RECT 203.14 14.47 203.35 14.54 ;
    RECT 203.14 14.83 203.35 14.9 ;
    RECT 203.14 15.19 203.35 15.26 ;
    RECT 200.28 14.47 200.49 14.54 ;
    RECT 200.28 14.83 200.49 14.9 ;
    RECT 200.28 15.19 200.49 15.26 ;
    RECT 199.82 14.47 200.03 14.54 ;
    RECT 199.82 14.83 200.03 14.9 ;
    RECT 199.82 15.19 200.03 15.26 ;
    RECT 196.96 14.47 197.17 14.54 ;
    RECT 196.96 14.83 197.17 14.9 ;
    RECT 196.96 15.19 197.17 15.26 ;
    RECT 196.5 14.47 196.71 14.54 ;
    RECT 196.5 14.83 196.71 14.9 ;
    RECT 196.5 15.19 196.71 15.26 ;
    RECT 193.64 14.47 193.85 14.54 ;
    RECT 193.64 14.83 193.85 14.9 ;
    RECT 193.64 15.19 193.85 15.26 ;
    RECT 193.18 14.47 193.39 14.54 ;
    RECT 193.18 14.83 193.39 14.9 ;
    RECT 193.18 15.19 193.39 15.26 ;
    RECT 190.32 14.47 190.53 14.54 ;
    RECT 190.32 14.83 190.53 14.9 ;
    RECT 190.32 15.19 190.53 15.26 ;
    RECT 189.86 14.47 190.07 14.54 ;
    RECT 189.86 14.83 190.07 14.9 ;
    RECT 189.86 15.19 190.07 15.26 ;
    RECT 150.48 14.47 150.69 14.54 ;
    RECT 150.48 14.83 150.69 14.9 ;
    RECT 150.48 15.19 150.69 15.26 ;
    RECT 150.02 14.47 150.23 14.54 ;
    RECT 150.02 14.83 150.23 14.9 ;
    RECT 150.02 15.19 150.23 15.26 ;
    RECT 187.0 14.47 187.21 14.54 ;
    RECT 187.0 14.83 187.21 14.9 ;
    RECT 187.0 15.19 187.21 15.26 ;
    RECT 186.54 14.47 186.75 14.54 ;
    RECT 186.54 14.83 186.75 14.9 ;
    RECT 186.54 15.19 186.75 15.26 ;
    RECT 183.68 14.47 183.89 14.54 ;
    RECT 183.68 14.83 183.89 14.9 ;
    RECT 183.68 15.19 183.89 15.26 ;
    RECT 183.22 14.47 183.43 14.54 ;
    RECT 183.22 14.83 183.43 14.9 ;
    RECT 183.22 15.19 183.43 15.26 ;
    RECT 263.36 14.47 263.57 14.54 ;
    RECT 263.36 14.83 263.57 14.9 ;
    RECT 263.36 15.19 263.57 15.26 ;
    RECT 262.9 14.47 263.11 14.54 ;
    RECT 262.9 14.83 263.11 14.9 ;
    RECT 262.9 15.19 263.11 15.26 ;
    RECT 260.04 14.47 260.25 14.54 ;
    RECT 260.04 14.83 260.25 14.9 ;
    RECT 260.04 15.19 260.25 15.26 ;
    RECT 259.58 14.47 259.79 14.54 ;
    RECT 259.58 14.83 259.79 14.9 ;
    RECT 259.58 15.19 259.79 15.26 ;
    RECT 256.72 14.47 256.93 14.54 ;
    RECT 256.72 14.83 256.93 14.9 ;
    RECT 256.72 15.19 256.93 15.26 ;
    RECT 256.26 14.47 256.47 14.54 ;
    RECT 256.26 14.83 256.47 14.9 ;
    RECT 256.26 15.19 256.47 15.26 ;
    RECT 253.4 14.47 253.61 14.54 ;
    RECT 253.4 14.83 253.61 14.9 ;
    RECT 253.4 15.19 253.61 15.26 ;
    RECT 252.94 14.47 253.15 14.54 ;
    RECT 252.94 14.83 253.15 14.9 ;
    RECT 252.94 15.19 253.15 15.26 ;
    RECT 250.08 89.37 250.29 89.44 ;
    RECT 250.08 89.73 250.29 89.8 ;
    RECT 250.08 90.09 250.29 90.16 ;
    RECT 249.62 89.37 249.83 89.44 ;
    RECT 249.62 89.73 249.83 89.8 ;
    RECT 249.62 90.09 249.83 90.16 ;
    RECT 246.76 89.37 246.97 89.44 ;
    RECT 246.76 89.73 246.97 89.8 ;
    RECT 246.76 90.09 246.97 90.16 ;
    RECT 246.3 89.37 246.51 89.44 ;
    RECT 246.3 89.73 246.51 89.8 ;
    RECT 246.3 90.09 246.51 90.16 ;
    RECT 243.44 89.37 243.65 89.44 ;
    RECT 243.44 89.73 243.65 89.8 ;
    RECT 243.44 90.09 243.65 90.16 ;
    RECT 242.98 89.37 243.19 89.44 ;
    RECT 242.98 89.73 243.19 89.8 ;
    RECT 242.98 90.09 243.19 90.16 ;
    RECT 240.12 89.37 240.33 89.44 ;
    RECT 240.12 89.73 240.33 89.8 ;
    RECT 240.12 90.09 240.33 90.16 ;
    RECT 239.66 89.37 239.87 89.44 ;
    RECT 239.66 89.73 239.87 89.8 ;
    RECT 239.66 90.09 239.87 90.16 ;
    RECT 236.8 89.37 237.01 89.44 ;
    RECT 236.8 89.73 237.01 89.8 ;
    RECT 236.8 90.09 237.01 90.16 ;
    RECT 236.34 89.37 236.55 89.44 ;
    RECT 236.34 89.73 236.55 89.8 ;
    RECT 236.34 90.09 236.55 90.16 ;
    RECT 233.48 89.37 233.69 89.44 ;
    RECT 233.48 89.73 233.69 89.8 ;
    RECT 233.48 90.09 233.69 90.16 ;
    RECT 233.02 89.37 233.23 89.44 ;
    RECT 233.02 89.73 233.23 89.8 ;
    RECT 233.02 90.09 233.23 90.16 ;
    RECT 230.16 89.37 230.37 89.44 ;
    RECT 230.16 89.73 230.37 89.8 ;
    RECT 230.16 90.09 230.37 90.16 ;
    RECT 229.7 89.37 229.91 89.44 ;
    RECT 229.7 89.73 229.91 89.8 ;
    RECT 229.7 90.09 229.91 90.16 ;
    RECT 226.84 89.37 227.05 89.44 ;
    RECT 226.84 89.73 227.05 89.8 ;
    RECT 226.84 90.09 227.05 90.16 ;
    RECT 226.38 89.37 226.59 89.44 ;
    RECT 226.38 89.73 226.59 89.8 ;
    RECT 226.38 90.09 226.59 90.16 ;
    RECT 223.52 89.37 223.73 89.44 ;
    RECT 223.52 89.73 223.73 89.8 ;
    RECT 223.52 90.09 223.73 90.16 ;
    RECT 223.06 89.37 223.27 89.44 ;
    RECT 223.06 89.73 223.27 89.8 ;
    RECT 223.06 90.09 223.27 90.16 ;
    RECT 220.2 89.37 220.41 89.44 ;
    RECT 220.2 89.73 220.41 89.8 ;
    RECT 220.2 90.09 220.41 90.16 ;
    RECT 219.74 89.37 219.95 89.44 ;
    RECT 219.74 89.73 219.95 89.8 ;
    RECT 219.74 90.09 219.95 90.16 ;
    RECT 216.88 89.37 217.09 89.44 ;
    RECT 216.88 89.73 217.09 89.8 ;
    RECT 216.88 90.09 217.09 90.16 ;
    RECT 216.42 89.37 216.63 89.44 ;
    RECT 216.42 89.73 216.63 89.8 ;
    RECT 216.42 90.09 216.63 90.16 ;
    RECT 267.91 89.73 267.98 89.8 ;
    RECT 180.36 89.37 180.57 89.44 ;
    RECT 180.36 89.73 180.57 89.8 ;
    RECT 180.36 90.09 180.57 90.16 ;
    RECT 179.9 89.37 180.11 89.44 ;
    RECT 179.9 89.73 180.11 89.8 ;
    RECT 179.9 90.09 180.11 90.16 ;
    RECT 177.04 89.37 177.25 89.44 ;
    RECT 177.04 89.73 177.25 89.8 ;
    RECT 177.04 90.09 177.25 90.16 ;
    RECT 176.58 89.37 176.79 89.44 ;
    RECT 176.58 89.73 176.79 89.8 ;
    RECT 176.58 90.09 176.79 90.16 ;
    RECT 173.72 89.37 173.93 89.44 ;
    RECT 173.72 89.73 173.93 89.8 ;
    RECT 173.72 90.09 173.93 90.16 ;
    RECT 173.26 89.37 173.47 89.44 ;
    RECT 173.26 89.73 173.47 89.8 ;
    RECT 173.26 90.09 173.47 90.16 ;
    RECT 170.4 89.37 170.61 89.44 ;
    RECT 170.4 89.73 170.61 89.8 ;
    RECT 170.4 90.09 170.61 90.16 ;
    RECT 169.94 89.37 170.15 89.44 ;
    RECT 169.94 89.73 170.15 89.8 ;
    RECT 169.94 90.09 170.15 90.16 ;
    RECT 167.08 89.37 167.29 89.44 ;
    RECT 167.08 89.73 167.29 89.8 ;
    RECT 167.08 90.09 167.29 90.16 ;
    RECT 166.62 89.37 166.83 89.44 ;
    RECT 166.62 89.73 166.83 89.8 ;
    RECT 166.62 90.09 166.83 90.16 ;
    RECT 163.76 89.37 163.97 89.44 ;
    RECT 163.76 89.73 163.97 89.8 ;
    RECT 163.76 90.09 163.97 90.16 ;
    RECT 163.3 89.37 163.51 89.44 ;
    RECT 163.3 89.73 163.51 89.8 ;
    RECT 163.3 90.09 163.51 90.16 ;
    RECT 160.44 89.37 160.65 89.44 ;
    RECT 160.44 89.73 160.65 89.8 ;
    RECT 160.44 90.09 160.65 90.16 ;
    RECT 159.98 89.37 160.19 89.44 ;
    RECT 159.98 89.73 160.19 89.8 ;
    RECT 159.98 90.09 160.19 90.16 ;
    RECT 157.12 89.37 157.33 89.44 ;
    RECT 157.12 89.73 157.33 89.8 ;
    RECT 157.12 90.09 157.33 90.16 ;
    RECT 156.66 89.37 156.87 89.44 ;
    RECT 156.66 89.73 156.87 89.8 ;
    RECT 156.66 90.09 156.87 90.16 ;
    RECT 153.8 89.37 154.01 89.44 ;
    RECT 153.8 89.73 154.01 89.8 ;
    RECT 153.8 90.09 154.01 90.16 ;
    RECT 153.34 89.37 153.55 89.44 ;
    RECT 153.34 89.73 153.55 89.8 ;
    RECT 153.34 90.09 153.55 90.16 ;
    RECT 150.48 89.37 150.69 89.44 ;
    RECT 150.48 89.73 150.69 89.8 ;
    RECT 150.48 90.09 150.69 90.16 ;
    RECT 150.02 89.37 150.23 89.44 ;
    RECT 150.02 89.73 150.23 89.8 ;
    RECT 150.02 90.09 150.23 90.16 ;
    RECT 213.56 89.37 213.77 89.44 ;
    RECT 213.56 89.73 213.77 89.8 ;
    RECT 213.56 90.09 213.77 90.16 ;
    RECT 213.1 89.37 213.31 89.44 ;
    RECT 213.1 89.73 213.31 89.8 ;
    RECT 213.1 90.09 213.31 90.16 ;
    RECT 210.24 89.37 210.45 89.44 ;
    RECT 210.24 89.73 210.45 89.8 ;
    RECT 210.24 90.09 210.45 90.16 ;
    RECT 209.78 89.37 209.99 89.44 ;
    RECT 209.78 89.73 209.99 89.8 ;
    RECT 209.78 90.09 209.99 90.16 ;
    RECT 206.92 89.37 207.13 89.44 ;
    RECT 206.92 89.73 207.13 89.8 ;
    RECT 206.92 90.09 207.13 90.16 ;
    RECT 206.46 89.37 206.67 89.44 ;
    RECT 206.46 89.73 206.67 89.8 ;
    RECT 206.46 90.09 206.67 90.16 ;
    RECT 203.6 89.37 203.81 89.44 ;
    RECT 203.6 89.73 203.81 89.8 ;
    RECT 203.6 90.09 203.81 90.16 ;
    RECT 203.14 89.37 203.35 89.44 ;
    RECT 203.14 89.73 203.35 89.8 ;
    RECT 203.14 90.09 203.35 90.16 ;
    RECT 200.28 89.37 200.49 89.44 ;
    RECT 200.28 89.73 200.49 89.8 ;
    RECT 200.28 90.09 200.49 90.16 ;
    RECT 199.82 89.37 200.03 89.44 ;
    RECT 199.82 89.73 200.03 89.8 ;
    RECT 199.82 90.09 200.03 90.16 ;
    RECT 196.96 89.37 197.17 89.44 ;
    RECT 196.96 89.73 197.17 89.8 ;
    RECT 196.96 90.09 197.17 90.16 ;
    RECT 196.5 89.37 196.71 89.44 ;
    RECT 196.5 89.73 196.71 89.8 ;
    RECT 196.5 90.09 196.71 90.16 ;
    RECT 193.64 89.37 193.85 89.44 ;
    RECT 193.64 89.73 193.85 89.8 ;
    RECT 193.64 90.09 193.85 90.16 ;
    RECT 193.18 89.37 193.39 89.44 ;
    RECT 193.18 89.73 193.39 89.8 ;
    RECT 193.18 90.09 193.39 90.16 ;
    RECT 190.32 89.37 190.53 89.44 ;
    RECT 190.32 89.73 190.53 89.8 ;
    RECT 190.32 90.09 190.53 90.16 ;
    RECT 189.86 89.37 190.07 89.44 ;
    RECT 189.86 89.73 190.07 89.8 ;
    RECT 189.86 90.09 190.07 90.16 ;
    RECT 187.0 89.37 187.21 89.44 ;
    RECT 187.0 89.73 187.21 89.8 ;
    RECT 187.0 90.09 187.21 90.16 ;
    RECT 186.54 89.37 186.75 89.44 ;
    RECT 186.54 89.73 186.75 89.8 ;
    RECT 186.54 90.09 186.75 90.16 ;
    RECT 183.68 89.37 183.89 89.44 ;
    RECT 183.68 89.73 183.89 89.8 ;
    RECT 183.68 90.09 183.89 90.16 ;
    RECT 183.22 89.37 183.43 89.44 ;
    RECT 183.22 89.73 183.43 89.8 ;
    RECT 183.22 90.09 183.43 90.16 ;
    RECT 147.485 89.73 147.555 89.8 ;
    RECT 266.68 89.37 266.89 89.44 ;
    RECT 266.68 89.73 266.89 89.8 ;
    RECT 266.68 90.09 266.89 90.16 ;
    RECT 266.22 89.37 266.43 89.44 ;
    RECT 266.22 89.73 266.43 89.8 ;
    RECT 266.22 90.09 266.43 90.16 ;
    RECT 263.36 89.37 263.57 89.44 ;
    RECT 263.36 89.73 263.57 89.8 ;
    RECT 263.36 90.09 263.57 90.16 ;
    RECT 262.9 89.37 263.11 89.44 ;
    RECT 262.9 89.73 263.11 89.8 ;
    RECT 262.9 90.09 263.11 90.16 ;
    RECT 260.04 89.37 260.25 89.44 ;
    RECT 260.04 89.73 260.25 89.8 ;
    RECT 260.04 90.09 260.25 90.16 ;
    RECT 259.58 89.37 259.79 89.44 ;
    RECT 259.58 89.73 259.79 89.8 ;
    RECT 259.58 90.09 259.79 90.16 ;
    RECT 256.72 89.37 256.93 89.44 ;
    RECT 256.72 89.73 256.93 89.8 ;
    RECT 256.72 90.09 256.93 90.16 ;
    RECT 256.26 89.37 256.47 89.44 ;
    RECT 256.26 89.73 256.47 89.8 ;
    RECT 256.26 90.09 256.47 90.16 ;
    RECT 253.4 89.37 253.61 89.44 ;
    RECT 253.4 89.73 253.61 89.8 ;
    RECT 253.4 90.09 253.61 90.16 ;
    RECT 252.94 89.37 253.15 89.44 ;
    RECT 252.94 89.73 253.15 89.8 ;
    RECT 252.94 90.09 253.15 90.16 ;
    RECT 250.08 52.63 250.29 52.7 ;
    RECT 250.08 52.99 250.29 53.06 ;
    RECT 250.08 53.35 250.29 53.42 ;
    RECT 249.62 52.63 249.83 52.7 ;
    RECT 249.62 52.99 249.83 53.06 ;
    RECT 249.62 53.35 249.83 53.42 ;
    RECT 246.76 52.63 246.97 52.7 ;
    RECT 246.76 52.99 246.97 53.06 ;
    RECT 246.76 53.35 246.97 53.42 ;
    RECT 246.3 52.63 246.51 52.7 ;
    RECT 246.3 52.99 246.51 53.06 ;
    RECT 246.3 53.35 246.51 53.42 ;
    RECT 243.44 52.63 243.65 52.7 ;
    RECT 243.44 52.99 243.65 53.06 ;
    RECT 243.44 53.35 243.65 53.42 ;
    RECT 242.98 52.63 243.19 52.7 ;
    RECT 242.98 52.99 243.19 53.06 ;
    RECT 242.98 53.35 243.19 53.42 ;
    RECT 240.12 52.63 240.33 52.7 ;
    RECT 240.12 52.99 240.33 53.06 ;
    RECT 240.12 53.35 240.33 53.42 ;
    RECT 239.66 52.63 239.87 52.7 ;
    RECT 239.66 52.99 239.87 53.06 ;
    RECT 239.66 53.35 239.87 53.42 ;
    RECT 236.8 52.63 237.01 52.7 ;
    RECT 236.8 52.99 237.01 53.06 ;
    RECT 236.8 53.35 237.01 53.42 ;
    RECT 236.34 52.63 236.55 52.7 ;
    RECT 236.34 52.99 236.55 53.06 ;
    RECT 236.34 53.35 236.55 53.42 ;
    RECT 233.48 52.63 233.69 52.7 ;
    RECT 233.48 52.99 233.69 53.06 ;
    RECT 233.48 53.35 233.69 53.42 ;
    RECT 233.02 52.63 233.23 52.7 ;
    RECT 233.02 52.99 233.23 53.06 ;
    RECT 233.02 53.35 233.23 53.42 ;
    RECT 230.16 52.63 230.37 52.7 ;
    RECT 230.16 52.99 230.37 53.06 ;
    RECT 230.16 53.35 230.37 53.42 ;
    RECT 229.7 52.63 229.91 52.7 ;
    RECT 229.7 52.99 229.91 53.06 ;
    RECT 229.7 53.35 229.91 53.42 ;
    RECT 226.84 52.63 227.05 52.7 ;
    RECT 226.84 52.99 227.05 53.06 ;
    RECT 226.84 53.35 227.05 53.42 ;
    RECT 226.38 52.63 226.59 52.7 ;
    RECT 226.38 52.99 226.59 53.06 ;
    RECT 226.38 53.35 226.59 53.42 ;
    RECT 223.52 52.63 223.73 52.7 ;
    RECT 223.52 52.99 223.73 53.06 ;
    RECT 223.52 53.35 223.73 53.42 ;
    RECT 223.06 52.63 223.27 52.7 ;
    RECT 223.06 52.99 223.27 53.06 ;
    RECT 223.06 53.35 223.27 53.42 ;
    RECT 220.2 52.63 220.41 52.7 ;
    RECT 220.2 52.99 220.41 53.06 ;
    RECT 220.2 53.35 220.41 53.42 ;
    RECT 219.74 52.63 219.95 52.7 ;
    RECT 219.74 52.99 219.95 53.06 ;
    RECT 219.74 53.35 219.95 53.42 ;
    RECT 216.88 52.63 217.09 52.7 ;
    RECT 216.88 52.99 217.09 53.06 ;
    RECT 216.88 53.35 217.09 53.42 ;
    RECT 216.42 52.63 216.63 52.7 ;
    RECT 216.42 52.99 216.63 53.06 ;
    RECT 216.42 53.35 216.63 53.42 ;
    RECT 267.91 52.99 267.98 53.06 ;
    RECT 180.36 52.63 180.57 52.7 ;
    RECT 180.36 52.99 180.57 53.06 ;
    RECT 180.36 53.35 180.57 53.42 ;
    RECT 179.9 52.63 180.11 52.7 ;
    RECT 179.9 52.99 180.11 53.06 ;
    RECT 179.9 53.35 180.11 53.42 ;
    RECT 177.04 52.63 177.25 52.7 ;
    RECT 177.04 52.99 177.25 53.06 ;
    RECT 177.04 53.35 177.25 53.42 ;
    RECT 176.58 52.63 176.79 52.7 ;
    RECT 176.58 52.99 176.79 53.06 ;
    RECT 176.58 53.35 176.79 53.42 ;
    RECT 173.72 52.63 173.93 52.7 ;
    RECT 173.72 52.99 173.93 53.06 ;
    RECT 173.72 53.35 173.93 53.42 ;
    RECT 173.26 52.63 173.47 52.7 ;
    RECT 173.26 52.99 173.47 53.06 ;
    RECT 173.26 53.35 173.47 53.42 ;
    RECT 170.4 52.63 170.61 52.7 ;
    RECT 170.4 52.99 170.61 53.06 ;
    RECT 170.4 53.35 170.61 53.42 ;
    RECT 169.94 52.63 170.15 52.7 ;
    RECT 169.94 52.99 170.15 53.06 ;
    RECT 169.94 53.35 170.15 53.42 ;
    RECT 167.08 52.63 167.29 52.7 ;
    RECT 167.08 52.99 167.29 53.06 ;
    RECT 167.08 53.35 167.29 53.42 ;
    RECT 166.62 52.63 166.83 52.7 ;
    RECT 166.62 52.99 166.83 53.06 ;
    RECT 166.62 53.35 166.83 53.42 ;
    RECT 163.76 52.63 163.97 52.7 ;
    RECT 163.76 52.99 163.97 53.06 ;
    RECT 163.76 53.35 163.97 53.42 ;
    RECT 163.3 52.63 163.51 52.7 ;
    RECT 163.3 52.99 163.51 53.06 ;
    RECT 163.3 53.35 163.51 53.42 ;
    RECT 160.44 52.63 160.65 52.7 ;
    RECT 160.44 52.99 160.65 53.06 ;
    RECT 160.44 53.35 160.65 53.42 ;
    RECT 159.98 52.63 160.19 52.7 ;
    RECT 159.98 52.99 160.19 53.06 ;
    RECT 159.98 53.35 160.19 53.42 ;
    RECT 157.12 52.63 157.33 52.7 ;
    RECT 157.12 52.99 157.33 53.06 ;
    RECT 157.12 53.35 157.33 53.42 ;
    RECT 156.66 52.63 156.87 52.7 ;
    RECT 156.66 52.99 156.87 53.06 ;
    RECT 156.66 53.35 156.87 53.42 ;
    RECT 153.8 52.63 154.01 52.7 ;
    RECT 153.8 52.99 154.01 53.06 ;
    RECT 153.8 53.35 154.01 53.42 ;
    RECT 153.34 52.63 153.55 52.7 ;
    RECT 153.34 52.99 153.55 53.06 ;
    RECT 153.34 53.35 153.55 53.42 ;
    RECT 150.48 52.63 150.69 52.7 ;
    RECT 150.48 52.99 150.69 53.06 ;
    RECT 150.48 53.35 150.69 53.42 ;
    RECT 150.02 52.63 150.23 52.7 ;
    RECT 150.02 52.99 150.23 53.06 ;
    RECT 150.02 53.35 150.23 53.42 ;
    RECT 213.56 52.63 213.77 52.7 ;
    RECT 213.56 52.99 213.77 53.06 ;
    RECT 213.56 53.35 213.77 53.42 ;
    RECT 213.1 52.63 213.31 52.7 ;
    RECT 213.1 52.99 213.31 53.06 ;
    RECT 213.1 53.35 213.31 53.42 ;
    RECT 210.24 52.63 210.45 52.7 ;
    RECT 210.24 52.99 210.45 53.06 ;
    RECT 210.24 53.35 210.45 53.42 ;
    RECT 209.78 52.63 209.99 52.7 ;
    RECT 209.78 52.99 209.99 53.06 ;
    RECT 209.78 53.35 209.99 53.42 ;
    RECT 206.92 52.63 207.13 52.7 ;
    RECT 206.92 52.99 207.13 53.06 ;
    RECT 206.92 53.35 207.13 53.42 ;
    RECT 206.46 52.63 206.67 52.7 ;
    RECT 206.46 52.99 206.67 53.06 ;
    RECT 206.46 53.35 206.67 53.42 ;
    RECT 203.6 52.63 203.81 52.7 ;
    RECT 203.6 52.99 203.81 53.06 ;
    RECT 203.6 53.35 203.81 53.42 ;
    RECT 203.14 52.63 203.35 52.7 ;
    RECT 203.14 52.99 203.35 53.06 ;
    RECT 203.14 53.35 203.35 53.42 ;
    RECT 200.28 52.63 200.49 52.7 ;
    RECT 200.28 52.99 200.49 53.06 ;
    RECT 200.28 53.35 200.49 53.42 ;
    RECT 199.82 52.63 200.03 52.7 ;
    RECT 199.82 52.99 200.03 53.06 ;
    RECT 199.82 53.35 200.03 53.42 ;
    RECT 196.96 52.63 197.17 52.7 ;
    RECT 196.96 52.99 197.17 53.06 ;
    RECT 196.96 53.35 197.17 53.42 ;
    RECT 196.5 52.63 196.71 52.7 ;
    RECT 196.5 52.99 196.71 53.06 ;
    RECT 196.5 53.35 196.71 53.42 ;
    RECT 193.64 52.63 193.85 52.7 ;
    RECT 193.64 52.99 193.85 53.06 ;
    RECT 193.64 53.35 193.85 53.42 ;
    RECT 193.18 52.63 193.39 52.7 ;
    RECT 193.18 52.99 193.39 53.06 ;
    RECT 193.18 53.35 193.39 53.42 ;
    RECT 190.32 52.63 190.53 52.7 ;
    RECT 190.32 52.99 190.53 53.06 ;
    RECT 190.32 53.35 190.53 53.42 ;
    RECT 189.86 52.63 190.07 52.7 ;
    RECT 189.86 52.99 190.07 53.06 ;
    RECT 189.86 53.35 190.07 53.42 ;
    RECT 187.0 52.63 187.21 52.7 ;
    RECT 187.0 52.99 187.21 53.06 ;
    RECT 187.0 53.35 187.21 53.42 ;
    RECT 186.54 52.63 186.75 52.7 ;
    RECT 186.54 52.99 186.75 53.06 ;
    RECT 186.54 53.35 186.75 53.42 ;
    RECT 183.68 52.63 183.89 52.7 ;
    RECT 183.68 52.99 183.89 53.06 ;
    RECT 183.68 53.35 183.89 53.42 ;
    RECT 183.22 52.63 183.43 52.7 ;
    RECT 183.22 52.99 183.43 53.06 ;
    RECT 183.22 53.35 183.43 53.42 ;
    RECT 147.485 52.99 147.555 53.06 ;
    RECT 266.68 52.63 266.89 52.7 ;
    RECT 266.68 52.99 266.89 53.06 ;
    RECT 266.68 53.35 266.89 53.42 ;
    RECT 266.22 52.63 266.43 52.7 ;
    RECT 266.22 52.99 266.43 53.06 ;
    RECT 266.22 53.35 266.43 53.42 ;
    RECT 263.36 52.63 263.57 52.7 ;
    RECT 263.36 52.99 263.57 53.06 ;
    RECT 263.36 53.35 263.57 53.42 ;
    RECT 262.9 52.63 263.11 52.7 ;
    RECT 262.9 52.99 263.11 53.06 ;
    RECT 262.9 53.35 263.11 53.42 ;
    RECT 260.04 52.63 260.25 52.7 ;
    RECT 260.04 52.99 260.25 53.06 ;
    RECT 260.04 53.35 260.25 53.42 ;
    RECT 259.58 52.63 259.79 52.7 ;
    RECT 259.58 52.99 259.79 53.06 ;
    RECT 259.58 53.35 259.79 53.42 ;
    RECT 256.72 52.63 256.93 52.7 ;
    RECT 256.72 52.99 256.93 53.06 ;
    RECT 256.72 53.35 256.93 53.42 ;
    RECT 256.26 52.63 256.47 52.7 ;
    RECT 256.26 52.99 256.47 53.06 ;
    RECT 256.26 53.35 256.47 53.42 ;
    RECT 253.4 52.63 253.61 52.7 ;
    RECT 253.4 52.99 253.61 53.06 ;
    RECT 253.4 53.35 253.61 53.42 ;
    RECT 252.94 52.63 253.15 52.7 ;
    RECT 252.94 52.99 253.15 53.06 ;
    RECT 252.94 53.35 253.15 53.42 ;
    RECT 250.08 88.65 250.29 88.72 ;
    RECT 250.08 89.01 250.29 89.08 ;
    RECT 250.08 89.37 250.29 89.44 ;
    RECT 249.62 88.65 249.83 88.72 ;
    RECT 249.62 89.01 249.83 89.08 ;
    RECT 249.62 89.37 249.83 89.44 ;
    RECT 246.76 88.65 246.97 88.72 ;
    RECT 246.76 89.01 246.97 89.08 ;
    RECT 246.76 89.37 246.97 89.44 ;
    RECT 246.3 88.65 246.51 88.72 ;
    RECT 246.3 89.01 246.51 89.08 ;
    RECT 246.3 89.37 246.51 89.44 ;
    RECT 243.44 88.65 243.65 88.72 ;
    RECT 243.44 89.01 243.65 89.08 ;
    RECT 243.44 89.37 243.65 89.44 ;
    RECT 242.98 88.65 243.19 88.72 ;
    RECT 242.98 89.01 243.19 89.08 ;
    RECT 242.98 89.37 243.19 89.44 ;
    RECT 240.12 88.65 240.33 88.72 ;
    RECT 240.12 89.01 240.33 89.08 ;
    RECT 240.12 89.37 240.33 89.44 ;
    RECT 239.66 88.65 239.87 88.72 ;
    RECT 239.66 89.01 239.87 89.08 ;
    RECT 239.66 89.37 239.87 89.44 ;
    RECT 236.8 88.65 237.01 88.72 ;
    RECT 236.8 89.01 237.01 89.08 ;
    RECT 236.8 89.37 237.01 89.44 ;
    RECT 236.34 88.65 236.55 88.72 ;
    RECT 236.34 89.01 236.55 89.08 ;
    RECT 236.34 89.37 236.55 89.44 ;
    RECT 233.48 88.65 233.69 88.72 ;
    RECT 233.48 89.01 233.69 89.08 ;
    RECT 233.48 89.37 233.69 89.44 ;
    RECT 233.02 88.65 233.23 88.72 ;
    RECT 233.02 89.01 233.23 89.08 ;
    RECT 233.02 89.37 233.23 89.44 ;
    RECT 230.16 88.65 230.37 88.72 ;
    RECT 230.16 89.01 230.37 89.08 ;
    RECT 230.16 89.37 230.37 89.44 ;
    RECT 229.7 88.65 229.91 88.72 ;
    RECT 229.7 89.01 229.91 89.08 ;
    RECT 229.7 89.37 229.91 89.44 ;
    RECT 226.84 88.65 227.05 88.72 ;
    RECT 226.84 89.01 227.05 89.08 ;
    RECT 226.84 89.37 227.05 89.44 ;
    RECT 226.38 88.65 226.59 88.72 ;
    RECT 226.38 89.01 226.59 89.08 ;
    RECT 226.38 89.37 226.59 89.44 ;
    RECT 223.52 88.65 223.73 88.72 ;
    RECT 223.52 89.01 223.73 89.08 ;
    RECT 223.52 89.37 223.73 89.44 ;
    RECT 223.06 88.65 223.27 88.72 ;
    RECT 223.06 89.01 223.27 89.08 ;
    RECT 223.06 89.37 223.27 89.44 ;
    RECT 220.2 88.65 220.41 88.72 ;
    RECT 220.2 89.01 220.41 89.08 ;
    RECT 220.2 89.37 220.41 89.44 ;
    RECT 219.74 88.65 219.95 88.72 ;
    RECT 219.74 89.01 219.95 89.08 ;
    RECT 219.74 89.37 219.95 89.44 ;
    RECT 216.88 88.65 217.09 88.72 ;
    RECT 216.88 89.01 217.09 89.08 ;
    RECT 216.88 89.37 217.09 89.44 ;
    RECT 216.42 88.65 216.63 88.72 ;
    RECT 216.42 89.01 216.63 89.08 ;
    RECT 216.42 89.37 216.63 89.44 ;
    RECT 267.91 89.01 267.98 89.08 ;
    RECT 180.36 88.65 180.57 88.72 ;
    RECT 180.36 89.01 180.57 89.08 ;
    RECT 180.36 89.37 180.57 89.44 ;
    RECT 179.9 88.65 180.11 88.72 ;
    RECT 179.9 89.01 180.11 89.08 ;
    RECT 179.9 89.37 180.11 89.44 ;
    RECT 177.04 88.65 177.25 88.72 ;
    RECT 177.04 89.01 177.25 89.08 ;
    RECT 177.04 89.37 177.25 89.44 ;
    RECT 176.58 88.65 176.79 88.72 ;
    RECT 176.58 89.01 176.79 89.08 ;
    RECT 176.58 89.37 176.79 89.44 ;
    RECT 173.72 88.65 173.93 88.72 ;
    RECT 173.72 89.01 173.93 89.08 ;
    RECT 173.72 89.37 173.93 89.44 ;
    RECT 173.26 88.65 173.47 88.72 ;
    RECT 173.26 89.01 173.47 89.08 ;
    RECT 173.26 89.37 173.47 89.44 ;
    RECT 170.4 88.65 170.61 88.72 ;
    RECT 170.4 89.01 170.61 89.08 ;
    RECT 170.4 89.37 170.61 89.44 ;
    RECT 169.94 88.65 170.15 88.72 ;
    RECT 169.94 89.01 170.15 89.08 ;
    RECT 169.94 89.37 170.15 89.44 ;
    RECT 167.08 88.65 167.29 88.72 ;
    RECT 167.08 89.01 167.29 89.08 ;
    RECT 167.08 89.37 167.29 89.44 ;
    RECT 166.62 88.65 166.83 88.72 ;
    RECT 166.62 89.01 166.83 89.08 ;
    RECT 166.62 89.37 166.83 89.44 ;
    RECT 163.76 88.65 163.97 88.72 ;
    RECT 163.76 89.01 163.97 89.08 ;
    RECT 163.76 89.37 163.97 89.44 ;
    RECT 163.3 88.65 163.51 88.72 ;
    RECT 163.3 89.01 163.51 89.08 ;
    RECT 163.3 89.37 163.51 89.44 ;
    RECT 160.44 88.65 160.65 88.72 ;
    RECT 160.44 89.01 160.65 89.08 ;
    RECT 160.44 89.37 160.65 89.44 ;
    RECT 159.98 88.65 160.19 88.72 ;
    RECT 159.98 89.01 160.19 89.08 ;
    RECT 159.98 89.37 160.19 89.44 ;
    RECT 157.12 88.65 157.33 88.72 ;
    RECT 157.12 89.01 157.33 89.08 ;
    RECT 157.12 89.37 157.33 89.44 ;
    RECT 156.66 88.65 156.87 88.72 ;
    RECT 156.66 89.01 156.87 89.08 ;
    RECT 156.66 89.37 156.87 89.44 ;
    RECT 153.8 88.65 154.01 88.72 ;
    RECT 153.8 89.01 154.01 89.08 ;
    RECT 153.8 89.37 154.01 89.44 ;
    RECT 153.34 88.65 153.55 88.72 ;
    RECT 153.34 89.01 153.55 89.08 ;
    RECT 153.34 89.37 153.55 89.44 ;
    RECT 150.48 88.65 150.69 88.72 ;
    RECT 150.48 89.01 150.69 89.08 ;
    RECT 150.48 89.37 150.69 89.44 ;
    RECT 150.02 88.65 150.23 88.72 ;
    RECT 150.02 89.01 150.23 89.08 ;
    RECT 150.02 89.37 150.23 89.44 ;
    RECT 213.56 88.65 213.77 88.72 ;
    RECT 213.56 89.01 213.77 89.08 ;
    RECT 213.56 89.37 213.77 89.44 ;
    RECT 213.1 88.65 213.31 88.72 ;
    RECT 213.1 89.01 213.31 89.08 ;
    RECT 213.1 89.37 213.31 89.44 ;
    RECT 210.24 88.65 210.45 88.72 ;
    RECT 210.24 89.01 210.45 89.08 ;
    RECT 210.24 89.37 210.45 89.44 ;
    RECT 209.78 88.65 209.99 88.72 ;
    RECT 209.78 89.01 209.99 89.08 ;
    RECT 209.78 89.37 209.99 89.44 ;
    RECT 206.92 88.65 207.13 88.72 ;
    RECT 206.92 89.01 207.13 89.08 ;
    RECT 206.92 89.37 207.13 89.44 ;
    RECT 206.46 88.65 206.67 88.72 ;
    RECT 206.46 89.01 206.67 89.08 ;
    RECT 206.46 89.37 206.67 89.44 ;
    RECT 203.6 88.65 203.81 88.72 ;
    RECT 203.6 89.01 203.81 89.08 ;
    RECT 203.6 89.37 203.81 89.44 ;
    RECT 203.14 88.65 203.35 88.72 ;
    RECT 203.14 89.01 203.35 89.08 ;
    RECT 203.14 89.37 203.35 89.44 ;
    RECT 200.28 88.65 200.49 88.72 ;
    RECT 200.28 89.01 200.49 89.08 ;
    RECT 200.28 89.37 200.49 89.44 ;
    RECT 199.82 88.65 200.03 88.72 ;
    RECT 199.82 89.01 200.03 89.08 ;
    RECT 199.82 89.37 200.03 89.44 ;
    RECT 196.96 88.65 197.17 88.72 ;
    RECT 196.96 89.01 197.17 89.08 ;
    RECT 196.96 89.37 197.17 89.44 ;
    RECT 196.5 88.65 196.71 88.72 ;
    RECT 196.5 89.01 196.71 89.08 ;
    RECT 196.5 89.37 196.71 89.44 ;
    RECT 193.64 88.65 193.85 88.72 ;
    RECT 193.64 89.01 193.85 89.08 ;
    RECT 193.64 89.37 193.85 89.44 ;
    RECT 193.18 88.65 193.39 88.72 ;
    RECT 193.18 89.01 193.39 89.08 ;
    RECT 193.18 89.37 193.39 89.44 ;
    RECT 190.32 88.65 190.53 88.72 ;
    RECT 190.32 89.01 190.53 89.08 ;
    RECT 190.32 89.37 190.53 89.44 ;
    RECT 189.86 88.65 190.07 88.72 ;
    RECT 189.86 89.01 190.07 89.08 ;
    RECT 189.86 89.37 190.07 89.44 ;
    RECT 187.0 88.65 187.21 88.72 ;
    RECT 187.0 89.01 187.21 89.08 ;
    RECT 187.0 89.37 187.21 89.44 ;
    RECT 186.54 88.65 186.75 88.72 ;
    RECT 186.54 89.01 186.75 89.08 ;
    RECT 186.54 89.37 186.75 89.44 ;
    RECT 183.68 88.65 183.89 88.72 ;
    RECT 183.68 89.01 183.89 89.08 ;
    RECT 183.68 89.37 183.89 89.44 ;
    RECT 183.22 88.65 183.43 88.72 ;
    RECT 183.22 89.01 183.43 89.08 ;
    RECT 183.22 89.37 183.43 89.44 ;
    RECT 147.485 89.01 147.555 89.08 ;
    RECT 266.68 88.65 266.89 88.72 ;
    RECT 266.68 89.01 266.89 89.08 ;
    RECT 266.68 89.37 266.89 89.44 ;
    RECT 266.22 88.65 266.43 88.72 ;
    RECT 266.22 89.01 266.43 89.08 ;
    RECT 266.22 89.37 266.43 89.44 ;
    RECT 263.36 88.65 263.57 88.72 ;
    RECT 263.36 89.01 263.57 89.08 ;
    RECT 263.36 89.37 263.57 89.44 ;
    RECT 262.9 88.65 263.11 88.72 ;
    RECT 262.9 89.01 263.11 89.08 ;
    RECT 262.9 89.37 263.11 89.44 ;
    RECT 260.04 88.65 260.25 88.72 ;
    RECT 260.04 89.01 260.25 89.08 ;
    RECT 260.04 89.37 260.25 89.44 ;
    RECT 259.58 88.65 259.79 88.72 ;
    RECT 259.58 89.01 259.79 89.08 ;
    RECT 259.58 89.37 259.79 89.44 ;
    RECT 256.72 88.65 256.93 88.72 ;
    RECT 256.72 89.01 256.93 89.08 ;
    RECT 256.72 89.37 256.93 89.44 ;
    RECT 256.26 88.65 256.47 88.72 ;
    RECT 256.26 89.01 256.47 89.08 ;
    RECT 256.26 89.37 256.47 89.44 ;
    RECT 253.4 88.65 253.61 88.72 ;
    RECT 253.4 89.01 253.61 89.08 ;
    RECT 253.4 89.37 253.61 89.44 ;
    RECT 252.94 88.65 253.15 88.72 ;
    RECT 252.94 89.01 253.15 89.08 ;
    RECT 252.94 89.37 253.15 89.44 ;
    RECT 250.08 51.91 250.29 51.98 ;
    RECT 250.08 52.27 250.29 52.34 ;
    RECT 250.08 52.63 250.29 52.7 ;
    RECT 249.62 51.91 249.83 51.98 ;
    RECT 249.62 52.27 249.83 52.34 ;
    RECT 249.62 52.63 249.83 52.7 ;
    RECT 246.76 51.91 246.97 51.98 ;
    RECT 246.76 52.27 246.97 52.34 ;
    RECT 246.76 52.63 246.97 52.7 ;
    RECT 246.3 51.91 246.51 51.98 ;
    RECT 246.3 52.27 246.51 52.34 ;
    RECT 246.3 52.63 246.51 52.7 ;
    RECT 243.44 51.91 243.65 51.98 ;
    RECT 243.44 52.27 243.65 52.34 ;
    RECT 243.44 52.63 243.65 52.7 ;
    RECT 242.98 51.91 243.19 51.98 ;
    RECT 242.98 52.27 243.19 52.34 ;
    RECT 242.98 52.63 243.19 52.7 ;
    RECT 240.12 51.91 240.33 51.98 ;
    RECT 240.12 52.27 240.33 52.34 ;
    RECT 240.12 52.63 240.33 52.7 ;
    RECT 239.66 51.91 239.87 51.98 ;
    RECT 239.66 52.27 239.87 52.34 ;
    RECT 239.66 52.63 239.87 52.7 ;
    RECT 236.8 51.91 237.01 51.98 ;
    RECT 236.8 52.27 237.01 52.34 ;
    RECT 236.8 52.63 237.01 52.7 ;
    RECT 236.34 51.91 236.55 51.98 ;
    RECT 236.34 52.27 236.55 52.34 ;
    RECT 236.34 52.63 236.55 52.7 ;
    RECT 233.48 51.91 233.69 51.98 ;
    RECT 233.48 52.27 233.69 52.34 ;
    RECT 233.48 52.63 233.69 52.7 ;
    RECT 233.02 51.91 233.23 51.98 ;
    RECT 233.02 52.27 233.23 52.34 ;
    RECT 233.02 52.63 233.23 52.7 ;
    RECT 230.16 51.91 230.37 51.98 ;
    RECT 230.16 52.27 230.37 52.34 ;
    RECT 230.16 52.63 230.37 52.7 ;
    RECT 229.7 51.91 229.91 51.98 ;
    RECT 229.7 52.27 229.91 52.34 ;
    RECT 229.7 52.63 229.91 52.7 ;
    RECT 226.84 51.91 227.05 51.98 ;
    RECT 226.84 52.27 227.05 52.34 ;
    RECT 226.84 52.63 227.05 52.7 ;
    RECT 226.38 51.91 226.59 51.98 ;
    RECT 226.38 52.27 226.59 52.34 ;
    RECT 226.38 52.63 226.59 52.7 ;
    RECT 223.52 51.91 223.73 51.98 ;
    RECT 223.52 52.27 223.73 52.34 ;
    RECT 223.52 52.63 223.73 52.7 ;
    RECT 223.06 51.91 223.27 51.98 ;
    RECT 223.06 52.27 223.27 52.34 ;
    RECT 223.06 52.63 223.27 52.7 ;
    RECT 220.2 51.91 220.41 51.98 ;
    RECT 220.2 52.27 220.41 52.34 ;
    RECT 220.2 52.63 220.41 52.7 ;
    RECT 219.74 51.91 219.95 51.98 ;
    RECT 219.74 52.27 219.95 52.34 ;
    RECT 219.74 52.63 219.95 52.7 ;
    RECT 216.88 51.91 217.09 51.98 ;
    RECT 216.88 52.27 217.09 52.34 ;
    RECT 216.88 52.63 217.09 52.7 ;
    RECT 216.42 51.91 216.63 51.98 ;
    RECT 216.42 52.27 216.63 52.34 ;
    RECT 216.42 52.63 216.63 52.7 ;
    RECT 267.91 52.27 267.98 52.34 ;
    RECT 180.36 51.91 180.57 51.98 ;
    RECT 180.36 52.27 180.57 52.34 ;
    RECT 180.36 52.63 180.57 52.7 ;
    RECT 179.9 51.91 180.11 51.98 ;
    RECT 179.9 52.27 180.11 52.34 ;
    RECT 179.9 52.63 180.11 52.7 ;
    RECT 177.04 51.91 177.25 51.98 ;
    RECT 177.04 52.27 177.25 52.34 ;
    RECT 177.04 52.63 177.25 52.7 ;
    RECT 176.58 51.91 176.79 51.98 ;
    RECT 176.58 52.27 176.79 52.34 ;
    RECT 176.58 52.63 176.79 52.7 ;
    RECT 173.72 51.91 173.93 51.98 ;
    RECT 173.72 52.27 173.93 52.34 ;
    RECT 173.72 52.63 173.93 52.7 ;
    RECT 173.26 51.91 173.47 51.98 ;
    RECT 173.26 52.27 173.47 52.34 ;
    RECT 173.26 52.63 173.47 52.7 ;
    RECT 170.4 51.91 170.61 51.98 ;
    RECT 170.4 52.27 170.61 52.34 ;
    RECT 170.4 52.63 170.61 52.7 ;
    RECT 169.94 51.91 170.15 51.98 ;
    RECT 169.94 52.27 170.15 52.34 ;
    RECT 169.94 52.63 170.15 52.7 ;
    RECT 167.08 51.91 167.29 51.98 ;
    RECT 167.08 52.27 167.29 52.34 ;
    RECT 167.08 52.63 167.29 52.7 ;
    RECT 166.62 51.91 166.83 51.98 ;
    RECT 166.62 52.27 166.83 52.34 ;
    RECT 166.62 52.63 166.83 52.7 ;
    RECT 163.76 51.91 163.97 51.98 ;
    RECT 163.76 52.27 163.97 52.34 ;
    RECT 163.76 52.63 163.97 52.7 ;
    RECT 163.3 51.91 163.51 51.98 ;
    RECT 163.3 52.27 163.51 52.34 ;
    RECT 163.3 52.63 163.51 52.7 ;
    RECT 160.44 51.91 160.65 51.98 ;
    RECT 160.44 52.27 160.65 52.34 ;
    RECT 160.44 52.63 160.65 52.7 ;
    RECT 159.98 51.91 160.19 51.98 ;
    RECT 159.98 52.27 160.19 52.34 ;
    RECT 159.98 52.63 160.19 52.7 ;
    RECT 157.12 51.91 157.33 51.98 ;
    RECT 157.12 52.27 157.33 52.34 ;
    RECT 157.12 52.63 157.33 52.7 ;
    RECT 156.66 51.91 156.87 51.98 ;
    RECT 156.66 52.27 156.87 52.34 ;
    RECT 156.66 52.63 156.87 52.7 ;
    RECT 153.8 51.91 154.01 51.98 ;
    RECT 153.8 52.27 154.01 52.34 ;
    RECT 153.8 52.63 154.01 52.7 ;
    RECT 153.34 51.91 153.55 51.98 ;
    RECT 153.34 52.27 153.55 52.34 ;
    RECT 153.34 52.63 153.55 52.7 ;
    RECT 150.48 51.91 150.69 51.98 ;
    RECT 150.48 52.27 150.69 52.34 ;
    RECT 150.48 52.63 150.69 52.7 ;
    RECT 150.02 51.91 150.23 51.98 ;
    RECT 150.02 52.27 150.23 52.34 ;
    RECT 150.02 52.63 150.23 52.7 ;
    RECT 213.56 51.91 213.77 51.98 ;
    RECT 213.56 52.27 213.77 52.34 ;
    RECT 213.56 52.63 213.77 52.7 ;
    RECT 213.1 51.91 213.31 51.98 ;
    RECT 213.1 52.27 213.31 52.34 ;
    RECT 213.1 52.63 213.31 52.7 ;
    RECT 210.24 51.91 210.45 51.98 ;
    RECT 210.24 52.27 210.45 52.34 ;
    RECT 210.24 52.63 210.45 52.7 ;
    RECT 209.78 51.91 209.99 51.98 ;
    RECT 209.78 52.27 209.99 52.34 ;
    RECT 209.78 52.63 209.99 52.7 ;
    RECT 206.92 51.91 207.13 51.98 ;
    RECT 206.92 52.27 207.13 52.34 ;
    RECT 206.92 52.63 207.13 52.7 ;
    RECT 206.46 51.91 206.67 51.98 ;
    RECT 206.46 52.27 206.67 52.34 ;
    RECT 206.46 52.63 206.67 52.7 ;
    RECT 203.6 51.91 203.81 51.98 ;
    RECT 203.6 52.27 203.81 52.34 ;
    RECT 203.6 52.63 203.81 52.7 ;
    RECT 203.14 51.91 203.35 51.98 ;
    RECT 203.14 52.27 203.35 52.34 ;
    RECT 203.14 52.63 203.35 52.7 ;
    RECT 200.28 51.91 200.49 51.98 ;
    RECT 200.28 52.27 200.49 52.34 ;
    RECT 200.28 52.63 200.49 52.7 ;
    RECT 199.82 51.91 200.03 51.98 ;
    RECT 199.82 52.27 200.03 52.34 ;
    RECT 199.82 52.63 200.03 52.7 ;
    RECT 196.96 51.91 197.17 51.98 ;
    RECT 196.96 52.27 197.17 52.34 ;
    RECT 196.96 52.63 197.17 52.7 ;
    RECT 196.5 51.91 196.71 51.98 ;
    RECT 196.5 52.27 196.71 52.34 ;
    RECT 196.5 52.63 196.71 52.7 ;
    RECT 193.64 51.91 193.85 51.98 ;
    RECT 193.64 52.27 193.85 52.34 ;
    RECT 193.64 52.63 193.85 52.7 ;
    RECT 193.18 51.91 193.39 51.98 ;
    RECT 193.18 52.27 193.39 52.34 ;
    RECT 193.18 52.63 193.39 52.7 ;
    RECT 190.32 51.91 190.53 51.98 ;
    RECT 190.32 52.27 190.53 52.34 ;
    RECT 190.32 52.63 190.53 52.7 ;
    RECT 189.86 51.91 190.07 51.98 ;
    RECT 189.86 52.27 190.07 52.34 ;
    RECT 189.86 52.63 190.07 52.7 ;
    RECT 187.0 51.91 187.21 51.98 ;
    RECT 187.0 52.27 187.21 52.34 ;
    RECT 187.0 52.63 187.21 52.7 ;
    RECT 186.54 51.91 186.75 51.98 ;
    RECT 186.54 52.27 186.75 52.34 ;
    RECT 186.54 52.63 186.75 52.7 ;
    RECT 183.68 51.91 183.89 51.98 ;
    RECT 183.68 52.27 183.89 52.34 ;
    RECT 183.68 52.63 183.89 52.7 ;
    RECT 183.22 51.91 183.43 51.98 ;
    RECT 183.22 52.27 183.43 52.34 ;
    RECT 183.22 52.63 183.43 52.7 ;
    RECT 147.485 52.27 147.555 52.34 ;
    RECT 266.68 51.91 266.89 51.98 ;
    RECT 266.68 52.27 266.89 52.34 ;
    RECT 266.68 52.63 266.89 52.7 ;
    RECT 266.22 51.91 266.43 51.98 ;
    RECT 266.22 52.27 266.43 52.34 ;
    RECT 266.22 52.63 266.43 52.7 ;
    RECT 263.36 51.91 263.57 51.98 ;
    RECT 263.36 52.27 263.57 52.34 ;
    RECT 263.36 52.63 263.57 52.7 ;
    RECT 262.9 51.91 263.11 51.98 ;
    RECT 262.9 52.27 263.11 52.34 ;
    RECT 262.9 52.63 263.11 52.7 ;
    RECT 260.04 51.91 260.25 51.98 ;
    RECT 260.04 52.27 260.25 52.34 ;
    RECT 260.04 52.63 260.25 52.7 ;
    RECT 259.58 51.91 259.79 51.98 ;
    RECT 259.58 52.27 259.79 52.34 ;
    RECT 259.58 52.63 259.79 52.7 ;
    RECT 256.72 51.91 256.93 51.98 ;
    RECT 256.72 52.27 256.93 52.34 ;
    RECT 256.72 52.63 256.93 52.7 ;
    RECT 256.26 51.91 256.47 51.98 ;
    RECT 256.26 52.27 256.47 52.34 ;
    RECT 256.26 52.63 256.47 52.7 ;
    RECT 253.4 51.91 253.61 51.98 ;
    RECT 253.4 52.27 253.61 52.34 ;
    RECT 253.4 52.63 253.61 52.7 ;
    RECT 252.94 51.91 253.15 51.98 ;
    RECT 252.94 52.27 253.15 52.34 ;
    RECT 252.94 52.63 253.15 52.7 ;
    RECT 250.08 87.93 250.29 88.0 ;
    RECT 250.08 88.29 250.29 88.36 ;
    RECT 250.08 88.65 250.29 88.72 ;
    RECT 249.62 87.93 249.83 88.0 ;
    RECT 249.62 88.29 249.83 88.36 ;
    RECT 249.62 88.65 249.83 88.72 ;
    RECT 246.76 87.93 246.97 88.0 ;
    RECT 246.76 88.29 246.97 88.36 ;
    RECT 246.76 88.65 246.97 88.72 ;
    RECT 246.3 87.93 246.51 88.0 ;
    RECT 246.3 88.29 246.51 88.36 ;
    RECT 246.3 88.65 246.51 88.72 ;
    RECT 243.44 87.93 243.65 88.0 ;
    RECT 243.44 88.29 243.65 88.36 ;
    RECT 243.44 88.65 243.65 88.72 ;
    RECT 242.98 87.93 243.19 88.0 ;
    RECT 242.98 88.29 243.19 88.36 ;
    RECT 242.98 88.65 243.19 88.72 ;
    RECT 240.12 87.93 240.33 88.0 ;
    RECT 240.12 88.29 240.33 88.36 ;
    RECT 240.12 88.65 240.33 88.72 ;
    RECT 239.66 87.93 239.87 88.0 ;
    RECT 239.66 88.29 239.87 88.36 ;
    RECT 239.66 88.65 239.87 88.72 ;
    RECT 236.8 87.93 237.01 88.0 ;
    RECT 236.8 88.29 237.01 88.36 ;
    RECT 236.8 88.65 237.01 88.72 ;
    RECT 236.34 87.93 236.55 88.0 ;
    RECT 236.34 88.29 236.55 88.36 ;
    RECT 236.34 88.65 236.55 88.72 ;
    RECT 233.48 87.93 233.69 88.0 ;
    RECT 233.48 88.29 233.69 88.36 ;
    RECT 233.48 88.65 233.69 88.72 ;
    RECT 233.02 87.93 233.23 88.0 ;
    RECT 233.02 88.29 233.23 88.36 ;
    RECT 233.02 88.65 233.23 88.72 ;
    RECT 230.16 87.93 230.37 88.0 ;
    RECT 230.16 88.29 230.37 88.36 ;
    RECT 230.16 88.65 230.37 88.72 ;
    RECT 229.7 87.93 229.91 88.0 ;
    RECT 229.7 88.29 229.91 88.36 ;
    RECT 229.7 88.65 229.91 88.72 ;
    RECT 226.84 87.93 227.05 88.0 ;
    RECT 226.84 88.29 227.05 88.36 ;
    RECT 226.84 88.65 227.05 88.72 ;
    RECT 226.38 87.93 226.59 88.0 ;
    RECT 226.38 88.29 226.59 88.36 ;
    RECT 226.38 88.65 226.59 88.72 ;
    RECT 223.52 87.93 223.73 88.0 ;
    RECT 223.52 88.29 223.73 88.36 ;
    RECT 223.52 88.65 223.73 88.72 ;
    RECT 223.06 87.93 223.27 88.0 ;
    RECT 223.06 88.29 223.27 88.36 ;
    RECT 223.06 88.65 223.27 88.72 ;
    RECT 220.2 87.93 220.41 88.0 ;
    RECT 220.2 88.29 220.41 88.36 ;
    RECT 220.2 88.65 220.41 88.72 ;
    RECT 219.74 87.93 219.95 88.0 ;
    RECT 219.74 88.29 219.95 88.36 ;
    RECT 219.74 88.65 219.95 88.72 ;
    RECT 216.88 87.93 217.09 88.0 ;
    RECT 216.88 88.29 217.09 88.36 ;
    RECT 216.88 88.65 217.09 88.72 ;
    RECT 216.42 87.93 216.63 88.0 ;
    RECT 216.42 88.29 216.63 88.36 ;
    RECT 216.42 88.65 216.63 88.72 ;
    RECT 267.91 88.29 267.98 88.36 ;
    RECT 180.36 87.93 180.57 88.0 ;
    RECT 180.36 88.29 180.57 88.36 ;
    RECT 180.36 88.65 180.57 88.72 ;
    RECT 179.9 87.93 180.11 88.0 ;
    RECT 179.9 88.29 180.11 88.36 ;
    RECT 179.9 88.65 180.11 88.72 ;
    RECT 177.04 87.93 177.25 88.0 ;
    RECT 177.04 88.29 177.25 88.36 ;
    RECT 177.04 88.65 177.25 88.72 ;
    RECT 176.58 87.93 176.79 88.0 ;
    RECT 176.58 88.29 176.79 88.36 ;
    RECT 176.58 88.65 176.79 88.72 ;
    RECT 173.72 87.93 173.93 88.0 ;
    RECT 173.72 88.29 173.93 88.36 ;
    RECT 173.72 88.65 173.93 88.72 ;
    RECT 173.26 87.93 173.47 88.0 ;
    RECT 173.26 88.29 173.47 88.36 ;
    RECT 173.26 88.65 173.47 88.72 ;
    RECT 170.4 87.93 170.61 88.0 ;
    RECT 170.4 88.29 170.61 88.36 ;
    RECT 170.4 88.65 170.61 88.72 ;
    RECT 169.94 87.93 170.15 88.0 ;
    RECT 169.94 88.29 170.15 88.36 ;
    RECT 169.94 88.65 170.15 88.72 ;
    RECT 167.08 87.93 167.29 88.0 ;
    RECT 167.08 88.29 167.29 88.36 ;
    RECT 167.08 88.65 167.29 88.72 ;
    RECT 166.62 87.93 166.83 88.0 ;
    RECT 166.62 88.29 166.83 88.36 ;
    RECT 166.62 88.65 166.83 88.72 ;
    RECT 163.76 87.93 163.97 88.0 ;
    RECT 163.76 88.29 163.97 88.36 ;
    RECT 163.76 88.65 163.97 88.72 ;
    RECT 163.3 87.93 163.51 88.0 ;
    RECT 163.3 88.29 163.51 88.36 ;
    RECT 163.3 88.65 163.51 88.72 ;
    RECT 160.44 87.93 160.65 88.0 ;
    RECT 160.44 88.29 160.65 88.36 ;
    RECT 160.44 88.65 160.65 88.72 ;
    RECT 159.98 87.93 160.19 88.0 ;
    RECT 159.98 88.29 160.19 88.36 ;
    RECT 159.98 88.65 160.19 88.72 ;
    RECT 157.12 87.93 157.33 88.0 ;
    RECT 157.12 88.29 157.33 88.36 ;
    RECT 157.12 88.65 157.33 88.72 ;
    RECT 156.66 87.93 156.87 88.0 ;
    RECT 156.66 88.29 156.87 88.36 ;
    RECT 156.66 88.65 156.87 88.72 ;
    RECT 153.8 87.93 154.01 88.0 ;
    RECT 153.8 88.29 154.01 88.36 ;
    RECT 153.8 88.65 154.01 88.72 ;
    RECT 153.34 87.93 153.55 88.0 ;
    RECT 153.34 88.29 153.55 88.36 ;
    RECT 153.34 88.65 153.55 88.72 ;
    RECT 150.48 87.93 150.69 88.0 ;
    RECT 150.48 88.29 150.69 88.36 ;
    RECT 150.48 88.65 150.69 88.72 ;
    RECT 150.02 87.93 150.23 88.0 ;
    RECT 150.02 88.29 150.23 88.36 ;
    RECT 150.02 88.65 150.23 88.72 ;
    RECT 213.56 87.93 213.77 88.0 ;
    RECT 213.56 88.29 213.77 88.36 ;
    RECT 213.56 88.65 213.77 88.72 ;
    RECT 213.1 87.93 213.31 88.0 ;
    RECT 213.1 88.29 213.31 88.36 ;
    RECT 213.1 88.65 213.31 88.72 ;
    RECT 210.24 87.93 210.45 88.0 ;
    RECT 210.24 88.29 210.45 88.36 ;
    RECT 210.24 88.65 210.45 88.72 ;
    RECT 209.78 87.93 209.99 88.0 ;
    RECT 209.78 88.29 209.99 88.36 ;
    RECT 209.78 88.65 209.99 88.72 ;
    RECT 206.92 87.93 207.13 88.0 ;
    RECT 206.92 88.29 207.13 88.36 ;
    RECT 206.92 88.65 207.13 88.72 ;
    RECT 206.46 87.93 206.67 88.0 ;
    RECT 206.46 88.29 206.67 88.36 ;
    RECT 206.46 88.65 206.67 88.72 ;
    RECT 203.6 87.93 203.81 88.0 ;
    RECT 203.6 88.29 203.81 88.36 ;
    RECT 203.6 88.65 203.81 88.72 ;
    RECT 203.14 87.93 203.35 88.0 ;
    RECT 203.14 88.29 203.35 88.36 ;
    RECT 203.14 88.65 203.35 88.72 ;
    RECT 200.28 87.93 200.49 88.0 ;
    RECT 200.28 88.29 200.49 88.36 ;
    RECT 200.28 88.65 200.49 88.72 ;
    RECT 199.82 87.93 200.03 88.0 ;
    RECT 199.82 88.29 200.03 88.36 ;
    RECT 199.82 88.65 200.03 88.72 ;
    RECT 196.96 87.93 197.17 88.0 ;
    RECT 196.96 88.29 197.17 88.36 ;
    RECT 196.96 88.65 197.17 88.72 ;
    RECT 196.5 87.93 196.71 88.0 ;
    RECT 196.5 88.29 196.71 88.36 ;
    RECT 196.5 88.65 196.71 88.72 ;
    RECT 193.64 87.93 193.85 88.0 ;
    RECT 193.64 88.29 193.85 88.36 ;
    RECT 193.64 88.65 193.85 88.72 ;
    RECT 193.18 87.93 193.39 88.0 ;
    RECT 193.18 88.29 193.39 88.36 ;
    RECT 193.18 88.65 193.39 88.72 ;
    RECT 190.32 87.93 190.53 88.0 ;
    RECT 190.32 88.29 190.53 88.36 ;
    RECT 190.32 88.65 190.53 88.72 ;
    RECT 189.86 87.93 190.07 88.0 ;
    RECT 189.86 88.29 190.07 88.36 ;
    RECT 189.86 88.65 190.07 88.72 ;
    RECT 187.0 87.93 187.21 88.0 ;
    RECT 187.0 88.29 187.21 88.36 ;
    RECT 187.0 88.65 187.21 88.72 ;
    RECT 186.54 87.93 186.75 88.0 ;
    RECT 186.54 88.29 186.75 88.36 ;
    RECT 186.54 88.65 186.75 88.72 ;
    RECT 183.68 87.93 183.89 88.0 ;
    RECT 183.68 88.29 183.89 88.36 ;
    RECT 183.68 88.65 183.89 88.72 ;
    RECT 183.22 87.93 183.43 88.0 ;
    RECT 183.22 88.29 183.43 88.36 ;
    RECT 183.22 88.65 183.43 88.72 ;
    RECT 147.485 88.29 147.555 88.36 ;
    RECT 266.68 87.93 266.89 88.0 ;
    RECT 266.68 88.29 266.89 88.36 ;
    RECT 266.68 88.65 266.89 88.72 ;
    RECT 266.22 87.93 266.43 88.0 ;
    RECT 266.22 88.29 266.43 88.36 ;
    RECT 266.22 88.65 266.43 88.72 ;
    RECT 263.36 87.93 263.57 88.0 ;
    RECT 263.36 88.29 263.57 88.36 ;
    RECT 263.36 88.65 263.57 88.72 ;
    RECT 262.9 87.93 263.11 88.0 ;
    RECT 262.9 88.29 263.11 88.36 ;
    RECT 262.9 88.65 263.11 88.72 ;
    RECT 260.04 87.93 260.25 88.0 ;
    RECT 260.04 88.29 260.25 88.36 ;
    RECT 260.04 88.65 260.25 88.72 ;
    RECT 259.58 87.93 259.79 88.0 ;
    RECT 259.58 88.29 259.79 88.36 ;
    RECT 259.58 88.65 259.79 88.72 ;
    RECT 256.72 87.93 256.93 88.0 ;
    RECT 256.72 88.29 256.93 88.36 ;
    RECT 256.72 88.65 256.93 88.72 ;
    RECT 256.26 87.93 256.47 88.0 ;
    RECT 256.26 88.29 256.47 88.36 ;
    RECT 256.26 88.65 256.47 88.72 ;
    RECT 253.4 87.93 253.61 88.0 ;
    RECT 253.4 88.29 253.61 88.36 ;
    RECT 253.4 88.65 253.61 88.72 ;
    RECT 252.94 87.93 253.15 88.0 ;
    RECT 252.94 88.29 253.15 88.36 ;
    RECT 252.94 88.65 253.15 88.72 ;
    RECT 250.08 51.19 250.29 51.26 ;
    RECT 250.08 51.55 250.29 51.62 ;
    RECT 250.08 51.91 250.29 51.98 ;
    RECT 249.62 51.19 249.83 51.26 ;
    RECT 249.62 51.55 249.83 51.62 ;
    RECT 249.62 51.91 249.83 51.98 ;
    RECT 246.76 51.19 246.97 51.26 ;
    RECT 246.76 51.55 246.97 51.62 ;
    RECT 246.76 51.91 246.97 51.98 ;
    RECT 246.3 51.19 246.51 51.26 ;
    RECT 246.3 51.55 246.51 51.62 ;
    RECT 246.3 51.91 246.51 51.98 ;
    RECT 243.44 51.19 243.65 51.26 ;
    RECT 243.44 51.55 243.65 51.62 ;
    RECT 243.44 51.91 243.65 51.98 ;
    RECT 242.98 51.19 243.19 51.26 ;
    RECT 242.98 51.55 243.19 51.62 ;
    RECT 242.98 51.91 243.19 51.98 ;
    RECT 240.12 51.19 240.33 51.26 ;
    RECT 240.12 51.55 240.33 51.62 ;
    RECT 240.12 51.91 240.33 51.98 ;
    RECT 239.66 51.19 239.87 51.26 ;
    RECT 239.66 51.55 239.87 51.62 ;
    RECT 239.66 51.91 239.87 51.98 ;
    RECT 236.8 51.19 237.01 51.26 ;
    RECT 236.8 51.55 237.01 51.62 ;
    RECT 236.8 51.91 237.01 51.98 ;
    RECT 236.34 51.19 236.55 51.26 ;
    RECT 236.34 51.55 236.55 51.62 ;
    RECT 236.34 51.91 236.55 51.98 ;
    RECT 233.48 51.19 233.69 51.26 ;
    RECT 233.48 51.55 233.69 51.62 ;
    RECT 233.48 51.91 233.69 51.98 ;
    RECT 233.02 51.19 233.23 51.26 ;
    RECT 233.02 51.55 233.23 51.62 ;
    RECT 233.02 51.91 233.23 51.98 ;
    RECT 230.16 51.19 230.37 51.26 ;
    RECT 230.16 51.55 230.37 51.62 ;
    RECT 230.16 51.91 230.37 51.98 ;
    RECT 229.7 51.19 229.91 51.26 ;
    RECT 229.7 51.55 229.91 51.62 ;
    RECT 229.7 51.91 229.91 51.98 ;
    RECT 226.84 51.19 227.05 51.26 ;
    RECT 226.84 51.55 227.05 51.62 ;
    RECT 226.84 51.91 227.05 51.98 ;
    RECT 226.38 51.19 226.59 51.26 ;
    RECT 226.38 51.55 226.59 51.62 ;
    RECT 226.38 51.91 226.59 51.98 ;
    RECT 223.52 51.19 223.73 51.26 ;
    RECT 223.52 51.55 223.73 51.62 ;
    RECT 223.52 51.91 223.73 51.98 ;
    RECT 223.06 51.19 223.27 51.26 ;
    RECT 223.06 51.55 223.27 51.62 ;
    RECT 223.06 51.91 223.27 51.98 ;
    RECT 220.2 51.19 220.41 51.26 ;
    RECT 220.2 51.55 220.41 51.62 ;
    RECT 220.2 51.91 220.41 51.98 ;
    RECT 219.74 51.19 219.95 51.26 ;
    RECT 219.74 51.55 219.95 51.62 ;
    RECT 219.74 51.91 219.95 51.98 ;
    RECT 216.88 51.19 217.09 51.26 ;
    RECT 216.88 51.55 217.09 51.62 ;
    RECT 216.88 51.91 217.09 51.98 ;
    RECT 216.42 51.19 216.63 51.26 ;
    RECT 216.42 51.55 216.63 51.62 ;
    RECT 216.42 51.91 216.63 51.98 ;
    RECT 267.91 51.55 267.98 51.62 ;
    RECT 180.36 51.19 180.57 51.26 ;
    RECT 180.36 51.55 180.57 51.62 ;
    RECT 180.36 51.91 180.57 51.98 ;
    RECT 179.9 51.19 180.11 51.26 ;
    RECT 179.9 51.55 180.11 51.62 ;
    RECT 179.9 51.91 180.11 51.98 ;
    RECT 177.04 51.19 177.25 51.26 ;
    RECT 177.04 51.55 177.25 51.62 ;
    RECT 177.04 51.91 177.25 51.98 ;
    RECT 176.58 51.19 176.79 51.26 ;
    RECT 176.58 51.55 176.79 51.62 ;
    RECT 176.58 51.91 176.79 51.98 ;
    RECT 173.72 51.19 173.93 51.26 ;
    RECT 173.72 51.55 173.93 51.62 ;
    RECT 173.72 51.91 173.93 51.98 ;
    RECT 173.26 51.19 173.47 51.26 ;
    RECT 173.26 51.55 173.47 51.62 ;
    RECT 173.26 51.91 173.47 51.98 ;
    RECT 170.4 51.19 170.61 51.26 ;
    RECT 170.4 51.55 170.61 51.62 ;
    RECT 170.4 51.91 170.61 51.98 ;
    RECT 169.94 51.19 170.15 51.26 ;
    RECT 169.94 51.55 170.15 51.62 ;
    RECT 169.94 51.91 170.15 51.98 ;
    RECT 167.08 51.19 167.29 51.26 ;
    RECT 167.08 51.55 167.29 51.62 ;
    RECT 167.08 51.91 167.29 51.98 ;
    RECT 166.62 51.19 166.83 51.26 ;
    RECT 166.62 51.55 166.83 51.62 ;
    RECT 166.62 51.91 166.83 51.98 ;
    RECT 163.76 51.19 163.97 51.26 ;
    RECT 163.76 51.55 163.97 51.62 ;
    RECT 163.76 51.91 163.97 51.98 ;
    RECT 163.3 51.19 163.51 51.26 ;
    RECT 163.3 51.55 163.51 51.62 ;
    RECT 163.3 51.91 163.51 51.98 ;
    RECT 160.44 51.19 160.65 51.26 ;
    RECT 160.44 51.55 160.65 51.62 ;
    RECT 160.44 51.91 160.65 51.98 ;
    RECT 159.98 51.19 160.19 51.26 ;
    RECT 159.98 51.55 160.19 51.62 ;
    RECT 159.98 51.91 160.19 51.98 ;
    RECT 157.12 51.19 157.33 51.26 ;
    RECT 157.12 51.55 157.33 51.62 ;
    RECT 157.12 51.91 157.33 51.98 ;
    RECT 156.66 51.19 156.87 51.26 ;
    RECT 156.66 51.55 156.87 51.62 ;
    RECT 156.66 51.91 156.87 51.98 ;
    RECT 153.8 51.19 154.01 51.26 ;
    RECT 153.8 51.55 154.01 51.62 ;
    RECT 153.8 51.91 154.01 51.98 ;
    RECT 153.34 51.19 153.55 51.26 ;
    RECT 153.34 51.55 153.55 51.62 ;
    RECT 153.34 51.91 153.55 51.98 ;
    RECT 150.48 51.19 150.69 51.26 ;
    RECT 150.48 51.55 150.69 51.62 ;
    RECT 150.48 51.91 150.69 51.98 ;
    RECT 150.02 51.19 150.23 51.26 ;
    RECT 150.02 51.55 150.23 51.62 ;
    RECT 150.02 51.91 150.23 51.98 ;
    RECT 213.56 51.19 213.77 51.26 ;
    RECT 213.56 51.55 213.77 51.62 ;
    RECT 213.56 51.91 213.77 51.98 ;
    RECT 213.1 51.19 213.31 51.26 ;
    RECT 213.1 51.55 213.31 51.62 ;
    RECT 213.1 51.91 213.31 51.98 ;
    RECT 210.24 51.19 210.45 51.26 ;
    RECT 210.24 51.55 210.45 51.62 ;
    RECT 210.24 51.91 210.45 51.98 ;
    RECT 209.78 51.19 209.99 51.26 ;
    RECT 209.78 51.55 209.99 51.62 ;
    RECT 209.78 51.91 209.99 51.98 ;
    RECT 206.92 51.19 207.13 51.26 ;
    RECT 206.92 51.55 207.13 51.62 ;
    RECT 206.92 51.91 207.13 51.98 ;
    RECT 206.46 51.19 206.67 51.26 ;
    RECT 206.46 51.55 206.67 51.62 ;
    RECT 206.46 51.91 206.67 51.98 ;
    RECT 203.6 51.19 203.81 51.26 ;
    RECT 203.6 51.55 203.81 51.62 ;
    RECT 203.6 51.91 203.81 51.98 ;
    RECT 203.14 51.19 203.35 51.26 ;
    RECT 203.14 51.55 203.35 51.62 ;
    RECT 203.14 51.91 203.35 51.98 ;
    RECT 200.28 51.19 200.49 51.26 ;
    RECT 200.28 51.55 200.49 51.62 ;
    RECT 200.28 51.91 200.49 51.98 ;
    RECT 199.82 51.19 200.03 51.26 ;
    RECT 199.82 51.55 200.03 51.62 ;
    RECT 199.82 51.91 200.03 51.98 ;
    RECT 196.96 51.19 197.17 51.26 ;
    RECT 196.96 51.55 197.17 51.62 ;
    RECT 196.96 51.91 197.17 51.98 ;
    RECT 196.5 51.19 196.71 51.26 ;
    RECT 196.5 51.55 196.71 51.62 ;
    RECT 196.5 51.91 196.71 51.98 ;
    RECT 193.64 51.19 193.85 51.26 ;
    RECT 193.64 51.55 193.85 51.62 ;
    RECT 193.64 51.91 193.85 51.98 ;
    RECT 193.18 51.19 193.39 51.26 ;
    RECT 193.18 51.55 193.39 51.62 ;
    RECT 193.18 51.91 193.39 51.98 ;
    RECT 190.32 51.19 190.53 51.26 ;
    RECT 190.32 51.55 190.53 51.62 ;
    RECT 190.32 51.91 190.53 51.98 ;
    RECT 189.86 51.19 190.07 51.26 ;
    RECT 189.86 51.55 190.07 51.62 ;
    RECT 189.86 51.91 190.07 51.98 ;
    RECT 187.0 51.19 187.21 51.26 ;
    RECT 187.0 51.55 187.21 51.62 ;
    RECT 187.0 51.91 187.21 51.98 ;
    RECT 186.54 51.19 186.75 51.26 ;
    RECT 186.54 51.55 186.75 51.62 ;
    RECT 186.54 51.91 186.75 51.98 ;
    RECT 183.68 51.19 183.89 51.26 ;
    RECT 183.68 51.55 183.89 51.62 ;
    RECT 183.68 51.91 183.89 51.98 ;
    RECT 183.22 51.19 183.43 51.26 ;
    RECT 183.22 51.55 183.43 51.62 ;
    RECT 183.22 51.91 183.43 51.98 ;
    RECT 147.485 51.55 147.555 51.62 ;
    RECT 266.68 51.19 266.89 51.26 ;
    RECT 266.68 51.55 266.89 51.62 ;
    RECT 266.68 51.91 266.89 51.98 ;
    RECT 266.22 51.19 266.43 51.26 ;
    RECT 266.22 51.55 266.43 51.62 ;
    RECT 266.22 51.91 266.43 51.98 ;
    RECT 263.36 51.19 263.57 51.26 ;
    RECT 263.36 51.55 263.57 51.62 ;
    RECT 263.36 51.91 263.57 51.98 ;
    RECT 262.9 51.19 263.11 51.26 ;
    RECT 262.9 51.55 263.11 51.62 ;
    RECT 262.9 51.91 263.11 51.98 ;
    RECT 260.04 51.19 260.25 51.26 ;
    RECT 260.04 51.55 260.25 51.62 ;
    RECT 260.04 51.91 260.25 51.98 ;
    RECT 259.58 51.19 259.79 51.26 ;
    RECT 259.58 51.55 259.79 51.62 ;
    RECT 259.58 51.91 259.79 51.98 ;
    RECT 256.72 51.19 256.93 51.26 ;
    RECT 256.72 51.55 256.93 51.62 ;
    RECT 256.72 51.91 256.93 51.98 ;
    RECT 256.26 51.19 256.47 51.26 ;
    RECT 256.26 51.55 256.47 51.62 ;
    RECT 256.26 51.91 256.47 51.98 ;
    RECT 253.4 51.19 253.61 51.26 ;
    RECT 253.4 51.55 253.61 51.62 ;
    RECT 253.4 51.91 253.61 51.98 ;
    RECT 252.94 51.19 253.15 51.26 ;
    RECT 252.94 51.55 253.15 51.62 ;
    RECT 252.94 51.91 253.15 51.98 ;
    RECT 250.08 87.21 250.29 87.28 ;
    RECT 250.08 87.57 250.29 87.64 ;
    RECT 250.08 87.93 250.29 88.0 ;
    RECT 249.62 87.21 249.83 87.28 ;
    RECT 249.62 87.57 249.83 87.64 ;
    RECT 249.62 87.93 249.83 88.0 ;
    RECT 246.76 87.21 246.97 87.28 ;
    RECT 246.76 87.57 246.97 87.64 ;
    RECT 246.76 87.93 246.97 88.0 ;
    RECT 246.3 87.21 246.51 87.28 ;
    RECT 246.3 87.57 246.51 87.64 ;
    RECT 246.3 87.93 246.51 88.0 ;
    RECT 243.44 87.21 243.65 87.28 ;
    RECT 243.44 87.57 243.65 87.64 ;
    RECT 243.44 87.93 243.65 88.0 ;
    RECT 242.98 87.21 243.19 87.28 ;
    RECT 242.98 87.57 243.19 87.64 ;
    RECT 242.98 87.93 243.19 88.0 ;
    RECT 240.12 87.21 240.33 87.28 ;
    RECT 240.12 87.57 240.33 87.64 ;
    RECT 240.12 87.93 240.33 88.0 ;
    RECT 239.66 87.21 239.87 87.28 ;
    RECT 239.66 87.57 239.87 87.64 ;
    RECT 239.66 87.93 239.87 88.0 ;
    RECT 236.8 87.21 237.01 87.28 ;
    RECT 236.8 87.57 237.01 87.64 ;
    RECT 236.8 87.93 237.01 88.0 ;
    RECT 236.34 87.21 236.55 87.28 ;
    RECT 236.34 87.57 236.55 87.64 ;
    RECT 236.34 87.93 236.55 88.0 ;
    RECT 233.48 87.21 233.69 87.28 ;
    RECT 233.48 87.57 233.69 87.64 ;
    RECT 233.48 87.93 233.69 88.0 ;
    RECT 233.02 87.21 233.23 87.28 ;
    RECT 233.02 87.57 233.23 87.64 ;
    RECT 233.02 87.93 233.23 88.0 ;
    RECT 230.16 87.21 230.37 87.28 ;
    RECT 230.16 87.57 230.37 87.64 ;
    RECT 230.16 87.93 230.37 88.0 ;
    RECT 229.7 87.21 229.91 87.28 ;
    RECT 229.7 87.57 229.91 87.64 ;
    RECT 229.7 87.93 229.91 88.0 ;
    RECT 226.84 87.21 227.05 87.28 ;
    RECT 226.84 87.57 227.05 87.64 ;
    RECT 226.84 87.93 227.05 88.0 ;
    RECT 226.38 87.21 226.59 87.28 ;
    RECT 226.38 87.57 226.59 87.64 ;
    RECT 226.38 87.93 226.59 88.0 ;
    RECT 223.52 87.21 223.73 87.28 ;
    RECT 223.52 87.57 223.73 87.64 ;
    RECT 223.52 87.93 223.73 88.0 ;
    RECT 223.06 87.21 223.27 87.28 ;
    RECT 223.06 87.57 223.27 87.64 ;
    RECT 223.06 87.93 223.27 88.0 ;
    RECT 220.2 87.21 220.41 87.28 ;
    RECT 220.2 87.57 220.41 87.64 ;
    RECT 220.2 87.93 220.41 88.0 ;
    RECT 219.74 87.21 219.95 87.28 ;
    RECT 219.74 87.57 219.95 87.64 ;
    RECT 219.74 87.93 219.95 88.0 ;
    RECT 216.88 87.21 217.09 87.28 ;
    RECT 216.88 87.57 217.09 87.64 ;
    RECT 216.88 87.93 217.09 88.0 ;
    RECT 216.42 87.21 216.63 87.28 ;
    RECT 216.42 87.57 216.63 87.64 ;
    RECT 216.42 87.93 216.63 88.0 ;
    RECT 267.91 87.57 267.98 87.64 ;
    RECT 180.36 87.21 180.57 87.28 ;
    RECT 180.36 87.57 180.57 87.64 ;
    RECT 180.36 87.93 180.57 88.0 ;
    RECT 179.9 87.21 180.11 87.28 ;
    RECT 179.9 87.57 180.11 87.64 ;
    RECT 179.9 87.93 180.11 88.0 ;
    RECT 177.04 87.21 177.25 87.28 ;
    RECT 177.04 87.57 177.25 87.64 ;
    RECT 177.04 87.93 177.25 88.0 ;
    RECT 176.58 87.21 176.79 87.28 ;
    RECT 176.58 87.57 176.79 87.64 ;
    RECT 176.58 87.93 176.79 88.0 ;
    RECT 173.72 87.21 173.93 87.28 ;
    RECT 173.72 87.57 173.93 87.64 ;
    RECT 173.72 87.93 173.93 88.0 ;
    RECT 173.26 87.21 173.47 87.28 ;
    RECT 173.26 87.57 173.47 87.64 ;
    RECT 173.26 87.93 173.47 88.0 ;
    RECT 170.4 87.21 170.61 87.28 ;
    RECT 170.4 87.57 170.61 87.64 ;
    RECT 170.4 87.93 170.61 88.0 ;
    RECT 169.94 87.21 170.15 87.28 ;
    RECT 169.94 87.57 170.15 87.64 ;
    RECT 169.94 87.93 170.15 88.0 ;
    RECT 167.08 87.21 167.29 87.28 ;
    RECT 167.08 87.57 167.29 87.64 ;
    RECT 167.08 87.93 167.29 88.0 ;
    RECT 166.62 87.21 166.83 87.28 ;
    RECT 166.62 87.57 166.83 87.64 ;
    RECT 166.62 87.93 166.83 88.0 ;
    RECT 163.76 87.21 163.97 87.28 ;
    RECT 163.76 87.57 163.97 87.64 ;
    RECT 163.76 87.93 163.97 88.0 ;
    RECT 163.3 87.21 163.51 87.28 ;
    RECT 163.3 87.57 163.51 87.64 ;
    RECT 163.3 87.93 163.51 88.0 ;
    RECT 160.44 87.21 160.65 87.28 ;
    RECT 160.44 87.57 160.65 87.64 ;
    RECT 160.44 87.93 160.65 88.0 ;
    RECT 159.98 87.21 160.19 87.28 ;
    RECT 159.98 87.57 160.19 87.64 ;
    RECT 159.98 87.93 160.19 88.0 ;
    RECT 157.12 87.21 157.33 87.28 ;
    RECT 157.12 87.57 157.33 87.64 ;
    RECT 157.12 87.93 157.33 88.0 ;
    RECT 156.66 87.21 156.87 87.28 ;
    RECT 156.66 87.57 156.87 87.64 ;
    RECT 156.66 87.93 156.87 88.0 ;
    RECT 153.8 87.21 154.01 87.28 ;
    RECT 153.8 87.57 154.01 87.64 ;
    RECT 153.8 87.93 154.01 88.0 ;
    RECT 153.34 87.21 153.55 87.28 ;
    RECT 153.34 87.57 153.55 87.64 ;
    RECT 153.34 87.93 153.55 88.0 ;
    RECT 150.48 87.21 150.69 87.28 ;
    RECT 150.48 87.57 150.69 87.64 ;
    RECT 150.48 87.93 150.69 88.0 ;
    RECT 150.02 87.21 150.23 87.28 ;
    RECT 150.02 87.57 150.23 87.64 ;
    RECT 150.02 87.93 150.23 88.0 ;
    RECT 213.56 87.21 213.77 87.28 ;
    RECT 213.56 87.57 213.77 87.64 ;
    RECT 213.56 87.93 213.77 88.0 ;
    RECT 213.1 87.21 213.31 87.28 ;
    RECT 213.1 87.57 213.31 87.64 ;
    RECT 213.1 87.93 213.31 88.0 ;
    RECT 210.24 87.21 210.45 87.28 ;
    RECT 210.24 87.57 210.45 87.64 ;
    RECT 210.24 87.93 210.45 88.0 ;
    RECT 209.78 87.21 209.99 87.28 ;
    RECT 209.78 87.57 209.99 87.64 ;
    RECT 209.78 87.93 209.99 88.0 ;
    RECT 206.92 87.21 207.13 87.28 ;
    RECT 206.92 87.57 207.13 87.64 ;
    RECT 206.92 87.93 207.13 88.0 ;
    RECT 206.46 87.21 206.67 87.28 ;
    RECT 206.46 87.57 206.67 87.64 ;
    RECT 206.46 87.93 206.67 88.0 ;
    RECT 203.6 87.21 203.81 87.28 ;
    RECT 203.6 87.57 203.81 87.64 ;
    RECT 203.6 87.93 203.81 88.0 ;
    RECT 203.14 87.21 203.35 87.28 ;
    RECT 203.14 87.57 203.35 87.64 ;
    RECT 203.14 87.93 203.35 88.0 ;
    RECT 200.28 87.21 200.49 87.28 ;
    RECT 200.28 87.57 200.49 87.64 ;
    RECT 200.28 87.93 200.49 88.0 ;
    RECT 199.82 87.21 200.03 87.28 ;
    RECT 199.82 87.57 200.03 87.64 ;
    RECT 199.82 87.93 200.03 88.0 ;
    RECT 196.96 87.21 197.17 87.28 ;
    RECT 196.96 87.57 197.17 87.64 ;
    RECT 196.96 87.93 197.17 88.0 ;
    RECT 196.5 87.21 196.71 87.28 ;
    RECT 196.5 87.57 196.71 87.64 ;
    RECT 196.5 87.93 196.71 88.0 ;
    RECT 193.64 87.21 193.85 87.28 ;
    RECT 193.64 87.57 193.85 87.64 ;
    RECT 193.64 87.93 193.85 88.0 ;
    RECT 193.18 87.21 193.39 87.28 ;
    RECT 193.18 87.57 193.39 87.64 ;
    RECT 193.18 87.93 193.39 88.0 ;
    RECT 190.32 87.21 190.53 87.28 ;
    RECT 190.32 87.57 190.53 87.64 ;
    RECT 190.32 87.93 190.53 88.0 ;
    RECT 189.86 87.21 190.07 87.28 ;
    RECT 189.86 87.57 190.07 87.64 ;
    RECT 189.86 87.93 190.07 88.0 ;
    RECT 187.0 87.21 187.21 87.28 ;
    RECT 187.0 87.57 187.21 87.64 ;
    RECT 187.0 87.93 187.21 88.0 ;
    RECT 186.54 87.21 186.75 87.28 ;
    RECT 186.54 87.57 186.75 87.64 ;
    RECT 186.54 87.93 186.75 88.0 ;
    RECT 183.68 87.21 183.89 87.28 ;
    RECT 183.68 87.57 183.89 87.64 ;
    RECT 183.68 87.93 183.89 88.0 ;
    RECT 183.22 87.21 183.43 87.28 ;
    RECT 183.22 87.57 183.43 87.64 ;
    RECT 183.22 87.93 183.43 88.0 ;
    RECT 147.485 87.57 147.555 87.64 ;
    RECT 266.68 87.21 266.89 87.28 ;
    RECT 266.68 87.57 266.89 87.64 ;
    RECT 266.68 87.93 266.89 88.0 ;
    RECT 266.22 87.21 266.43 87.28 ;
    RECT 266.22 87.57 266.43 87.64 ;
    RECT 266.22 87.93 266.43 88.0 ;
    RECT 263.36 87.21 263.57 87.28 ;
    RECT 263.36 87.57 263.57 87.64 ;
    RECT 263.36 87.93 263.57 88.0 ;
    RECT 262.9 87.21 263.11 87.28 ;
    RECT 262.9 87.57 263.11 87.64 ;
    RECT 262.9 87.93 263.11 88.0 ;
    RECT 260.04 87.21 260.25 87.28 ;
    RECT 260.04 87.57 260.25 87.64 ;
    RECT 260.04 87.93 260.25 88.0 ;
    RECT 259.58 87.21 259.79 87.28 ;
    RECT 259.58 87.57 259.79 87.64 ;
    RECT 259.58 87.93 259.79 88.0 ;
    RECT 256.72 87.21 256.93 87.28 ;
    RECT 256.72 87.57 256.93 87.64 ;
    RECT 256.72 87.93 256.93 88.0 ;
    RECT 256.26 87.21 256.47 87.28 ;
    RECT 256.26 87.57 256.47 87.64 ;
    RECT 256.26 87.93 256.47 88.0 ;
    RECT 253.4 87.21 253.61 87.28 ;
    RECT 253.4 87.57 253.61 87.64 ;
    RECT 253.4 87.93 253.61 88.0 ;
    RECT 252.94 87.21 253.15 87.28 ;
    RECT 252.94 87.57 253.15 87.64 ;
    RECT 252.94 87.93 253.15 88.0 ;
    RECT 250.08 50.47 250.29 50.54 ;
    RECT 250.08 50.83 250.29 50.9 ;
    RECT 250.08 51.19 250.29 51.26 ;
    RECT 249.62 50.47 249.83 50.54 ;
    RECT 249.62 50.83 249.83 50.9 ;
    RECT 249.62 51.19 249.83 51.26 ;
    RECT 246.76 50.47 246.97 50.54 ;
    RECT 246.76 50.83 246.97 50.9 ;
    RECT 246.76 51.19 246.97 51.26 ;
    RECT 246.3 50.47 246.51 50.54 ;
    RECT 246.3 50.83 246.51 50.9 ;
    RECT 246.3 51.19 246.51 51.26 ;
    RECT 243.44 50.47 243.65 50.54 ;
    RECT 243.44 50.83 243.65 50.9 ;
    RECT 243.44 51.19 243.65 51.26 ;
    RECT 242.98 50.47 243.19 50.54 ;
    RECT 242.98 50.83 243.19 50.9 ;
    RECT 242.98 51.19 243.19 51.26 ;
    RECT 240.12 50.47 240.33 50.54 ;
    RECT 240.12 50.83 240.33 50.9 ;
    RECT 240.12 51.19 240.33 51.26 ;
    RECT 239.66 50.47 239.87 50.54 ;
    RECT 239.66 50.83 239.87 50.9 ;
    RECT 239.66 51.19 239.87 51.26 ;
    RECT 236.8 50.47 237.01 50.54 ;
    RECT 236.8 50.83 237.01 50.9 ;
    RECT 236.8 51.19 237.01 51.26 ;
    RECT 236.34 50.47 236.55 50.54 ;
    RECT 236.34 50.83 236.55 50.9 ;
    RECT 236.34 51.19 236.55 51.26 ;
    RECT 233.48 50.47 233.69 50.54 ;
    RECT 233.48 50.83 233.69 50.9 ;
    RECT 233.48 51.19 233.69 51.26 ;
    RECT 233.02 50.47 233.23 50.54 ;
    RECT 233.02 50.83 233.23 50.9 ;
    RECT 233.02 51.19 233.23 51.26 ;
    RECT 230.16 50.47 230.37 50.54 ;
    RECT 230.16 50.83 230.37 50.9 ;
    RECT 230.16 51.19 230.37 51.26 ;
    RECT 229.7 50.47 229.91 50.54 ;
    RECT 229.7 50.83 229.91 50.9 ;
    RECT 229.7 51.19 229.91 51.26 ;
    RECT 226.84 50.47 227.05 50.54 ;
    RECT 226.84 50.83 227.05 50.9 ;
    RECT 226.84 51.19 227.05 51.26 ;
    RECT 226.38 50.47 226.59 50.54 ;
    RECT 226.38 50.83 226.59 50.9 ;
    RECT 226.38 51.19 226.59 51.26 ;
    RECT 223.52 50.47 223.73 50.54 ;
    RECT 223.52 50.83 223.73 50.9 ;
    RECT 223.52 51.19 223.73 51.26 ;
    RECT 223.06 50.47 223.27 50.54 ;
    RECT 223.06 50.83 223.27 50.9 ;
    RECT 223.06 51.19 223.27 51.26 ;
    RECT 220.2 50.47 220.41 50.54 ;
    RECT 220.2 50.83 220.41 50.9 ;
    RECT 220.2 51.19 220.41 51.26 ;
    RECT 219.74 50.47 219.95 50.54 ;
    RECT 219.74 50.83 219.95 50.9 ;
    RECT 219.74 51.19 219.95 51.26 ;
    RECT 216.88 50.47 217.09 50.54 ;
    RECT 216.88 50.83 217.09 50.9 ;
    RECT 216.88 51.19 217.09 51.26 ;
    RECT 216.42 50.47 216.63 50.54 ;
    RECT 216.42 50.83 216.63 50.9 ;
    RECT 216.42 51.19 216.63 51.26 ;
    RECT 267.91 50.83 267.98 50.9 ;
    RECT 180.36 50.47 180.57 50.54 ;
    RECT 180.36 50.83 180.57 50.9 ;
    RECT 180.36 51.19 180.57 51.26 ;
    RECT 179.9 50.47 180.11 50.54 ;
    RECT 179.9 50.83 180.11 50.9 ;
    RECT 179.9 51.19 180.11 51.26 ;
    RECT 177.04 50.47 177.25 50.54 ;
    RECT 177.04 50.83 177.25 50.9 ;
    RECT 177.04 51.19 177.25 51.26 ;
    RECT 176.58 50.47 176.79 50.54 ;
    RECT 176.58 50.83 176.79 50.9 ;
    RECT 176.58 51.19 176.79 51.26 ;
    RECT 173.72 50.47 173.93 50.54 ;
    RECT 173.72 50.83 173.93 50.9 ;
    RECT 173.72 51.19 173.93 51.26 ;
    RECT 173.26 50.47 173.47 50.54 ;
    RECT 173.26 50.83 173.47 50.9 ;
    RECT 173.26 51.19 173.47 51.26 ;
    RECT 170.4 50.47 170.61 50.54 ;
    RECT 170.4 50.83 170.61 50.9 ;
    RECT 170.4 51.19 170.61 51.26 ;
    RECT 169.94 50.47 170.15 50.54 ;
    RECT 169.94 50.83 170.15 50.9 ;
    RECT 169.94 51.19 170.15 51.26 ;
    RECT 167.08 50.47 167.29 50.54 ;
    RECT 167.08 50.83 167.29 50.9 ;
    RECT 167.08 51.19 167.29 51.26 ;
    RECT 166.62 50.47 166.83 50.54 ;
    RECT 166.62 50.83 166.83 50.9 ;
    RECT 166.62 51.19 166.83 51.26 ;
    RECT 163.76 50.47 163.97 50.54 ;
    RECT 163.76 50.83 163.97 50.9 ;
    RECT 163.76 51.19 163.97 51.26 ;
    RECT 163.3 50.47 163.51 50.54 ;
    RECT 163.3 50.83 163.51 50.9 ;
    RECT 163.3 51.19 163.51 51.26 ;
    RECT 160.44 50.47 160.65 50.54 ;
    RECT 160.44 50.83 160.65 50.9 ;
    RECT 160.44 51.19 160.65 51.26 ;
    RECT 159.98 50.47 160.19 50.54 ;
    RECT 159.98 50.83 160.19 50.9 ;
    RECT 159.98 51.19 160.19 51.26 ;
    RECT 157.12 50.47 157.33 50.54 ;
    RECT 157.12 50.83 157.33 50.9 ;
    RECT 157.12 51.19 157.33 51.26 ;
    RECT 156.66 50.47 156.87 50.54 ;
    RECT 156.66 50.83 156.87 50.9 ;
    RECT 156.66 51.19 156.87 51.26 ;
    RECT 153.8 50.47 154.01 50.54 ;
    RECT 153.8 50.83 154.01 50.9 ;
    RECT 153.8 51.19 154.01 51.26 ;
    RECT 153.34 50.47 153.55 50.54 ;
    RECT 153.34 50.83 153.55 50.9 ;
    RECT 153.34 51.19 153.55 51.26 ;
    RECT 150.48 50.47 150.69 50.54 ;
    RECT 150.48 50.83 150.69 50.9 ;
    RECT 150.48 51.19 150.69 51.26 ;
    RECT 150.02 50.47 150.23 50.54 ;
    RECT 150.02 50.83 150.23 50.9 ;
    RECT 150.02 51.19 150.23 51.26 ;
    RECT 213.56 50.47 213.77 50.54 ;
    RECT 213.56 50.83 213.77 50.9 ;
    RECT 213.56 51.19 213.77 51.26 ;
    RECT 213.1 50.47 213.31 50.54 ;
    RECT 213.1 50.83 213.31 50.9 ;
    RECT 213.1 51.19 213.31 51.26 ;
    RECT 210.24 50.47 210.45 50.54 ;
    RECT 210.24 50.83 210.45 50.9 ;
    RECT 210.24 51.19 210.45 51.26 ;
    RECT 209.78 50.47 209.99 50.54 ;
    RECT 209.78 50.83 209.99 50.9 ;
    RECT 209.78 51.19 209.99 51.26 ;
    RECT 206.92 50.47 207.13 50.54 ;
    RECT 206.92 50.83 207.13 50.9 ;
    RECT 206.92 51.19 207.13 51.26 ;
    RECT 206.46 50.47 206.67 50.54 ;
    RECT 206.46 50.83 206.67 50.9 ;
    RECT 206.46 51.19 206.67 51.26 ;
    RECT 203.6 50.47 203.81 50.54 ;
    RECT 203.6 50.83 203.81 50.9 ;
    RECT 203.6 51.19 203.81 51.26 ;
    RECT 203.14 50.47 203.35 50.54 ;
    RECT 203.14 50.83 203.35 50.9 ;
    RECT 203.14 51.19 203.35 51.26 ;
    RECT 200.28 50.47 200.49 50.54 ;
    RECT 200.28 50.83 200.49 50.9 ;
    RECT 200.28 51.19 200.49 51.26 ;
    RECT 199.82 50.47 200.03 50.54 ;
    RECT 199.82 50.83 200.03 50.9 ;
    RECT 199.82 51.19 200.03 51.26 ;
    RECT 196.96 50.47 197.17 50.54 ;
    RECT 196.96 50.83 197.17 50.9 ;
    RECT 196.96 51.19 197.17 51.26 ;
    RECT 196.5 50.47 196.71 50.54 ;
    RECT 196.5 50.83 196.71 50.9 ;
    RECT 196.5 51.19 196.71 51.26 ;
    RECT 193.64 50.47 193.85 50.54 ;
    RECT 193.64 50.83 193.85 50.9 ;
    RECT 193.64 51.19 193.85 51.26 ;
    RECT 193.18 50.47 193.39 50.54 ;
    RECT 193.18 50.83 193.39 50.9 ;
    RECT 193.18 51.19 193.39 51.26 ;
    RECT 190.32 50.47 190.53 50.54 ;
    RECT 190.32 50.83 190.53 50.9 ;
    RECT 190.32 51.19 190.53 51.26 ;
    RECT 189.86 50.47 190.07 50.54 ;
    RECT 189.86 50.83 190.07 50.9 ;
    RECT 189.86 51.19 190.07 51.26 ;
    RECT 187.0 50.47 187.21 50.54 ;
    RECT 187.0 50.83 187.21 50.9 ;
    RECT 187.0 51.19 187.21 51.26 ;
    RECT 186.54 50.47 186.75 50.54 ;
    RECT 186.54 50.83 186.75 50.9 ;
    RECT 186.54 51.19 186.75 51.26 ;
    RECT 183.68 50.47 183.89 50.54 ;
    RECT 183.68 50.83 183.89 50.9 ;
    RECT 183.68 51.19 183.89 51.26 ;
    RECT 183.22 50.47 183.43 50.54 ;
    RECT 183.22 50.83 183.43 50.9 ;
    RECT 183.22 51.19 183.43 51.26 ;
    RECT 147.485 50.83 147.555 50.9 ;
    RECT 266.68 50.47 266.89 50.54 ;
    RECT 266.68 50.83 266.89 50.9 ;
    RECT 266.68 51.19 266.89 51.26 ;
    RECT 266.22 50.47 266.43 50.54 ;
    RECT 266.22 50.83 266.43 50.9 ;
    RECT 266.22 51.19 266.43 51.26 ;
    RECT 263.36 50.47 263.57 50.54 ;
    RECT 263.36 50.83 263.57 50.9 ;
    RECT 263.36 51.19 263.57 51.26 ;
    RECT 262.9 50.47 263.11 50.54 ;
    RECT 262.9 50.83 263.11 50.9 ;
    RECT 262.9 51.19 263.11 51.26 ;
    RECT 260.04 50.47 260.25 50.54 ;
    RECT 260.04 50.83 260.25 50.9 ;
    RECT 260.04 51.19 260.25 51.26 ;
    RECT 259.58 50.47 259.79 50.54 ;
    RECT 259.58 50.83 259.79 50.9 ;
    RECT 259.58 51.19 259.79 51.26 ;
    RECT 256.72 50.47 256.93 50.54 ;
    RECT 256.72 50.83 256.93 50.9 ;
    RECT 256.72 51.19 256.93 51.26 ;
    RECT 256.26 50.47 256.47 50.54 ;
    RECT 256.26 50.83 256.47 50.9 ;
    RECT 256.26 51.19 256.47 51.26 ;
    RECT 253.4 50.47 253.61 50.54 ;
    RECT 253.4 50.83 253.61 50.9 ;
    RECT 253.4 51.19 253.61 51.26 ;
    RECT 252.94 50.47 253.15 50.54 ;
    RECT 252.94 50.83 253.15 50.9 ;
    RECT 252.94 51.19 253.15 51.26 ;
    RECT 250.08 49.75 250.29 49.82 ;
    RECT 250.08 50.11 250.29 50.18 ;
    RECT 250.08 50.47 250.29 50.54 ;
    RECT 249.62 49.75 249.83 49.82 ;
    RECT 249.62 50.11 249.83 50.18 ;
    RECT 249.62 50.47 249.83 50.54 ;
    RECT 246.76 49.75 246.97 49.82 ;
    RECT 246.76 50.11 246.97 50.18 ;
    RECT 246.76 50.47 246.97 50.54 ;
    RECT 246.3 49.75 246.51 49.82 ;
    RECT 246.3 50.11 246.51 50.18 ;
    RECT 246.3 50.47 246.51 50.54 ;
    RECT 243.44 49.75 243.65 49.82 ;
    RECT 243.44 50.11 243.65 50.18 ;
    RECT 243.44 50.47 243.65 50.54 ;
    RECT 242.98 49.75 243.19 49.82 ;
    RECT 242.98 50.11 243.19 50.18 ;
    RECT 242.98 50.47 243.19 50.54 ;
    RECT 240.12 49.75 240.33 49.82 ;
    RECT 240.12 50.11 240.33 50.18 ;
    RECT 240.12 50.47 240.33 50.54 ;
    RECT 239.66 49.75 239.87 49.82 ;
    RECT 239.66 50.11 239.87 50.18 ;
    RECT 239.66 50.47 239.87 50.54 ;
    RECT 236.8 49.75 237.01 49.82 ;
    RECT 236.8 50.11 237.01 50.18 ;
    RECT 236.8 50.47 237.01 50.54 ;
    RECT 236.34 49.75 236.55 49.82 ;
    RECT 236.34 50.11 236.55 50.18 ;
    RECT 236.34 50.47 236.55 50.54 ;
    RECT 233.48 49.75 233.69 49.82 ;
    RECT 233.48 50.11 233.69 50.18 ;
    RECT 233.48 50.47 233.69 50.54 ;
    RECT 233.02 49.75 233.23 49.82 ;
    RECT 233.02 50.11 233.23 50.18 ;
    RECT 233.02 50.47 233.23 50.54 ;
    RECT 230.16 49.75 230.37 49.82 ;
    RECT 230.16 50.11 230.37 50.18 ;
    RECT 230.16 50.47 230.37 50.54 ;
    RECT 229.7 49.75 229.91 49.82 ;
    RECT 229.7 50.11 229.91 50.18 ;
    RECT 229.7 50.47 229.91 50.54 ;
    RECT 226.84 49.75 227.05 49.82 ;
    RECT 226.84 50.11 227.05 50.18 ;
    RECT 226.84 50.47 227.05 50.54 ;
    RECT 226.38 49.75 226.59 49.82 ;
    RECT 226.38 50.11 226.59 50.18 ;
    RECT 226.38 50.47 226.59 50.54 ;
    RECT 223.52 49.75 223.73 49.82 ;
    RECT 223.52 50.11 223.73 50.18 ;
    RECT 223.52 50.47 223.73 50.54 ;
    RECT 223.06 49.75 223.27 49.82 ;
    RECT 223.06 50.11 223.27 50.18 ;
    RECT 223.06 50.47 223.27 50.54 ;
    RECT 220.2 49.75 220.41 49.82 ;
    RECT 220.2 50.11 220.41 50.18 ;
    RECT 220.2 50.47 220.41 50.54 ;
    RECT 219.74 49.75 219.95 49.82 ;
    RECT 219.74 50.11 219.95 50.18 ;
    RECT 219.74 50.47 219.95 50.54 ;
    RECT 216.88 49.75 217.09 49.82 ;
    RECT 216.88 50.11 217.09 50.18 ;
    RECT 216.88 50.47 217.09 50.54 ;
    RECT 216.42 49.75 216.63 49.82 ;
    RECT 216.42 50.11 216.63 50.18 ;
    RECT 216.42 50.47 216.63 50.54 ;
    RECT 267.91 50.11 267.98 50.18 ;
    RECT 180.36 49.75 180.57 49.82 ;
    RECT 180.36 50.11 180.57 50.18 ;
    RECT 180.36 50.47 180.57 50.54 ;
    RECT 179.9 49.75 180.11 49.82 ;
    RECT 179.9 50.11 180.11 50.18 ;
    RECT 179.9 50.47 180.11 50.54 ;
    RECT 177.04 49.75 177.25 49.82 ;
    RECT 177.04 50.11 177.25 50.18 ;
    RECT 177.04 50.47 177.25 50.54 ;
    RECT 176.58 49.75 176.79 49.82 ;
    RECT 176.58 50.11 176.79 50.18 ;
    RECT 176.58 50.47 176.79 50.54 ;
    RECT 173.72 49.75 173.93 49.82 ;
    RECT 173.72 50.11 173.93 50.18 ;
    RECT 173.72 50.47 173.93 50.54 ;
    RECT 173.26 49.75 173.47 49.82 ;
    RECT 173.26 50.11 173.47 50.18 ;
    RECT 173.26 50.47 173.47 50.54 ;
    RECT 170.4 49.75 170.61 49.82 ;
    RECT 170.4 50.11 170.61 50.18 ;
    RECT 170.4 50.47 170.61 50.54 ;
    RECT 169.94 49.75 170.15 49.82 ;
    RECT 169.94 50.11 170.15 50.18 ;
    RECT 169.94 50.47 170.15 50.54 ;
    RECT 167.08 49.75 167.29 49.82 ;
    RECT 167.08 50.11 167.29 50.18 ;
    RECT 167.08 50.47 167.29 50.54 ;
    RECT 166.62 49.75 166.83 49.82 ;
    RECT 166.62 50.11 166.83 50.18 ;
    RECT 166.62 50.47 166.83 50.54 ;
    RECT 163.76 49.75 163.97 49.82 ;
    RECT 163.76 50.11 163.97 50.18 ;
    RECT 163.76 50.47 163.97 50.54 ;
    RECT 163.3 49.75 163.51 49.82 ;
    RECT 163.3 50.11 163.51 50.18 ;
    RECT 163.3 50.47 163.51 50.54 ;
    RECT 160.44 49.75 160.65 49.82 ;
    RECT 160.44 50.11 160.65 50.18 ;
    RECT 160.44 50.47 160.65 50.54 ;
    RECT 159.98 49.75 160.19 49.82 ;
    RECT 159.98 50.11 160.19 50.18 ;
    RECT 159.98 50.47 160.19 50.54 ;
    RECT 157.12 49.75 157.33 49.82 ;
    RECT 157.12 50.11 157.33 50.18 ;
    RECT 157.12 50.47 157.33 50.54 ;
    RECT 156.66 49.75 156.87 49.82 ;
    RECT 156.66 50.11 156.87 50.18 ;
    RECT 156.66 50.47 156.87 50.54 ;
    RECT 153.8 49.75 154.01 49.82 ;
    RECT 153.8 50.11 154.01 50.18 ;
    RECT 153.8 50.47 154.01 50.54 ;
    RECT 153.34 49.75 153.55 49.82 ;
    RECT 153.34 50.11 153.55 50.18 ;
    RECT 153.34 50.47 153.55 50.54 ;
    RECT 150.48 49.75 150.69 49.82 ;
    RECT 150.48 50.11 150.69 50.18 ;
    RECT 150.48 50.47 150.69 50.54 ;
    RECT 150.02 49.75 150.23 49.82 ;
    RECT 150.02 50.11 150.23 50.18 ;
    RECT 150.02 50.47 150.23 50.54 ;
    RECT 213.56 49.75 213.77 49.82 ;
    RECT 213.56 50.11 213.77 50.18 ;
    RECT 213.56 50.47 213.77 50.54 ;
    RECT 213.1 49.75 213.31 49.82 ;
    RECT 213.1 50.11 213.31 50.18 ;
    RECT 213.1 50.47 213.31 50.54 ;
    RECT 210.24 49.75 210.45 49.82 ;
    RECT 210.24 50.11 210.45 50.18 ;
    RECT 210.24 50.47 210.45 50.54 ;
    RECT 209.78 49.75 209.99 49.82 ;
    RECT 209.78 50.11 209.99 50.18 ;
    RECT 209.78 50.47 209.99 50.54 ;
    RECT 206.92 49.75 207.13 49.82 ;
    RECT 206.92 50.11 207.13 50.18 ;
    RECT 206.92 50.47 207.13 50.54 ;
    RECT 206.46 49.75 206.67 49.82 ;
    RECT 206.46 50.11 206.67 50.18 ;
    RECT 206.46 50.47 206.67 50.54 ;
    RECT 203.6 49.75 203.81 49.82 ;
    RECT 203.6 50.11 203.81 50.18 ;
    RECT 203.6 50.47 203.81 50.54 ;
    RECT 203.14 49.75 203.35 49.82 ;
    RECT 203.14 50.11 203.35 50.18 ;
    RECT 203.14 50.47 203.35 50.54 ;
    RECT 200.28 49.75 200.49 49.82 ;
    RECT 200.28 50.11 200.49 50.18 ;
    RECT 200.28 50.47 200.49 50.54 ;
    RECT 199.82 49.75 200.03 49.82 ;
    RECT 199.82 50.11 200.03 50.18 ;
    RECT 199.82 50.47 200.03 50.54 ;
    RECT 196.96 49.75 197.17 49.82 ;
    RECT 196.96 50.11 197.17 50.18 ;
    RECT 196.96 50.47 197.17 50.54 ;
    RECT 196.5 49.75 196.71 49.82 ;
    RECT 196.5 50.11 196.71 50.18 ;
    RECT 196.5 50.47 196.71 50.54 ;
    RECT 193.64 49.75 193.85 49.82 ;
    RECT 193.64 50.11 193.85 50.18 ;
    RECT 193.64 50.47 193.85 50.54 ;
    RECT 193.18 49.75 193.39 49.82 ;
    RECT 193.18 50.11 193.39 50.18 ;
    RECT 193.18 50.47 193.39 50.54 ;
    RECT 190.32 49.75 190.53 49.82 ;
    RECT 190.32 50.11 190.53 50.18 ;
    RECT 190.32 50.47 190.53 50.54 ;
    RECT 189.86 49.75 190.07 49.82 ;
    RECT 189.86 50.11 190.07 50.18 ;
    RECT 189.86 50.47 190.07 50.54 ;
    RECT 187.0 49.75 187.21 49.82 ;
    RECT 187.0 50.11 187.21 50.18 ;
    RECT 187.0 50.47 187.21 50.54 ;
    RECT 186.54 49.75 186.75 49.82 ;
    RECT 186.54 50.11 186.75 50.18 ;
    RECT 186.54 50.47 186.75 50.54 ;
    RECT 183.68 49.75 183.89 49.82 ;
    RECT 183.68 50.11 183.89 50.18 ;
    RECT 183.68 50.47 183.89 50.54 ;
    RECT 183.22 49.75 183.43 49.82 ;
    RECT 183.22 50.11 183.43 50.18 ;
    RECT 183.22 50.47 183.43 50.54 ;
    RECT 147.485 50.11 147.555 50.18 ;
    RECT 266.68 49.75 266.89 49.82 ;
    RECT 266.68 50.11 266.89 50.18 ;
    RECT 266.68 50.47 266.89 50.54 ;
    RECT 266.22 49.75 266.43 49.82 ;
    RECT 266.22 50.11 266.43 50.18 ;
    RECT 266.22 50.47 266.43 50.54 ;
    RECT 263.36 49.75 263.57 49.82 ;
    RECT 263.36 50.11 263.57 50.18 ;
    RECT 263.36 50.47 263.57 50.54 ;
    RECT 262.9 49.75 263.11 49.82 ;
    RECT 262.9 50.11 263.11 50.18 ;
    RECT 262.9 50.47 263.11 50.54 ;
    RECT 260.04 49.75 260.25 49.82 ;
    RECT 260.04 50.11 260.25 50.18 ;
    RECT 260.04 50.47 260.25 50.54 ;
    RECT 259.58 49.75 259.79 49.82 ;
    RECT 259.58 50.11 259.79 50.18 ;
    RECT 259.58 50.47 259.79 50.54 ;
    RECT 256.72 49.75 256.93 49.82 ;
    RECT 256.72 50.11 256.93 50.18 ;
    RECT 256.72 50.47 256.93 50.54 ;
    RECT 256.26 49.75 256.47 49.82 ;
    RECT 256.26 50.11 256.47 50.18 ;
    RECT 256.26 50.47 256.47 50.54 ;
    RECT 253.4 49.75 253.61 49.82 ;
    RECT 253.4 50.11 253.61 50.18 ;
    RECT 253.4 50.47 253.61 50.54 ;
    RECT 252.94 49.75 253.15 49.82 ;
    RECT 252.94 50.11 253.15 50.18 ;
    RECT 252.94 50.47 253.15 50.54 ;
    RECT 250.08 49.03 250.29 49.1 ;
    RECT 250.08 49.39 250.29 49.46 ;
    RECT 250.08 49.75 250.29 49.82 ;
    RECT 249.62 49.03 249.83 49.1 ;
    RECT 249.62 49.39 249.83 49.46 ;
    RECT 249.62 49.75 249.83 49.82 ;
    RECT 246.76 49.03 246.97 49.1 ;
    RECT 246.76 49.39 246.97 49.46 ;
    RECT 246.76 49.75 246.97 49.82 ;
    RECT 246.3 49.03 246.51 49.1 ;
    RECT 246.3 49.39 246.51 49.46 ;
    RECT 246.3 49.75 246.51 49.82 ;
    RECT 243.44 49.03 243.65 49.1 ;
    RECT 243.44 49.39 243.65 49.46 ;
    RECT 243.44 49.75 243.65 49.82 ;
    RECT 242.98 49.03 243.19 49.1 ;
    RECT 242.98 49.39 243.19 49.46 ;
    RECT 242.98 49.75 243.19 49.82 ;
    RECT 240.12 49.03 240.33 49.1 ;
    RECT 240.12 49.39 240.33 49.46 ;
    RECT 240.12 49.75 240.33 49.82 ;
    RECT 239.66 49.03 239.87 49.1 ;
    RECT 239.66 49.39 239.87 49.46 ;
    RECT 239.66 49.75 239.87 49.82 ;
    RECT 236.8 49.03 237.01 49.1 ;
    RECT 236.8 49.39 237.01 49.46 ;
    RECT 236.8 49.75 237.01 49.82 ;
    RECT 236.34 49.03 236.55 49.1 ;
    RECT 236.34 49.39 236.55 49.46 ;
    RECT 236.34 49.75 236.55 49.82 ;
    RECT 233.48 49.03 233.69 49.1 ;
    RECT 233.48 49.39 233.69 49.46 ;
    RECT 233.48 49.75 233.69 49.82 ;
    RECT 233.02 49.03 233.23 49.1 ;
    RECT 233.02 49.39 233.23 49.46 ;
    RECT 233.02 49.75 233.23 49.82 ;
    RECT 230.16 49.03 230.37 49.1 ;
    RECT 230.16 49.39 230.37 49.46 ;
    RECT 230.16 49.75 230.37 49.82 ;
    RECT 229.7 49.03 229.91 49.1 ;
    RECT 229.7 49.39 229.91 49.46 ;
    RECT 229.7 49.75 229.91 49.82 ;
    RECT 226.84 49.03 227.05 49.1 ;
    RECT 226.84 49.39 227.05 49.46 ;
    RECT 226.84 49.75 227.05 49.82 ;
    RECT 226.38 49.03 226.59 49.1 ;
    RECT 226.38 49.39 226.59 49.46 ;
    RECT 226.38 49.75 226.59 49.82 ;
    RECT 223.52 49.03 223.73 49.1 ;
    RECT 223.52 49.39 223.73 49.46 ;
    RECT 223.52 49.75 223.73 49.82 ;
    RECT 223.06 49.03 223.27 49.1 ;
    RECT 223.06 49.39 223.27 49.46 ;
    RECT 223.06 49.75 223.27 49.82 ;
    RECT 220.2 49.03 220.41 49.1 ;
    RECT 220.2 49.39 220.41 49.46 ;
    RECT 220.2 49.75 220.41 49.82 ;
    RECT 219.74 49.03 219.95 49.1 ;
    RECT 219.74 49.39 219.95 49.46 ;
    RECT 219.74 49.75 219.95 49.82 ;
    RECT 216.88 49.03 217.09 49.1 ;
    RECT 216.88 49.39 217.09 49.46 ;
    RECT 216.88 49.75 217.09 49.82 ;
    RECT 216.42 49.03 216.63 49.1 ;
    RECT 216.42 49.39 216.63 49.46 ;
    RECT 216.42 49.75 216.63 49.82 ;
    RECT 267.91 49.39 267.98 49.46 ;
    RECT 180.36 49.03 180.57 49.1 ;
    RECT 180.36 49.39 180.57 49.46 ;
    RECT 180.36 49.75 180.57 49.82 ;
    RECT 179.9 49.03 180.11 49.1 ;
    RECT 179.9 49.39 180.11 49.46 ;
    RECT 179.9 49.75 180.11 49.82 ;
    RECT 177.04 49.03 177.25 49.1 ;
    RECT 177.04 49.39 177.25 49.46 ;
    RECT 177.04 49.75 177.25 49.82 ;
    RECT 176.58 49.03 176.79 49.1 ;
    RECT 176.58 49.39 176.79 49.46 ;
    RECT 176.58 49.75 176.79 49.82 ;
    RECT 173.72 49.03 173.93 49.1 ;
    RECT 173.72 49.39 173.93 49.46 ;
    RECT 173.72 49.75 173.93 49.82 ;
    RECT 173.26 49.03 173.47 49.1 ;
    RECT 173.26 49.39 173.47 49.46 ;
    RECT 173.26 49.75 173.47 49.82 ;
    RECT 170.4 49.03 170.61 49.1 ;
    RECT 170.4 49.39 170.61 49.46 ;
    RECT 170.4 49.75 170.61 49.82 ;
    RECT 169.94 49.03 170.15 49.1 ;
    RECT 169.94 49.39 170.15 49.46 ;
    RECT 169.94 49.75 170.15 49.82 ;
    RECT 167.08 49.03 167.29 49.1 ;
    RECT 167.08 49.39 167.29 49.46 ;
    RECT 167.08 49.75 167.29 49.82 ;
    RECT 166.62 49.03 166.83 49.1 ;
    RECT 166.62 49.39 166.83 49.46 ;
    RECT 166.62 49.75 166.83 49.82 ;
    RECT 163.76 49.03 163.97 49.1 ;
    RECT 163.76 49.39 163.97 49.46 ;
    RECT 163.76 49.75 163.97 49.82 ;
    RECT 163.3 49.03 163.51 49.1 ;
    RECT 163.3 49.39 163.51 49.46 ;
    RECT 163.3 49.75 163.51 49.82 ;
    RECT 160.44 49.03 160.65 49.1 ;
    RECT 160.44 49.39 160.65 49.46 ;
    RECT 160.44 49.75 160.65 49.82 ;
    RECT 159.98 49.03 160.19 49.1 ;
    RECT 159.98 49.39 160.19 49.46 ;
    RECT 159.98 49.75 160.19 49.82 ;
    RECT 157.12 49.03 157.33 49.1 ;
    RECT 157.12 49.39 157.33 49.46 ;
    RECT 157.12 49.75 157.33 49.82 ;
    RECT 156.66 49.03 156.87 49.1 ;
    RECT 156.66 49.39 156.87 49.46 ;
    RECT 156.66 49.75 156.87 49.82 ;
    RECT 153.8 49.03 154.01 49.1 ;
    RECT 153.8 49.39 154.01 49.46 ;
    RECT 153.8 49.75 154.01 49.82 ;
    RECT 153.34 49.03 153.55 49.1 ;
    RECT 153.34 49.39 153.55 49.46 ;
    RECT 153.34 49.75 153.55 49.82 ;
    RECT 150.48 49.03 150.69 49.1 ;
    RECT 150.48 49.39 150.69 49.46 ;
    RECT 150.48 49.75 150.69 49.82 ;
    RECT 150.02 49.03 150.23 49.1 ;
    RECT 150.02 49.39 150.23 49.46 ;
    RECT 150.02 49.75 150.23 49.82 ;
    RECT 213.56 49.03 213.77 49.1 ;
    RECT 213.56 49.39 213.77 49.46 ;
    RECT 213.56 49.75 213.77 49.82 ;
    RECT 213.1 49.03 213.31 49.1 ;
    RECT 213.1 49.39 213.31 49.46 ;
    RECT 213.1 49.75 213.31 49.82 ;
    RECT 210.24 49.03 210.45 49.1 ;
    RECT 210.24 49.39 210.45 49.46 ;
    RECT 210.24 49.75 210.45 49.82 ;
    RECT 209.78 49.03 209.99 49.1 ;
    RECT 209.78 49.39 209.99 49.46 ;
    RECT 209.78 49.75 209.99 49.82 ;
    RECT 206.92 49.03 207.13 49.1 ;
    RECT 206.92 49.39 207.13 49.46 ;
    RECT 206.92 49.75 207.13 49.82 ;
    RECT 206.46 49.03 206.67 49.1 ;
    RECT 206.46 49.39 206.67 49.46 ;
    RECT 206.46 49.75 206.67 49.82 ;
    RECT 203.6 49.03 203.81 49.1 ;
    RECT 203.6 49.39 203.81 49.46 ;
    RECT 203.6 49.75 203.81 49.82 ;
    RECT 203.14 49.03 203.35 49.1 ;
    RECT 203.14 49.39 203.35 49.46 ;
    RECT 203.14 49.75 203.35 49.82 ;
    RECT 200.28 49.03 200.49 49.1 ;
    RECT 200.28 49.39 200.49 49.46 ;
    RECT 200.28 49.75 200.49 49.82 ;
    RECT 199.82 49.03 200.03 49.1 ;
    RECT 199.82 49.39 200.03 49.46 ;
    RECT 199.82 49.75 200.03 49.82 ;
    RECT 196.96 49.03 197.17 49.1 ;
    RECT 196.96 49.39 197.17 49.46 ;
    RECT 196.96 49.75 197.17 49.82 ;
    RECT 196.5 49.03 196.71 49.1 ;
    RECT 196.5 49.39 196.71 49.46 ;
    RECT 196.5 49.75 196.71 49.82 ;
    RECT 193.64 49.03 193.85 49.1 ;
    RECT 193.64 49.39 193.85 49.46 ;
    RECT 193.64 49.75 193.85 49.82 ;
    RECT 193.18 49.03 193.39 49.1 ;
    RECT 193.18 49.39 193.39 49.46 ;
    RECT 193.18 49.75 193.39 49.82 ;
    RECT 190.32 49.03 190.53 49.1 ;
    RECT 190.32 49.39 190.53 49.46 ;
    RECT 190.32 49.75 190.53 49.82 ;
    RECT 189.86 49.03 190.07 49.1 ;
    RECT 189.86 49.39 190.07 49.46 ;
    RECT 189.86 49.75 190.07 49.82 ;
    RECT 187.0 49.03 187.21 49.1 ;
    RECT 187.0 49.39 187.21 49.46 ;
    RECT 187.0 49.75 187.21 49.82 ;
    RECT 186.54 49.03 186.75 49.1 ;
    RECT 186.54 49.39 186.75 49.46 ;
    RECT 186.54 49.75 186.75 49.82 ;
    RECT 183.68 49.03 183.89 49.1 ;
    RECT 183.68 49.39 183.89 49.46 ;
    RECT 183.68 49.75 183.89 49.82 ;
    RECT 183.22 49.03 183.43 49.1 ;
    RECT 183.22 49.39 183.43 49.46 ;
    RECT 183.22 49.75 183.43 49.82 ;
    RECT 147.485 49.39 147.555 49.46 ;
    RECT 266.68 49.03 266.89 49.1 ;
    RECT 266.68 49.39 266.89 49.46 ;
    RECT 266.68 49.75 266.89 49.82 ;
    RECT 266.22 49.03 266.43 49.1 ;
    RECT 266.22 49.39 266.43 49.46 ;
    RECT 266.22 49.75 266.43 49.82 ;
    RECT 263.36 49.03 263.57 49.1 ;
    RECT 263.36 49.39 263.57 49.46 ;
    RECT 263.36 49.75 263.57 49.82 ;
    RECT 262.9 49.03 263.11 49.1 ;
    RECT 262.9 49.39 263.11 49.46 ;
    RECT 262.9 49.75 263.11 49.82 ;
    RECT 260.04 49.03 260.25 49.1 ;
    RECT 260.04 49.39 260.25 49.46 ;
    RECT 260.04 49.75 260.25 49.82 ;
    RECT 259.58 49.03 259.79 49.1 ;
    RECT 259.58 49.39 259.79 49.46 ;
    RECT 259.58 49.75 259.79 49.82 ;
    RECT 256.72 49.03 256.93 49.1 ;
    RECT 256.72 49.39 256.93 49.46 ;
    RECT 256.72 49.75 256.93 49.82 ;
    RECT 256.26 49.03 256.47 49.1 ;
    RECT 256.26 49.39 256.47 49.46 ;
    RECT 256.26 49.75 256.47 49.82 ;
    RECT 253.4 49.03 253.61 49.1 ;
    RECT 253.4 49.39 253.61 49.46 ;
    RECT 253.4 49.75 253.61 49.82 ;
    RECT 252.94 49.03 253.15 49.1 ;
    RECT 252.94 49.39 253.15 49.46 ;
    RECT 252.94 49.75 253.15 49.82 ;
    RECT 250.08 48.31 250.29 48.38 ;
    RECT 250.08 48.67 250.29 48.74 ;
    RECT 250.08 49.03 250.29 49.1 ;
    RECT 249.62 48.31 249.83 48.38 ;
    RECT 249.62 48.67 249.83 48.74 ;
    RECT 249.62 49.03 249.83 49.1 ;
    RECT 246.76 48.31 246.97 48.38 ;
    RECT 246.76 48.67 246.97 48.74 ;
    RECT 246.76 49.03 246.97 49.1 ;
    RECT 246.3 48.31 246.51 48.38 ;
    RECT 246.3 48.67 246.51 48.74 ;
    RECT 246.3 49.03 246.51 49.1 ;
    RECT 243.44 48.31 243.65 48.38 ;
    RECT 243.44 48.67 243.65 48.74 ;
    RECT 243.44 49.03 243.65 49.1 ;
    RECT 242.98 48.31 243.19 48.38 ;
    RECT 242.98 48.67 243.19 48.74 ;
    RECT 242.98 49.03 243.19 49.1 ;
    RECT 240.12 48.31 240.33 48.38 ;
    RECT 240.12 48.67 240.33 48.74 ;
    RECT 240.12 49.03 240.33 49.1 ;
    RECT 239.66 48.31 239.87 48.38 ;
    RECT 239.66 48.67 239.87 48.74 ;
    RECT 239.66 49.03 239.87 49.1 ;
    RECT 236.8 48.31 237.01 48.38 ;
    RECT 236.8 48.67 237.01 48.74 ;
    RECT 236.8 49.03 237.01 49.1 ;
    RECT 236.34 48.31 236.55 48.38 ;
    RECT 236.34 48.67 236.55 48.74 ;
    RECT 236.34 49.03 236.55 49.1 ;
    RECT 233.48 48.31 233.69 48.38 ;
    RECT 233.48 48.67 233.69 48.74 ;
    RECT 233.48 49.03 233.69 49.1 ;
    RECT 233.02 48.31 233.23 48.38 ;
    RECT 233.02 48.67 233.23 48.74 ;
    RECT 233.02 49.03 233.23 49.1 ;
    RECT 230.16 48.31 230.37 48.38 ;
    RECT 230.16 48.67 230.37 48.74 ;
    RECT 230.16 49.03 230.37 49.1 ;
    RECT 229.7 48.31 229.91 48.38 ;
    RECT 229.7 48.67 229.91 48.74 ;
    RECT 229.7 49.03 229.91 49.1 ;
    RECT 226.84 48.31 227.05 48.38 ;
    RECT 226.84 48.67 227.05 48.74 ;
    RECT 226.84 49.03 227.05 49.1 ;
    RECT 226.38 48.31 226.59 48.38 ;
    RECT 226.38 48.67 226.59 48.74 ;
    RECT 226.38 49.03 226.59 49.1 ;
    RECT 223.52 48.31 223.73 48.38 ;
    RECT 223.52 48.67 223.73 48.74 ;
    RECT 223.52 49.03 223.73 49.1 ;
    RECT 223.06 48.31 223.27 48.38 ;
    RECT 223.06 48.67 223.27 48.74 ;
    RECT 223.06 49.03 223.27 49.1 ;
    RECT 220.2 48.31 220.41 48.38 ;
    RECT 220.2 48.67 220.41 48.74 ;
    RECT 220.2 49.03 220.41 49.1 ;
    RECT 219.74 48.31 219.95 48.38 ;
    RECT 219.74 48.67 219.95 48.74 ;
    RECT 219.74 49.03 219.95 49.1 ;
    RECT 216.88 48.31 217.09 48.38 ;
    RECT 216.88 48.67 217.09 48.74 ;
    RECT 216.88 49.03 217.09 49.1 ;
    RECT 216.42 48.31 216.63 48.38 ;
    RECT 216.42 48.67 216.63 48.74 ;
    RECT 216.42 49.03 216.63 49.1 ;
    RECT 267.91 48.67 267.98 48.74 ;
    RECT 180.36 48.31 180.57 48.38 ;
    RECT 180.36 48.67 180.57 48.74 ;
    RECT 180.36 49.03 180.57 49.1 ;
    RECT 179.9 48.31 180.11 48.38 ;
    RECT 179.9 48.67 180.11 48.74 ;
    RECT 179.9 49.03 180.11 49.1 ;
    RECT 177.04 48.31 177.25 48.38 ;
    RECT 177.04 48.67 177.25 48.74 ;
    RECT 177.04 49.03 177.25 49.1 ;
    RECT 176.58 48.31 176.79 48.38 ;
    RECT 176.58 48.67 176.79 48.74 ;
    RECT 176.58 49.03 176.79 49.1 ;
    RECT 173.72 48.31 173.93 48.38 ;
    RECT 173.72 48.67 173.93 48.74 ;
    RECT 173.72 49.03 173.93 49.1 ;
    RECT 173.26 48.31 173.47 48.38 ;
    RECT 173.26 48.67 173.47 48.74 ;
    RECT 173.26 49.03 173.47 49.1 ;
    RECT 170.4 48.31 170.61 48.38 ;
    RECT 170.4 48.67 170.61 48.74 ;
    RECT 170.4 49.03 170.61 49.1 ;
    RECT 169.94 48.31 170.15 48.38 ;
    RECT 169.94 48.67 170.15 48.74 ;
    RECT 169.94 49.03 170.15 49.1 ;
    RECT 167.08 48.31 167.29 48.38 ;
    RECT 167.08 48.67 167.29 48.74 ;
    RECT 167.08 49.03 167.29 49.1 ;
    RECT 166.62 48.31 166.83 48.38 ;
    RECT 166.62 48.67 166.83 48.74 ;
    RECT 166.62 49.03 166.83 49.1 ;
    RECT 163.76 48.31 163.97 48.38 ;
    RECT 163.76 48.67 163.97 48.74 ;
    RECT 163.76 49.03 163.97 49.1 ;
    RECT 163.3 48.31 163.51 48.38 ;
    RECT 163.3 48.67 163.51 48.74 ;
    RECT 163.3 49.03 163.51 49.1 ;
    RECT 160.44 48.31 160.65 48.38 ;
    RECT 160.44 48.67 160.65 48.74 ;
    RECT 160.44 49.03 160.65 49.1 ;
    RECT 159.98 48.31 160.19 48.38 ;
    RECT 159.98 48.67 160.19 48.74 ;
    RECT 159.98 49.03 160.19 49.1 ;
    RECT 157.12 48.31 157.33 48.38 ;
    RECT 157.12 48.67 157.33 48.74 ;
    RECT 157.12 49.03 157.33 49.1 ;
    RECT 156.66 48.31 156.87 48.38 ;
    RECT 156.66 48.67 156.87 48.74 ;
    RECT 156.66 49.03 156.87 49.1 ;
    RECT 153.8 48.31 154.01 48.38 ;
    RECT 153.8 48.67 154.01 48.74 ;
    RECT 153.8 49.03 154.01 49.1 ;
    RECT 153.34 48.31 153.55 48.38 ;
    RECT 153.34 48.67 153.55 48.74 ;
    RECT 153.34 49.03 153.55 49.1 ;
    RECT 150.48 48.31 150.69 48.38 ;
    RECT 150.48 48.67 150.69 48.74 ;
    RECT 150.48 49.03 150.69 49.1 ;
    RECT 150.02 48.31 150.23 48.38 ;
    RECT 150.02 48.67 150.23 48.74 ;
    RECT 150.02 49.03 150.23 49.1 ;
    RECT 213.56 48.31 213.77 48.38 ;
    RECT 213.56 48.67 213.77 48.74 ;
    RECT 213.56 49.03 213.77 49.1 ;
    RECT 213.1 48.31 213.31 48.38 ;
    RECT 213.1 48.67 213.31 48.74 ;
    RECT 213.1 49.03 213.31 49.1 ;
    RECT 210.24 48.31 210.45 48.38 ;
    RECT 210.24 48.67 210.45 48.74 ;
    RECT 210.24 49.03 210.45 49.1 ;
    RECT 209.78 48.31 209.99 48.38 ;
    RECT 209.78 48.67 209.99 48.74 ;
    RECT 209.78 49.03 209.99 49.1 ;
    RECT 206.92 48.31 207.13 48.38 ;
    RECT 206.92 48.67 207.13 48.74 ;
    RECT 206.92 49.03 207.13 49.1 ;
    RECT 206.46 48.31 206.67 48.38 ;
    RECT 206.46 48.67 206.67 48.74 ;
    RECT 206.46 49.03 206.67 49.1 ;
    RECT 203.6 48.31 203.81 48.38 ;
    RECT 203.6 48.67 203.81 48.74 ;
    RECT 203.6 49.03 203.81 49.1 ;
    RECT 203.14 48.31 203.35 48.38 ;
    RECT 203.14 48.67 203.35 48.74 ;
    RECT 203.14 49.03 203.35 49.1 ;
    RECT 200.28 48.31 200.49 48.38 ;
    RECT 200.28 48.67 200.49 48.74 ;
    RECT 200.28 49.03 200.49 49.1 ;
    RECT 199.82 48.31 200.03 48.38 ;
    RECT 199.82 48.67 200.03 48.74 ;
    RECT 199.82 49.03 200.03 49.1 ;
    RECT 196.96 48.31 197.17 48.38 ;
    RECT 196.96 48.67 197.17 48.74 ;
    RECT 196.96 49.03 197.17 49.1 ;
    RECT 196.5 48.31 196.71 48.38 ;
    RECT 196.5 48.67 196.71 48.74 ;
    RECT 196.5 49.03 196.71 49.1 ;
    RECT 193.64 48.31 193.85 48.38 ;
    RECT 193.64 48.67 193.85 48.74 ;
    RECT 193.64 49.03 193.85 49.1 ;
    RECT 193.18 48.31 193.39 48.38 ;
    RECT 193.18 48.67 193.39 48.74 ;
    RECT 193.18 49.03 193.39 49.1 ;
    RECT 190.32 48.31 190.53 48.38 ;
    RECT 190.32 48.67 190.53 48.74 ;
    RECT 190.32 49.03 190.53 49.1 ;
    RECT 189.86 48.31 190.07 48.38 ;
    RECT 189.86 48.67 190.07 48.74 ;
    RECT 189.86 49.03 190.07 49.1 ;
    RECT 187.0 48.31 187.21 48.38 ;
    RECT 187.0 48.67 187.21 48.74 ;
    RECT 187.0 49.03 187.21 49.1 ;
    RECT 186.54 48.31 186.75 48.38 ;
    RECT 186.54 48.67 186.75 48.74 ;
    RECT 186.54 49.03 186.75 49.1 ;
    RECT 183.68 48.31 183.89 48.38 ;
    RECT 183.68 48.67 183.89 48.74 ;
    RECT 183.68 49.03 183.89 49.1 ;
    RECT 183.22 48.31 183.43 48.38 ;
    RECT 183.22 48.67 183.43 48.74 ;
    RECT 183.22 49.03 183.43 49.1 ;
    RECT 147.485 48.67 147.555 48.74 ;
    RECT 266.68 48.31 266.89 48.38 ;
    RECT 266.68 48.67 266.89 48.74 ;
    RECT 266.68 49.03 266.89 49.1 ;
    RECT 266.22 48.31 266.43 48.38 ;
    RECT 266.22 48.67 266.43 48.74 ;
    RECT 266.22 49.03 266.43 49.1 ;
    RECT 263.36 48.31 263.57 48.38 ;
    RECT 263.36 48.67 263.57 48.74 ;
    RECT 263.36 49.03 263.57 49.1 ;
    RECT 262.9 48.31 263.11 48.38 ;
    RECT 262.9 48.67 263.11 48.74 ;
    RECT 262.9 49.03 263.11 49.1 ;
    RECT 260.04 48.31 260.25 48.38 ;
    RECT 260.04 48.67 260.25 48.74 ;
    RECT 260.04 49.03 260.25 49.1 ;
    RECT 259.58 48.31 259.79 48.38 ;
    RECT 259.58 48.67 259.79 48.74 ;
    RECT 259.58 49.03 259.79 49.1 ;
    RECT 256.72 48.31 256.93 48.38 ;
    RECT 256.72 48.67 256.93 48.74 ;
    RECT 256.72 49.03 256.93 49.1 ;
    RECT 256.26 48.31 256.47 48.38 ;
    RECT 256.26 48.67 256.47 48.74 ;
    RECT 256.26 49.03 256.47 49.1 ;
    RECT 253.4 48.31 253.61 48.38 ;
    RECT 253.4 48.67 253.61 48.74 ;
    RECT 253.4 49.03 253.61 49.1 ;
    RECT 252.94 48.31 253.15 48.38 ;
    RECT 252.94 48.67 253.15 48.74 ;
    RECT 252.94 49.03 253.15 49.1 ;
    RECT 250.08 47.59 250.29 47.66 ;
    RECT 250.08 47.95 250.29 48.02 ;
    RECT 250.08 48.31 250.29 48.38 ;
    RECT 249.62 47.59 249.83 47.66 ;
    RECT 249.62 47.95 249.83 48.02 ;
    RECT 249.62 48.31 249.83 48.38 ;
    RECT 246.76 47.59 246.97 47.66 ;
    RECT 246.76 47.95 246.97 48.02 ;
    RECT 246.76 48.31 246.97 48.38 ;
    RECT 246.3 47.59 246.51 47.66 ;
    RECT 246.3 47.95 246.51 48.02 ;
    RECT 246.3 48.31 246.51 48.38 ;
    RECT 243.44 47.59 243.65 47.66 ;
    RECT 243.44 47.95 243.65 48.02 ;
    RECT 243.44 48.31 243.65 48.38 ;
    RECT 242.98 47.59 243.19 47.66 ;
    RECT 242.98 47.95 243.19 48.02 ;
    RECT 242.98 48.31 243.19 48.38 ;
    RECT 240.12 47.59 240.33 47.66 ;
    RECT 240.12 47.95 240.33 48.02 ;
    RECT 240.12 48.31 240.33 48.38 ;
    RECT 239.66 47.59 239.87 47.66 ;
    RECT 239.66 47.95 239.87 48.02 ;
    RECT 239.66 48.31 239.87 48.38 ;
    RECT 236.8 47.59 237.01 47.66 ;
    RECT 236.8 47.95 237.01 48.02 ;
    RECT 236.8 48.31 237.01 48.38 ;
    RECT 236.34 47.59 236.55 47.66 ;
    RECT 236.34 47.95 236.55 48.02 ;
    RECT 236.34 48.31 236.55 48.38 ;
    RECT 233.48 47.59 233.69 47.66 ;
    RECT 233.48 47.95 233.69 48.02 ;
    RECT 233.48 48.31 233.69 48.38 ;
    RECT 233.02 47.59 233.23 47.66 ;
    RECT 233.02 47.95 233.23 48.02 ;
    RECT 233.02 48.31 233.23 48.38 ;
    RECT 230.16 47.59 230.37 47.66 ;
    RECT 230.16 47.95 230.37 48.02 ;
    RECT 230.16 48.31 230.37 48.38 ;
    RECT 229.7 47.59 229.91 47.66 ;
    RECT 229.7 47.95 229.91 48.02 ;
    RECT 229.7 48.31 229.91 48.38 ;
    RECT 226.84 47.59 227.05 47.66 ;
    RECT 226.84 47.95 227.05 48.02 ;
    RECT 226.84 48.31 227.05 48.38 ;
    RECT 226.38 47.59 226.59 47.66 ;
    RECT 226.38 47.95 226.59 48.02 ;
    RECT 226.38 48.31 226.59 48.38 ;
    RECT 223.52 47.59 223.73 47.66 ;
    RECT 223.52 47.95 223.73 48.02 ;
    RECT 223.52 48.31 223.73 48.38 ;
    RECT 223.06 47.59 223.27 47.66 ;
    RECT 223.06 47.95 223.27 48.02 ;
    RECT 223.06 48.31 223.27 48.38 ;
    RECT 220.2 47.59 220.41 47.66 ;
    RECT 220.2 47.95 220.41 48.02 ;
    RECT 220.2 48.31 220.41 48.38 ;
    RECT 219.74 47.59 219.95 47.66 ;
    RECT 219.74 47.95 219.95 48.02 ;
    RECT 219.74 48.31 219.95 48.38 ;
    RECT 216.88 47.59 217.09 47.66 ;
    RECT 216.88 47.95 217.09 48.02 ;
    RECT 216.88 48.31 217.09 48.38 ;
    RECT 216.42 47.59 216.63 47.66 ;
    RECT 216.42 47.95 216.63 48.02 ;
    RECT 216.42 48.31 216.63 48.38 ;
    RECT 267.91 47.95 267.98 48.02 ;
    RECT 180.36 47.59 180.57 47.66 ;
    RECT 180.36 47.95 180.57 48.02 ;
    RECT 180.36 48.31 180.57 48.38 ;
    RECT 179.9 47.59 180.11 47.66 ;
    RECT 179.9 47.95 180.11 48.02 ;
    RECT 179.9 48.31 180.11 48.38 ;
    RECT 177.04 47.59 177.25 47.66 ;
    RECT 177.04 47.95 177.25 48.02 ;
    RECT 177.04 48.31 177.25 48.38 ;
    RECT 176.58 47.59 176.79 47.66 ;
    RECT 176.58 47.95 176.79 48.02 ;
    RECT 176.58 48.31 176.79 48.38 ;
    RECT 173.72 47.59 173.93 47.66 ;
    RECT 173.72 47.95 173.93 48.02 ;
    RECT 173.72 48.31 173.93 48.38 ;
    RECT 173.26 47.59 173.47 47.66 ;
    RECT 173.26 47.95 173.47 48.02 ;
    RECT 173.26 48.31 173.47 48.38 ;
    RECT 170.4 47.59 170.61 47.66 ;
    RECT 170.4 47.95 170.61 48.02 ;
    RECT 170.4 48.31 170.61 48.38 ;
    RECT 169.94 47.59 170.15 47.66 ;
    RECT 169.94 47.95 170.15 48.02 ;
    RECT 169.94 48.31 170.15 48.38 ;
    RECT 167.08 47.59 167.29 47.66 ;
    RECT 167.08 47.95 167.29 48.02 ;
    RECT 167.08 48.31 167.29 48.38 ;
    RECT 166.62 47.59 166.83 47.66 ;
    RECT 166.62 47.95 166.83 48.02 ;
    RECT 166.62 48.31 166.83 48.38 ;
    RECT 163.76 47.59 163.97 47.66 ;
    RECT 163.76 47.95 163.97 48.02 ;
    RECT 163.76 48.31 163.97 48.38 ;
    RECT 163.3 47.59 163.51 47.66 ;
    RECT 163.3 47.95 163.51 48.02 ;
    RECT 163.3 48.31 163.51 48.38 ;
    RECT 160.44 47.59 160.65 47.66 ;
    RECT 160.44 47.95 160.65 48.02 ;
    RECT 160.44 48.31 160.65 48.38 ;
    RECT 159.98 47.59 160.19 47.66 ;
    RECT 159.98 47.95 160.19 48.02 ;
    RECT 159.98 48.31 160.19 48.38 ;
    RECT 157.12 47.59 157.33 47.66 ;
    RECT 157.12 47.95 157.33 48.02 ;
    RECT 157.12 48.31 157.33 48.38 ;
    RECT 156.66 47.59 156.87 47.66 ;
    RECT 156.66 47.95 156.87 48.02 ;
    RECT 156.66 48.31 156.87 48.38 ;
    RECT 153.8 47.59 154.01 47.66 ;
    RECT 153.8 47.95 154.01 48.02 ;
    RECT 153.8 48.31 154.01 48.38 ;
    RECT 153.34 47.59 153.55 47.66 ;
    RECT 153.34 47.95 153.55 48.02 ;
    RECT 153.34 48.31 153.55 48.38 ;
    RECT 150.48 47.59 150.69 47.66 ;
    RECT 150.48 47.95 150.69 48.02 ;
    RECT 150.48 48.31 150.69 48.38 ;
    RECT 150.02 47.59 150.23 47.66 ;
    RECT 150.02 47.95 150.23 48.02 ;
    RECT 150.02 48.31 150.23 48.38 ;
    RECT 213.56 47.59 213.77 47.66 ;
    RECT 213.56 47.95 213.77 48.02 ;
    RECT 213.56 48.31 213.77 48.38 ;
    RECT 213.1 47.59 213.31 47.66 ;
    RECT 213.1 47.95 213.31 48.02 ;
    RECT 213.1 48.31 213.31 48.38 ;
    RECT 210.24 47.59 210.45 47.66 ;
    RECT 210.24 47.95 210.45 48.02 ;
    RECT 210.24 48.31 210.45 48.38 ;
    RECT 209.78 47.59 209.99 47.66 ;
    RECT 209.78 47.95 209.99 48.02 ;
    RECT 209.78 48.31 209.99 48.38 ;
    RECT 206.92 47.59 207.13 47.66 ;
    RECT 206.92 47.95 207.13 48.02 ;
    RECT 206.92 48.31 207.13 48.38 ;
    RECT 206.46 47.59 206.67 47.66 ;
    RECT 206.46 47.95 206.67 48.02 ;
    RECT 206.46 48.31 206.67 48.38 ;
    RECT 203.6 47.59 203.81 47.66 ;
    RECT 203.6 47.95 203.81 48.02 ;
    RECT 203.6 48.31 203.81 48.38 ;
    RECT 203.14 47.59 203.35 47.66 ;
    RECT 203.14 47.95 203.35 48.02 ;
    RECT 203.14 48.31 203.35 48.38 ;
    RECT 200.28 47.59 200.49 47.66 ;
    RECT 200.28 47.95 200.49 48.02 ;
    RECT 200.28 48.31 200.49 48.38 ;
    RECT 199.82 47.59 200.03 47.66 ;
    RECT 199.82 47.95 200.03 48.02 ;
    RECT 199.82 48.31 200.03 48.38 ;
    RECT 196.96 47.59 197.17 47.66 ;
    RECT 196.96 47.95 197.17 48.02 ;
    RECT 196.96 48.31 197.17 48.38 ;
    RECT 196.5 47.59 196.71 47.66 ;
    RECT 196.5 47.95 196.71 48.02 ;
    RECT 196.5 48.31 196.71 48.38 ;
    RECT 193.64 47.59 193.85 47.66 ;
    RECT 193.64 47.95 193.85 48.02 ;
    RECT 193.64 48.31 193.85 48.38 ;
    RECT 193.18 47.59 193.39 47.66 ;
    RECT 193.18 47.95 193.39 48.02 ;
    RECT 193.18 48.31 193.39 48.38 ;
    RECT 190.32 47.59 190.53 47.66 ;
    RECT 190.32 47.95 190.53 48.02 ;
    RECT 190.32 48.31 190.53 48.38 ;
    RECT 189.86 47.59 190.07 47.66 ;
    RECT 189.86 47.95 190.07 48.02 ;
    RECT 189.86 48.31 190.07 48.38 ;
    RECT 187.0 47.59 187.21 47.66 ;
    RECT 187.0 47.95 187.21 48.02 ;
    RECT 187.0 48.31 187.21 48.38 ;
    RECT 186.54 47.59 186.75 47.66 ;
    RECT 186.54 47.95 186.75 48.02 ;
    RECT 186.54 48.31 186.75 48.38 ;
    RECT 183.68 47.59 183.89 47.66 ;
    RECT 183.68 47.95 183.89 48.02 ;
    RECT 183.68 48.31 183.89 48.38 ;
    RECT 183.22 47.59 183.43 47.66 ;
    RECT 183.22 47.95 183.43 48.02 ;
    RECT 183.22 48.31 183.43 48.38 ;
    RECT 147.485 47.95 147.555 48.02 ;
    RECT 266.68 47.59 266.89 47.66 ;
    RECT 266.68 47.95 266.89 48.02 ;
    RECT 266.68 48.31 266.89 48.38 ;
    RECT 266.22 47.59 266.43 47.66 ;
    RECT 266.22 47.95 266.43 48.02 ;
    RECT 266.22 48.31 266.43 48.38 ;
    RECT 263.36 47.59 263.57 47.66 ;
    RECT 263.36 47.95 263.57 48.02 ;
    RECT 263.36 48.31 263.57 48.38 ;
    RECT 262.9 47.59 263.11 47.66 ;
    RECT 262.9 47.95 263.11 48.02 ;
    RECT 262.9 48.31 263.11 48.38 ;
    RECT 260.04 47.59 260.25 47.66 ;
    RECT 260.04 47.95 260.25 48.02 ;
    RECT 260.04 48.31 260.25 48.38 ;
    RECT 259.58 47.59 259.79 47.66 ;
    RECT 259.58 47.95 259.79 48.02 ;
    RECT 259.58 48.31 259.79 48.38 ;
    RECT 256.72 47.59 256.93 47.66 ;
    RECT 256.72 47.95 256.93 48.02 ;
    RECT 256.72 48.31 256.93 48.38 ;
    RECT 256.26 47.59 256.47 47.66 ;
    RECT 256.26 47.95 256.47 48.02 ;
    RECT 256.26 48.31 256.47 48.38 ;
    RECT 253.4 47.59 253.61 47.66 ;
    RECT 253.4 47.95 253.61 48.02 ;
    RECT 253.4 48.31 253.61 48.38 ;
    RECT 252.94 47.59 253.15 47.66 ;
    RECT 252.94 47.95 253.15 48.02 ;
    RECT 252.94 48.31 253.15 48.38 ;
    RECT 250.08 46.87 250.29 46.94 ;
    RECT 250.08 47.23 250.29 47.3 ;
    RECT 250.08 47.59 250.29 47.66 ;
    RECT 249.62 46.87 249.83 46.94 ;
    RECT 249.62 47.23 249.83 47.3 ;
    RECT 249.62 47.59 249.83 47.66 ;
    RECT 246.76 46.87 246.97 46.94 ;
    RECT 246.76 47.23 246.97 47.3 ;
    RECT 246.76 47.59 246.97 47.66 ;
    RECT 246.3 46.87 246.51 46.94 ;
    RECT 246.3 47.23 246.51 47.3 ;
    RECT 246.3 47.59 246.51 47.66 ;
    RECT 243.44 46.87 243.65 46.94 ;
    RECT 243.44 47.23 243.65 47.3 ;
    RECT 243.44 47.59 243.65 47.66 ;
    RECT 242.98 46.87 243.19 46.94 ;
    RECT 242.98 47.23 243.19 47.3 ;
    RECT 242.98 47.59 243.19 47.66 ;
    RECT 240.12 46.87 240.33 46.94 ;
    RECT 240.12 47.23 240.33 47.3 ;
    RECT 240.12 47.59 240.33 47.66 ;
    RECT 239.66 46.87 239.87 46.94 ;
    RECT 239.66 47.23 239.87 47.3 ;
    RECT 239.66 47.59 239.87 47.66 ;
    RECT 236.8 46.87 237.01 46.94 ;
    RECT 236.8 47.23 237.01 47.3 ;
    RECT 236.8 47.59 237.01 47.66 ;
    RECT 236.34 46.87 236.55 46.94 ;
    RECT 236.34 47.23 236.55 47.3 ;
    RECT 236.34 47.59 236.55 47.66 ;
    RECT 233.48 46.87 233.69 46.94 ;
    RECT 233.48 47.23 233.69 47.3 ;
    RECT 233.48 47.59 233.69 47.66 ;
    RECT 233.02 46.87 233.23 46.94 ;
    RECT 233.02 47.23 233.23 47.3 ;
    RECT 233.02 47.59 233.23 47.66 ;
    RECT 230.16 46.87 230.37 46.94 ;
    RECT 230.16 47.23 230.37 47.3 ;
    RECT 230.16 47.59 230.37 47.66 ;
    RECT 229.7 46.87 229.91 46.94 ;
    RECT 229.7 47.23 229.91 47.3 ;
    RECT 229.7 47.59 229.91 47.66 ;
    RECT 226.84 46.87 227.05 46.94 ;
    RECT 226.84 47.23 227.05 47.3 ;
    RECT 226.84 47.59 227.05 47.66 ;
    RECT 226.38 46.87 226.59 46.94 ;
    RECT 226.38 47.23 226.59 47.3 ;
    RECT 226.38 47.59 226.59 47.66 ;
    RECT 223.52 46.87 223.73 46.94 ;
    RECT 223.52 47.23 223.73 47.3 ;
    RECT 223.52 47.59 223.73 47.66 ;
    RECT 223.06 46.87 223.27 46.94 ;
    RECT 223.06 47.23 223.27 47.3 ;
    RECT 223.06 47.59 223.27 47.66 ;
    RECT 220.2 46.87 220.41 46.94 ;
    RECT 220.2 47.23 220.41 47.3 ;
    RECT 220.2 47.59 220.41 47.66 ;
    RECT 219.74 46.87 219.95 46.94 ;
    RECT 219.74 47.23 219.95 47.3 ;
    RECT 219.74 47.59 219.95 47.66 ;
    RECT 216.88 46.87 217.09 46.94 ;
    RECT 216.88 47.23 217.09 47.3 ;
    RECT 216.88 47.59 217.09 47.66 ;
    RECT 216.42 46.87 216.63 46.94 ;
    RECT 216.42 47.23 216.63 47.3 ;
    RECT 216.42 47.59 216.63 47.66 ;
    RECT 267.91 47.23 267.98 47.3 ;
    RECT 180.36 46.87 180.57 46.94 ;
    RECT 180.36 47.23 180.57 47.3 ;
    RECT 180.36 47.59 180.57 47.66 ;
    RECT 179.9 46.87 180.11 46.94 ;
    RECT 179.9 47.23 180.11 47.3 ;
    RECT 179.9 47.59 180.11 47.66 ;
    RECT 177.04 46.87 177.25 46.94 ;
    RECT 177.04 47.23 177.25 47.3 ;
    RECT 177.04 47.59 177.25 47.66 ;
    RECT 176.58 46.87 176.79 46.94 ;
    RECT 176.58 47.23 176.79 47.3 ;
    RECT 176.58 47.59 176.79 47.66 ;
    RECT 173.72 46.87 173.93 46.94 ;
    RECT 173.72 47.23 173.93 47.3 ;
    RECT 173.72 47.59 173.93 47.66 ;
    RECT 173.26 46.87 173.47 46.94 ;
    RECT 173.26 47.23 173.47 47.3 ;
    RECT 173.26 47.59 173.47 47.66 ;
    RECT 170.4 46.87 170.61 46.94 ;
    RECT 170.4 47.23 170.61 47.3 ;
    RECT 170.4 47.59 170.61 47.66 ;
    RECT 169.94 46.87 170.15 46.94 ;
    RECT 169.94 47.23 170.15 47.3 ;
    RECT 169.94 47.59 170.15 47.66 ;
    RECT 167.08 46.87 167.29 46.94 ;
    RECT 167.08 47.23 167.29 47.3 ;
    RECT 167.08 47.59 167.29 47.66 ;
    RECT 166.62 46.87 166.83 46.94 ;
    RECT 166.62 47.23 166.83 47.3 ;
    RECT 166.62 47.59 166.83 47.66 ;
    RECT 163.76 46.87 163.97 46.94 ;
    RECT 163.76 47.23 163.97 47.3 ;
    RECT 163.76 47.59 163.97 47.66 ;
    RECT 163.3 46.87 163.51 46.94 ;
    RECT 163.3 47.23 163.51 47.3 ;
    RECT 163.3 47.59 163.51 47.66 ;
    RECT 160.44 46.87 160.65 46.94 ;
    RECT 160.44 47.23 160.65 47.3 ;
    RECT 160.44 47.59 160.65 47.66 ;
    RECT 159.98 46.87 160.19 46.94 ;
    RECT 159.98 47.23 160.19 47.3 ;
    RECT 159.98 47.59 160.19 47.66 ;
    RECT 157.12 46.87 157.33 46.94 ;
    RECT 157.12 47.23 157.33 47.3 ;
    RECT 157.12 47.59 157.33 47.66 ;
    RECT 156.66 46.87 156.87 46.94 ;
    RECT 156.66 47.23 156.87 47.3 ;
    RECT 156.66 47.59 156.87 47.66 ;
    RECT 153.8 46.87 154.01 46.94 ;
    RECT 153.8 47.23 154.01 47.3 ;
    RECT 153.8 47.59 154.01 47.66 ;
    RECT 153.34 46.87 153.55 46.94 ;
    RECT 153.34 47.23 153.55 47.3 ;
    RECT 153.34 47.59 153.55 47.66 ;
    RECT 150.48 46.87 150.69 46.94 ;
    RECT 150.48 47.23 150.69 47.3 ;
    RECT 150.48 47.59 150.69 47.66 ;
    RECT 150.02 46.87 150.23 46.94 ;
    RECT 150.02 47.23 150.23 47.3 ;
    RECT 150.02 47.59 150.23 47.66 ;
    RECT 213.56 46.87 213.77 46.94 ;
    RECT 213.56 47.23 213.77 47.3 ;
    RECT 213.56 47.59 213.77 47.66 ;
    RECT 213.1 46.87 213.31 46.94 ;
    RECT 213.1 47.23 213.31 47.3 ;
    RECT 213.1 47.59 213.31 47.66 ;
    RECT 210.24 46.87 210.45 46.94 ;
    RECT 210.24 47.23 210.45 47.3 ;
    RECT 210.24 47.59 210.45 47.66 ;
    RECT 209.78 46.87 209.99 46.94 ;
    RECT 209.78 47.23 209.99 47.3 ;
    RECT 209.78 47.59 209.99 47.66 ;
    RECT 206.92 46.87 207.13 46.94 ;
    RECT 206.92 47.23 207.13 47.3 ;
    RECT 206.92 47.59 207.13 47.66 ;
    RECT 206.46 46.87 206.67 46.94 ;
    RECT 206.46 47.23 206.67 47.3 ;
    RECT 206.46 47.59 206.67 47.66 ;
    RECT 203.6 46.87 203.81 46.94 ;
    RECT 203.6 47.23 203.81 47.3 ;
    RECT 203.6 47.59 203.81 47.66 ;
    RECT 203.14 46.87 203.35 46.94 ;
    RECT 203.14 47.23 203.35 47.3 ;
    RECT 203.14 47.59 203.35 47.66 ;
    RECT 200.28 46.87 200.49 46.94 ;
    RECT 200.28 47.23 200.49 47.3 ;
    RECT 200.28 47.59 200.49 47.66 ;
    RECT 199.82 46.87 200.03 46.94 ;
    RECT 199.82 47.23 200.03 47.3 ;
    RECT 199.82 47.59 200.03 47.66 ;
    RECT 196.96 46.87 197.17 46.94 ;
    RECT 196.96 47.23 197.17 47.3 ;
    RECT 196.96 47.59 197.17 47.66 ;
    RECT 196.5 46.87 196.71 46.94 ;
    RECT 196.5 47.23 196.71 47.3 ;
    RECT 196.5 47.59 196.71 47.66 ;
    RECT 193.64 46.87 193.85 46.94 ;
    RECT 193.64 47.23 193.85 47.3 ;
    RECT 193.64 47.59 193.85 47.66 ;
    RECT 193.18 46.87 193.39 46.94 ;
    RECT 193.18 47.23 193.39 47.3 ;
    RECT 193.18 47.59 193.39 47.66 ;
    RECT 190.32 46.87 190.53 46.94 ;
    RECT 190.32 47.23 190.53 47.3 ;
    RECT 190.32 47.59 190.53 47.66 ;
    RECT 189.86 46.87 190.07 46.94 ;
    RECT 189.86 47.23 190.07 47.3 ;
    RECT 189.86 47.59 190.07 47.66 ;
    RECT 187.0 46.87 187.21 46.94 ;
    RECT 187.0 47.23 187.21 47.3 ;
    RECT 187.0 47.59 187.21 47.66 ;
    RECT 186.54 46.87 186.75 46.94 ;
    RECT 186.54 47.23 186.75 47.3 ;
    RECT 186.54 47.59 186.75 47.66 ;
    RECT 183.68 46.87 183.89 46.94 ;
    RECT 183.68 47.23 183.89 47.3 ;
    RECT 183.68 47.59 183.89 47.66 ;
    RECT 183.22 46.87 183.43 46.94 ;
    RECT 183.22 47.23 183.43 47.3 ;
    RECT 183.22 47.59 183.43 47.66 ;
    RECT 147.485 47.23 147.555 47.3 ;
    RECT 266.68 46.87 266.89 46.94 ;
    RECT 266.68 47.23 266.89 47.3 ;
    RECT 266.68 47.59 266.89 47.66 ;
    RECT 266.22 46.87 266.43 46.94 ;
    RECT 266.22 47.23 266.43 47.3 ;
    RECT 266.22 47.59 266.43 47.66 ;
    RECT 263.36 46.87 263.57 46.94 ;
    RECT 263.36 47.23 263.57 47.3 ;
    RECT 263.36 47.59 263.57 47.66 ;
    RECT 262.9 46.87 263.11 46.94 ;
    RECT 262.9 47.23 263.11 47.3 ;
    RECT 262.9 47.59 263.11 47.66 ;
    RECT 260.04 46.87 260.25 46.94 ;
    RECT 260.04 47.23 260.25 47.3 ;
    RECT 260.04 47.59 260.25 47.66 ;
    RECT 259.58 46.87 259.79 46.94 ;
    RECT 259.58 47.23 259.79 47.3 ;
    RECT 259.58 47.59 259.79 47.66 ;
    RECT 256.72 46.87 256.93 46.94 ;
    RECT 256.72 47.23 256.93 47.3 ;
    RECT 256.72 47.59 256.93 47.66 ;
    RECT 256.26 46.87 256.47 46.94 ;
    RECT 256.26 47.23 256.47 47.3 ;
    RECT 256.26 47.59 256.47 47.66 ;
    RECT 253.4 46.87 253.61 46.94 ;
    RECT 253.4 47.23 253.61 47.3 ;
    RECT 253.4 47.59 253.61 47.66 ;
    RECT 252.94 46.87 253.15 46.94 ;
    RECT 252.94 47.23 253.15 47.3 ;
    RECT 252.94 47.59 253.15 47.66 ;
    RECT 250.08 86.49 250.29 86.56 ;
    RECT 250.08 86.85 250.29 86.92 ;
    RECT 250.08 87.21 250.29 87.28 ;
    RECT 249.62 86.49 249.83 86.56 ;
    RECT 249.62 86.85 249.83 86.92 ;
    RECT 249.62 87.21 249.83 87.28 ;
    RECT 246.76 86.49 246.97 86.56 ;
    RECT 246.76 86.85 246.97 86.92 ;
    RECT 246.76 87.21 246.97 87.28 ;
    RECT 246.3 86.49 246.51 86.56 ;
    RECT 246.3 86.85 246.51 86.92 ;
    RECT 246.3 87.21 246.51 87.28 ;
    RECT 243.44 86.49 243.65 86.56 ;
    RECT 243.44 86.85 243.65 86.92 ;
    RECT 243.44 87.21 243.65 87.28 ;
    RECT 242.98 86.49 243.19 86.56 ;
    RECT 242.98 86.85 243.19 86.92 ;
    RECT 242.98 87.21 243.19 87.28 ;
    RECT 240.12 86.49 240.33 86.56 ;
    RECT 240.12 86.85 240.33 86.92 ;
    RECT 240.12 87.21 240.33 87.28 ;
    RECT 239.66 86.49 239.87 86.56 ;
    RECT 239.66 86.85 239.87 86.92 ;
    RECT 239.66 87.21 239.87 87.28 ;
    RECT 236.8 86.49 237.01 86.56 ;
    RECT 236.8 86.85 237.01 86.92 ;
    RECT 236.8 87.21 237.01 87.28 ;
    RECT 236.34 86.49 236.55 86.56 ;
    RECT 236.34 86.85 236.55 86.92 ;
    RECT 236.34 87.21 236.55 87.28 ;
    RECT 233.48 86.49 233.69 86.56 ;
    RECT 233.48 86.85 233.69 86.92 ;
    RECT 233.48 87.21 233.69 87.28 ;
    RECT 233.02 86.49 233.23 86.56 ;
    RECT 233.02 86.85 233.23 86.92 ;
    RECT 233.02 87.21 233.23 87.28 ;
    RECT 230.16 86.49 230.37 86.56 ;
    RECT 230.16 86.85 230.37 86.92 ;
    RECT 230.16 87.21 230.37 87.28 ;
    RECT 229.7 86.49 229.91 86.56 ;
    RECT 229.7 86.85 229.91 86.92 ;
    RECT 229.7 87.21 229.91 87.28 ;
    RECT 226.84 86.49 227.05 86.56 ;
    RECT 226.84 86.85 227.05 86.92 ;
    RECT 226.84 87.21 227.05 87.28 ;
    RECT 226.38 86.49 226.59 86.56 ;
    RECT 226.38 86.85 226.59 86.92 ;
    RECT 226.38 87.21 226.59 87.28 ;
    RECT 223.52 86.49 223.73 86.56 ;
    RECT 223.52 86.85 223.73 86.92 ;
    RECT 223.52 87.21 223.73 87.28 ;
    RECT 223.06 86.49 223.27 86.56 ;
    RECT 223.06 86.85 223.27 86.92 ;
    RECT 223.06 87.21 223.27 87.28 ;
    RECT 220.2 86.49 220.41 86.56 ;
    RECT 220.2 86.85 220.41 86.92 ;
    RECT 220.2 87.21 220.41 87.28 ;
    RECT 219.74 86.49 219.95 86.56 ;
    RECT 219.74 86.85 219.95 86.92 ;
    RECT 219.74 87.21 219.95 87.28 ;
    RECT 216.88 86.49 217.09 86.56 ;
    RECT 216.88 86.85 217.09 86.92 ;
    RECT 216.88 87.21 217.09 87.28 ;
    RECT 216.42 86.49 216.63 86.56 ;
    RECT 216.42 86.85 216.63 86.92 ;
    RECT 216.42 87.21 216.63 87.28 ;
    RECT 267.91 86.85 267.98 86.92 ;
    RECT 180.36 86.49 180.57 86.56 ;
    RECT 180.36 86.85 180.57 86.92 ;
    RECT 180.36 87.21 180.57 87.28 ;
    RECT 179.9 86.49 180.11 86.56 ;
    RECT 179.9 86.85 180.11 86.92 ;
    RECT 179.9 87.21 180.11 87.28 ;
    RECT 177.04 86.49 177.25 86.56 ;
    RECT 177.04 86.85 177.25 86.92 ;
    RECT 177.04 87.21 177.25 87.28 ;
    RECT 176.58 86.49 176.79 86.56 ;
    RECT 176.58 86.85 176.79 86.92 ;
    RECT 176.58 87.21 176.79 87.28 ;
    RECT 173.72 86.49 173.93 86.56 ;
    RECT 173.72 86.85 173.93 86.92 ;
    RECT 173.72 87.21 173.93 87.28 ;
    RECT 173.26 86.49 173.47 86.56 ;
    RECT 173.26 86.85 173.47 86.92 ;
    RECT 173.26 87.21 173.47 87.28 ;
    RECT 170.4 86.49 170.61 86.56 ;
    RECT 170.4 86.85 170.61 86.92 ;
    RECT 170.4 87.21 170.61 87.28 ;
    RECT 169.94 86.49 170.15 86.56 ;
    RECT 169.94 86.85 170.15 86.92 ;
    RECT 169.94 87.21 170.15 87.28 ;
    RECT 167.08 86.49 167.29 86.56 ;
    RECT 167.08 86.85 167.29 86.92 ;
    RECT 167.08 87.21 167.29 87.28 ;
    RECT 166.62 86.49 166.83 86.56 ;
    RECT 166.62 86.85 166.83 86.92 ;
    RECT 166.62 87.21 166.83 87.28 ;
    RECT 163.76 86.49 163.97 86.56 ;
    RECT 163.76 86.85 163.97 86.92 ;
    RECT 163.76 87.21 163.97 87.28 ;
    RECT 163.3 86.49 163.51 86.56 ;
    RECT 163.3 86.85 163.51 86.92 ;
    RECT 163.3 87.21 163.51 87.28 ;
    RECT 160.44 86.49 160.65 86.56 ;
    RECT 160.44 86.85 160.65 86.92 ;
    RECT 160.44 87.21 160.65 87.28 ;
    RECT 159.98 86.49 160.19 86.56 ;
    RECT 159.98 86.85 160.19 86.92 ;
    RECT 159.98 87.21 160.19 87.28 ;
    RECT 157.12 86.49 157.33 86.56 ;
    RECT 157.12 86.85 157.33 86.92 ;
    RECT 157.12 87.21 157.33 87.28 ;
    RECT 156.66 86.49 156.87 86.56 ;
    RECT 156.66 86.85 156.87 86.92 ;
    RECT 156.66 87.21 156.87 87.28 ;
    RECT 153.8 86.49 154.01 86.56 ;
    RECT 153.8 86.85 154.01 86.92 ;
    RECT 153.8 87.21 154.01 87.28 ;
    RECT 153.34 86.49 153.55 86.56 ;
    RECT 153.34 86.85 153.55 86.92 ;
    RECT 153.34 87.21 153.55 87.28 ;
    RECT 150.48 86.49 150.69 86.56 ;
    RECT 150.48 86.85 150.69 86.92 ;
    RECT 150.48 87.21 150.69 87.28 ;
    RECT 150.02 86.49 150.23 86.56 ;
    RECT 150.02 86.85 150.23 86.92 ;
    RECT 150.02 87.21 150.23 87.28 ;
    RECT 213.56 86.49 213.77 86.56 ;
    RECT 213.56 86.85 213.77 86.92 ;
    RECT 213.56 87.21 213.77 87.28 ;
    RECT 213.1 86.49 213.31 86.56 ;
    RECT 213.1 86.85 213.31 86.92 ;
    RECT 213.1 87.21 213.31 87.28 ;
    RECT 210.24 86.49 210.45 86.56 ;
    RECT 210.24 86.85 210.45 86.92 ;
    RECT 210.24 87.21 210.45 87.28 ;
    RECT 209.78 86.49 209.99 86.56 ;
    RECT 209.78 86.85 209.99 86.92 ;
    RECT 209.78 87.21 209.99 87.28 ;
    RECT 206.92 86.49 207.13 86.56 ;
    RECT 206.92 86.85 207.13 86.92 ;
    RECT 206.92 87.21 207.13 87.28 ;
    RECT 206.46 86.49 206.67 86.56 ;
    RECT 206.46 86.85 206.67 86.92 ;
    RECT 206.46 87.21 206.67 87.28 ;
    RECT 203.6 86.49 203.81 86.56 ;
    RECT 203.6 86.85 203.81 86.92 ;
    RECT 203.6 87.21 203.81 87.28 ;
    RECT 203.14 86.49 203.35 86.56 ;
    RECT 203.14 86.85 203.35 86.92 ;
    RECT 203.14 87.21 203.35 87.28 ;
    RECT 200.28 86.49 200.49 86.56 ;
    RECT 200.28 86.85 200.49 86.92 ;
    RECT 200.28 87.21 200.49 87.28 ;
    RECT 199.82 86.49 200.03 86.56 ;
    RECT 199.82 86.85 200.03 86.92 ;
    RECT 199.82 87.21 200.03 87.28 ;
    RECT 196.96 86.49 197.17 86.56 ;
    RECT 196.96 86.85 197.17 86.92 ;
    RECT 196.96 87.21 197.17 87.28 ;
    RECT 196.5 86.49 196.71 86.56 ;
    RECT 196.5 86.85 196.71 86.92 ;
    RECT 196.5 87.21 196.71 87.28 ;
    RECT 193.64 86.49 193.85 86.56 ;
    RECT 193.64 86.85 193.85 86.92 ;
    RECT 193.64 87.21 193.85 87.28 ;
    RECT 193.18 86.49 193.39 86.56 ;
    RECT 193.18 86.85 193.39 86.92 ;
    RECT 193.18 87.21 193.39 87.28 ;
    RECT 190.32 86.49 190.53 86.56 ;
    RECT 190.32 86.85 190.53 86.92 ;
    RECT 190.32 87.21 190.53 87.28 ;
    RECT 189.86 86.49 190.07 86.56 ;
    RECT 189.86 86.85 190.07 86.92 ;
    RECT 189.86 87.21 190.07 87.28 ;
    RECT 187.0 86.49 187.21 86.56 ;
    RECT 187.0 86.85 187.21 86.92 ;
    RECT 187.0 87.21 187.21 87.28 ;
    RECT 186.54 86.49 186.75 86.56 ;
    RECT 186.54 86.85 186.75 86.92 ;
    RECT 186.54 87.21 186.75 87.28 ;
    RECT 183.68 86.49 183.89 86.56 ;
    RECT 183.68 86.85 183.89 86.92 ;
    RECT 183.68 87.21 183.89 87.28 ;
    RECT 183.22 86.49 183.43 86.56 ;
    RECT 183.22 86.85 183.43 86.92 ;
    RECT 183.22 87.21 183.43 87.28 ;
    RECT 147.485 86.85 147.555 86.92 ;
    RECT 266.68 86.49 266.89 86.56 ;
    RECT 266.68 86.85 266.89 86.92 ;
    RECT 266.68 87.21 266.89 87.28 ;
    RECT 266.22 86.49 266.43 86.56 ;
    RECT 266.22 86.85 266.43 86.92 ;
    RECT 266.22 87.21 266.43 87.28 ;
    RECT 263.36 86.49 263.57 86.56 ;
    RECT 263.36 86.85 263.57 86.92 ;
    RECT 263.36 87.21 263.57 87.28 ;
    RECT 262.9 86.49 263.11 86.56 ;
    RECT 262.9 86.85 263.11 86.92 ;
    RECT 262.9 87.21 263.11 87.28 ;
    RECT 260.04 86.49 260.25 86.56 ;
    RECT 260.04 86.85 260.25 86.92 ;
    RECT 260.04 87.21 260.25 87.28 ;
    RECT 259.58 86.49 259.79 86.56 ;
    RECT 259.58 86.85 259.79 86.92 ;
    RECT 259.58 87.21 259.79 87.28 ;
    RECT 256.72 86.49 256.93 86.56 ;
    RECT 256.72 86.85 256.93 86.92 ;
    RECT 256.72 87.21 256.93 87.28 ;
    RECT 256.26 86.49 256.47 86.56 ;
    RECT 256.26 86.85 256.47 86.92 ;
    RECT 256.26 87.21 256.47 87.28 ;
    RECT 253.4 86.49 253.61 86.56 ;
    RECT 253.4 86.85 253.61 86.92 ;
    RECT 253.4 87.21 253.61 87.28 ;
    RECT 252.94 86.49 253.15 86.56 ;
    RECT 252.94 86.85 253.15 86.92 ;
    RECT 252.94 87.21 253.15 87.28 ;
    RECT 250.08 46.15 250.29 46.22 ;
    RECT 250.08 46.51 250.29 46.58 ;
    RECT 250.08 46.87 250.29 46.94 ;
    RECT 249.62 46.15 249.83 46.22 ;
    RECT 249.62 46.51 249.83 46.58 ;
    RECT 249.62 46.87 249.83 46.94 ;
    RECT 246.76 46.15 246.97 46.22 ;
    RECT 246.76 46.51 246.97 46.58 ;
    RECT 246.76 46.87 246.97 46.94 ;
    RECT 246.3 46.15 246.51 46.22 ;
    RECT 246.3 46.51 246.51 46.58 ;
    RECT 246.3 46.87 246.51 46.94 ;
    RECT 243.44 46.15 243.65 46.22 ;
    RECT 243.44 46.51 243.65 46.58 ;
    RECT 243.44 46.87 243.65 46.94 ;
    RECT 242.98 46.15 243.19 46.22 ;
    RECT 242.98 46.51 243.19 46.58 ;
    RECT 242.98 46.87 243.19 46.94 ;
    RECT 240.12 46.15 240.33 46.22 ;
    RECT 240.12 46.51 240.33 46.58 ;
    RECT 240.12 46.87 240.33 46.94 ;
    RECT 239.66 46.15 239.87 46.22 ;
    RECT 239.66 46.51 239.87 46.58 ;
    RECT 239.66 46.87 239.87 46.94 ;
    RECT 236.8 46.15 237.01 46.22 ;
    RECT 236.8 46.51 237.01 46.58 ;
    RECT 236.8 46.87 237.01 46.94 ;
    RECT 236.34 46.15 236.55 46.22 ;
    RECT 236.34 46.51 236.55 46.58 ;
    RECT 236.34 46.87 236.55 46.94 ;
    RECT 233.48 46.15 233.69 46.22 ;
    RECT 233.48 46.51 233.69 46.58 ;
    RECT 233.48 46.87 233.69 46.94 ;
    RECT 233.02 46.15 233.23 46.22 ;
    RECT 233.02 46.51 233.23 46.58 ;
    RECT 233.02 46.87 233.23 46.94 ;
    RECT 230.16 46.15 230.37 46.22 ;
    RECT 230.16 46.51 230.37 46.58 ;
    RECT 230.16 46.87 230.37 46.94 ;
    RECT 229.7 46.15 229.91 46.22 ;
    RECT 229.7 46.51 229.91 46.58 ;
    RECT 229.7 46.87 229.91 46.94 ;
    RECT 226.84 46.15 227.05 46.22 ;
    RECT 226.84 46.51 227.05 46.58 ;
    RECT 226.84 46.87 227.05 46.94 ;
    RECT 226.38 46.15 226.59 46.22 ;
    RECT 226.38 46.51 226.59 46.58 ;
    RECT 226.38 46.87 226.59 46.94 ;
    RECT 223.52 46.15 223.73 46.22 ;
    RECT 223.52 46.51 223.73 46.58 ;
    RECT 223.52 46.87 223.73 46.94 ;
    RECT 223.06 46.15 223.27 46.22 ;
    RECT 223.06 46.51 223.27 46.58 ;
    RECT 223.06 46.87 223.27 46.94 ;
    RECT 220.2 46.15 220.41 46.22 ;
    RECT 220.2 46.51 220.41 46.58 ;
    RECT 220.2 46.87 220.41 46.94 ;
    RECT 219.74 46.15 219.95 46.22 ;
    RECT 219.74 46.51 219.95 46.58 ;
    RECT 219.74 46.87 219.95 46.94 ;
    RECT 216.88 46.15 217.09 46.22 ;
    RECT 216.88 46.51 217.09 46.58 ;
    RECT 216.88 46.87 217.09 46.94 ;
    RECT 216.42 46.15 216.63 46.22 ;
    RECT 216.42 46.51 216.63 46.58 ;
    RECT 216.42 46.87 216.63 46.94 ;
    RECT 267.91 46.51 267.98 46.58 ;
    RECT 180.36 46.15 180.57 46.22 ;
    RECT 180.36 46.51 180.57 46.58 ;
    RECT 180.36 46.87 180.57 46.94 ;
    RECT 179.9 46.15 180.11 46.22 ;
    RECT 179.9 46.51 180.11 46.58 ;
    RECT 179.9 46.87 180.11 46.94 ;
    RECT 177.04 46.15 177.25 46.22 ;
    RECT 177.04 46.51 177.25 46.58 ;
    RECT 177.04 46.87 177.25 46.94 ;
    RECT 176.58 46.15 176.79 46.22 ;
    RECT 176.58 46.51 176.79 46.58 ;
    RECT 176.58 46.87 176.79 46.94 ;
    RECT 173.72 46.15 173.93 46.22 ;
    RECT 173.72 46.51 173.93 46.58 ;
    RECT 173.72 46.87 173.93 46.94 ;
    RECT 173.26 46.15 173.47 46.22 ;
    RECT 173.26 46.51 173.47 46.58 ;
    RECT 173.26 46.87 173.47 46.94 ;
    RECT 170.4 46.15 170.61 46.22 ;
    RECT 170.4 46.51 170.61 46.58 ;
    RECT 170.4 46.87 170.61 46.94 ;
    RECT 169.94 46.15 170.15 46.22 ;
    RECT 169.94 46.51 170.15 46.58 ;
    RECT 169.94 46.87 170.15 46.94 ;
    RECT 167.08 46.15 167.29 46.22 ;
    RECT 167.08 46.51 167.29 46.58 ;
    RECT 167.08 46.87 167.29 46.94 ;
    RECT 166.62 46.15 166.83 46.22 ;
    RECT 166.62 46.51 166.83 46.58 ;
    RECT 166.62 46.87 166.83 46.94 ;
    RECT 163.76 46.15 163.97 46.22 ;
    RECT 163.76 46.51 163.97 46.58 ;
    RECT 163.76 46.87 163.97 46.94 ;
    RECT 163.3 46.15 163.51 46.22 ;
    RECT 163.3 46.51 163.51 46.58 ;
    RECT 163.3 46.87 163.51 46.94 ;
    RECT 160.44 46.15 160.65 46.22 ;
    RECT 160.44 46.51 160.65 46.58 ;
    RECT 160.44 46.87 160.65 46.94 ;
    RECT 159.98 46.15 160.19 46.22 ;
    RECT 159.98 46.51 160.19 46.58 ;
    RECT 159.98 46.87 160.19 46.94 ;
    RECT 157.12 46.15 157.33 46.22 ;
    RECT 157.12 46.51 157.33 46.58 ;
    RECT 157.12 46.87 157.33 46.94 ;
    RECT 156.66 46.15 156.87 46.22 ;
    RECT 156.66 46.51 156.87 46.58 ;
    RECT 156.66 46.87 156.87 46.94 ;
    RECT 153.8 46.15 154.01 46.22 ;
    RECT 153.8 46.51 154.01 46.58 ;
    RECT 153.8 46.87 154.01 46.94 ;
    RECT 153.34 46.15 153.55 46.22 ;
    RECT 153.34 46.51 153.55 46.58 ;
    RECT 153.34 46.87 153.55 46.94 ;
    RECT 150.48 46.15 150.69 46.22 ;
    RECT 150.48 46.51 150.69 46.58 ;
    RECT 150.48 46.87 150.69 46.94 ;
    RECT 150.02 46.15 150.23 46.22 ;
    RECT 150.02 46.51 150.23 46.58 ;
    RECT 150.02 46.87 150.23 46.94 ;
    RECT 213.56 46.15 213.77 46.22 ;
    RECT 213.56 46.51 213.77 46.58 ;
    RECT 213.56 46.87 213.77 46.94 ;
    RECT 213.1 46.15 213.31 46.22 ;
    RECT 213.1 46.51 213.31 46.58 ;
    RECT 213.1 46.87 213.31 46.94 ;
    RECT 210.24 46.15 210.45 46.22 ;
    RECT 210.24 46.51 210.45 46.58 ;
    RECT 210.24 46.87 210.45 46.94 ;
    RECT 209.78 46.15 209.99 46.22 ;
    RECT 209.78 46.51 209.99 46.58 ;
    RECT 209.78 46.87 209.99 46.94 ;
    RECT 206.92 46.15 207.13 46.22 ;
    RECT 206.92 46.51 207.13 46.58 ;
    RECT 206.92 46.87 207.13 46.94 ;
    RECT 206.46 46.15 206.67 46.22 ;
    RECT 206.46 46.51 206.67 46.58 ;
    RECT 206.46 46.87 206.67 46.94 ;
    RECT 203.6 46.15 203.81 46.22 ;
    RECT 203.6 46.51 203.81 46.58 ;
    RECT 203.6 46.87 203.81 46.94 ;
    RECT 203.14 46.15 203.35 46.22 ;
    RECT 203.14 46.51 203.35 46.58 ;
    RECT 203.14 46.87 203.35 46.94 ;
    RECT 200.28 46.15 200.49 46.22 ;
    RECT 200.28 46.51 200.49 46.58 ;
    RECT 200.28 46.87 200.49 46.94 ;
    RECT 199.82 46.15 200.03 46.22 ;
    RECT 199.82 46.51 200.03 46.58 ;
    RECT 199.82 46.87 200.03 46.94 ;
    RECT 196.96 46.15 197.17 46.22 ;
    RECT 196.96 46.51 197.17 46.58 ;
    RECT 196.96 46.87 197.17 46.94 ;
    RECT 196.5 46.15 196.71 46.22 ;
    RECT 196.5 46.51 196.71 46.58 ;
    RECT 196.5 46.87 196.71 46.94 ;
    RECT 193.64 46.15 193.85 46.22 ;
    RECT 193.64 46.51 193.85 46.58 ;
    RECT 193.64 46.87 193.85 46.94 ;
    RECT 193.18 46.15 193.39 46.22 ;
    RECT 193.18 46.51 193.39 46.58 ;
    RECT 193.18 46.87 193.39 46.94 ;
    RECT 190.32 46.15 190.53 46.22 ;
    RECT 190.32 46.51 190.53 46.58 ;
    RECT 190.32 46.87 190.53 46.94 ;
    RECT 189.86 46.15 190.07 46.22 ;
    RECT 189.86 46.51 190.07 46.58 ;
    RECT 189.86 46.87 190.07 46.94 ;
    RECT 187.0 46.15 187.21 46.22 ;
    RECT 187.0 46.51 187.21 46.58 ;
    RECT 187.0 46.87 187.21 46.94 ;
    RECT 186.54 46.15 186.75 46.22 ;
    RECT 186.54 46.51 186.75 46.58 ;
    RECT 186.54 46.87 186.75 46.94 ;
    RECT 183.68 46.15 183.89 46.22 ;
    RECT 183.68 46.51 183.89 46.58 ;
    RECT 183.68 46.87 183.89 46.94 ;
    RECT 183.22 46.15 183.43 46.22 ;
    RECT 183.22 46.51 183.43 46.58 ;
    RECT 183.22 46.87 183.43 46.94 ;
    RECT 147.485 46.51 147.555 46.58 ;
    RECT 266.68 46.15 266.89 46.22 ;
    RECT 266.68 46.51 266.89 46.58 ;
    RECT 266.68 46.87 266.89 46.94 ;
    RECT 266.22 46.15 266.43 46.22 ;
    RECT 266.22 46.51 266.43 46.58 ;
    RECT 266.22 46.87 266.43 46.94 ;
    RECT 263.36 46.15 263.57 46.22 ;
    RECT 263.36 46.51 263.57 46.58 ;
    RECT 263.36 46.87 263.57 46.94 ;
    RECT 262.9 46.15 263.11 46.22 ;
    RECT 262.9 46.51 263.11 46.58 ;
    RECT 262.9 46.87 263.11 46.94 ;
    RECT 260.04 46.15 260.25 46.22 ;
    RECT 260.04 46.51 260.25 46.58 ;
    RECT 260.04 46.87 260.25 46.94 ;
    RECT 259.58 46.15 259.79 46.22 ;
    RECT 259.58 46.51 259.79 46.58 ;
    RECT 259.58 46.87 259.79 46.94 ;
    RECT 256.72 46.15 256.93 46.22 ;
    RECT 256.72 46.51 256.93 46.58 ;
    RECT 256.72 46.87 256.93 46.94 ;
    RECT 256.26 46.15 256.47 46.22 ;
    RECT 256.26 46.51 256.47 46.58 ;
    RECT 256.26 46.87 256.47 46.94 ;
    RECT 253.4 46.15 253.61 46.22 ;
    RECT 253.4 46.51 253.61 46.58 ;
    RECT 253.4 46.87 253.61 46.94 ;
    RECT 252.94 46.15 253.15 46.22 ;
    RECT 252.94 46.51 253.15 46.58 ;
    RECT 252.94 46.87 253.15 46.94 ;
    RECT 250.08 85.77 250.29 85.84 ;
    RECT 250.08 86.13 250.29 86.2 ;
    RECT 250.08 86.49 250.29 86.56 ;
    RECT 249.62 85.77 249.83 85.84 ;
    RECT 249.62 86.13 249.83 86.2 ;
    RECT 249.62 86.49 249.83 86.56 ;
    RECT 246.76 85.77 246.97 85.84 ;
    RECT 246.76 86.13 246.97 86.2 ;
    RECT 246.76 86.49 246.97 86.56 ;
    RECT 246.3 85.77 246.51 85.84 ;
    RECT 246.3 86.13 246.51 86.2 ;
    RECT 246.3 86.49 246.51 86.56 ;
    RECT 243.44 85.77 243.65 85.84 ;
    RECT 243.44 86.13 243.65 86.2 ;
    RECT 243.44 86.49 243.65 86.56 ;
    RECT 242.98 85.77 243.19 85.84 ;
    RECT 242.98 86.13 243.19 86.2 ;
    RECT 242.98 86.49 243.19 86.56 ;
    RECT 240.12 85.77 240.33 85.84 ;
    RECT 240.12 86.13 240.33 86.2 ;
    RECT 240.12 86.49 240.33 86.56 ;
    RECT 239.66 85.77 239.87 85.84 ;
    RECT 239.66 86.13 239.87 86.2 ;
    RECT 239.66 86.49 239.87 86.56 ;
    RECT 236.8 85.77 237.01 85.84 ;
    RECT 236.8 86.13 237.01 86.2 ;
    RECT 236.8 86.49 237.01 86.56 ;
    RECT 236.34 85.77 236.55 85.84 ;
    RECT 236.34 86.13 236.55 86.2 ;
    RECT 236.34 86.49 236.55 86.56 ;
    RECT 233.48 85.77 233.69 85.84 ;
    RECT 233.48 86.13 233.69 86.2 ;
    RECT 233.48 86.49 233.69 86.56 ;
    RECT 233.02 85.77 233.23 85.84 ;
    RECT 233.02 86.13 233.23 86.2 ;
    RECT 233.02 86.49 233.23 86.56 ;
    RECT 230.16 85.77 230.37 85.84 ;
    RECT 230.16 86.13 230.37 86.2 ;
    RECT 230.16 86.49 230.37 86.56 ;
    RECT 229.7 85.77 229.91 85.84 ;
    RECT 229.7 86.13 229.91 86.2 ;
    RECT 229.7 86.49 229.91 86.56 ;
    RECT 226.84 85.77 227.05 85.84 ;
    RECT 226.84 86.13 227.05 86.2 ;
    RECT 226.84 86.49 227.05 86.56 ;
    RECT 226.38 85.77 226.59 85.84 ;
    RECT 226.38 86.13 226.59 86.2 ;
    RECT 226.38 86.49 226.59 86.56 ;
    RECT 223.52 85.77 223.73 85.84 ;
    RECT 223.52 86.13 223.73 86.2 ;
    RECT 223.52 86.49 223.73 86.56 ;
    RECT 223.06 85.77 223.27 85.84 ;
    RECT 223.06 86.13 223.27 86.2 ;
    RECT 223.06 86.49 223.27 86.56 ;
    RECT 220.2 85.77 220.41 85.84 ;
    RECT 220.2 86.13 220.41 86.2 ;
    RECT 220.2 86.49 220.41 86.56 ;
    RECT 219.74 85.77 219.95 85.84 ;
    RECT 219.74 86.13 219.95 86.2 ;
    RECT 219.74 86.49 219.95 86.56 ;
    RECT 216.88 85.77 217.09 85.84 ;
    RECT 216.88 86.13 217.09 86.2 ;
    RECT 216.88 86.49 217.09 86.56 ;
    RECT 216.42 85.77 216.63 85.84 ;
    RECT 216.42 86.13 216.63 86.2 ;
    RECT 216.42 86.49 216.63 86.56 ;
    RECT 267.91 86.13 267.98 86.2 ;
    RECT 180.36 85.77 180.57 85.84 ;
    RECT 180.36 86.13 180.57 86.2 ;
    RECT 180.36 86.49 180.57 86.56 ;
    RECT 179.9 85.77 180.11 85.84 ;
    RECT 179.9 86.13 180.11 86.2 ;
    RECT 179.9 86.49 180.11 86.56 ;
    RECT 177.04 85.77 177.25 85.84 ;
    RECT 177.04 86.13 177.25 86.2 ;
    RECT 177.04 86.49 177.25 86.56 ;
    RECT 176.58 85.77 176.79 85.84 ;
    RECT 176.58 86.13 176.79 86.2 ;
    RECT 176.58 86.49 176.79 86.56 ;
    RECT 173.72 85.77 173.93 85.84 ;
    RECT 173.72 86.13 173.93 86.2 ;
    RECT 173.72 86.49 173.93 86.56 ;
    RECT 173.26 85.77 173.47 85.84 ;
    RECT 173.26 86.13 173.47 86.2 ;
    RECT 173.26 86.49 173.47 86.56 ;
    RECT 170.4 85.77 170.61 85.84 ;
    RECT 170.4 86.13 170.61 86.2 ;
    RECT 170.4 86.49 170.61 86.56 ;
    RECT 169.94 85.77 170.15 85.84 ;
    RECT 169.94 86.13 170.15 86.2 ;
    RECT 169.94 86.49 170.15 86.56 ;
    RECT 167.08 85.77 167.29 85.84 ;
    RECT 167.08 86.13 167.29 86.2 ;
    RECT 167.08 86.49 167.29 86.56 ;
    RECT 166.62 85.77 166.83 85.84 ;
    RECT 166.62 86.13 166.83 86.2 ;
    RECT 166.62 86.49 166.83 86.56 ;
    RECT 163.76 85.77 163.97 85.84 ;
    RECT 163.76 86.13 163.97 86.2 ;
    RECT 163.76 86.49 163.97 86.56 ;
    RECT 163.3 85.77 163.51 85.84 ;
    RECT 163.3 86.13 163.51 86.2 ;
    RECT 163.3 86.49 163.51 86.56 ;
    RECT 160.44 85.77 160.65 85.84 ;
    RECT 160.44 86.13 160.65 86.2 ;
    RECT 160.44 86.49 160.65 86.56 ;
    RECT 159.98 85.77 160.19 85.84 ;
    RECT 159.98 86.13 160.19 86.2 ;
    RECT 159.98 86.49 160.19 86.56 ;
    RECT 157.12 85.77 157.33 85.84 ;
    RECT 157.12 86.13 157.33 86.2 ;
    RECT 157.12 86.49 157.33 86.56 ;
    RECT 156.66 85.77 156.87 85.84 ;
    RECT 156.66 86.13 156.87 86.2 ;
    RECT 156.66 86.49 156.87 86.56 ;
    RECT 153.8 85.77 154.01 85.84 ;
    RECT 153.8 86.13 154.01 86.2 ;
    RECT 153.8 86.49 154.01 86.56 ;
    RECT 153.34 85.77 153.55 85.84 ;
    RECT 153.34 86.13 153.55 86.2 ;
    RECT 153.34 86.49 153.55 86.56 ;
    RECT 150.48 85.77 150.69 85.84 ;
    RECT 150.48 86.13 150.69 86.2 ;
    RECT 150.48 86.49 150.69 86.56 ;
    RECT 150.02 85.77 150.23 85.84 ;
    RECT 150.02 86.13 150.23 86.2 ;
    RECT 150.02 86.49 150.23 86.56 ;
    RECT 213.56 85.77 213.77 85.84 ;
    RECT 213.56 86.13 213.77 86.2 ;
    RECT 213.56 86.49 213.77 86.56 ;
    RECT 213.1 85.77 213.31 85.84 ;
    RECT 213.1 86.13 213.31 86.2 ;
    RECT 213.1 86.49 213.31 86.56 ;
    RECT 210.24 85.77 210.45 85.84 ;
    RECT 210.24 86.13 210.45 86.2 ;
    RECT 210.24 86.49 210.45 86.56 ;
    RECT 209.78 85.77 209.99 85.84 ;
    RECT 209.78 86.13 209.99 86.2 ;
    RECT 209.78 86.49 209.99 86.56 ;
    RECT 206.92 85.77 207.13 85.84 ;
    RECT 206.92 86.13 207.13 86.2 ;
    RECT 206.92 86.49 207.13 86.56 ;
    RECT 206.46 85.77 206.67 85.84 ;
    RECT 206.46 86.13 206.67 86.2 ;
    RECT 206.46 86.49 206.67 86.56 ;
    RECT 203.6 85.77 203.81 85.84 ;
    RECT 203.6 86.13 203.81 86.2 ;
    RECT 203.6 86.49 203.81 86.56 ;
    RECT 203.14 85.77 203.35 85.84 ;
    RECT 203.14 86.13 203.35 86.2 ;
    RECT 203.14 86.49 203.35 86.56 ;
    RECT 200.28 85.77 200.49 85.84 ;
    RECT 200.28 86.13 200.49 86.2 ;
    RECT 200.28 86.49 200.49 86.56 ;
    RECT 199.82 85.77 200.03 85.84 ;
    RECT 199.82 86.13 200.03 86.2 ;
    RECT 199.82 86.49 200.03 86.56 ;
    RECT 196.96 85.77 197.17 85.84 ;
    RECT 196.96 86.13 197.17 86.2 ;
    RECT 196.96 86.49 197.17 86.56 ;
    RECT 196.5 85.77 196.71 85.84 ;
    RECT 196.5 86.13 196.71 86.2 ;
    RECT 196.5 86.49 196.71 86.56 ;
    RECT 193.64 85.77 193.85 85.84 ;
    RECT 193.64 86.13 193.85 86.2 ;
    RECT 193.64 86.49 193.85 86.56 ;
    RECT 193.18 85.77 193.39 85.84 ;
    RECT 193.18 86.13 193.39 86.2 ;
    RECT 193.18 86.49 193.39 86.56 ;
    RECT 190.32 85.77 190.53 85.84 ;
    RECT 190.32 86.13 190.53 86.2 ;
    RECT 190.32 86.49 190.53 86.56 ;
    RECT 189.86 85.77 190.07 85.84 ;
    RECT 189.86 86.13 190.07 86.2 ;
    RECT 189.86 86.49 190.07 86.56 ;
    RECT 187.0 85.77 187.21 85.84 ;
    RECT 187.0 86.13 187.21 86.2 ;
    RECT 187.0 86.49 187.21 86.56 ;
    RECT 186.54 85.77 186.75 85.84 ;
    RECT 186.54 86.13 186.75 86.2 ;
    RECT 186.54 86.49 186.75 86.56 ;
    RECT 183.68 85.77 183.89 85.84 ;
    RECT 183.68 86.13 183.89 86.2 ;
    RECT 183.68 86.49 183.89 86.56 ;
    RECT 183.22 85.77 183.43 85.84 ;
    RECT 183.22 86.13 183.43 86.2 ;
    RECT 183.22 86.49 183.43 86.56 ;
    RECT 147.485 86.13 147.555 86.2 ;
    RECT 266.68 85.77 266.89 85.84 ;
    RECT 266.68 86.13 266.89 86.2 ;
    RECT 266.68 86.49 266.89 86.56 ;
    RECT 266.22 85.77 266.43 85.84 ;
    RECT 266.22 86.13 266.43 86.2 ;
    RECT 266.22 86.49 266.43 86.56 ;
    RECT 263.36 85.77 263.57 85.84 ;
    RECT 263.36 86.13 263.57 86.2 ;
    RECT 263.36 86.49 263.57 86.56 ;
    RECT 262.9 85.77 263.11 85.84 ;
    RECT 262.9 86.13 263.11 86.2 ;
    RECT 262.9 86.49 263.11 86.56 ;
    RECT 260.04 85.77 260.25 85.84 ;
    RECT 260.04 86.13 260.25 86.2 ;
    RECT 260.04 86.49 260.25 86.56 ;
    RECT 259.58 85.77 259.79 85.84 ;
    RECT 259.58 86.13 259.79 86.2 ;
    RECT 259.58 86.49 259.79 86.56 ;
    RECT 256.72 85.77 256.93 85.84 ;
    RECT 256.72 86.13 256.93 86.2 ;
    RECT 256.72 86.49 256.93 86.56 ;
    RECT 256.26 85.77 256.47 85.84 ;
    RECT 256.26 86.13 256.47 86.2 ;
    RECT 256.26 86.49 256.47 86.56 ;
    RECT 253.4 85.77 253.61 85.84 ;
    RECT 253.4 86.13 253.61 86.2 ;
    RECT 253.4 86.49 253.61 86.56 ;
    RECT 252.94 85.77 253.15 85.84 ;
    RECT 252.94 86.13 253.15 86.2 ;
    RECT 252.94 86.49 253.15 86.56 ;
    RECT 250.08 45.43 250.29 45.5 ;
    RECT 250.08 45.79 250.29 45.86 ;
    RECT 250.08 46.15 250.29 46.22 ;
    RECT 249.62 45.43 249.83 45.5 ;
    RECT 249.62 45.79 249.83 45.86 ;
    RECT 249.62 46.15 249.83 46.22 ;
    RECT 246.76 45.43 246.97 45.5 ;
    RECT 246.76 45.79 246.97 45.86 ;
    RECT 246.76 46.15 246.97 46.22 ;
    RECT 246.3 45.43 246.51 45.5 ;
    RECT 246.3 45.79 246.51 45.86 ;
    RECT 246.3 46.15 246.51 46.22 ;
    RECT 243.44 45.43 243.65 45.5 ;
    RECT 243.44 45.79 243.65 45.86 ;
    RECT 243.44 46.15 243.65 46.22 ;
    RECT 242.98 45.43 243.19 45.5 ;
    RECT 242.98 45.79 243.19 45.86 ;
    RECT 242.98 46.15 243.19 46.22 ;
    RECT 240.12 45.43 240.33 45.5 ;
    RECT 240.12 45.79 240.33 45.86 ;
    RECT 240.12 46.15 240.33 46.22 ;
    RECT 239.66 45.43 239.87 45.5 ;
    RECT 239.66 45.79 239.87 45.86 ;
    RECT 239.66 46.15 239.87 46.22 ;
    RECT 236.8 45.43 237.01 45.5 ;
    RECT 236.8 45.79 237.01 45.86 ;
    RECT 236.8 46.15 237.01 46.22 ;
    RECT 236.34 45.43 236.55 45.5 ;
    RECT 236.34 45.79 236.55 45.86 ;
    RECT 236.34 46.15 236.55 46.22 ;
    RECT 233.48 45.43 233.69 45.5 ;
    RECT 233.48 45.79 233.69 45.86 ;
    RECT 233.48 46.15 233.69 46.22 ;
    RECT 233.02 45.43 233.23 45.5 ;
    RECT 233.02 45.79 233.23 45.86 ;
    RECT 233.02 46.15 233.23 46.22 ;
    RECT 230.16 45.43 230.37 45.5 ;
    RECT 230.16 45.79 230.37 45.86 ;
    RECT 230.16 46.15 230.37 46.22 ;
    RECT 229.7 45.43 229.91 45.5 ;
    RECT 229.7 45.79 229.91 45.86 ;
    RECT 229.7 46.15 229.91 46.22 ;
    RECT 226.84 45.43 227.05 45.5 ;
    RECT 226.84 45.79 227.05 45.86 ;
    RECT 226.84 46.15 227.05 46.22 ;
    RECT 226.38 45.43 226.59 45.5 ;
    RECT 226.38 45.79 226.59 45.86 ;
    RECT 226.38 46.15 226.59 46.22 ;
    RECT 223.52 45.43 223.73 45.5 ;
    RECT 223.52 45.79 223.73 45.86 ;
    RECT 223.52 46.15 223.73 46.22 ;
    RECT 223.06 45.43 223.27 45.5 ;
    RECT 223.06 45.79 223.27 45.86 ;
    RECT 223.06 46.15 223.27 46.22 ;
    RECT 220.2 45.43 220.41 45.5 ;
    RECT 220.2 45.79 220.41 45.86 ;
    RECT 220.2 46.15 220.41 46.22 ;
    RECT 219.74 45.43 219.95 45.5 ;
    RECT 219.74 45.79 219.95 45.86 ;
    RECT 219.74 46.15 219.95 46.22 ;
    RECT 216.88 45.43 217.09 45.5 ;
    RECT 216.88 45.79 217.09 45.86 ;
    RECT 216.88 46.15 217.09 46.22 ;
    RECT 216.42 45.43 216.63 45.5 ;
    RECT 216.42 45.79 216.63 45.86 ;
    RECT 216.42 46.15 216.63 46.22 ;
    RECT 267.91 45.79 267.98 45.86 ;
    RECT 180.36 45.43 180.57 45.5 ;
    RECT 180.36 45.79 180.57 45.86 ;
    RECT 180.36 46.15 180.57 46.22 ;
    RECT 179.9 45.43 180.11 45.5 ;
    RECT 179.9 45.79 180.11 45.86 ;
    RECT 179.9 46.15 180.11 46.22 ;
    RECT 177.04 45.43 177.25 45.5 ;
    RECT 177.04 45.79 177.25 45.86 ;
    RECT 177.04 46.15 177.25 46.22 ;
    RECT 176.58 45.43 176.79 45.5 ;
    RECT 176.58 45.79 176.79 45.86 ;
    RECT 176.58 46.15 176.79 46.22 ;
    RECT 173.72 45.43 173.93 45.5 ;
    RECT 173.72 45.79 173.93 45.86 ;
    RECT 173.72 46.15 173.93 46.22 ;
    RECT 173.26 45.43 173.47 45.5 ;
    RECT 173.26 45.79 173.47 45.86 ;
    RECT 173.26 46.15 173.47 46.22 ;
    RECT 170.4 45.43 170.61 45.5 ;
    RECT 170.4 45.79 170.61 45.86 ;
    RECT 170.4 46.15 170.61 46.22 ;
    RECT 169.94 45.43 170.15 45.5 ;
    RECT 169.94 45.79 170.15 45.86 ;
    RECT 169.94 46.15 170.15 46.22 ;
    RECT 167.08 45.43 167.29 45.5 ;
    RECT 167.08 45.79 167.29 45.86 ;
    RECT 167.08 46.15 167.29 46.22 ;
    RECT 166.62 45.43 166.83 45.5 ;
    RECT 166.62 45.79 166.83 45.86 ;
    RECT 166.62 46.15 166.83 46.22 ;
    RECT 163.76 45.43 163.97 45.5 ;
    RECT 163.76 45.79 163.97 45.86 ;
    RECT 163.76 46.15 163.97 46.22 ;
    RECT 163.3 45.43 163.51 45.5 ;
    RECT 163.3 45.79 163.51 45.86 ;
    RECT 163.3 46.15 163.51 46.22 ;
    RECT 160.44 45.43 160.65 45.5 ;
    RECT 160.44 45.79 160.65 45.86 ;
    RECT 160.44 46.15 160.65 46.22 ;
    RECT 159.98 45.43 160.19 45.5 ;
    RECT 159.98 45.79 160.19 45.86 ;
    RECT 159.98 46.15 160.19 46.22 ;
    RECT 157.12 45.43 157.33 45.5 ;
    RECT 157.12 45.79 157.33 45.86 ;
    RECT 157.12 46.15 157.33 46.22 ;
    RECT 156.66 45.43 156.87 45.5 ;
    RECT 156.66 45.79 156.87 45.86 ;
    RECT 156.66 46.15 156.87 46.22 ;
    RECT 153.8 45.43 154.01 45.5 ;
    RECT 153.8 45.79 154.01 45.86 ;
    RECT 153.8 46.15 154.01 46.22 ;
    RECT 153.34 45.43 153.55 45.5 ;
    RECT 153.34 45.79 153.55 45.86 ;
    RECT 153.34 46.15 153.55 46.22 ;
    RECT 150.48 45.43 150.69 45.5 ;
    RECT 150.48 45.79 150.69 45.86 ;
    RECT 150.48 46.15 150.69 46.22 ;
    RECT 150.02 45.43 150.23 45.5 ;
    RECT 150.02 45.79 150.23 45.86 ;
    RECT 150.02 46.15 150.23 46.22 ;
    RECT 213.56 45.43 213.77 45.5 ;
    RECT 213.56 45.79 213.77 45.86 ;
    RECT 213.56 46.15 213.77 46.22 ;
    RECT 213.1 45.43 213.31 45.5 ;
    RECT 213.1 45.79 213.31 45.86 ;
    RECT 213.1 46.15 213.31 46.22 ;
    RECT 210.24 45.43 210.45 45.5 ;
    RECT 210.24 45.79 210.45 45.86 ;
    RECT 210.24 46.15 210.45 46.22 ;
    RECT 209.78 45.43 209.99 45.5 ;
    RECT 209.78 45.79 209.99 45.86 ;
    RECT 209.78 46.15 209.99 46.22 ;
    RECT 206.92 45.43 207.13 45.5 ;
    RECT 206.92 45.79 207.13 45.86 ;
    RECT 206.92 46.15 207.13 46.22 ;
    RECT 206.46 45.43 206.67 45.5 ;
    RECT 206.46 45.79 206.67 45.86 ;
    RECT 206.46 46.15 206.67 46.22 ;
    RECT 203.6 45.43 203.81 45.5 ;
    RECT 203.6 45.79 203.81 45.86 ;
    RECT 203.6 46.15 203.81 46.22 ;
    RECT 203.14 45.43 203.35 45.5 ;
    RECT 203.14 45.79 203.35 45.86 ;
    RECT 203.14 46.15 203.35 46.22 ;
    RECT 200.28 45.43 200.49 45.5 ;
    RECT 200.28 45.79 200.49 45.86 ;
    RECT 200.28 46.15 200.49 46.22 ;
    RECT 199.82 45.43 200.03 45.5 ;
    RECT 199.82 45.79 200.03 45.86 ;
    RECT 199.82 46.15 200.03 46.22 ;
    RECT 196.96 45.43 197.17 45.5 ;
    RECT 196.96 45.79 197.17 45.86 ;
    RECT 196.96 46.15 197.17 46.22 ;
    RECT 196.5 45.43 196.71 45.5 ;
    RECT 196.5 45.79 196.71 45.86 ;
    RECT 196.5 46.15 196.71 46.22 ;
    RECT 193.64 45.43 193.85 45.5 ;
    RECT 193.64 45.79 193.85 45.86 ;
    RECT 193.64 46.15 193.85 46.22 ;
    RECT 193.18 45.43 193.39 45.5 ;
    RECT 193.18 45.79 193.39 45.86 ;
    RECT 193.18 46.15 193.39 46.22 ;
    RECT 190.32 45.43 190.53 45.5 ;
    RECT 190.32 45.79 190.53 45.86 ;
    RECT 190.32 46.15 190.53 46.22 ;
    RECT 189.86 45.43 190.07 45.5 ;
    RECT 189.86 45.79 190.07 45.86 ;
    RECT 189.86 46.15 190.07 46.22 ;
    RECT 187.0 45.43 187.21 45.5 ;
    RECT 187.0 45.79 187.21 45.86 ;
    RECT 187.0 46.15 187.21 46.22 ;
    RECT 186.54 45.43 186.75 45.5 ;
    RECT 186.54 45.79 186.75 45.86 ;
    RECT 186.54 46.15 186.75 46.22 ;
    RECT 183.68 45.43 183.89 45.5 ;
    RECT 183.68 45.79 183.89 45.86 ;
    RECT 183.68 46.15 183.89 46.22 ;
    RECT 183.22 45.43 183.43 45.5 ;
    RECT 183.22 45.79 183.43 45.86 ;
    RECT 183.22 46.15 183.43 46.22 ;
    RECT 147.485 45.79 147.555 45.86 ;
    RECT 266.68 45.43 266.89 45.5 ;
    RECT 266.68 45.79 266.89 45.86 ;
    RECT 266.68 46.15 266.89 46.22 ;
    RECT 266.22 45.43 266.43 45.5 ;
    RECT 266.22 45.79 266.43 45.86 ;
    RECT 266.22 46.15 266.43 46.22 ;
    RECT 263.36 45.43 263.57 45.5 ;
    RECT 263.36 45.79 263.57 45.86 ;
    RECT 263.36 46.15 263.57 46.22 ;
    RECT 262.9 45.43 263.11 45.5 ;
    RECT 262.9 45.79 263.11 45.86 ;
    RECT 262.9 46.15 263.11 46.22 ;
    RECT 260.04 45.43 260.25 45.5 ;
    RECT 260.04 45.79 260.25 45.86 ;
    RECT 260.04 46.15 260.25 46.22 ;
    RECT 259.58 45.43 259.79 45.5 ;
    RECT 259.58 45.79 259.79 45.86 ;
    RECT 259.58 46.15 259.79 46.22 ;
    RECT 256.72 45.43 256.93 45.5 ;
    RECT 256.72 45.79 256.93 45.86 ;
    RECT 256.72 46.15 256.93 46.22 ;
    RECT 256.26 45.43 256.47 45.5 ;
    RECT 256.26 45.79 256.47 45.86 ;
    RECT 256.26 46.15 256.47 46.22 ;
    RECT 253.4 45.43 253.61 45.5 ;
    RECT 253.4 45.79 253.61 45.86 ;
    RECT 253.4 46.15 253.61 46.22 ;
    RECT 252.94 45.43 253.15 45.5 ;
    RECT 252.94 45.79 253.15 45.86 ;
    RECT 252.94 46.15 253.15 46.22 ;
    RECT 250.08 85.05 250.29 85.12 ;
    RECT 250.08 85.41 250.29 85.48 ;
    RECT 250.08 85.77 250.29 85.84 ;
    RECT 249.62 85.05 249.83 85.12 ;
    RECT 249.62 85.41 249.83 85.48 ;
    RECT 249.62 85.77 249.83 85.84 ;
    RECT 246.76 85.05 246.97 85.12 ;
    RECT 246.76 85.41 246.97 85.48 ;
    RECT 246.76 85.77 246.97 85.84 ;
    RECT 246.3 85.05 246.51 85.12 ;
    RECT 246.3 85.41 246.51 85.48 ;
    RECT 246.3 85.77 246.51 85.84 ;
    RECT 243.44 85.05 243.65 85.12 ;
    RECT 243.44 85.41 243.65 85.48 ;
    RECT 243.44 85.77 243.65 85.84 ;
    RECT 242.98 85.05 243.19 85.12 ;
    RECT 242.98 85.41 243.19 85.48 ;
    RECT 242.98 85.77 243.19 85.84 ;
    RECT 240.12 85.05 240.33 85.12 ;
    RECT 240.12 85.41 240.33 85.48 ;
    RECT 240.12 85.77 240.33 85.84 ;
    RECT 239.66 85.05 239.87 85.12 ;
    RECT 239.66 85.41 239.87 85.48 ;
    RECT 239.66 85.77 239.87 85.84 ;
    RECT 236.8 85.05 237.01 85.12 ;
    RECT 236.8 85.41 237.01 85.48 ;
    RECT 236.8 85.77 237.01 85.84 ;
    RECT 236.34 85.05 236.55 85.12 ;
    RECT 236.34 85.41 236.55 85.48 ;
    RECT 236.34 85.77 236.55 85.84 ;
    RECT 233.48 85.05 233.69 85.12 ;
    RECT 233.48 85.41 233.69 85.48 ;
    RECT 233.48 85.77 233.69 85.84 ;
    RECT 233.02 85.05 233.23 85.12 ;
    RECT 233.02 85.41 233.23 85.48 ;
    RECT 233.02 85.77 233.23 85.84 ;
    RECT 230.16 85.05 230.37 85.12 ;
    RECT 230.16 85.41 230.37 85.48 ;
    RECT 230.16 85.77 230.37 85.84 ;
    RECT 229.7 85.05 229.91 85.12 ;
    RECT 229.7 85.41 229.91 85.48 ;
    RECT 229.7 85.77 229.91 85.84 ;
    RECT 226.84 85.05 227.05 85.12 ;
    RECT 226.84 85.41 227.05 85.48 ;
    RECT 226.84 85.77 227.05 85.84 ;
    RECT 226.38 85.05 226.59 85.12 ;
    RECT 226.38 85.41 226.59 85.48 ;
    RECT 226.38 85.77 226.59 85.84 ;
    RECT 223.52 85.05 223.73 85.12 ;
    RECT 223.52 85.41 223.73 85.48 ;
    RECT 223.52 85.77 223.73 85.84 ;
    RECT 223.06 85.05 223.27 85.12 ;
    RECT 223.06 85.41 223.27 85.48 ;
    RECT 223.06 85.77 223.27 85.84 ;
    RECT 220.2 85.05 220.41 85.12 ;
    RECT 220.2 85.41 220.41 85.48 ;
    RECT 220.2 85.77 220.41 85.84 ;
    RECT 219.74 85.05 219.95 85.12 ;
    RECT 219.74 85.41 219.95 85.48 ;
    RECT 219.74 85.77 219.95 85.84 ;
    RECT 216.88 85.05 217.09 85.12 ;
    RECT 216.88 85.41 217.09 85.48 ;
    RECT 216.88 85.77 217.09 85.84 ;
    RECT 216.42 85.05 216.63 85.12 ;
    RECT 216.42 85.41 216.63 85.48 ;
    RECT 216.42 85.77 216.63 85.84 ;
    RECT 267.91 85.41 267.98 85.48 ;
    RECT 180.36 85.05 180.57 85.12 ;
    RECT 180.36 85.41 180.57 85.48 ;
    RECT 180.36 85.77 180.57 85.84 ;
    RECT 179.9 85.05 180.11 85.12 ;
    RECT 179.9 85.41 180.11 85.48 ;
    RECT 179.9 85.77 180.11 85.84 ;
    RECT 177.04 85.05 177.25 85.12 ;
    RECT 177.04 85.41 177.25 85.48 ;
    RECT 177.04 85.77 177.25 85.84 ;
    RECT 176.58 85.05 176.79 85.12 ;
    RECT 176.58 85.41 176.79 85.48 ;
    RECT 176.58 85.77 176.79 85.84 ;
    RECT 173.72 85.05 173.93 85.12 ;
    RECT 173.72 85.41 173.93 85.48 ;
    RECT 173.72 85.77 173.93 85.84 ;
    RECT 173.26 85.05 173.47 85.12 ;
    RECT 173.26 85.41 173.47 85.48 ;
    RECT 173.26 85.77 173.47 85.84 ;
    RECT 170.4 85.05 170.61 85.12 ;
    RECT 170.4 85.41 170.61 85.48 ;
    RECT 170.4 85.77 170.61 85.84 ;
    RECT 169.94 85.05 170.15 85.12 ;
    RECT 169.94 85.41 170.15 85.48 ;
    RECT 169.94 85.77 170.15 85.84 ;
    RECT 167.08 85.05 167.29 85.12 ;
    RECT 167.08 85.41 167.29 85.48 ;
    RECT 167.08 85.77 167.29 85.84 ;
    RECT 166.62 85.05 166.83 85.12 ;
    RECT 166.62 85.41 166.83 85.48 ;
    RECT 166.62 85.77 166.83 85.84 ;
    RECT 163.76 85.05 163.97 85.12 ;
    RECT 163.76 85.41 163.97 85.48 ;
    RECT 163.76 85.77 163.97 85.84 ;
    RECT 163.3 85.05 163.51 85.12 ;
    RECT 163.3 85.41 163.51 85.48 ;
    RECT 163.3 85.77 163.51 85.84 ;
    RECT 160.44 85.05 160.65 85.12 ;
    RECT 160.44 85.41 160.65 85.48 ;
    RECT 160.44 85.77 160.65 85.84 ;
    RECT 159.98 85.05 160.19 85.12 ;
    RECT 159.98 85.41 160.19 85.48 ;
    RECT 159.98 85.77 160.19 85.84 ;
    RECT 157.12 85.05 157.33 85.12 ;
    RECT 157.12 85.41 157.33 85.48 ;
    RECT 157.12 85.77 157.33 85.84 ;
    RECT 156.66 85.05 156.87 85.12 ;
    RECT 156.66 85.41 156.87 85.48 ;
    RECT 156.66 85.77 156.87 85.84 ;
    RECT 153.8 85.05 154.01 85.12 ;
    RECT 153.8 85.41 154.01 85.48 ;
    RECT 153.8 85.77 154.01 85.84 ;
    RECT 153.34 85.05 153.55 85.12 ;
    RECT 153.34 85.41 153.55 85.48 ;
    RECT 153.34 85.77 153.55 85.84 ;
    RECT 150.48 85.05 150.69 85.12 ;
    RECT 150.48 85.41 150.69 85.48 ;
    RECT 150.48 85.77 150.69 85.84 ;
    RECT 150.02 85.05 150.23 85.12 ;
    RECT 150.02 85.41 150.23 85.48 ;
    RECT 150.02 85.77 150.23 85.84 ;
    RECT 213.56 85.05 213.77 85.12 ;
    RECT 213.56 85.41 213.77 85.48 ;
    RECT 213.56 85.77 213.77 85.84 ;
    RECT 213.1 85.05 213.31 85.12 ;
    RECT 213.1 85.41 213.31 85.48 ;
    RECT 213.1 85.77 213.31 85.84 ;
    RECT 210.24 85.05 210.45 85.12 ;
    RECT 210.24 85.41 210.45 85.48 ;
    RECT 210.24 85.77 210.45 85.84 ;
    RECT 209.78 85.05 209.99 85.12 ;
    RECT 209.78 85.41 209.99 85.48 ;
    RECT 209.78 85.77 209.99 85.84 ;
    RECT 206.92 85.05 207.13 85.12 ;
    RECT 206.92 85.41 207.13 85.48 ;
    RECT 206.92 85.77 207.13 85.84 ;
    RECT 206.46 85.05 206.67 85.12 ;
    RECT 206.46 85.41 206.67 85.48 ;
    RECT 206.46 85.77 206.67 85.84 ;
    RECT 203.6 85.05 203.81 85.12 ;
    RECT 203.6 85.41 203.81 85.48 ;
    RECT 203.6 85.77 203.81 85.84 ;
    RECT 203.14 85.05 203.35 85.12 ;
    RECT 203.14 85.41 203.35 85.48 ;
    RECT 203.14 85.77 203.35 85.84 ;
    RECT 200.28 85.05 200.49 85.12 ;
    RECT 200.28 85.41 200.49 85.48 ;
    RECT 200.28 85.77 200.49 85.84 ;
    RECT 199.82 85.05 200.03 85.12 ;
    RECT 199.82 85.41 200.03 85.48 ;
    RECT 199.82 85.77 200.03 85.84 ;
    RECT 196.96 85.05 197.17 85.12 ;
    RECT 196.96 85.41 197.17 85.48 ;
    RECT 196.96 85.77 197.17 85.84 ;
    RECT 196.5 85.05 196.71 85.12 ;
    RECT 196.5 85.41 196.71 85.48 ;
    RECT 196.5 85.77 196.71 85.84 ;
    RECT 193.64 85.05 193.85 85.12 ;
    RECT 193.64 85.41 193.85 85.48 ;
    RECT 193.64 85.77 193.85 85.84 ;
    RECT 193.18 85.05 193.39 85.12 ;
    RECT 193.18 85.41 193.39 85.48 ;
    RECT 193.18 85.77 193.39 85.84 ;
    RECT 190.32 85.05 190.53 85.12 ;
    RECT 190.32 85.41 190.53 85.48 ;
    RECT 190.32 85.77 190.53 85.84 ;
    RECT 189.86 85.05 190.07 85.12 ;
    RECT 189.86 85.41 190.07 85.48 ;
    RECT 189.86 85.77 190.07 85.84 ;
    RECT 187.0 85.05 187.21 85.12 ;
    RECT 187.0 85.41 187.21 85.48 ;
    RECT 187.0 85.77 187.21 85.84 ;
    RECT 186.54 85.05 186.75 85.12 ;
    RECT 186.54 85.41 186.75 85.48 ;
    RECT 186.54 85.77 186.75 85.84 ;
    RECT 183.68 85.05 183.89 85.12 ;
    RECT 183.68 85.41 183.89 85.48 ;
    RECT 183.68 85.77 183.89 85.84 ;
    RECT 183.22 85.05 183.43 85.12 ;
    RECT 183.22 85.41 183.43 85.48 ;
    RECT 183.22 85.77 183.43 85.84 ;
    RECT 147.485 85.41 147.555 85.48 ;
    RECT 266.68 85.05 266.89 85.12 ;
    RECT 266.68 85.41 266.89 85.48 ;
    RECT 266.68 85.77 266.89 85.84 ;
    RECT 266.22 85.05 266.43 85.12 ;
    RECT 266.22 85.41 266.43 85.48 ;
    RECT 266.22 85.77 266.43 85.84 ;
    RECT 263.36 85.05 263.57 85.12 ;
    RECT 263.36 85.41 263.57 85.48 ;
    RECT 263.36 85.77 263.57 85.84 ;
    RECT 262.9 85.05 263.11 85.12 ;
    RECT 262.9 85.41 263.11 85.48 ;
    RECT 262.9 85.77 263.11 85.84 ;
    RECT 260.04 85.05 260.25 85.12 ;
    RECT 260.04 85.41 260.25 85.48 ;
    RECT 260.04 85.77 260.25 85.84 ;
    RECT 259.58 85.05 259.79 85.12 ;
    RECT 259.58 85.41 259.79 85.48 ;
    RECT 259.58 85.77 259.79 85.84 ;
    RECT 256.72 85.05 256.93 85.12 ;
    RECT 256.72 85.41 256.93 85.48 ;
    RECT 256.72 85.77 256.93 85.84 ;
    RECT 256.26 85.05 256.47 85.12 ;
    RECT 256.26 85.41 256.47 85.48 ;
    RECT 256.26 85.77 256.47 85.84 ;
    RECT 253.4 85.05 253.61 85.12 ;
    RECT 253.4 85.41 253.61 85.48 ;
    RECT 253.4 85.77 253.61 85.84 ;
    RECT 252.94 85.05 253.15 85.12 ;
    RECT 252.94 85.41 253.15 85.48 ;
    RECT 252.94 85.77 253.15 85.84 ;
    RECT 250.08 44.71 250.29 44.78 ;
    RECT 250.08 45.07 250.29 45.14 ;
    RECT 250.08 45.43 250.29 45.5 ;
    RECT 249.62 44.71 249.83 44.78 ;
    RECT 249.62 45.07 249.83 45.14 ;
    RECT 249.62 45.43 249.83 45.5 ;
    RECT 246.76 44.71 246.97 44.78 ;
    RECT 246.76 45.07 246.97 45.14 ;
    RECT 246.76 45.43 246.97 45.5 ;
    RECT 246.3 44.71 246.51 44.78 ;
    RECT 246.3 45.07 246.51 45.14 ;
    RECT 246.3 45.43 246.51 45.5 ;
    RECT 243.44 44.71 243.65 44.78 ;
    RECT 243.44 45.07 243.65 45.14 ;
    RECT 243.44 45.43 243.65 45.5 ;
    RECT 242.98 44.71 243.19 44.78 ;
    RECT 242.98 45.07 243.19 45.14 ;
    RECT 242.98 45.43 243.19 45.5 ;
    RECT 240.12 44.71 240.33 44.78 ;
    RECT 240.12 45.07 240.33 45.14 ;
    RECT 240.12 45.43 240.33 45.5 ;
    RECT 239.66 44.71 239.87 44.78 ;
    RECT 239.66 45.07 239.87 45.14 ;
    RECT 239.66 45.43 239.87 45.5 ;
    RECT 236.8 44.71 237.01 44.78 ;
    RECT 236.8 45.07 237.01 45.14 ;
    RECT 236.8 45.43 237.01 45.5 ;
    RECT 236.34 44.71 236.55 44.78 ;
    RECT 236.34 45.07 236.55 45.14 ;
    RECT 236.34 45.43 236.55 45.5 ;
    RECT 233.48 44.71 233.69 44.78 ;
    RECT 233.48 45.07 233.69 45.14 ;
    RECT 233.48 45.43 233.69 45.5 ;
    RECT 233.02 44.71 233.23 44.78 ;
    RECT 233.02 45.07 233.23 45.14 ;
    RECT 233.02 45.43 233.23 45.5 ;
    RECT 230.16 44.71 230.37 44.78 ;
    RECT 230.16 45.07 230.37 45.14 ;
    RECT 230.16 45.43 230.37 45.5 ;
    RECT 229.7 44.71 229.91 44.78 ;
    RECT 229.7 45.07 229.91 45.14 ;
    RECT 229.7 45.43 229.91 45.5 ;
    RECT 226.84 44.71 227.05 44.78 ;
    RECT 226.84 45.07 227.05 45.14 ;
    RECT 226.84 45.43 227.05 45.5 ;
    RECT 226.38 44.71 226.59 44.78 ;
    RECT 226.38 45.07 226.59 45.14 ;
    RECT 226.38 45.43 226.59 45.5 ;
    RECT 223.52 44.71 223.73 44.78 ;
    RECT 223.52 45.07 223.73 45.14 ;
    RECT 223.52 45.43 223.73 45.5 ;
    RECT 223.06 44.71 223.27 44.78 ;
    RECT 223.06 45.07 223.27 45.14 ;
    RECT 223.06 45.43 223.27 45.5 ;
    RECT 220.2 44.71 220.41 44.78 ;
    RECT 220.2 45.07 220.41 45.14 ;
    RECT 220.2 45.43 220.41 45.5 ;
    RECT 219.74 44.71 219.95 44.78 ;
    RECT 219.74 45.07 219.95 45.14 ;
    RECT 219.74 45.43 219.95 45.5 ;
    RECT 216.88 44.71 217.09 44.78 ;
    RECT 216.88 45.07 217.09 45.14 ;
    RECT 216.88 45.43 217.09 45.5 ;
    RECT 216.42 44.71 216.63 44.78 ;
    RECT 216.42 45.07 216.63 45.14 ;
    RECT 216.42 45.43 216.63 45.5 ;
    RECT 267.91 45.07 267.98 45.14 ;
    RECT 180.36 44.71 180.57 44.78 ;
    RECT 180.36 45.07 180.57 45.14 ;
    RECT 180.36 45.43 180.57 45.5 ;
    RECT 179.9 44.71 180.11 44.78 ;
    RECT 179.9 45.07 180.11 45.14 ;
    RECT 179.9 45.43 180.11 45.5 ;
    RECT 177.04 44.71 177.25 44.78 ;
    RECT 177.04 45.07 177.25 45.14 ;
    RECT 177.04 45.43 177.25 45.5 ;
    RECT 176.58 44.71 176.79 44.78 ;
    RECT 176.58 45.07 176.79 45.14 ;
    RECT 176.58 45.43 176.79 45.5 ;
    RECT 173.72 44.71 173.93 44.78 ;
    RECT 173.72 45.07 173.93 45.14 ;
    RECT 173.72 45.43 173.93 45.5 ;
    RECT 173.26 44.71 173.47 44.78 ;
    RECT 173.26 45.07 173.47 45.14 ;
    RECT 173.26 45.43 173.47 45.5 ;
    RECT 170.4 44.71 170.61 44.78 ;
    RECT 170.4 45.07 170.61 45.14 ;
    RECT 170.4 45.43 170.61 45.5 ;
    RECT 169.94 44.71 170.15 44.78 ;
    RECT 169.94 45.07 170.15 45.14 ;
    RECT 169.94 45.43 170.15 45.5 ;
    RECT 167.08 44.71 167.29 44.78 ;
    RECT 167.08 45.07 167.29 45.14 ;
    RECT 167.08 45.43 167.29 45.5 ;
    RECT 166.62 44.71 166.83 44.78 ;
    RECT 166.62 45.07 166.83 45.14 ;
    RECT 166.62 45.43 166.83 45.5 ;
    RECT 163.76 44.71 163.97 44.78 ;
    RECT 163.76 45.07 163.97 45.14 ;
    RECT 163.76 45.43 163.97 45.5 ;
    RECT 163.3 44.71 163.51 44.78 ;
    RECT 163.3 45.07 163.51 45.14 ;
    RECT 163.3 45.43 163.51 45.5 ;
    RECT 160.44 44.71 160.65 44.78 ;
    RECT 160.44 45.07 160.65 45.14 ;
    RECT 160.44 45.43 160.65 45.5 ;
    RECT 159.98 44.71 160.19 44.78 ;
    RECT 159.98 45.07 160.19 45.14 ;
    RECT 159.98 45.43 160.19 45.5 ;
    RECT 157.12 44.71 157.33 44.78 ;
    RECT 157.12 45.07 157.33 45.14 ;
    RECT 157.12 45.43 157.33 45.5 ;
    RECT 156.66 44.71 156.87 44.78 ;
    RECT 156.66 45.07 156.87 45.14 ;
    RECT 156.66 45.43 156.87 45.5 ;
    RECT 153.8 44.71 154.01 44.78 ;
    RECT 153.8 45.07 154.01 45.14 ;
    RECT 153.8 45.43 154.01 45.5 ;
    RECT 153.34 44.71 153.55 44.78 ;
    RECT 153.34 45.07 153.55 45.14 ;
    RECT 153.34 45.43 153.55 45.5 ;
    RECT 150.48 44.71 150.69 44.78 ;
    RECT 150.48 45.07 150.69 45.14 ;
    RECT 150.48 45.43 150.69 45.5 ;
    RECT 150.02 44.71 150.23 44.78 ;
    RECT 150.02 45.07 150.23 45.14 ;
    RECT 150.02 45.43 150.23 45.5 ;
    RECT 213.56 44.71 213.77 44.78 ;
    RECT 213.56 45.07 213.77 45.14 ;
    RECT 213.56 45.43 213.77 45.5 ;
    RECT 213.1 44.71 213.31 44.78 ;
    RECT 213.1 45.07 213.31 45.14 ;
    RECT 213.1 45.43 213.31 45.5 ;
    RECT 210.24 44.71 210.45 44.78 ;
    RECT 210.24 45.07 210.45 45.14 ;
    RECT 210.24 45.43 210.45 45.5 ;
    RECT 209.78 44.71 209.99 44.78 ;
    RECT 209.78 45.07 209.99 45.14 ;
    RECT 209.78 45.43 209.99 45.5 ;
    RECT 206.92 44.71 207.13 44.78 ;
    RECT 206.92 45.07 207.13 45.14 ;
    RECT 206.92 45.43 207.13 45.5 ;
    RECT 206.46 44.71 206.67 44.78 ;
    RECT 206.46 45.07 206.67 45.14 ;
    RECT 206.46 45.43 206.67 45.5 ;
    RECT 203.6 44.71 203.81 44.78 ;
    RECT 203.6 45.07 203.81 45.14 ;
    RECT 203.6 45.43 203.81 45.5 ;
    RECT 203.14 44.71 203.35 44.78 ;
    RECT 203.14 45.07 203.35 45.14 ;
    RECT 203.14 45.43 203.35 45.5 ;
    RECT 200.28 44.71 200.49 44.78 ;
    RECT 200.28 45.07 200.49 45.14 ;
    RECT 200.28 45.43 200.49 45.5 ;
    RECT 199.82 44.71 200.03 44.78 ;
    RECT 199.82 45.07 200.03 45.14 ;
    RECT 199.82 45.43 200.03 45.5 ;
    RECT 196.96 44.71 197.17 44.78 ;
    RECT 196.96 45.07 197.17 45.14 ;
    RECT 196.96 45.43 197.17 45.5 ;
    RECT 196.5 44.71 196.71 44.78 ;
    RECT 196.5 45.07 196.71 45.14 ;
    RECT 196.5 45.43 196.71 45.5 ;
    RECT 193.64 44.71 193.85 44.78 ;
    RECT 193.64 45.07 193.85 45.14 ;
    RECT 193.64 45.43 193.85 45.5 ;
    RECT 193.18 44.71 193.39 44.78 ;
    RECT 193.18 45.07 193.39 45.14 ;
    RECT 193.18 45.43 193.39 45.5 ;
    RECT 190.32 44.71 190.53 44.78 ;
    RECT 190.32 45.07 190.53 45.14 ;
    RECT 190.32 45.43 190.53 45.5 ;
    RECT 189.86 44.71 190.07 44.78 ;
    RECT 189.86 45.07 190.07 45.14 ;
    RECT 189.86 45.43 190.07 45.5 ;
    RECT 187.0 44.71 187.21 44.78 ;
    RECT 187.0 45.07 187.21 45.14 ;
    RECT 187.0 45.43 187.21 45.5 ;
    RECT 186.54 44.71 186.75 44.78 ;
    RECT 186.54 45.07 186.75 45.14 ;
    RECT 186.54 45.43 186.75 45.5 ;
    RECT 183.68 44.71 183.89 44.78 ;
    RECT 183.68 45.07 183.89 45.14 ;
    RECT 183.68 45.43 183.89 45.5 ;
    RECT 183.22 44.71 183.43 44.78 ;
    RECT 183.22 45.07 183.43 45.14 ;
    RECT 183.22 45.43 183.43 45.5 ;
    RECT 147.485 45.07 147.555 45.14 ;
    RECT 266.68 44.71 266.89 44.78 ;
    RECT 266.68 45.07 266.89 45.14 ;
    RECT 266.68 45.43 266.89 45.5 ;
    RECT 266.22 44.71 266.43 44.78 ;
    RECT 266.22 45.07 266.43 45.14 ;
    RECT 266.22 45.43 266.43 45.5 ;
    RECT 263.36 44.71 263.57 44.78 ;
    RECT 263.36 45.07 263.57 45.14 ;
    RECT 263.36 45.43 263.57 45.5 ;
    RECT 262.9 44.71 263.11 44.78 ;
    RECT 262.9 45.07 263.11 45.14 ;
    RECT 262.9 45.43 263.11 45.5 ;
    RECT 260.04 44.71 260.25 44.78 ;
    RECT 260.04 45.07 260.25 45.14 ;
    RECT 260.04 45.43 260.25 45.5 ;
    RECT 259.58 44.71 259.79 44.78 ;
    RECT 259.58 45.07 259.79 45.14 ;
    RECT 259.58 45.43 259.79 45.5 ;
    RECT 256.72 44.71 256.93 44.78 ;
    RECT 256.72 45.07 256.93 45.14 ;
    RECT 256.72 45.43 256.93 45.5 ;
    RECT 256.26 44.71 256.47 44.78 ;
    RECT 256.26 45.07 256.47 45.14 ;
    RECT 256.26 45.43 256.47 45.5 ;
    RECT 253.4 44.71 253.61 44.78 ;
    RECT 253.4 45.07 253.61 45.14 ;
    RECT 253.4 45.43 253.61 45.5 ;
    RECT 252.94 44.71 253.15 44.78 ;
    RECT 252.94 45.07 253.15 45.14 ;
    RECT 252.94 45.43 253.15 45.5 ;
    RECT 250.08 84.33 250.29 84.4 ;
    RECT 250.08 84.69 250.29 84.76 ;
    RECT 250.08 85.05 250.29 85.12 ;
    RECT 249.62 84.33 249.83 84.4 ;
    RECT 249.62 84.69 249.83 84.76 ;
    RECT 249.62 85.05 249.83 85.12 ;
    RECT 246.76 84.33 246.97 84.4 ;
    RECT 246.76 84.69 246.97 84.76 ;
    RECT 246.76 85.05 246.97 85.12 ;
    RECT 246.3 84.33 246.51 84.4 ;
    RECT 246.3 84.69 246.51 84.76 ;
    RECT 246.3 85.05 246.51 85.12 ;
    RECT 243.44 84.33 243.65 84.4 ;
    RECT 243.44 84.69 243.65 84.76 ;
    RECT 243.44 85.05 243.65 85.12 ;
    RECT 242.98 84.33 243.19 84.4 ;
    RECT 242.98 84.69 243.19 84.76 ;
    RECT 242.98 85.05 243.19 85.12 ;
    RECT 240.12 84.33 240.33 84.4 ;
    RECT 240.12 84.69 240.33 84.76 ;
    RECT 240.12 85.05 240.33 85.12 ;
    RECT 239.66 84.33 239.87 84.4 ;
    RECT 239.66 84.69 239.87 84.76 ;
    RECT 239.66 85.05 239.87 85.12 ;
    RECT 236.8 84.33 237.01 84.4 ;
    RECT 236.8 84.69 237.01 84.76 ;
    RECT 236.8 85.05 237.01 85.12 ;
    RECT 236.34 84.33 236.55 84.4 ;
    RECT 236.34 84.69 236.55 84.76 ;
    RECT 236.34 85.05 236.55 85.12 ;
    RECT 233.48 84.33 233.69 84.4 ;
    RECT 233.48 84.69 233.69 84.76 ;
    RECT 233.48 85.05 233.69 85.12 ;
    RECT 233.02 84.33 233.23 84.4 ;
    RECT 233.02 84.69 233.23 84.76 ;
    RECT 233.02 85.05 233.23 85.12 ;
    RECT 230.16 84.33 230.37 84.4 ;
    RECT 230.16 84.69 230.37 84.76 ;
    RECT 230.16 85.05 230.37 85.12 ;
    RECT 229.7 84.33 229.91 84.4 ;
    RECT 229.7 84.69 229.91 84.76 ;
    RECT 229.7 85.05 229.91 85.12 ;
    RECT 226.84 84.33 227.05 84.4 ;
    RECT 226.84 84.69 227.05 84.76 ;
    RECT 226.84 85.05 227.05 85.12 ;
    RECT 226.38 84.33 226.59 84.4 ;
    RECT 226.38 84.69 226.59 84.76 ;
    RECT 226.38 85.05 226.59 85.12 ;
    RECT 223.52 84.33 223.73 84.4 ;
    RECT 223.52 84.69 223.73 84.76 ;
    RECT 223.52 85.05 223.73 85.12 ;
    RECT 223.06 84.33 223.27 84.4 ;
    RECT 223.06 84.69 223.27 84.76 ;
    RECT 223.06 85.05 223.27 85.12 ;
    RECT 220.2 84.33 220.41 84.4 ;
    RECT 220.2 84.69 220.41 84.76 ;
    RECT 220.2 85.05 220.41 85.12 ;
    RECT 219.74 84.33 219.95 84.4 ;
    RECT 219.74 84.69 219.95 84.76 ;
    RECT 219.74 85.05 219.95 85.12 ;
    RECT 216.88 84.33 217.09 84.4 ;
    RECT 216.88 84.69 217.09 84.76 ;
    RECT 216.88 85.05 217.09 85.12 ;
    RECT 216.42 84.33 216.63 84.4 ;
    RECT 216.42 84.69 216.63 84.76 ;
    RECT 216.42 85.05 216.63 85.12 ;
    RECT 267.91 84.69 267.98 84.76 ;
    RECT 180.36 84.33 180.57 84.4 ;
    RECT 180.36 84.69 180.57 84.76 ;
    RECT 180.36 85.05 180.57 85.12 ;
    RECT 179.9 84.33 180.11 84.4 ;
    RECT 179.9 84.69 180.11 84.76 ;
    RECT 179.9 85.05 180.11 85.12 ;
    RECT 177.04 84.33 177.25 84.4 ;
    RECT 177.04 84.69 177.25 84.76 ;
    RECT 177.04 85.05 177.25 85.12 ;
    RECT 176.58 84.33 176.79 84.4 ;
    RECT 176.58 84.69 176.79 84.76 ;
    RECT 176.58 85.05 176.79 85.12 ;
    RECT 173.72 84.33 173.93 84.4 ;
    RECT 173.72 84.69 173.93 84.76 ;
    RECT 173.72 85.05 173.93 85.12 ;
    RECT 173.26 84.33 173.47 84.4 ;
    RECT 173.26 84.69 173.47 84.76 ;
    RECT 173.26 85.05 173.47 85.12 ;
    RECT 170.4 84.33 170.61 84.4 ;
    RECT 170.4 84.69 170.61 84.76 ;
    RECT 170.4 85.05 170.61 85.12 ;
    RECT 169.94 84.33 170.15 84.4 ;
    RECT 169.94 84.69 170.15 84.76 ;
    RECT 169.94 85.05 170.15 85.12 ;
    RECT 167.08 84.33 167.29 84.4 ;
    RECT 167.08 84.69 167.29 84.76 ;
    RECT 167.08 85.05 167.29 85.12 ;
    RECT 166.62 84.33 166.83 84.4 ;
    RECT 166.62 84.69 166.83 84.76 ;
    RECT 166.62 85.05 166.83 85.12 ;
    RECT 163.76 84.33 163.97 84.4 ;
    RECT 163.76 84.69 163.97 84.76 ;
    RECT 163.76 85.05 163.97 85.12 ;
    RECT 163.3 84.33 163.51 84.4 ;
    RECT 163.3 84.69 163.51 84.76 ;
    RECT 163.3 85.05 163.51 85.12 ;
    RECT 160.44 84.33 160.65 84.4 ;
    RECT 160.44 84.69 160.65 84.76 ;
    RECT 160.44 85.05 160.65 85.12 ;
    RECT 159.98 84.33 160.19 84.4 ;
    RECT 159.98 84.69 160.19 84.76 ;
    RECT 159.98 85.05 160.19 85.12 ;
    RECT 157.12 84.33 157.33 84.4 ;
    RECT 157.12 84.69 157.33 84.76 ;
    RECT 157.12 85.05 157.33 85.12 ;
    RECT 156.66 84.33 156.87 84.4 ;
    RECT 156.66 84.69 156.87 84.76 ;
    RECT 156.66 85.05 156.87 85.12 ;
    RECT 153.8 84.33 154.01 84.4 ;
    RECT 153.8 84.69 154.01 84.76 ;
    RECT 153.8 85.05 154.01 85.12 ;
    RECT 153.34 84.33 153.55 84.4 ;
    RECT 153.34 84.69 153.55 84.76 ;
    RECT 153.34 85.05 153.55 85.12 ;
    RECT 150.48 84.33 150.69 84.4 ;
    RECT 150.48 84.69 150.69 84.76 ;
    RECT 150.48 85.05 150.69 85.12 ;
    RECT 150.02 84.33 150.23 84.4 ;
    RECT 150.02 84.69 150.23 84.76 ;
    RECT 150.02 85.05 150.23 85.12 ;
    RECT 213.56 84.33 213.77 84.4 ;
    RECT 213.56 84.69 213.77 84.76 ;
    RECT 213.56 85.05 213.77 85.12 ;
    RECT 213.1 84.33 213.31 84.4 ;
    RECT 213.1 84.69 213.31 84.76 ;
    RECT 213.1 85.05 213.31 85.12 ;
    RECT 210.24 84.33 210.45 84.4 ;
    RECT 210.24 84.69 210.45 84.76 ;
    RECT 210.24 85.05 210.45 85.12 ;
    RECT 209.78 84.33 209.99 84.4 ;
    RECT 209.78 84.69 209.99 84.76 ;
    RECT 209.78 85.05 209.99 85.12 ;
    RECT 206.92 84.33 207.13 84.4 ;
    RECT 206.92 84.69 207.13 84.76 ;
    RECT 206.92 85.05 207.13 85.12 ;
    RECT 206.46 84.33 206.67 84.4 ;
    RECT 206.46 84.69 206.67 84.76 ;
    RECT 206.46 85.05 206.67 85.12 ;
    RECT 203.6 84.33 203.81 84.4 ;
    RECT 203.6 84.69 203.81 84.76 ;
    RECT 203.6 85.05 203.81 85.12 ;
    RECT 203.14 84.33 203.35 84.4 ;
    RECT 203.14 84.69 203.35 84.76 ;
    RECT 203.14 85.05 203.35 85.12 ;
    RECT 200.28 84.33 200.49 84.4 ;
    RECT 200.28 84.69 200.49 84.76 ;
    RECT 200.28 85.05 200.49 85.12 ;
    RECT 199.82 84.33 200.03 84.4 ;
    RECT 199.82 84.69 200.03 84.76 ;
    RECT 199.82 85.05 200.03 85.12 ;
    RECT 196.96 84.33 197.17 84.4 ;
    RECT 196.96 84.69 197.17 84.76 ;
    RECT 196.96 85.05 197.17 85.12 ;
    RECT 196.5 84.33 196.71 84.4 ;
    RECT 196.5 84.69 196.71 84.76 ;
    RECT 196.5 85.05 196.71 85.12 ;
    RECT 193.64 84.33 193.85 84.4 ;
    RECT 193.64 84.69 193.85 84.76 ;
    RECT 193.64 85.05 193.85 85.12 ;
    RECT 193.18 84.33 193.39 84.4 ;
    RECT 193.18 84.69 193.39 84.76 ;
    RECT 193.18 85.05 193.39 85.12 ;
    RECT 190.32 84.33 190.53 84.4 ;
    RECT 190.32 84.69 190.53 84.76 ;
    RECT 190.32 85.05 190.53 85.12 ;
    RECT 189.86 84.33 190.07 84.4 ;
    RECT 189.86 84.69 190.07 84.76 ;
    RECT 189.86 85.05 190.07 85.12 ;
    RECT 187.0 84.33 187.21 84.4 ;
    RECT 187.0 84.69 187.21 84.76 ;
    RECT 187.0 85.05 187.21 85.12 ;
    RECT 186.54 84.33 186.75 84.4 ;
    RECT 186.54 84.69 186.75 84.76 ;
    RECT 186.54 85.05 186.75 85.12 ;
    RECT 183.68 84.33 183.89 84.4 ;
    RECT 183.68 84.69 183.89 84.76 ;
    RECT 183.68 85.05 183.89 85.12 ;
    RECT 183.22 84.33 183.43 84.4 ;
    RECT 183.22 84.69 183.43 84.76 ;
    RECT 183.22 85.05 183.43 85.12 ;
    RECT 147.485 84.69 147.555 84.76 ;
    RECT 266.68 84.33 266.89 84.4 ;
    RECT 266.68 84.69 266.89 84.76 ;
    RECT 266.68 85.05 266.89 85.12 ;
    RECT 266.22 84.33 266.43 84.4 ;
    RECT 266.22 84.69 266.43 84.76 ;
    RECT 266.22 85.05 266.43 85.12 ;
    RECT 263.36 84.33 263.57 84.4 ;
    RECT 263.36 84.69 263.57 84.76 ;
    RECT 263.36 85.05 263.57 85.12 ;
    RECT 262.9 84.33 263.11 84.4 ;
    RECT 262.9 84.69 263.11 84.76 ;
    RECT 262.9 85.05 263.11 85.12 ;
    RECT 260.04 84.33 260.25 84.4 ;
    RECT 260.04 84.69 260.25 84.76 ;
    RECT 260.04 85.05 260.25 85.12 ;
    RECT 259.58 84.33 259.79 84.4 ;
    RECT 259.58 84.69 259.79 84.76 ;
    RECT 259.58 85.05 259.79 85.12 ;
    RECT 256.72 84.33 256.93 84.4 ;
    RECT 256.72 84.69 256.93 84.76 ;
    RECT 256.72 85.05 256.93 85.12 ;
    RECT 256.26 84.33 256.47 84.4 ;
    RECT 256.26 84.69 256.47 84.76 ;
    RECT 256.26 85.05 256.47 85.12 ;
    RECT 253.4 84.33 253.61 84.4 ;
    RECT 253.4 84.69 253.61 84.76 ;
    RECT 253.4 85.05 253.61 85.12 ;
    RECT 252.94 84.33 253.15 84.4 ;
    RECT 252.94 84.69 253.15 84.76 ;
    RECT 252.94 85.05 253.15 85.12 ;
    RECT 250.08 43.99 250.29 44.06 ;
    RECT 250.08 44.35 250.29 44.42 ;
    RECT 250.08 44.71 250.29 44.78 ;
    RECT 249.62 43.99 249.83 44.06 ;
    RECT 249.62 44.35 249.83 44.42 ;
    RECT 249.62 44.71 249.83 44.78 ;
    RECT 246.76 43.99 246.97 44.06 ;
    RECT 246.76 44.35 246.97 44.42 ;
    RECT 246.76 44.71 246.97 44.78 ;
    RECT 246.3 43.99 246.51 44.06 ;
    RECT 246.3 44.35 246.51 44.42 ;
    RECT 246.3 44.71 246.51 44.78 ;
    RECT 243.44 43.99 243.65 44.06 ;
    RECT 243.44 44.35 243.65 44.42 ;
    RECT 243.44 44.71 243.65 44.78 ;
    RECT 242.98 43.99 243.19 44.06 ;
    RECT 242.98 44.35 243.19 44.42 ;
    RECT 242.98 44.71 243.19 44.78 ;
    RECT 240.12 43.99 240.33 44.06 ;
    RECT 240.12 44.35 240.33 44.42 ;
    RECT 240.12 44.71 240.33 44.78 ;
    RECT 239.66 43.99 239.87 44.06 ;
    RECT 239.66 44.35 239.87 44.42 ;
    RECT 239.66 44.71 239.87 44.78 ;
    RECT 236.8 43.99 237.01 44.06 ;
    RECT 236.8 44.35 237.01 44.42 ;
    RECT 236.8 44.71 237.01 44.78 ;
    RECT 236.34 43.99 236.55 44.06 ;
    RECT 236.34 44.35 236.55 44.42 ;
    RECT 236.34 44.71 236.55 44.78 ;
    RECT 233.48 43.99 233.69 44.06 ;
    RECT 233.48 44.35 233.69 44.42 ;
    RECT 233.48 44.71 233.69 44.78 ;
    RECT 233.02 43.99 233.23 44.06 ;
    RECT 233.02 44.35 233.23 44.42 ;
    RECT 233.02 44.71 233.23 44.78 ;
    RECT 230.16 43.99 230.37 44.06 ;
    RECT 230.16 44.35 230.37 44.42 ;
    RECT 230.16 44.71 230.37 44.78 ;
    RECT 229.7 43.99 229.91 44.06 ;
    RECT 229.7 44.35 229.91 44.42 ;
    RECT 229.7 44.71 229.91 44.78 ;
    RECT 226.84 43.99 227.05 44.06 ;
    RECT 226.84 44.35 227.05 44.42 ;
    RECT 226.84 44.71 227.05 44.78 ;
    RECT 226.38 43.99 226.59 44.06 ;
    RECT 226.38 44.35 226.59 44.42 ;
    RECT 226.38 44.71 226.59 44.78 ;
    RECT 223.52 43.99 223.73 44.06 ;
    RECT 223.52 44.35 223.73 44.42 ;
    RECT 223.52 44.71 223.73 44.78 ;
    RECT 223.06 43.99 223.27 44.06 ;
    RECT 223.06 44.35 223.27 44.42 ;
    RECT 223.06 44.71 223.27 44.78 ;
    RECT 220.2 43.99 220.41 44.06 ;
    RECT 220.2 44.35 220.41 44.42 ;
    RECT 220.2 44.71 220.41 44.78 ;
    RECT 219.74 43.99 219.95 44.06 ;
    RECT 219.74 44.35 219.95 44.42 ;
    RECT 219.74 44.71 219.95 44.78 ;
    RECT 216.88 43.99 217.09 44.06 ;
    RECT 216.88 44.35 217.09 44.42 ;
    RECT 216.88 44.71 217.09 44.78 ;
    RECT 216.42 43.99 216.63 44.06 ;
    RECT 216.42 44.35 216.63 44.42 ;
    RECT 216.42 44.71 216.63 44.78 ;
    RECT 267.91 44.35 267.98 44.42 ;
    RECT 180.36 43.99 180.57 44.06 ;
    RECT 180.36 44.35 180.57 44.42 ;
    RECT 180.36 44.71 180.57 44.78 ;
    RECT 179.9 43.99 180.11 44.06 ;
    RECT 179.9 44.35 180.11 44.42 ;
    RECT 179.9 44.71 180.11 44.78 ;
    RECT 177.04 43.99 177.25 44.06 ;
    RECT 177.04 44.35 177.25 44.42 ;
    RECT 177.04 44.71 177.25 44.78 ;
    RECT 176.58 43.99 176.79 44.06 ;
    RECT 176.58 44.35 176.79 44.42 ;
    RECT 176.58 44.71 176.79 44.78 ;
    RECT 173.72 43.99 173.93 44.06 ;
    RECT 173.72 44.35 173.93 44.42 ;
    RECT 173.72 44.71 173.93 44.78 ;
    RECT 173.26 43.99 173.47 44.06 ;
    RECT 173.26 44.35 173.47 44.42 ;
    RECT 173.26 44.71 173.47 44.78 ;
    RECT 170.4 43.99 170.61 44.06 ;
    RECT 170.4 44.35 170.61 44.42 ;
    RECT 170.4 44.71 170.61 44.78 ;
    RECT 169.94 43.99 170.15 44.06 ;
    RECT 169.94 44.35 170.15 44.42 ;
    RECT 169.94 44.71 170.15 44.78 ;
    RECT 167.08 43.99 167.29 44.06 ;
    RECT 167.08 44.35 167.29 44.42 ;
    RECT 167.08 44.71 167.29 44.78 ;
    RECT 166.62 43.99 166.83 44.06 ;
    RECT 166.62 44.35 166.83 44.42 ;
    RECT 166.62 44.71 166.83 44.78 ;
    RECT 163.76 43.99 163.97 44.06 ;
    RECT 163.76 44.35 163.97 44.42 ;
    RECT 163.76 44.71 163.97 44.78 ;
    RECT 163.3 43.99 163.51 44.06 ;
    RECT 163.3 44.35 163.51 44.42 ;
    RECT 163.3 44.71 163.51 44.78 ;
    RECT 160.44 43.99 160.65 44.06 ;
    RECT 160.44 44.35 160.65 44.42 ;
    RECT 160.44 44.71 160.65 44.78 ;
    RECT 159.98 43.99 160.19 44.06 ;
    RECT 159.98 44.35 160.19 44.42 ;
    RECT 159.98 44.71 160.19 44.78 ;
    RECT 157.12 43.99 157.33 44.06 ;
    RECT 157.12 44.35 157.33 44.42 ;
    RECT 157.12 44.71 157.33 44.78 ;
    RECT 156.66 43.99 156.87 44.06 ;
    RECT 156.66 44.35 156.87 44.42 ;
    RECT 156.66 44.71 156.87 44.78 ;
    RECT 153.8 43.99 154.01 44.06 ;
    RECT 153.8 44.35 154.01 44.42 ;
    RECT 153.8 44.71 154.01 44.78 ;
    RECT 153.34 43.99 153.55 44.06 ;
    RECT 153.34 44.35 153.55 44.42 ;
    RECT 153.34 44.71 153.55 44.78 ;
    RECT 150.48 43.99 150.69 44.06 ;
    RECT 150.48 44.35 150.69 44.42 ;
    RECT 150.48 44.71 150.69 44.78 ;
    RECT 150.02 43.99 150.23 44.06 ;
    RECT 150.02 44.35 150.23 44.42 ;
    RECT 150.02 44.71 150.23 44.78 ;
    RECT 213.56 43.99 213.77 44.06 ;
    RECT 213.56 44.35 213.77 44.42 ;
    RECT 213.56 44.71 213.77 44.78 ;
    RECT 213.1 43.99 213.31 44.06 ;
    RECT 213.1 44.35 213.31 44.42 ;
    RECT 213.1 44.71 213.31 44.78 ;
    RECT 210.24 43.99 210.45 44.06 ;
    RECT 210.24 44.35 210.45 44.42 ;
    RECT 210.24 44.71 210.45 44.78 ;
    RECT 209.78 43.99 209.99 44.06 ;
    RECT 209.78 44.35 209.99 44.42 ;
    RECT 209.78 44.71 209.99 44.78 ;
    RECT 206.92 43.99 207.13 44.06 ;
    RECT 206.92 44.35 207.13 44.42 ;
    RECT 206.92 44.71 207.13 44.78 ;
    RECT 206.46 43.99 206.67 44.06 ;
    RECT 206.46 44.35 206.67 44.42 ;
    RECT 206.46 44.71 206.67 44.78 ;
    RECT 203.6 43.99 203.81 44.06 ;
    RECT 203.6 44.35 203.81 44.42 ;
    RECT 203.6 44.71 203.81 44.78 ;
    RECT 203.14 43.99 203.35 44.06 ;
    RECT 203.14 44.35 203.35 44.42 ;
    RECT 203.14 44.71 203.35 44.78 ;
    RECT 200.28 43.99 200.49 44.06 ;
    RECT 200.28 44.35 200.49 44.42 ;
    RECT 200.28 44.71 200.49 44.78 ;
    RECT 199.82 43.99 200.03 44.06 ;
    RECT 199.82 44.35 200.03 44.42 ;
    RECT 199.82 44.71 200.03 44.78 ;
    RECT 196.96 43.99 197.17 44.06 ;
    RECT 196.96 44.35 197.17 44.42 ;
    RECT 196.96 44.71 197.17 44.78 ;
    RECT 196.5 43.99 196.71 44.06 ;
    RECT 196.5 44.35 196.71 44.42 ;
    RECT 196.5 44.71 196.71 44.78 ;
    RECT 193.64 43.99 193.85 44.06 ;
    RECT 193.64 44.35 193.85 44.42 ;
    RECT 193.64 44.71 193.85 44.78 ;
    RECT 193.18 43.99 193.39 44.06 ;
    RECT 193.18 44.35 193.39 44.42 ;
    RECT 193.18 44.71 193.39 44.78 ;
    RECT 190.32 43.99 190.53 44.06 ;
    RECT 190.32 44.35 190.53 44.42 ;
    RECT 190.32 44.71 190.53 44.78 ;
    RECT 189.86 43.99 190.07 44.06 ;
    RECT 189.86 44.35 190.07 44.42 ;
    RECT 189.86 44.71 190.07 44.78 ;
    RECT 187.0 43.99 187.21 44.06 ;
    RECT 187.0 44.35 187.21 44.42 ;
    RECT 187.0 44.71 187.21 44.78 ;
    RECT 186.54 43.99 186.75 44.06 ;
    RECT 186.54 44.35 186.75 44.42 ;
    RECT 186.54 44.71 186.75 44.78 ;
    RECT 183.68 43.99 183.89 44.06 ;
    RECT 183.68 44.35 183.89 44.42 ;
    RECT 183.68 44.71 183.89 44.78 ;
    RECT 183.22 43.99 183.43 44.06 ;
    RECT 183.22 44.35 183.43 44.42 ;
    RECT 183.22 44.71 183.43 44.78 ;
    RECT 147.485 44.35 147.555 44.42 ;
    RECT 266.68 43.99 266.89 44.06 ;
    RECT 266.68 44.35 266.89 44.42 ;
    RECT 266.68 44.71 266.89 44.78 ;
    RECT 266.22 43.99 266.43 44.06 ;
    RECT 266.22 44.35 266.43 44.42 ;
    RECT 266.22 44.71 266.43 44.78 ;
    RECT 263.36 43.99 263.57 44.06 ;
    RECT 263.36 44.35 263.57 44.42 ;
    RECT 263.36 44.71 263.57 44.78 ;
    RECT 262.9 43.99 263.11 44.06 ;
    RECT 262.9 44.35 263.11 44.42 ;
    RECT 262.9 44.71 263.11 44.78 ;
    RECT 260.04 43.99 260.25 44.06 ;
    RECT 260.04 44.35 260.25 44.42 ;
    RECT 260.04 44.71 260.25 44.78 ;
    RECT 259.58 43.99 259.79 44.06 ;
    RECT 259.58 44.35 259.79 44.42 ;
    RECT 259.58 44.71 259.79 44.78 ;
    RECT 256.72 43.99 256.93 44.06 ;
    RECT 256.72 44.35 256.93 44.42 ;
    RECT 256.72 44.71 256.93 44.78 ;
    RECT 256.26 43.99 256.47 44.06 ;
    RECT 256.26 44.35 256.47 44.42 ;
    RECT 256.26 44.71 256.47 44.78 ;
    RECT 253.4 43.99 253.61 44.06 ;
    RECT 253.4 44.35 253.61 44.42 ;
    RECT 253.4 44.71 253.61 44.78 ;
    RECT 252.94 43.99 253.15 44.06 ;
    RECT 252.94 44.35 253.15 44.42 ;
    RECT 252.94 44.71 253.15 44.78 ;
    RECT 250.08 83.61 250.29 83.68 ;
    RECT 250.08 83.97 250.29 84.04 ;
    RECT 250.08 84.33 250.29 84.4 ;
    RECT 249.62 83.61 249.83 83.68 ;
    RECT 249.62 83.97 249.83 84.04 ;
    RECT 249.62 84.33 249.83 84.4 ;
    RECT 246.76 83.61 246.97 83.68 ;
    RECT 246.76 83.97 246.97 84.04 ;
    RECT 246.76 84.33 246.97 84.4 ;
    RECT 246.3 83.61 246.51 83.68 ;
    RECT 246.3 83.97 246.51 84.04 ;
    RECT 246.3 84.33 246.51 84.4 ;
    RECT 243.44 83.61 243.65 83.68 ;
    RECT 243.44 83.97 243.65 84.04 ;
    RECT 243.44 84.33 243.65 84.4 ;
    RECT 242.98 83.61 243.19 83.68 ;
    RECT 242.98 83.97 243.19 84.04 ;
    RECT 242.98 84.33 243.19 84.4 ;
    RECT 240.12 83.61 240.33 83.68 ;
    RECT 240.12 83.97 240.33 84.04 ;
    RECT 240.12 84.33 240.33 84.4 ;
    RECT 239.66 83.61 239.87 83.68 ;
    RECT 239.66 83.97 239.87 84.04 ;
    RECT 239.66 84.33 239.87 84.4 ;
    RECT 236.8 83.61 237.01 83.68 ;
    RECT 236.8 83.97 237.01 84.04 ;
    RECT 236.8 84.33 237.01 84.4 ;
    RECT 236.34 83.61 236.55 83.68 ;
    RECT 236.34 83.97 236.55 84.04 ;
    RECT 236.34 84.33 236.55 84.4 ;
    RECT 233.48 83.61 233.69 83.68 ;
    RECT 233.48 83.97 233.69 84.04 ;
    RECT 233.48 84.33 233.69 84.4 ;
    RECT 233.02 83.61 233.23 83.68 ;
    RECT 233.02 83.97 233.23 84.04 ;
    RECT 233.02 84.33 233.23 84.4 ;
    RECT 230.16 83.61 230.37 83.68 ;
    RECT 230.16 83.97 230.37 84.04 ;
    RECT 230.16 84.33 230.37 84.4 ;
    RECT 229.7 83.61 229.91 83.68 ;
    RECT 229.7 83.97 229.91 84.04 ;
    RECT 229.7 84.33 229.91 84.4 ;
    RECT 226.84 83.61 227.05 83.68 ;
    RECT 226.84 83.97 227.05 84.04 ;
    RECT 226.84 84.33 227.05 84.4 ;
    RECT 226.38 83.61 226.59 83.68 ;
    RECT 226.38 83.97 226.59 84.04 ;
    RECT 226.38 84.33 226.59 84.4 ;
    RECT 223.52 83.61 223.73 83.68 ;
    RECT 223.52 83.97 223.73 84.04 ;
    RECT 223.52 84.33 223.73 84.4 ;
    RECT 223.06 83.61 223.27 83.68 ;
    RECT 223.06 83.97 223.27 84.04 ;
    RECT 223.06 84.33 223.27 84.4 ;
    RECT 220.2 83.61 220.41 83.68 ;
    RECT 220.2 83.97 220.41 84.04 ;
    RECT 220.2 84.33 220.41 84.4 ;
    RECT 219.74 83.61 219.95 83.68 ;
    RECT 219.74 83.97 219.95 84.04 ;
    RECT 219.74 84.33 219.95 84.4 ;
    RECT 216.88 83.61 217.09 83.68 ;
    RECT 216.88 83.97 217.09 84.04 ;
    RECT 216.88 84.33 217.09 84.4 ;
    RECT 216.42 83.61 216.63 83.68 ;
    RECT 216.42 83.97 216.63 84.04 ;
    RECT 216.42 84.33 216.63 84.4 ;
    RECT 267.91 83.97 267.98 84.04 ;
    RECT 180.36 83.61 180.57 83.68 ;
    RECT 180.36 83.97 180.57 84.04 ;
    RECT 180.36 84.33 180.57 84.4 ;
    RECT 179.9 83.61 180.11 83.68 ;
    RECT 179.9 83.97 180.11 84.04 ;
    RECT 179.9 84.33 180.11 84.4 ;
    RECT 177.04 83.61 177.25 83.68 ;
    RECT 177.04 83.97 177.25 84.04 ;
    RECT 177.04 84.33 177.25 84.4 ;
    RECT 176.58 83.61 176.79 83.68 ;
    RECT 176.58 83.97 176.79 84.04 ;
    RECT 176.58 84.33 176.79 84.4 ;
    RECT 173.72 83.61 173.93 83.68 ;
    RECT 173.72 83.97 173.93 84.04 ;
    RECT 173.72 84.33 173.93 84.4 ;
    RECT 173.26 83.61 173.47 83.68 ;
    RECT 173.26 83.97 173.47 84.04 ;
    RECT 173.26 84.33 173.47 84.4 ;
    RECT 170.4 83.61 170.61 83.68 ;
    RECT 170.4 83.97 170.61 84.04 ;
    RECT 170.4 84.33 170.61 84.4 ;
    RECT 169.94 83.61 170.15 83.68 ;
    RECT 169.94 83.97 170.15 84.04 ;
    RECT 169.94 84.33 170.15 84.4 ;
    RECT 167.08 83.61 167.29 83.68 ;
    RECT 167.08 83.97 167.29 84.04 ;
    RECT 167.08 84.33 167.29 84.4 ;
    RECT 166.62 83.61 166.83 83.68 ;
    RECT 166.62 83.97 166.83 84.04 ;
    RECT 166.62 84.33 166.83 84.4 ;
    RECT 163.76 83.61 163.97 83.68 ;
    RECT 163.76 83.97 163.97 84.04 ;
    RECT 163.76 84.33 163.97 84.4 ;
    RECT 163.3 83.61 163.51 83.68 ;
    RECT 163.3 83.97 163.51 84.04 ;
    RECT 163.3 84.33 163.51 84.4 ;
    RECT 160.44 83.61 160.65 83.68 ;
    RECT 160.44 83.97 160.65 84.04 ;
    RECT 160.44 84.33 160.65 84.4 ;
    RECT 159.98 83.61 160.19 83.68 ;
    RECT 159.98 83.97 160.19 84.04 ;
    RECT 159.98 84.33 160.19 84.4 ;
    RECT 157.12 83.61 157.33 83.68 ;
    RECT 157.12 83.97 157.33 84.04 ;
    RECT 157.12 84.33 157.33 84.4 ;
    RECT 156.66 83.61 156.87 83.68 ;
    RECT 156.66 83.97 156.87 84.04 ;
    RECT 156.66 84.33 156.87 84.4 ;
    RECT 153.8 83.61 154.01 83.68 ;
    RECT 153.8 83.97 154.01 84.04 ;
    RECT 153.8 84.33 154.01 84.4 ;
    RECT 153.34 83.61 153.55 83.68 ;
    RECT 153.34 83.97 153.55 84.04 ;
    RECT 153.34 84.33 153.55 84.4 ;
    RECT 150.48 83.61 150.69 83.68 ;
    RECT 150.48 83.97 150.69 84.04 ;
    RECT 150.48 84.33 150.69 84.4 ;
    RECT 150.02 83.61 150.23 83.68 ;
    RECT 150.02 83.97 150.23 84.04 ;
    RECT 150.02 84.33 150.23 84.4 ;
    RECT 213.56 83.61 213.77 83.68 ;
    RECT 213.56 83.97 213.77 84.04 ;
    RECT 213.56 84.33 213.77 84.4 ;
    RECT 213.1 83.61 213.31 83.68 ;
    RECT 213.1 83.97 213.31 84.04 ;
    RECT 213.1 84.33 213.31 84.4 ;
    RECT 210.24 83.61 210.45 83.68 ;
    RECT 210.24 83.97 210.45 84.04 ;
    RECT 210.24 84.33 210.45 84.4 ;
    RECT 209.78 83.61 209.99 83.68 ;
    RECT 209.78 83.97 209.99 84.04 ;
    RECT 209.78 84.33 209.99 84.4 ;
    RECT 206.92 83.61 207.13 83.68 ;
    RECT 206.92 83.97 207.13 84.04 ;
    RECT 206.92 84.33 207.13 84.4 ;
    RECT 206.46 83.61 206.67 83.68 ;
    RECT 206.46 83.97 206.67 84.04 ;
    RECT 206.46 84.33 206.67 84.4 ;
    RECT 203.6 83.61 203.81 83.68 ;
    RECT 203.6 83.97 203.81 84.04 ;
    RECT 203.6 84.33 203.81 84.4 ;
    RECT 203.14 83.61 203.35 83.68 ;
    RECT 203.14 83.97 203.35 84.04 ;
    RECT 203.14 84.33 203.35 84.4 ;
    RECT 200.28 83.61 200.49 83.68 ;
    RECT 200.28 83.97 200.49 84.04 ;
    RECT 200.28 84.33 200.49 84.4 ;
    RECT 199.82 83.61 200.03 83.68 ;
    RECT 199.82 83.97 200.03 84.04 ;
    RECT 199.82 84.33 200.03 84.4 ;
    RECT 196.96 83.61 197.17 83.68 ;
    RECT 196.96 83.97 197.17 84.04 ;
    RECT 196.96 84.33 197.17 84.4 ;
    RECT 196.5 83.61 196.71 83.68 ;
    RECT 196.5 83.97 196.71 84.04 ;
    RECT 196.5 84.33 196.71 84.4 ;
    RECT 193.64 83.61 193.85 83.68 ;
    RECT 193.64 83.97 193.85 84.04 ;
    RECT 193.64 84.33 193.85 84.4 ;
    RECT 193.18 83.61 193.39 83.68 ;
    RECT 193.18 83.97 193.39 84.04 ;
    RECT 193.18 84.33 193.39 84.4 ;
    RECT 190.32 83.61 190.53 83.68 ;
    RECT 190.32 83.97 190.53 84.04 ;
    RECT 190.32 84.33 190.53 84.4 ;
    RECT 189.86 83.61 190.07 83.68 ;
    RECT 189.86 83.97 190.07 84.04 ;
    RECT 189.86 84.33 190.07 84.4 ;
    RECT 187.0 83.61 187.21 83.68 ;
    RECT 187.0 83.97 187.21 84.04 ;
    RECT 187.0 84.33 187.21 84.4 ;
    RECT 186.54 83.61 186.75 83.68 ;
    RECT 186.54 83.97 186.75 84.04 ;
    RECT 186.54 84.33 186.75 84.4 ;
    RECT 183.68 83.61 183.89 83.68 ;
    RECT 183.68 83.97 183.89 84.04 ;
    RECT 183.68 84.33 183.89 84.4 ;
    RECT 183.22 83.61 183.43 83.68 ;
    RECT 183.22 83.97 183.43 84.04 ;
    RECT 183.22 84.33 183.43 84.4 ;
    RECT 147.485 83.97 147.555 84.04 ;
    RECT 266.68 83.61 266.89 83.68 ;
    RECT 266.68 83.97 266.89 84.04 ;
    RECT 266.68 84.33 266.89 84.4 ;
    RECT 266.22 83.61 266.43 83.68 ;
    RECT 266.22 83.97 266.43 84.04 ;
    RECT 266.22 84.33 266.43 84.4 ;
    RECT 263.36 83.61 263.57 83.68 ;
    RECT 263.36 83.97 263.57 84.04 ;
    RECT 263.36 84.33 263.57 84.4 ;
    RECT 262.9 83.61 263.11 83.68 ;
    RECT 262.9 83.97 263.11 84.04 ;
    RECT 262.9 84.33 263.11 84.4 ;
    RECT 260.04 83.61 260.25 83.68 ;
    RECT 260.04 83.97 260.25 84.04 ;
    RECT 260.04 84.33 260.25 84.4 ;
    RECT 259.58 83.61 259.79 83.68 ;
    RECT 259.58 83.97 259.79 84.04 ;
    RECT 259.58 84.33 259.79 84.4 ;
    RECT 256.72 83.61 256.93 83.68 ;
    RECT 256.72 83.97 256.93 84.04 ;
    RECT 256.72 84.33 256.93 84.4 ;
    RECT 256.26 83.61 256.47 83.68 ;
    RECT 256.26 83.97 256.47 84.04 ;
    RECT 256.26 84.33 256.47 84.4 ;
    RECT 253.4 83.61 253.61 83.68 ;
    RECT 253.4 83.97 253.61 84.04 ;
    RECT 253.4 84.33 253.61 84.4 ;
    RECT 252.94 83.61 253.15 83.68 ;
    RECT 252.94 83.97 253.15 84.04 ;
    RECT 252.94 84.33 253.15 84.4 ;
    RECT 250.08 43.27 250.29 43.34 ;
    RECT 250.08 43.63 250.29 43.7 ;
    RECT 250.08 43.99 250.29 44.06 ;
    RECT 249.62 43.27 249.83 43.34 ;
    RECT 249.62 43.63 249.83 43.7 ;
    RECT 249.62 43.99 249.83 44.06 ;
    RECT 246.76 43.27 246.97 43.34 ;
    RECT 246.76 43.63 246.97 43.7 ;
    RECT 246.76 43.99 246.97 44.06 ;
    RECT 246.3 43.27 246.51 43.34 ;
    RECT 246.3 43.63 246.51 43.7 ;
    RECT 246.3 43.99 246.51 44.06 ;
    RECT 243.44 43.27 243.65 43.34 ;
    RECT 243.44 43.63 243.65 43.7 ;
    RECT 243.44 43.99 243.65 44.06 ;
    RECT 242.98 43.27 243.19 43.34 ;
    RECT 242.98 43.63 243.19 43.7 ;
    RECT 242.98 43.99 243.19 44.06 ;
    RECT 240.12 43.27 240.33 43.34 ;
    RECT 240.12 43.63 240.33 43.7 ;
    RECT 240.12 43.99 240.33 44.06 ;
    RECT 239.66 43.27 239.87 43.34 ;
    RECT 239.66 43.63 239.87 43.7 ;
    RECT 239.66 43.99 239.87 44.06 ;
    RECT 236.8 43.27 237.01 43.34 ;
    RECT 236.8 43.63 237.01 43.7 ;
    RECT 236.8 43.99 237.01 44.06 ;
    RECT 236.34 43.27 236.55 43.34 ;
    RECT 236.34 43.63 236.55 43.7 ;
    RECT 236.34 43.99 236.55 44.06 ;
    RECT 233.48 43.27 233.69 43.34 ;
    RECT 233.48 43.63 233.69 43.7 ;
    RECT 233.48 43.99 233.69 44.06 ;
    RECT 233.02 43.27 233.23 43.34 ;
    RECT 233.02 43.63 233.23 43.7 ;
    RECT 233.02 43.99 233.23 44.06 ;
    RECT 230.16 43.27 230.37 43.34 ;
    RECT 230.16 43.63 230.37 43.7 ;
    RECT 230.16 43.99 230.37 44.06 ;
    RECT 229.7 43.27 229.91 43.34 ;
    RECT 229.7 43.63 229.91 43.7 ;
    RECT 229.7 43.99 229.91 44.06 ;
    RECT 226.84 43.27 227.05 43.34 ;
    RECT 226.84 43.63 227.05 43.7 ;
    RECT 226.84 43.99 227.05 44.06 ;
    RECT 226.38 43.27 226.59 43.34 ;
    RECT 226.38 43.63 226.59 43.7 ;
    RECT 226.38 43.99 226.59 44.06 ;
    RECT 223.52 43.27 223.73 43.34 ;
    RECT 223.52 43.63 223.73 43.7 ;
    RECT 223.52 43.99 223.73 44.06 ;
    RECT 223.06 43.27 223.27 43.34 ;
    RECT 223.06 43.63 223.27 43.7 ;
    RECT 223.06 43.99 223.27 44.06 ;
    RECT 220.2 43.27 220.41 43.34 ;
    RECT 220.2 43.63 220.41 43.7 ;
    RECT 220.2 43.99 220.41 44.06 ;
    RECT 219.74 43.27 219.95 43.34 ;
    RECT 219.74 43.63 219.95 43.7 ;
    RECT 219.74 43.99 219.95 44.06 ;
    RECT 216.88 43.27 217.09 43.34 ;
    RECT 216.88 43.63 217.09 43.7 ;
    RECT 216.88 43.99 217.09 44.06 ;
    RECT 216.42 43.27 216.63 43.34 ;
    RECT 216.42 43.63 216.63 43.7 ;
    RECT 216.42 43.99 216.63 44.06 ;
    RECT 267.91 43.63 267.98 43.7 ;
    RECT 180.36 43.27 180.57 43.34 ;
    RECT 180.36 43.63 180.57 43.7 ;
    RECT 180.36 43.99 180.57 44.06 ;
    RECT 179.9 43.27 180.11 43.34 ;
    RECT 179.9 43.63 180.11 43.7 ;
    RECT 179.9 43.99 180.11 44.06 ;
    RECT 177.04 43.27 177.25 43.34 ;
    RECT 177.04 43.63 177.25 43.7 ;
    RECT 177.04 43.99 177.25 44.06 ;
    RECT 176.58 43.27 176.79 43.34 ;
    RECT 176.58 43.63 176.79 43.7 ;
    RECT 176.58 43.99 176.79 44.06 ;
    RECT 173.72 43.27 173.93 43.34 ;
    RECT 173.72 43.63 173.93 43.7 ;
    RECT 173.72 43.99 173.93 44.06 ;
    RECT 173.26 43.27 173.47 43.34 ;
    RECT 173.26 43.63 173.47 43.7 ;
    RECT 173.26 43.99 173.47 44.06 ;
    RECT 170.4 43.27 170.61 43.34 ;
    RECT 170.4 43.63 170.61 43.7 ;
    RECT 170.4 43.99 170.61 44.06 ;
    RECT 169.94 43.27 170.15 43.34 ;
    RECT 169.94 43.63 170.15 43.7 ;
    RECT 169.94 43.99 170.15 44.06 ;
    RECT 167.08 43.27 167.29 43.34 ;
    RECT 167.08 43.63 167.29 43.7 ;
    RECT 167.08 43.99 167.29 44.06 ;
    RECT 166.62 43.27 166.83 43.34 ;
    RECT 166.62 43.63 166.83 43.7 ;
    RECT 166.62 43.99 166.83 44.06 ;
    RECT 163.76 43.27 163.97 43.34 ;
    RECT 163.76 43.63 163.97 43.7 ;
    RECT 163.76 43.99 163.97 44.06 ;
    RECT 163.3 43.27 163.51 43.34 ;
    RECT 163.3 43.63 163.51 43.7 ;
    RECT 163.3 43.99 163.51 44.06 ;
    RECT 160.44 43.27 160.65 43.34 ;
    RECT 160.44 43.63 160.65 43.7 ;
    RECT 160.44 43.99 160.65 44.06 ;
    RECT 159.98 43.27 160.19 43.34 ;
    RECT 159.98 43.63 160.19 43.7 ;
    RECT 159.98 43.99 160.19 44.06 ;
    RECT 157.12 43.27 157.33 43.34 ;
    RECT 157.12 43.63 157.33 43.7 ;
    RECT 157.12 43.99 157.33 44.06 ;
    RECT 156.66 43.27 156.87 43.34 ;
    RECT 156.66 43.63 156.87 43.7 ;
    RECT 156.66 43.99 156.87 44.06 ;
    RECT 153.8 43.27 154.01 43.34 ;
    RECT 153.8 43.63 154.01 43.7 ;
    RECT 153.8 43.99 154.01 44.06 ;
    RECT 153.34 43.27 153.55 43.34 ;
    RECT 153.34 43.63 153.55 43.7 ;
    RECT 153.34 43.99 153.55 44.06 ;
    RECT 150.48 43.27 150.69 43.34 ;
    RECT 150.48 43.63 150.69 43.7 ;
    RECT 150.48 43.99 150.69 44.06 ;
    RECT 150.02 43.27 150.23 43.34 ;
    RECT 150.02 43.63 150.23 43.7 ;
    RECT 150.02 43.99 150.23 44.06 ;
    RECT 213.56 43.27 213.77 43.34 ;
    RECT 213.56 43.63 213.77 43.7 ;
    RECT 213.56 43.99 213.77 44.06 ;
    RECT 213.1 43.27 213.31 43.34 ;
    RECT 213.1 43.63 213.31 43.7 ;
    RECT 213.1 43.99 213.31 44.06 ;
    RECT 210.24 43.27 210.45 43.34 ;
    RECT 210.24 43.63 210.45 43.7 ;
    RECT 210.24 43.99 210.45 44.06 ;
    RECT 209.78 43.27 209.99 43.34 ;
    RECT 209.78 43.63 209.99 43.7 ;
    RECT 209.78 43.99 209.99 44.06 ;
    RECT 206.92 43.27 207.13 43.34 ;
    RECT 206.92 43.63 207.13 43.7 ;
    RECT 206.92 43.99 207.13 44.06 ;
    RECT 206.46 43.27 206.67 43.34 ;
    RECT 206.46 43.63 206.67 43.7 ;
    RECT 206.46 43.99 206.67 44.06 ;
    RECT 203.6 43.27 203.81 43.34 ;
    RECT 203.6 43.63 203.81 43.7 ;
    RECT 203.6 43.99 203.81 44.06 ;
    RECT 203.14 43.27 203.35 43.34 ;
    RECT 203.14 43.63 203.35 43.7 ;
    RECT 203.14 43.99 203.35 44.06 ;
    RECT 200.28 43.27 200.49 43.34 ;
    RECT 200.28 43.63 200.49 43.7 ;
    RECT 200.28 43.99 200.49 44.06 ;
    RECT 199.82 43.27 200.03 43.34 ;
    RECT 199.82 43.63 200.03 43.7 ;
    RECT 199.82 43.99 200.03 44.06 ;
    RECT 196.96 43.27 197.17 43.34 ;
    RECT 196.96 43.63 197.17 43.7 ;
    RECT 196.96 43.99 197.17 44.06 ;
    RECT 196.5 43.27 196.71 43.34 ;
    RECT 196.5 43.63 196.71 43.7 ;
    RECT 196.5 43.99 196.71 44.06 ;
    RECT 193.64 43.27 193.85 43.34 ;
    RECT 193.64 43.63 193.85 43.7 ;
    RECT 193.64 43.99 193.85 44.06 ;
    RECT 193.18 43.27 193.39 43.34 ;
    RECT 193.18 43.63 193.39 43.7 ;
    RECT 193.18 43.99 193.39 44.06 ;
    RECT 190.32 43.27 190.53 43.34 ;
    RECT 190.32 43.63 190.53 43.7 ;
    RECT 190.32 43.99 190.53 44.06 ;
    RECT 189.86 43.27 190.07 43.34 ;
    RECT 189.86 43.63 190.07 43.7 ;
    RECT 189.86 43.99 190.07 44.06 ;
    RECT 187.0 43.27 187.21 43.34 ;
    RECT 187.0 43.63 187.21 43.7 ;
    RECT 187.0 43.99 187.21 44.06 ;
    RECT 186.54 43.27 186.75 43.34 ;
    RECT 186.54 43.63 186.75 43.7 ;
    RECT 186.54 43.99 186.75 44.06 ;
    RECT 183.68 43.27 183.89 43.34 ;
    RECT 183.68 43.63 183.89 43.7 ;
    RECT 183.68 43.99 183.89 44.06 ;
    RECT 183.22 43.27 183.43 43.34 ;
    RECT 183.22 43.63 183.43 43.7 ;
    RECT 183.22 43.99 183.43 44.06 ;
    RECT 147.485 43.63 147.555 43.7 ;
    RECT 266.68 43.27 266.89 43.34 ;
    RECT 266.68 43.63 266.89 43.7 ;
    RECT 266.68 43.99 266.89 44.06 ;
    RECT 266.22 43.27 266.43 43.34 ;
    RECT 266.22 43.63 266.43 43.7 ;
    RECT 266.22 43.99 266.43 44.06 ;
    RECT 263.36 43.27 263.57 43.34 ;
    RECT 263.36 43.63 263.57 43.7 ;
    RECT 263.36 43.99 263.57 44.06 ;
    RECT 262.9 43.27 263.11 43.34 ;
    RECT 262.9 43.63 263.11 43.7 ;
    RECT 262.9 43.99 263.11 44.06 ;
    RECT 260.04 43.27 260.25 43.34 ;
    RECT 260.04 43.63 260.25 43.7 ;
    RECT 260.04 43.99 260.25 44.06 ;
    RECT 259.58 43.27 259.79 43.34 ;
    RECT 259.58 43.63 259.79 43.7 ;
    RECT 259.58 43.99 259.79 44.06 ;
    RECT 256.72 43.27 256.93 43.34 ;
    RECT 256.72 43.63 256.93 43.7 ;
    RECT 256.72 43.99 256.93 44.06 ;
    RECT 256.26 43.27 256.47 43.34 ;
    RECT 256.26 43.63 256.47 43.7 ;
    RECT 256.26 43.99 256.47 44.06 ;
    RECT 253.4 43.27 253.61 43.34 ;
    RECT 253.4 43.63 253.61 43.7 ;
    RECT 253.4 43.99 253.61 44.06 ;
    RECT 252.94 43.27 253.15 43.34 ;
    RECT 252.94 43.63 253.15 43.7 ;
    RECT 252.94 43.99 253.15 44.06 ;
    RECT 250.08 82.89 250.29 82.96 ;
    RECT 250.08 83.25 250.29 83.32 ;
    RECT 250.08 83.61 250.29 83.68 ;
    RECT 249.62 82.89 249.83 82.96 ;
    RECT 249.62 83.25 249.83 83.32 ;
    RECT 249.62 83.61 249.83 83.68 ;
    RECT 246.76 82.89 246.97 82.96 ;
    RECT 246.76 83.25 246.97 83.32 ;
    RECT 246.76 83.61 246.97 83.68 ;
    RECT 246.3 82.89 246.51 82.96 ;
    RECT 246.3 83.25 246.51 83.32 ;
    RECT 246.3 83.61 246.51 83.68 ;
    RECT 243.44 82.89 243.65 82.96 ;
    RECT 243.44 83.25 243.65 83.32 ;
    RECT 243.44 83.61 243.65 83.68 ;
    RECT 242.98 82.89 243.19 82.96 ;
    RECT 242.98 83.25 243.19 83.32 ;
    RECT 242.98 83.61 243.19 83.68 ;
    RECT 240.12 82.89 240.33 82.96 ;
    RECT 240.12 83.25 240.33 83.32 ;
    RECT 240.12 83.61 240.33 83.68 ;
    RECT 239.66 82.89 239.87 82.96 ;
    RECT 239.66 83.25 239.87 83.32 ;
    RECT 239.66 83.61 239.87 83.68 ;
    RECT 236.8 82.89 237.01 82.96 ;
    RECT 236.8 83.25 237.01 83.32 ;
    RECT 236.8 83.61 237.01 83.68 ;
    RECT 236.34 82.89 236.55 82.96 ;
    RECT 236.34 83.25 236.55 83.32 ;
    RECT 236.34 83.61 236.55 83.68 ;
    RECT 233.48 82.89 233.69 82.96 ;
    RECT 233.48 83.25 233.69 83.32 ;
    RECT 233.48 83.61 233.69 83.68 ;
    RECT 233.02 82.89 233.23 82.96 ;
    RECT 233.02 83.25 233.23 83.32 ;
    RECT 233.02 83.61 233.23 83.68 ;
    RECT 230.16 82.89 230.37 82.96 ;
    RECT 230.16 83.25 230.37 83.32 ;
    RECT 230.16 83.61 230.37 83.68 ;
    RECT 229.7 82.89 229.91 82.96 ;
    RECT 229.7 83.25 229.91 83.32 ;
    RECT 229.7 83.61 229.91 83.68 ;
    RECT 226.84 82.89 227.05 82.96 ;
    RECT 226.84 83.25 227.05 83.32 ;
    RECT 226.84 83.61 227.05 83.68 ;
    RECT 226.38 82.89 226.59 82.96 ;
    RECT 226.38 83.25 226.59 83.32 ;
    RECT 226.38 83.61 226.59 83.68 ;
    RECT 223.52 82.89 223.73 82.96 ;
    RECT 223.52 83.25 223.73 83.32 ;
    RECT 223.52 83.61 223.73 83.68 ;
    RECT 223.06 82.89 223.27 82.96 ;
    RECT 223.06 83.25 223.27 83.32 ;
    RECT 223.06 83.61 223.27 83.68 ;
    RECT 220.2 82.89 220.41 82.96 ;
    RECT 220.2 83.25 220.41 83.32 ;
    RECT 220.2 83.61 220.41 83.68 ;
    RECT 219.74 82.89 219.95 82.96 ;
    RECT 219.74 83.25 219.95 83.32 ;
    RECT 219.74 83.61 219.95 83.68 ;
    RECT 216.88 82.89 217.09 82.96 ;
    RECT 216.88 83.25 217.09 83.32 ;
    RECT 216.88 83.61 217.09 83.68 ;
    RECT 216.42 82.89 216.63 82.96 ;
    RECT 216.42 83.25 216.63 83.32 ;
    RECT 216.42 83.61 216.63 83.68 ;
    RECT 267.91 83.25 267.98 83.32 ;
    RECT 180.36 82.89 180.57 82.96 ;
    RECT 180.36 83.25 180.57 83.32 ;
    RECT 180.36 83.61 180.57 83.68 ;
    RECT 179.9 82.89 180.11 82.96 ;
    RECT 179.9 83.25 180.11 83.32 ;
    RECT 179.9 83.61 180.11 83.68 ;
    RECT 177.04 82.89 177.25 82.96 ;
    RECT 177.04 83.25 177.25 83.32 ;
    RECT 177.04 83.61 177.25 83.68 ;
    RECT 176.58 82.89 176.79 82.96 ;
    RECT 176.58 83.25 176.79 83.32 ;
    RECT 176.58 83.61 176.79 83.68 ;
    RECT 173.72 82.89 173.93 82.96 ;
    RECT 173.72 83.25 173.93 83.32 ;
    RECT 173.72 83.61 173.93 83.68 ;
    RECT 173.26 82.89 173.47 82.96 ;
    RECT 173.26 83.25 173.47 83.32 ;
    RECT 173.26 83.61 173.47 83.68 ;
    RECT 170.4 82.89 170.61 82.96 ;
    RECT 170.4 83.25 170.61 83.32 ;
    RECT 170.4 83.61 170.61 83.68 ;
    RECT 169.94 82.89 170.15 82.96 ;
    RECT 169.94 83.25 170.15 83.32 ;
    RECT 169.94 83.61 170.15 83.68 ;
    RECT 167.08 82.89 167.29 82.96 ;
    RECT 167.08 83.25 167.29 83.32 ;
    RECT 167.08 83.61 167.29 83.68 ;
    RECT 166.62 82.89 166.83 82.96 ;
    RECT 166.62 83.25 166.83 83.32 ;
    RECT 166.62 83.61 166.83 83.68 ;
    RECT 163.76 82.89 163.97 82.96 ;
    RECT 163.76 83.25 163.97 83.32 ;
    RECT 163.76 83.61 163.97 83.68 ;
    RECT 163.3 82.89 163.51 82.96 ;
    RECT 163.3 83.25 163.51 83.32 ;
    RECT 163.3 83.61 163.51 83.68 ;
    RECT 160.44 82.89 160.65 82.96 ;
    RECT 160.44 83.25 160.65 83.32 ;
    RECT 160.44 83.61 160.65 83.68 ;
    RECT 159.98 82.89 160.19 82.96 ;
    RECT 159.98 83.25 160.19 83.32 ;
    RECT 159.98 83.61 160.19 83.68 ;
    RECT 157.12 82.89 157.33 82.96 ;
    RECT 157.12 83.25 157.33 83.32 ;
    RECT 157.12 83.61 157.33 83.68 ;
    RECT 156.66 82.89 156.87 82.96 ;
    RECT 156.66 83.25 156.87 83.32 ;
    RECT 156.66 83.61 156.87 83.68 ;
    RECT 153.8 82.89 154.01 82.96 ;
    RECT 153.8 83.25 154.01 83.32 ;
    RECT 153.8 83.61 154.01 83.68 ;
    RECT 153.34 82.89 153.55 82.96 ;
    RECT 153.34 83.25 153.55 83.32 ;
    RECT 153.34 83.61 153.55 83.68 ;
    RECT 150.48 82.89 150.69 82.96 ;
    RECT 150.48 83.25 150.69 83.32 ;
    RECT 150.48 83.61 150.69 83.68 ;
    RECT 150.02 82.89 150.23 82.96 ;
    RECT 150.02 83.25 150.23 83.32 ;
    RECT 150.02 83.61 150.23 83.68 ;
    RECT 213.56 82.89 213.77 82.96 ;
    RECT 213.56 83.25 213.77 83.32 ;
    RECT 213.56 83.61 213.77 83.68 ;
    RECT 213.1 82.89 213.31 82.96 ;
    RECT 213.1 83.25 213.31 83.32 ;
    RECT 213.1 83.61 213.31 83.68 ;
    RECT 210.24 82.89 210.45 82.96 ;
    RECT 210.24 83.25 210.45 83.32 ;
    RECT 210.24 83.61 210.45 83.68 ;
    RECT 209.78 82.89 209.99 82.96 ;
    RECT 209.78 83.25 209.99 83.32 ;
    RECT 209.78 83.61 209.99 83.68 ;
    RECT 206.92 82.89 207.13 82.96 ;
    RECT 206.92 83.25 207.13 83.32 ;
    RECT 206.92 83.61 207.13 83.68 ;
    RECT 206.46 82.89 206.67 82.96 ;
    RECT 206.46 83.25 206.67 83.32 ;
    RECT 206.46 83.61 206.67 83.68 ;
    RECT 203.6 82.89 203.81 82.96 ;
    RECT 203.6 83.25 203.81 83.32 ;
    RECT 203.6 83.61 203.81 83.68 ;
    RECT 203.14 82.89 203.35 82.96 ;
    RECT 203.14 83.25 203.35 83.32 ;
    RECT 203.14 83.61 203.35 83.68 ;
    RECT 200.28 82.89 200.49 82.96 ;
    RECT 200.28 83.25 200.49 83.32 ;
    RECT 200.28 83.61 200.49 83.68 ;
    RECT 199.82 82.89 200.03 82.96 ;
    RECT 199.82 83.25 200.03 83.32 ;
    RECT 199.82 83.61 200.03 83.68 ;
    RECT 196.96 82.89 197.17 82.96 ;
    RECT 196.96 83.25 197.17 83.32 ;
    RECT 196.96 83.61 197.17 83.68 ;
    RECT 196.5 82.89 196.71 82.96 ;
    RECT 196.5 83.25 196.71 83.32 ;
    RECT 196.5 83.61 196.71 83.68 ;
    RECT 193.64 82.89 193.85 82.96 ;
    RECT 193.64 83.25 193.85 83.32 ;
    RECT 193.64 83.61 193.85 83.68 ;
    RECT 193.18 82.89 193.39 82.96 ;
    RECT 193.18 83.25 193.39 83.32 ;
    RECT 193.18 83.61 193.39 83.68 ;
    RECT 190.32 82.89 190.53 82.96 ;
    RECT 190.32 83.25 190.53 83.32 ;
    RECT 190.32 83.61 190.53 83.68 ;
    RECT 189.86 82.89 190.07 82.96 ;
    RECT 189.86 83.25 190.07 83.32 ;
    RECT 189.86 83.61 190.07 83.68 ;
    RECT 187.0 82.89 187.21 82.96 ;
    RECT 187.0 83.25 187.21 83.32 ;
    RECT 187.0 83.61 187.21 83.68 ;
    RECT 186.54 82.89 186.75 82.96 ;
    RECT 186.54 83.25 186.75 83.32 ;
    RECT 186.54 83.61 186.75 83.68 ;
    RECT 183.68 82.89 183.89 82.96 ;
    RECT 183.68 83.25 183.89 83.32 ;
    RECT 183.68 83.61 183.89 83.68 ;
    RECT 183.22 82.89 183.43 82.96 ;
    RECT 183.22 83.25 183.43 83.32 ;
    RECT 183.22 83.61 183.43 83.68 ;
    RECT 147.485 83.25 147.555 83.32 ;
    RECT 266.68 82.89 266.89 82.96 ;
    RECT 266.68 83.25 266.89 83.32 ;
    RECT 266.68 83.61 266.89 83.68 ;
    RECT 266.22 82.89 266.43 82.96 ;
    RECT 266.22 83.25 266.43 83.32 ;
    RECT 266.22 83.61 266.43 83.68 ;
    RECT 263.36 82.89 263.57 82.96 ;
    RECT 263.36 83.25 263.57 83.32 ;
    RECT 263.36 83.61 263.57 83.68 ;
    RECT 262.9 82.89 263.11 82.96 ;
    RECT 262.9 83.25 263.11 83.32 ;
    RECT 262.9 83.61 263.11 83.68 ;
    RECT 260.04 82.89 260.25 82.96 ;
    RECT 260.04 83.25 260.25 83.32 ;
    RECT 260.04 83.61 260.25 83.68 ;
    RECT 259.58 82.89 259.79 82.96 ;
    RECT 259.58 83.25 259.79 83.32 ;
    RECT 259.58 83.61 259.79 83.68 ;
    RECT 256.72 82.89 256.93 82.96 ;
    RECT 256.72 83.25 256.93 83.32 ;
    RECT 256.72 83.61 256.93 83.68 ;
    RECT 256.26 82.89 256.47 82.96 ;
    RECT 256.26 83.25 256.47 83.32 ;
    RECT 256.26 83.61 256.47 83.68 ;
    RECT 253.4 82.89 253.61 82.96 ;
    RECT 253.4 83.25 253.61 83.32 ;
    RECT 253.4 83.61 253.61 83.68 ;
    RECT 252.94 82.89 253.15 82.96 ;
    RECT 252.94 83.25 253.15 83.32 ;
    RECT 252.94 83.61 253.15 83.68 ;
    RECT 250.08 82.17 250.29 82.24 ;
    RECT 250.08 82.53 250.29 82.6 ;
    RECT 250.08 82.89 250.29 82.96 ;
    RECT 249.62 82.17 249.83 82.24 ;
    RECT 249.62 82.53 249.83 82.6 ;
    RECT 249.62 82.89 249.83 82.96 ;
    RECT 246.76 82.17 246.97 82.24 ;
    RECT 246.76 82.53 246.97 82.6 ;
    RECT 246.76 82.89 246.97 82.96 ;
    RECT 246.3 82.17 246.51 82.24 ;
    RECT 246.3 82.53 246.51 82.6 ;
    RECT 246.3 82.89 246.51 82.96 ;
    RECT 243.44 82.17 243.65 82.24 ;
    RECT 243.44 82.53 243.65 82.6 ;
    RECT 243.44 82.89 243.65 82.96 ;
    RECT 242.98 82.17 243.19 82.24 ;
    RECT 242.98 82.53 243.19 82.6 ;
    RECT 242.98 82.89 243.19 82.96 ;
    RECT 240.12 82.17 240.33 82.24 ;
    RECT 240.12 82.53 240.33 82.6 ;
    RECT 240.12 82.89 240.33 82.96 ;
    RECT 239.66 82.17 239.87 82.24 ;
    RECT 239.66 82.53 239.87 82.6 ;
    RECT 239.66 82.89 239.87 82.96 ;
    RECT 236.8 82.17 237.01 82.24 ;
    RECT 236.8 82.53 237.01 82.6 ;
    RECT 236.8 82.89 237.01 82.96 ;
    RECT 236.34 82.17 236.55 82.24 ;
    RECT 236.34 82.53 236.55 82.6 ;
    RECT 236.34 82.89 236.55 82.96 ;
    RECT 233.48 82.17 233.69 82.24 ;
    RECT 233.48 82.53 233.69 82.6 ;
    RECT 233.48 82.89 233.69 82.96 ;
    RECT 233.02 82.17 233.23 82.24 ;
    RECT 233.02 82.53 233.23 82.6 ;
    RECT 233.02 82.89 233.23 82.96 ;
    RECT 230.16 82.17 230.37 82.24 ;
    RECT 230.16 82.53 230.37 82.6 ;
    RECT 230.16 82.89 230.37 82.96 ;
    RECT 229.7 82.17 229.91 82.24 ;
    RECT 229.7 82.53 229.91 82.6 ;
    RECT 229.7 82.89 229.91 82.96 ;
    RECT 226.84 82.17 227.05 82.24 ;
    RECT 226.84 82.53 227.05 82.6 ;
    RECT 226.84 82.89 227.05 82.96 ;
    RECT 226.38 82.17 226.59 82.24 ;
    RECT 226.38 82.53 226.59 82.6 ;
    RECT 226.38 82.89 226.59 82.96 ;
    RECT 223.52 82.17 223.73 82.24 ;
    RECT 223.52 82.53 223.73 82.6 ;
    RECT 223.52 82.89 223.73 82.96 ;
    RECT 223.06 82.17 223.27 82.24 ;
    RECT 223.06 82.53 223.27 82.6 ;
    RECT 223.06 82.89 223.27 82.96 ;
    RECT 220.2 82.17 220.41 82.24 ;
    RECT 220.2 82.53 220.41 82.6 ;
    RECT 220.2 82.89 220.41 82.96 ;
    RECT 219.74 82.17 219.95 82.24 ;
    RECT 219.74 82.53 219.95 82.6 ;
    RECT 219.74 82.89 219.95 82.96 ;
    RECT 216.88 82.17 217.09 82.24 ;
    RECT 216.88 82.53 217.09 82.6 ;
    RECT 216.88 82.89 217.09 82.96 ;
    RECT 216.42 82.17 216.63 82.24 ;
    RECT 216.42 82.53 216.63 82.6 ;
    RECT 216.42 82.89 216.63 82.96 ;
    RECT 267.91 82.53 267.98 82.6 ;
    RECT 180.36 82.17 180.57 82.24 ;
    RECT 180.36 82.53 180.57 82.6 ;
    RECT 180.36 82.89 180.57 82.96 ;
    RECT 179.9 82.17 180.11 82.24 ;
    RECT 179.9 82.53 180.11 82.6 ;
    RECT 179.9 82.89 180.11 82.96 ;
    RECT 177.04 82.17 177.25 82.24 ;
    RECT 177.04 82.53 177.25 82.6 ;
    RECT 177.04 82.89 177.25 82.96 ;
    RECT 176.58 82.17 176.79 82.24 ;
    RECT 176.58 82.53 176.79 82.6 ;
    RECT 176.58 82.89 176.79 82.96 ;
    RECT 173.72 82.17 173.93 82.24 ;
    RECT 173.72 82.53 173.93 82.6 ;
    RECT 173.72 82.89 173.93 82.96 ;
    RECT 173.26 82.17 173.47 82.24 ;
    RECT 173.26 82.53 173.47 82.6 ;
    RECT 173.26 82.89 173.47 82.96 ;
    RECT 170.4 82.17 170.61 82.24 ;
    RECT 170.4 82.53 170.61 82.6 ;
    RECT 170.4 82.89 170.61 82.96 ;
    RECT 169.94 82.17 170.15 82.24 ;
    RECT 169.94 82.53 170.15 82.6 ;
    RECT 169.94 82.89 170.15 82.96 ;
    RECT 167.08 82.17 167.29 82.24 ;
    RECT 167.08 82.53 167.29 82.6 ;
    RECT 167.08 82.89 167.29 82.96 ;
    RECT 166.62 82.17 166.83 82.24 ;
    RECT 166.62 82.53 166.83 82.6 ;
    RECT 166.62 82.89 166.83 82.96 ;
    RECT 163.76 82.17 163.97 82.24 ;
    RECT 163.76 82.53 163.97 82.6 ;
    RECT 163.76 82.89 163.97 82.96 ;
    RECT 163.3 82.17 163.51 82.24 ;
    RECT 163.3 82.53 163.51 82.6 ;
    RECT 163.3 82.89 163.51 82.96 ;
    RECT 160.44 82.17 160.65 82.24 ;
    RECT 160.44 82.53 160.65 82.6 ;
    RECT 160.44 82.89 160.65 82.96 ;
    RECT 159.98 82.17 160.19 82.24 ;
    RECT 159.98 82.53 160.19 82.6 ;
    RECT 159.98 82.89 160.19 82.96 ;
    RECT 157.12 82.17 157.33 82.24 ;
    RECT 157.12 82.53 157.33 82.6 ;
    RECT 157.12 82.89 157.33 82.96 ;
    RECT 156.66 82.17 156.87 82.24 ;
    RECT 156.66 82.53 156.87 82.6 ;
    RECT 156.66 82.89 156.87 82.96 ;
    RECT 153.8 82.17 154.01 82.24 ;
    RECT 153.8 82.53 154.01 82.6 ;
    RECT 153.8 82.89 154.01 82.96 ;
    RECT 153.34 82.17 153.55 82.24 ;
    RECT 153.34 82.53 153.55 82.6 ;
    RECT 153.34 82.89 153.55 82.96 ;
    RECT 150.48 82.17 150.69 82.24 ;
    RECT 150.48 82.53 150.69 82.6 ;
    RECT 150.48 82.89 150.69 82.96 ;
    RECT 150.02 82.17 150.23 82.24 ;
    RECT 150.02 82.53 150.23 82.6 ;
    RECT 150.02 82.89 150.23 82.96 ;
    RECT 213.56 82.17 213.77 82.24 ;
    RECT 213.56 82.53 213.77 82.6 ;
    RECT 213.56 82.89 213.77 82.96 ;
    RECT 213.1 82.17 213.31 82.24 ;
    RECT 213.1 82.53 213.31 82.6 ;
    RECT 213.1 82.89 213.31 82.96 ;
    RECT 210.24 82.17 210.45 82.24 ;
    RECT 210.24 82.53 210.45 82.6 ;
    RECT 210.24 82.89 210.45 82.96 ;
    RECT 209.78 82.17 209.99 82.24 ;
    RECT 209.78 82.53 209.99 82.6 ;
    RECT 209.78 82.89 209.99 82.96 ;
    RECT 206.92 82.17 207.13 82.24 ;
    RECT 206.92 82.53 207.13 82.6 ;
    RECT 206.92 82.89 207.13 82.96 ;
    RECT 206.46 82.17 206.67 82.24 ;
    RECT 206.46 82.53 206.67 82.6 ;
    RECT 206.46 82.89 206.67 82.96 ;
    RECT 203.6 82.17 203.81 82.24 ;
    RECT 203.6 82.53 203.81 82.6 ;
    RECT 203.6 82.89 203.81 82.96 ;
    RECT 203.14 82.17 203.35 82.24 ;
    RECT 203.14 82.53 203.35 82.6 ;
    RECT 203.14 82.89 203.35 82.96 ;
    RECT 200.28 82.17 200.49 82.24 ;
    RECT 200.28 82.53 200.49 82.6 ;
    RECT 200.28 82.89 200.49 82.96 ;
    RECT 199.82 82.17 200.03 82.24 ;
    RECT 199.82 82.53 200.03 82.6 ;
    RECT 199.82 82.89 200.03 82.96 ;
    RECT 196.96 82.17 197.17 82.24 ;
    RECT 196.96 82.53 197.17 82.6 ;
    RECT 196.96 82.89 197.17 82.96 ;
    RECT 196.5 82.17 196.71 82.24 ;
    RECT 196.5 82.53 196.71 82.6 ;
    RECT 196.5 82.89 196.71 82.96 ;
    RECT 193.64 82.17 193.85 82.24 ;
    RECT 193.64 82.53 193.85 82.6 ;
    RECT 193.64 82.89 193.85 82.96 ;
    RECT 193.18 82.17 193.39 82.24 ;
    RECT 193.18 82.53 193.39 82.6 ;
    RECT 193.18 82.89 193.39 82.96 ;
    RECT 190.32 82.17 190.53 82.24 ;
    RECT 190.32 82.53 190.53 82.6 ;
    RECT 190.32 82.89 190.53 82.96 ;
    RECT 189.86 82.17 190.07 82.24 ;
    RECT 189.86 82.53 190.07 82.6 ;
    RECT 189.86 82.89 190.07 82.96 ;
    RECT 187.0 82.17 187.21 82.24 ;
    RECT 187.0 82.53 187.21 82.6 ;
    RECT 187.0 82.89 187.21 82.96 ;
    RECT 186.54 82.17 186.75 82.24 ;
    RECT 186.54 82.53 186.75 82.6 ;
    RECT 186.54 82.89 186.75 82.96 ;
    RECT 183.68 82.17 183.89 82.24 ;
    RECT 183.68 82.53 183.89 82.6 ;
    RECT 183.68 82.89 183.89 82.96 ;
    RECT 183.22 82.17 183.43 82.24 ;
    RECT 183.22 82.53 183.43 82.6 ;
    RECT 183.22 82.89 183.43 82.96 ;
    RECT 147.485 82.53 147.555 82.6 ;
    RECT 266.68 82.17 266.89 82.24 ;
    RECT 266.68 82.53 266.89 82.6 ;
    RECT 266.68 82.89 266.89 82.96 ;
    RECT 266.22 82.17 266.43 82.24 ;
    RECT 266.22 82.53 266.43 82.6 ;
    RECT 266.22 82.89 266.43 82.96 ;
    RECT 263.36 82.17 263.57 82.24 ;
    RECT 263.36 82.53 263.57 82.6 ;
    RECT 263.36 82.89 263.57 82.96 ;
    RECT 262.9 82.17 263.11 82.24 ;
    RECT 262.9 82.53 263.11 82.6 ;
    RECT 262.9 82.89 263.11 82.96 ;
    RECT 260.04 82.17 260.25 82.24 ;
    RECT 260.04 82.53 260.25 82.6 ;
    RECT 260.04 82.89 260.25 82.96 ;
    RECT 259.58 82.17 259.79 82.24 ;
    RECT 259.58 82.53 259.79 82.6 ;
    RECT 259.58 82.89 259.79 82.96 ;
    RECT 256.72 82.17 256.93 82.24 ;
    RECT 256.72 82.53 256.93 82.6 ;
    RECT 256.72 82.89 256.93 82.96 ;
    RECT 256.26 82.17 256.47 82.24 ;
    RECT 256.26 82.53 256.47 82.6 ;
    RECT 256.26 82.89 256.47 82.96 ;
    RECT 253.4 82.17 253.61 82.24 ;
    RECT 253.4 82.53 253.61 82.6 ;
    RECT 253.4 82.89 253.61 82.96 ;
    RECT 252.94 82.17 253.15 82.24 ;
    RECT 252.94 82.53 253.15 82.6 ;
    RECT 252.94 82.89 253.15 82.96 ;
    RECT 250.08 81.45 250.29 81.52 ;
    RECT 250.08 81.81 250.29 81.88 ;
    RECT 250.08 82.17 250.29 82.24 ;
    RECT 249.62 81.45 249.83 81.52 ;
    RECT 249.62 81.81 249.83 81.88 ;
    RECT 249.62 82.17 249.83 82.24 ;
    RECT 246.76 81.45 246.97 81.52 ;
    RECT 246.76 81.81 246.97 81.88 ;
    RECT 246.76 82.17 246.97 82.24 ;
    RECT 246.3 81.45 246.51 81.52 ;
    RECT 246.3 81.81 246.51 81.88 ;
    RECT 246.3 82.17 246.51 82.24 ;
    RECT 243.44 81.45 243.65 81.52 ;
    RECT 243.44 81.81 243.65 81.88 ;
    RECT 243.44 82.17 243.65 82.24 ;
    RECT 242.98 81.45 243.19 81.52 ;
    RECT 242.98 81.81 243.19 81.88 ;
    RECT 242.98 82.17 243.19 82.24 ;
    RECT 240.12 81.45 240.33 81.52 ;
    RECT 240.12 81.81 240.33 81.88 ;
    RECT 240.12 82.17 240.33 82.24 ;
    RECT 239.66 81.45 239.87 81.52 ;
    RECT 239.66 81.81 239.87 81.88 ;
    RECT 239.66 82.17 239.87 82.24 ;
    RECT 236.8 81.45 237.01 81.52 ;
    RECT 236.8 81.81 237.01 81.88 ;
    RECT 236.8 82.17 237.01 82.24 ;
    RECT 236.34 81.45 236.55 81.52 ;
    RECT 236.34 81.81 236.55 81.88 ;
    RECT 236.34 82.17 236.55 82.24 ;
    RECT 233.48 81.45 233.69 81.52 ;
    RECT 233.48 81.81 233.69 81.88 ;
    RECT 233.48 82.17 233.69 82.24 ;
    RECT 233.02 81.45 233.23 81.52 ;
    RECT 233.02 81.81 233.23 81.88 ;
    RECT 233.02 82.17 233.23 82.24 ;
    RECT 230.16 81.45 230.37 81.52 ;
    RECT 230.16 81.81 230.37 81.88 ;
    RECT 230.16 82.17 230.37 82.24 ;
    RECT 229.7 81.45 229.91 81.52 ;
    RECT 229.7 81.81 229.91 81.88 ;
    RECT 229.7 82.17 229.91 82.24 ;
    RECT 226.84 81.45 227.05 81.52 ;
    RECT 226.84 81.81 227.05 81.88 ;
    RECT 226.84 82.17 227.05 82.24 ;
    RECT 226.38 81.45 226.59 81.52 ;
    RECT 226.38 81.81 226.59 81.88 ;
    RECT 226.38 82.17 226.59 82.24 ;
    RECT 223.52 81.45 223.73 81.52 ;
    RECT 223.52 81.81 223.73 81.88 ;
    RECT 223.52 82.17 223.73 82.24 ;
    RECT 223.06 81.45 223.27 81.52 ;
    RECT 223.06 81.81 223.27 81.88 ;
    RECT 223.06 82.17 223.27 82.24 ;
    RECT 220.2 81.45 220.41 81.52 ;
    RECT 220.2 81.81 220.41 81.88 ;
    RECT 220.2 82.17 220.41 82.24 ;
    RECT 219.74 81.45 219.95 81.52 ;
    RECT 219.74 81.81 219.95 81.88 ;
    RECT 219.74 82.17 219.95 82.24 ;
    RECT 216.88 81.45 217.09 81.52 ;
    RECT 216.88 81.81 217.09 81.88 ;
    RECT 216.88 82.17 217.09 82.24 ;
    RECT 216.42 81.45 216.63 81.52 ;
    RECT 216.42 81.81 216.63 81.88 ;
    RECT 216.42 82.17 216.63 82.24 ;
    RECT 267.91 81.81 267.98 81.88 ;
    RECT 180.36 81.45 180.57 81.52 ;
    RECT 180.36 81.81 180.57 81.88 ;
    RECT 180.36 82.17 180.57 82.24 ;
    RECT 179.9 81.45 180.11 81.52 ;
    RECT 179.9 81.81 180.11 81.88 ;
    RECT 179.9 82.17 180.11 82.24 ;
    RECT 177.04 81.45 177.25 81.52 ;
    RECT 177.04 81.81 177.25 81.88 ;
    RECT 177.04 82.17 177.25 82.24 ;
    RECT 176.58 81.45 176.79 81.52 ;
    RECT 176.58 81.81 176.79 81.88 ;
    RECT 176.58 82.17 176.79 82.24 ;
    RECT 173.72 81.45 173.93 81.52 ;
    RECT 173.72 81.81 173.93 81.88 ;
    RECT 173.72 82.17 173.93 82.24 ;
    RECT 173.26 81.45 173.47 81.52 ;
    RECT 173.26 81.81 173.47 81.88 ;
    RECT 173.26 82.17 173.47 82.24 ;
    RECT 170.4 81.45 170.61 81.52 ;
    RECT 170.4 81.81 170.61 81.88 ;
    RECT 170.4 82.17 170.61 82.24 ;
    RECT 169.94 81.45 170.15 81.52 ;
    RECT 169.94 81.81 170.15 81.88 ;
    RECT 169.94 82.17 170.15 82.24 ;
    RECT 167.08 81.45 167.29 81.52 ;
    RECT 167.08 81.81 167.29 81.88 ;
    RECT 167.08 82.17 167.29 82.24 ;
    RECT 166.62 81.45 166.83 81.52 ;
    RECT 166.62 81.81 166.83 81.88 ;
    RECT 166.62 82.17 166.83 82.24 ;
    RECT 163.76 81.45 163.97 81.52 ;
    RECT 163.76 81.81 163.97 81.88 ;
    RECT 163.76 82.17 163.97 82.24 ;
    RECT 163.3 81.45 163.51 81.52 ;
    RECT 163.3 81.81 163.51 81.88 ;
    RECT 163.3 82.17 163.51 82.24 ;
    RECT 160.44 81.45 160.65 81.52 ;
    RECT 160.44 81.81 160.65 81.88 ;
    RECT 160.44 82.17 160.65 82.24 ;
    RECT 159.98 81.45 160.19 81.52 ;
    RECT 159.98 81.81 160.19 81.88 ;
    RECT 159.98 82.17 160.19 82.24 ;
    RECT 157.12 81.45 157.33 81.52 ;
    RECT 157.12 81.81 157.33 81.88 ;
    RECT 157.12 82.17 157.33 82.24 ;
    RECT 156.66 81.45 156.87 81.52 ;
    RECT 156.66 81.81 156.87 81.88 ;
    RECT 156.66 82.17 156.87 82.24 ;
    RECT 153.8 81.45 154.01 81.52 ;
    RECT 153.8 81.81 154.01 81.88 ;
    RECT 153.8 82.17 154.01 82.24 ;
    RECT 153.34 81.45 153.55 81.52 ;
    RECT 153.34 81.81 153.55 81.88 ;
    RECT 153.34 82.17 153.55 82.24 ;
    RECT 150.48 81.45 150.69 81.52 ;
    RECT 150.48 81.81 150.69 81.88 ;
    RECT 150.48 82.17 150.69 82.24 ;
    RECT 150.02 81.45 150.23 81.52 ;
    RECT 150.02 81.81 150.23 81.88 ;
    RECT 150.02 82.17 150.23 82.24 ;
    RECT 213.56 81.45 213.77 81.52 ;
    RECT 213.56 81.81 213.77 81.88 ;
    RECT 213.56 82.17 213.77 82.24 ;
    RECT 213.1 81.45 213.31 81.52 ;
    RECT 213.1 81.81 213.31 81.88 ;
    RECT 213.1 82.17 213.31 82.24 ;
    RECT 210.24 81.45 210.45 81.52 ;
    RECT 210.24 81.81 210.45 81.88 ;
    RECT 210.24 82.17 210.45 82.24 ;
    RECT 209.78 81.45 209.99 81.52 ;
    RECT 209.78 81.81 209.99 81.88 ;
    RECT 209.78 82.17 209.99 82.24 ;
    RECT 206.92 81.45 207.13 81.52 ;
    RECT 206.92 81.81 207.13 81.88 ;
    RECT 206.92 82.17 207.13 82.24 ;
    RECT 206.46 81.45 206.67 81.52 ;
    RECT 206.46 81.81 206.67 81.88 ;
    RECT 206.46 82.17 206.67 82.24 ;
    RECT 203.6 81.45 203.81 81.52 ;
    RECT 203.6 81.81 203.81 81.88 ;
    RECT 203.6 82.17 203.81 82.24 ;
    RECT 203.14 81.45 203.35 81.52 ;
    RECT 203.14 81.81 203.35 81.88 ;
    RECT 203.14 82.17 203.35 82.24 ;
    RECT 200.28 81.45 200.49 81.52 ;
    RECT 200.28 81.81 200.49 81.88 ;
    RECT 200.28 82.17 200.49 82.24 ;
    RECT 199.82 81.45 200.03 81.52 ;
    RECT 199.82 81.81 200.03 81.88 ;
    RECT 199.82 82.17 200.03 82.24 ;
    RECT 196.96 81.45 197.17 81.52 ;
    RECT 196.96 81.81 197.17 81.88 ;
    RECT 196.96 82.17 197.17 82.24 ;
    RECT 196.5 81.45 196.71 81.52 ;
    RECT 196.5 81.81 196.71 81.88 ;
    RECT 196.5 82.17 196.71 82.24 ;
    RECT 193.64 81.45 193.85 81.52 ;
    RECT 193.64 81.81 193.85 81.88 ;
    RECT 193.64 82.17 193.85 82.24 ;
    RECT 193.18 81.45 193.39 81.52 ;
    RECT 193.18 81.81 193.39 81.88 ;
    RECT 193.18 82.17 193.39 82.24 ;
    RECT 190.32 81.45 190.53 81.52 ;
    RECT 190.32 81.81 190.53 81.88 ;
    RECT 190.32 82.17 190.53 82.24 ;
    RECT 189.86 81.45 190.07 81.52 ;
    RECT 189.86 81.81 190.07 81.88 ;
    RECT 189.86 82.17 190.07 82.24 ;
    RECT 187.0 81.45 187.21 81.52 ;
    RECT 187.0 81.81 187.21 81.88 ;
    RECT 187.0 82.17 187.21 82.24 ;
    RECT 186.54 81.45 186.75 81.52 ;
    RECT 186.54 81.81 186.75 81.88 ;
    RECT 186.54 82.17 186.75 82.24 ;
    RECT 183.68 81.45 183.89 81.52 ;
    RECT 183.68 81.81 183.89 81.88 ;
    RECT 183.68 82.17 183.89 82.24 ;
    RECT 183.22 81.45 183.43 81.52 ;
    RECT 183.22 81.81 183.43 81.88 ;
    RECT 183.22 82.17 183.43 82.24 ;
    RECT 147.485 81.81 147.555 81.88 ;
    RECT 266.68 81.45 266.89 81.52 ;
    RECT 266.68 81.81 266.89 81.88 ;
    RECT 266.68 82.17 266.89 82.24 ;
    RECT 266.22 81.45 266.43 81.52 ;
    RECT 266.22 81.81 266.43 81.88 ;
    RECT 266.22 82.17 266.43 82.24 ;
    RECT 263.36 81.45 263.57 81.52 ;
    RECT 263.36 81.81 263.57 81.88 ;
    RECT 263.36 82.17 263.57 82.24 ;
    RECT 262.9 81.45 263.11 81.52 ;
    RECT 262.9 81.81 263.11 81.88 ;
    RECT 262.9 82.17 263.11 82.24 ;
    RECT 260.04 81.45 260.25 81.52 ;
    RECT 260.04 81.81 260.25 81.88 ;
    RECT 260.04 82.17 260.25 82.24 ;
    RECT 259.58 81.45 259.79 81.52 ;
    RECT 259.58 81.81 259.79 81.88 ;
    RECT 259.58 82.17 259.79 82.24 ;
    RECT 256.72 81.45 256.93 81.52 ;
    RECT 256.72 81.81 256.93 81.88 ;
    RECT 256.72 82.17 256.93 82.24 ;
    RECT 256.26 81.45 256.47 81.52 ;
    RECT 256.26 81.81 256.47 81.88 ;
    RECT 256.26 82.17 256.47 82.24 ;
    RECT 253.4 81.45 253.61 81.52 ;
    RECT 253.4 81.81 253.61 81.88 ;
    RECT 253.4 82.17 253.61 82.24 ;
    RECT 252.94 81.45 253.15 81.52 ;
    RECT 252.94 81.81 253.15 81.88 ;
    RECT 252.94 82.17 253.15 82.24 ;
    RECT 250.08 98.01 250.29 98.08 ;
    RECT 250.08 98.37 250.29 98.44 ;
    RECT 250.08 98.73 250.29 98.8 ;
    RECT 249.62 98.01 249.83 98.08 ;
    RECT 249.62 98.37 249.83 98.44 ;
    RECT 249.62 98.73 249.83 98.8 ;
    RECT 267.91 98.37 267.98 98.44 ;
    RECT 246.76 98.01 246.97 98.08 ;
    RECT 246.76 98.37 246.97 98.44 ;
    RECT 246.76 98.73 246.97 98.8 ;
    RECT 246.3 98.01 246.51 98.08 ;
    RECT 246.3 98.37 246.51 98.44 ;
    RECT 246.3 98.73 246.51 98.8 ;
    RECT 243.44 98.01 243.65 98.08 ;
    RECT 243.44 98.37 243.65 98.44 ;
    RECT 243.44 98.73 243.65 98.8 ;
    RECT 242.98 98.01 243.19 98.08 ;
    RECT 242.98 98.37 243.19 98.44 ;
    RECT 242.98 98.73 243.19 98.8 ;
    RECT 240.12 98.01 240.33 98.08 ;
    RECT 240.12 98.37 240.33 98.44 ;
    RECT 240.12 98.73 240.33 98.8 ;
    RECT 239.66 98.01 239.87 98.08 ;
    RECT 239.66 98.37 239.87 98.44 ;
    RECT 239.66 98.73 239.87 98.8 ;
    RECT 236.8 98.01 237.01 98.08 ;
    RECT 236.8 98.37 237.01 98.44 ;
    RECT 236.8 98.73 237.01 98.8 ;
    RECT 236.34 98.01 236.55 98.08 ;
    RECT 236.34 98.37 236.55 98.44 ;
    RECT 236.34 98.73 236.55 98.8 ;
    RECT 233.48 98.01 233.69 98.08 ;
    RECT 233.48 98.37 233.69 98.44 ;
    RECT 233.48 98.73 233.69 98.8 ;
    RECT 233.02 98.01 233.23 98.08 ;
    RECT 233.02 98.37 233.23 98.44 ;
    RECT 233.02 98.73 233.23 98.8 ;
    RECT 230.16 98.01 230.37 98.08 ;
    RECT 230.16 98.37 230.37 98.44 ;
    RECT 230.16 98.73 230.37 98.8 ;
    RECT 229.7 98.01 229.91 98.08 ;
    RECT 229.7 98.37 229.91 98.44 ;
    RECT 229.7 98.73 229.91 98.8 ;
    RECT 226.84 98.01 227.05 98.08 ;
    RECT 226.84 98.37 227.05 98.44 ;
    RECT 226.84 98.73 227.05 98.8 ;
    RECT 226.38 98.01 226.59 98.08 ;
    RECT 226.38 98.37 226.59 98.44 ;
    RECT 226.38 98.73 226.59 98.8 ;
    RECT 223.52 98.01 223.73 98.08 ;
    RECT 223.52 98.37 223.73 98.44 ;
    RECT 223.52 98.73 223.73 98.8 ;
    RECT 223.06 98.01 223.27 98.08 ;
    RECT 223.06 98.37 223.27 98.44 ;
    RECT 223.06 98.73 223.27 98.8 ;
    RECT 220.2 98.01 220.41 98.08 ;
    RECT 220.2 98.37 220.41 98.44 ;
    RECT 220.2 98.73 220.41 98.8 ;
    RECT 219.74 98.01 219.95 98.08 ;
    RECT 219.74 98.37 219.95 98.44 ;
    RECT 219.74 98.73 219.95 98.8 ;
    RECT 216.88 98.01 217.09 98.08 ;
    RECT 216.88 98.37 217.09 98.44 ;
    RECT 216.88 98.73 217.09 98.8 ;
    RECT 216.42 98.01 216.63 98.08 ;
    RECT 216.42 98.37 216.63 98.44 ;
    RECT 216.42 98.73 216.63 98.8 ;
    RECT 180.36 98.01 180.57 98.08 ;
    RECT 180.36 98.37 180.57 98.44 ;
    RECT 180.36 98.73 180.57 98.8 ;
    RECT 179.9 98.01 180.11 98.08 ;
    RECT 179.9 98.37 180.11 98.44 ;
    RECT 179.9 98.73 180.11 98.8 ;
    RECT 177.04 98.01 177.25 98.08 ;
    RECT 177.04 98.37 177.25 98.44 ;
    RECT 177.04 98.73 177.25 98.8 ;
    RECT 176.58 98.01 176.79 98.08 ;
    RECT 176.58 98.37 176.79 98.44 ;
    RECT 176.58 98.73 176.79 98.8 ;
    RECT 173.72 98.01 173.93 98.08 ;
    RECT 173.72 98.37 173.93 98.44 ;
    RECT 173.72 98.73 173.93 98.8 ;
    RECT 173.26 98.01 173.47 98.08 ;
    RECT 173.26 98.37 173.47 98.44 ;
    RECT 173.26 98.73 173.47 98.8 ;
    RECT 170.4 98.01 170.61 98.08 ;
    RECT 170.4 98.37 170.61 98.44 ;
    RECT 170.4 98.73 170.61 98.8 ;
    RECT 169.94 98.01 170.15 98.08 ;
    RECT 169.94 98.37 170.15 98.44 ;
    RECT 169.94 98.73 170.15 98.8 ;
    RECT 167.08 98.01 167.29 98.08 ;
    RECT 167.08 98.37 167.29 98.44 ;
    RECT 167.08 98.73 167.29 98.8 ;
    RECT 166.62 98.01 166.83 98.08 ;
    RECT 166.62 98.37 166.83 98.44 ;
    RECT 166.62 98.73 166.83 98.8 ;
    RECT 163.76 98.01 163.97 98.08 ;
    RECT 163.76 98.37 163.97 98.44 ;
    RECT 163.76 98.73 163.97 98.8 ;
    RECT 163.3 98.01 163.51 98.08 ;
    RECT 163.3 98.37 163.51 98.44 ;
    RECT 163.3 98.73 163.51 98.8 ;
    RECT 160.44 98.01 160.65 98.08 ;
    RECT 160.44 98.37 160.65 98.44 ;
    RECT 160.44 98.73 160.65 98.8 ;
    RECT 159.98 98.01 160.19 98.08 ;
    RECT 159.98 98.37 160.19 98.44 ;
    RECT 159.98 98.73 160.19 98.8 ;
    RECT 157.12 98.01 157.33 98.08 ;
    RECT 157.12 98.37 157.33 98.44 ;
    RECT 157.12 98.73 157.33 98.8 ;
    RECT 156.66 98.01 156.87 98.08 ;
    RECT 156.66 98.37 156.87 98.44 ;
    RECT 156.66 98.73 156.87 98.8 ;
    RECT 153.8 98.01 154.01 98.08 ;
    RECT 153.8 98.37 154.01 98.44 ;
    RECT 153.8 98.73 154.01 98.8 ;
    RECT 153.34 98.01 153.55 98.08 ;
    RECT 153.34 98.37 153.55 98.44 ;
    RECT 153.34 98.73 153.55 98.8 ;
    RECT 147.485 98.37 147.555 98.44 ;
    RECT 213.56 98.01 213.77 98.08 ;
    RECT 213.56 98.37 213.77 98.44 ;
    RECT 213.56 98.73 213.77 98.8 ;
    RECT 213.1 98.01 213.31 98.08 ;
    RECT 213.1 98.37 213.31 98.44 ;
    RECT 213.1 98.73 213.31 98.8 ;
    RECT 210.24 98.01 210.45 98.08 ;
    RECT 210.24 98.37 210.45 98.44 ;
    RECT 210.24 98.73 210.45 98.8 ;
    RECT 209.78 98.01 209.99 98.08 ;
    RECT 209.78 98.37 209.99 98.44 ;
    RECT 209.78 98.73 209.99 98.8 ;
    RECT 206.92 98.01 207.13 98.08 ;
    RECT 206.92 98.37 207.13 98.44 ;
    RECT 206.92 98.73 207.13 98.8 ;
    RECT 206.46 98.01 206.67 98.08 ;
    RECT 206.46 98.37 206.67 98.44 ;
    RECT 206.46 98.73 206.67 98.8 ;
    RECT 203.6 98.01 203.81 98.08 ;
    RECT 203.6 98.37 203.81 98.44 ;
    RECT 203.6 98.73 203.81 98.8 ;
    RECT 203.14 98.01 203.35 98.08 ;
    RECT 203.14 98.37 203.35 98.44 ;
    RECT 203.14 98.73 203.35 98.8 ;
    RECT 200.28 98.01 200.49 98.08 ;
    RECT 200.28 98.37 200.49 98.44 ;
    RECT 200.28 98.73 200.49 98.8 ;
    RECT 199.82 98.01 200.03 98.08 ;
    RECT 199.82 98.37 200.03 98.44 ;
    RECT 199.82 98.73 200.03 98.8 ;
    RECT 196.96 98.01 197.17 98.08 ;
    RECT 196.96 98.37 197.17 98.44 ;
    RECT 196.96 98.73 197.17 98.8 ;
    RECT 196.5 98.01 196.71 98.08 ;
    RECT 196.5 98.37 196.71 98.44 ;
    RECT 196.5 98.73 196.71 98.8 ;
    RECT 193.64 98.01 193.85 98.08 ;
    RECT 193.64 98.37 193.85 98.44 ;
    RECT 193.64 98.73 193.85 98.8 ;
    RECT 193.18 98.01 193.39 98.08 ;
    RECT 193.18 98.37 193.39 98.44 ;
    RECT 193.18 98.73 193.39 98.8 ;
    RECT 190.32 98.01 190.53 98.08 ;
    RECT 190.32 98.37 190.53 98.44 ;
    RECT 190.32 98.73 190.53 98.8 ;
    RECT 189.86 98.01 190.07 98.08 ;
    RECT 189.86 98.37 190.07 98.44 ;
    RECT 189.86 98.73 190.07 98.8 ;
    RECT 187.0 98.01 187.21 98.08 ;
    RECT 187.0 98.37 187.21 98.44 ;
    RECT 187.0 98.73 187.21 98.8 ;
    RECT 186.54 98.01 186.75 98.08 ;
    RECT 186.54 98.37 186.75 98.44 ;
    RECT 186.54 98.73 186.75 98.8 ;
    RECT 183.68 98.01 183.89 98.08 ;
    RECT 183.68 98.37 183.89 98.44 ;
    RECT 183.68 98.73 183.89 98.8 ;
    RECT 183.22 98.01 183.43 98.08 ;
    RECT 183.22 98.37 183.43 98.44 ;
    RECT 183.22 98.73 183.43 98.8 ;
    RECT 266.68 98.01 266.89 98.08 ;
    RECT 266.68 98.37 266.89 98.44 ;
    RECT 266.68 98.73 266.89 98.8 ;
    RECT 266.22 98.01 266.43 98.08 ;
    RECT 266.22 98.37 266.43 98.44 ;
    RECT 266.22 98.73 266.43 98.8 ;
    RECT 150.48 98.01 150.69 98.08 ;
    RECT 150.48 98.37 150.69 98.44 ;
    RECT 150.48 98.73 150.69 98.8 ;
    RECT 150.02 98.01 150.23 98.08 ;
    RECT 150.02 98.37 150.23 98.44 ;
    RECT 150.02 98.73 150.23 98.8 ;
    RECT 263.36 98.01 263.57 98.08 ;
    RECT 263.36 98.37 263.57 98.44 ;
    RECT 263.36 98.73 263.57 98.8 ;
    RECT 262.9 98.01 263.11 98.08 ;
    RECT 262.9 98.37 263.11 98.44 ;
    RECT 262.9 98.73 263.11 98.8 ;
    RECT 260.04 98.01 260.25 98.08 ;
    RECT 260.04 98.37 260.25 98.44 ;
    RECT 260.04 98.73 260.25 98.8 ;
    RECT 259.58 98.01 259.79 98.08 ;
    RECT 259.58 98.37 259.79 98.44 ;
    RECT 259.58 98.73 259.79 98.8 ;
    RECT 256.72 98.01 256.93 98.08 ;
    RECT 256.72 98.37 256.93 98.44 ;
    RECT 256.72 98.73 256.93 98.8 ;
    RECT 256.26 98.01 256.47 98.08 ;
    RECT 256.26 98.37 256.47 98.44 ;
    RECT 256.26 98.73 256.47 98.8 ;
    RECT 253.4 98.01 253.61 98.08 ;
    RECT 253.4 98.37 253.61 98.44 ;
    RECT 253.4 98.73 253.61 98.8 ;
    RECT 252.94 98.01 253.15 98.08 ;
    RECT 252.94 98.37 253.15 98.44 ;
    RECT 252.94 98.73 253.15 98.8 ;
    RECT 250.08 80.73 250.29 80.8 ;
    RECT 250.08 81.09 250.29 81.16 ;
    RECT 250.08 81.45 250.29 81.52 ;
    RECT 249.62 80.73 249.83 80.8 ;
    RECT 249.62 81.09 249.83 81.16 ;
    RECT 249.62 81.45 249.83 81.52 ;
    RECT 246.76 80.73 246.97 80.8 ;
    RECT 246.76 81.09 246.97 81.16 ;
    RECT 246.76 81.45 246.97 81.52 ;
    RECT 246.3 80.73 246.51 80.8 ;
    RECT 246.3 81.09 246.51 81.16 ;
    RECT 246.3 81.45 246.51 81.52 ;
    RECT 243.44 80.73 243.65 80.8 ;
    RECT 243.44 81.09 243.65 81.16 ;
    RECT 243.44 81.45 243.65 81.52 ;
    RECT 242.98 80.73 243.19 80.8 ;
    RECT 242.98 81.09 243.19 81.16 ;
    RECT 242.98 81.45 243.19 81.52 ;
    RECT 240.12 80.73 240.33 80.8 ;
    RECT 240.12 81.09 240.33 81.16 ;
    RECT 240.12 81.45 240.33 81.52 ;
    RECT 239.66 80.73 239.87 80.8 ;
    RECT 239.66 81.09 239.87 81.16 ;
    RECT 239.66 81.45 239.87 81.52 ;
    RECT 236.8 80.73 237.01 80.8 ;
    RECT 236.8 81.09 237.01 81.16 ;
    RECT 236.8 81.45 237.01 81.52 ;
    RECT 236.34 80.73 236.55 80.8 ;
    RECT 236.34 81.09 236.55 81.16 ;
    RECT 236.34 81.45 236.55 81.52 ;
    RECT 233.48 80.73 233.69 80.8 ;
    RECT 233.48 81.09 233.69 81.16 ;
    RECT 233.48 81.45 233.69 81.52 ;
    RECT 233.02 80.73 233.23 80.8 ;
    RECT 233.02 81.09 233.23 81.16 ;
    RECT 233.02 81.45 233.23 81.52 ;
    RECT 230.16 80.73 230.37 80.8 ;
    RECT 230.16 81.09 230.37 81.16 ;
    RECT 230.16 81.45 230.37 81.52 ;
    RECT 229.7 80.73 229.91 80.8 ;
    RECT 229.7 81.09 229.91 81.16 ;
    RECT 229.7 81.45 229.91 81.52 ;
    RECT 226.84 80.73 227.05 80.8 ;
    RECT 226.84 81.09 227.05 81.16 ;
    RECT 226.84 81.45 227.05 81.52 ;
    RECT 226.38 80.73 226.59 80.8 ;
    RECT 226.38 81.09 226.59 81.16 ;
    RECT 226.38 81.45 226.59 81.52 ;
    RECT 223.52 80.73 223.73 80.8 ;
    RECT 223.52 81.09 223.73 81.16 ;
    RECT 223.52 81.45 223.73 81.52 ;
    RECT 223.06 80.73 223.27 80.8 ;
    RECT 223.06 81.09 223.27 81.16 ;
    RECT 223.06 81.45 223.27 81.52 ;
    RECT 220.2 80.73 220.41 80.8 ;
    RECT 220.2 81.09 220.41 81.16 ;
    RECT 220.2 81.45 220.41 81.52 ;
    RECT 219.74 80.73 219.95 80.8 ;
    RECT 219.74 81.09 219.95 81.16 ;
    RECT 219.74 81.45 219.95 81.52 ;
    RECT 216.88 80.73 217.09 80.8 ;
    RECT 216.88 81.09 217.09 81.16 ;
    RECT 216.88 81.45 217.09 81.52 ;
    RECT 216.42 80.73 216.63 80.8 ;
    RECT 216.42 81.09 216.63 81.16 ;
    RECT 216.42 81.45 216.63 81.52 ;
    RECT 267.91 81.09 267.98 81.16 ;
    RECT 180.36 80.73 180.57 80.8 ;
    RECT 180.36 81.09 180.57 81.16 ;
    RECT 180.36 81.45 180.57 81.52 ;
    RECT 179.9 80.73 180.11 80.8 ;
    RECT 179.9 81.09 180.11 81.16 ;
    RECT 179.9 81.45 180.11 81.52 ;
    RECT 177.04 80.73 177.25 80.8 ;
    RECT 177.04 81.09 177.25 81.16 ;
    RECT 177.04 81.45 177.25 81.52 ;
    RECT 176.58 80.73 176.79 80.8 ;
    RECT 176.58 81.09 176.79 81.16 ;
    RECT 176.58 81.45 176.79 81.52 ;
    RECT 173.72 80.73 173.93 80.8 ;
    RECT 173.72 81.09 173.93 81.16 ;
    RECT 173.72 81.45 173.93 81.52 ;
    RECT 173.26 80.73 173.47 80.8 ;
    RECT 173.26 81.09 173.47 81.16 ;
    RECT 173.26 81.45 173.47 81.52 ;
    RECT 170.4 80.73 170.61 80.8 ;
    RECT 170.4 81.09 170.61 81.16 ;
    RECT 170.4 81.45 170.61 81.52 ;
    RECT 169.94 80.73 170.15 80.8 ;
    RECT 169.94 81.09 170.15 81.16 ;
    RECT 169.94 81.45 170.15 81.52 ;
    RECT 167.08 80.73 167.29 80.8 ;
    RECT 167.08 81.09 167.29 81.16 ;
    RECT 167.08 81.45 167.29 81.52 ;
    RECT 166.62 80.73 166.83 80.8 ;
    RECT 166.62 81.09 166.83 81.16 ;
    RECT 166.62 81.45 166.83 81.52 ;
    RECT 163.76 80.73 163.97 80.8 ;
    RECT 163.76 81.09 163.97 81.16 ;
    RECT 163.76 81.45 163.97 81.52 ;
    RECT 163.3 80.73 163.51 80.8 ;
    RECT 163.3 81.09 163.51 81.16 ;
    RECT 163.3 81.45 163.51 81.52 ;
    RECT 160.44 80.73 160.65 80.8 ;
    RECT 160.44 81.09 160.65 81.16 ;
    RECT 160.44 81.45 160.65 81.52 ;
    RECT 159.98 80.73 160.19 80.8 ;
    RECT 159.98 81.09 160.19 81.16 ;
    RECT 159.98 81.45 160.19 81.52 ;
    RECT 157.12 80.73 157.33 80.8 ;
    RECT 157.12 81.09 157.33 81.16 ;
    RECT 157.12 81.45 157.33 81.52 ;
    RECT 156.66 80.73 156.87 80.8 ;
    RECT 156.66 81.09 156.87 81.16 ;
    RECT 156.66 81.45 156.87 81.52 ;
    RECT 153.8 80.73 154.01 80.8 ;
    RECT 153.8 81.09 154.01 81.16 ;
    RECT 153.8 81.45 154.01 81.52 ;
    RECT 153.34 80.73 153.55 80.8 ;
    RECT 153.34 81.09 153.55 81.16 ;
    RECT 153.34 81.45 153.55 81.52 ;
    RECT 150.48 80.73 150.69 80.8 ;
    RECT 150.48 81.09 150.69 81.16 ;
    RECT 150.48 81.45 150.69 81.52 ;
    RECT 150.02 80.73 150.23 80.8 ;
    RECT 150.02 81.09 150.23 81.16 ;
    RECT 150.02 81.45 150.23 81.52 ;
    RECT 213.56 80.73 213.77 80.8 ;
    RECT 213.56 81.09 213.77 81.16 ;
    RECT 213.56 81.45 213.77 81.52 ;
    RECT 213.1 80.73 213.31 80.8 ;
    RECT 213.1 81.09 213.31 81.16 ;
    RECT 213.1 81.45 213.31 81.52 ;
    RECT 210.24 80.73 210.45 80.8 ;
    RECT 210.24 81.09 210.45 81.16 ;
    RECT 210.24 81.45 210.45 81.52 ;
    RECT 209.78 80.73 209.99 80.8 ;
    RECT 209.78 81.09 209.99 81.16 ;
    RECT 209.78 81.45 209.99 81.52 ;
    RECT 206.92 80.73 207.13 80.8 ;
    RECT 206.92 81.09 207.13 81.16 ;
    RECT 206.92 81.45 207.13 81.52 ;
    RECT 206.46 80.73 206.67 80.8 ;
    RECT 206.46 81.09 206.67 81.16 ;
    RECT 206.46 81.45 206.67 81.52 ;
    RECT 203.6 80.73 203.81 80.8 ;
    RECT 203.6 81.09 203.81 81.16 ;
    RECT 203.6 81.45 203.81 81.52 ;
    RECT 203.14 80.73 203.35 80.8 ;
    RECT 203.14 81.09 203.35 81.16 ;
    RECT 203.14 81.45 203.35 81.52 ;
    RECT 200.28 80.73 200.49 80.8 ;
    RECT 200.28 81.09 200.49 81.16 ;
    RECT 200.28 81.45 200.49 81.52 ;
    RECT 199.82 80.73 200.03 80.8 ;
    RECT 199.82 81.09 200.03 81.16 ;
    RECT 199.82 81.45 200.03 81.52 ;
    RECT 196.96 80.73 197.17 80.8 ;
    RECT 196.96 81.09 197.17 81.16 ;
    RECT 196.96 81.45 197.17 81.52 ;
    RECT 196.5 80.73 196.71 80.8 ;
    RECT 196.5 81.09 196.71 81.16 ;
    RECT 196.5 81.45 196.71 81.52 ;
    RECT 193.64 80.73 193.85 80.8 ;
    RECT 193.64 81.09 193.85 81.16 ;
    RECT 193.64 81.45 193.85 81.52 ;
    RECT 193.18 80.73 193.39 80.8 ;
    RECT 193.18 81.09 193.39 81.16 ;
    RECT 193.18 81.45 193.39 81.52 ;
    RECT 190.32 80.73 190.53 80.8 ;
    RECT 190.32 81.09 190.53 81.16 ;
    RECT 190.32 81.45 190.53 81.52 ;
    RECT 189.86 80.73 190.07 80.8 ;
    RECT 189.86 81.09 190.07 81.16 ;
    RECT 189.86 81.45 190.07 81.52 ;
    RECT 187.0 80.73 187.21 80.8 ;
    RECT 187.0 81.09 187.21 81.16 ;
    RECT 187.0 81.45 187.21 81.52 ;
    RECT 186.54 80.73 186.75 80.8 ;
    RECT 186.54 81.09 186.75 81.16 ;
    RECT 186.54 81.45 186.75 81.52 ;
    RECT 183.68 80.73 183.89 80.8 ;
    RECT 183.68 81.09 183.89 81.16 ;
    RECT 183.68 81.45 183.89 81.52 ;
    RECT 183.22 80.73 183.43 80.8 ;
    RECT 183.22 81.09 183.43 81.16 ;
    RECT 183.22 81.45 183.43 81.52 ;
    RECT 147.485 81.09 147.555 81.16 ;
    RECT 266.68 80.73 266.89 80.8 ;
    RECT 266.68 81.09 266.89 81.16 ;
    RECT 266.68 81.45 266.89 81.52 ;
    RECT 266.22 80.73 266.43 80.8 ;
    RECT 266.22 81.09 266.43 81.16 ;
    RECT 266.22 81.45 266.43 81.52 ;
    RECT 263.36 80.73 263.57 80.8 ;
    RECT 263.36 81.09 263.57 81.16 ;
    RECT 263.36 81.45 263.57 81.52 ;
    RECT 262.9 80.73 263.11 80.8 ;
    RECT 262.9 81.09 263.11 81.16 ;
    RECT 262.9 81.45 263.11 81.52 ;
    RECT 260.04 80.73 260.25 80.8 ;
    RECT 260.04 81.09 260.25 81.16 ;
    RECT 260.04 81.45 260.25 81.52 ;
    RECT 259.58 80.73 259.79 80.8 ;
    RECT 259.58 81.09 259.79 81.16 ;
    RECT 259.58 81.45 259.79 81.52 ;
    RECT 256.72 80.73 256.93 80.8 ;
    RECT 256.72 81.09 256.93 81.16 ;
    RECT 256.72 81.45 256.93 81.52 ;
    RECT 256.26 80.73 256.47 80.8 ;
    RECT 256.26 81.09 256.47 81.16 ;
    RECT 256.26 81.45 256.47 81.52 ;
    RECT 253.4 80.73 253.61 80.8 ;
    RECT 253.4 81.09 253.61 81.16 ;
    RECT 253.4 81.45 253.61 81.52 ;
    RECT 252.94 80.73 253.15 80.8 ;
    RECT 252.94 81.09 253.15 81.16 ;
    RECT 252.94 81.45 253.15 81.52 ;
    RECT 250.08 80.01 250.29 80.08 ;
    RECT 250.08 80.37 250.29 80.44 ;
    RECT 250.08 80.73 250.29 80.8 ;
    RECT 249.62 80.01 249.83 80.08 ;
    RECT 249.62 80.37 249.83 80.44 ;
    RECT 249.62 80.73 249.83 80.8 ;
    RECT 246.76 80.01 246.97 80.08 ;
    RECT 246.76 80.37 246.97 80.44 ;
    RECT 246.76 80.73 246.97 80.8 ;
    RECT 246.3 80.01 246.51 80.08 ;
    RECT 246.3 80.37 246.51 80.44 ;
    RECT 246.3 80.73 246.51 80.8 ;
    RECT 243.44 80.01 243.65 80.08 ;
    RECT 243.44 80.37 243.65 80.44 ;
    RECT 243.44 80.73 243.65 80.8 ;
    RECT 242.98 80.01 243.19 80.08 ;
    RECT 242.98 80.37 243.19 80.44 ;
    RECT 242.98 80.73 243.19 80.8 ;
    RECT 240.12 80.01 240.33 80.08 ;
    RECT 240.12 80.37 240.33 80.44 ;
    RECT 240.12 80.73 240.33 80.8 ;
    RECT 239.66 80.01 239.87 80.08 ;
    RECT 239.66 80.37 239.87 80.44 ;
    RECT 239.66 80.73 239.87 80.8 ;
    RECT 236.8 80.01 237.01 80.08 ;
    RECT 236.8 80.37 237.01 80.44 ;
    RECT 236.8 80.73 237.01 80.8 ;
    RECT 236.34 80.01 236.55 80.08 ;
    RECT 236.34 80.37 236.55 80.44 ;
    RECT 236.34 80.73 236.55 80.8 ;
    RECT 233.48 80.01 233.69 80.08 ;
    RECT 233.48 80.37 233.69 80.44 ;
    RECT 233.48 80.73 233.69 80.8 ;
    RECT 233.02 80.01 233.23 80.08 ;
    RECT 233.02 80.37 233.23 80.44 ;
    RECT 233.02 80.73 233.23 80.8 ;
    RECT 230.16 80.01 230.37 80.08 ;
    RECT 230.16 80.37 230.37 80.44 ;
    RECT 230.16 80.73 230.37 80.8 ;
    RECT 229.7 80.01 229.91 80.08 ;
    RECT 229.7 80.37 229.91 80.44 ;
    RECT 229.7 80.73 229.91 80.8 ;
    RECT 226.84 80.01 227.05 80.08 ;
    RECT 226.84 80.37 227.05 80.44 ;
    RECT 226.84 80.73 227.05 80.8 ;
    RECT 226.38 80.01 226.59 80.08 ;
    RECT 226.38 80.37 226.59 80.44 ;
    RECT 226.38 80.73 226.59 80.8 ;
    RECT 223.52 80.01 223.73 80.08 ;
    RECT 223.52 80.37 223.73 80.44 ;
    RECT 223.52 80.73 223.73 80.8 ;
    RECT 223.06 80.01 223.27 80.08 ;
    RECT 223.06 80.37 223.27 80.44 ;
    RECT 223.06 80.73 223.27 80.8 ;
    RECT 220.2 80.01 220.41 80.08 ;
    RECT 220.2 80.37 220.41 80.44 ;
    RECT 220.2 80.73 220.41 80.8 ;
    RECT 219.74 80.01 219.95 80.08 ;
    RECT 219.74 80.37 219.95 80.44 ;
    RECT 219.74 80.73 219.95 80.8 ;
    RECT 216.88 80.01 217.09 80.08 ;
    RECT 216.88 80.37 217.09 80.44 ;
    RECT 216.88 80.73 217.09 80.8 ;
    RECT 216.42 80.01 216.63 80.08 ;
    RECT 216.42 80.37 216.63 80.44 ;
    RECT 216.42 80.73 216.63 80.8 ;
    RECT 267.91 80.37 267.98 80.44 ;
    RECT 180.36 80.01 180.57 80.08 ;
    RECT 180.36 80.37 180.57 80.44 ;
    RECT 180.36 80.73 180.57 80.8 ;
    RECT 179.9 80.01 180.11 80.08 ;
    RECT 179.9 80.37 180.11 80.44 ;
    RECT 179.9 80.73 180.11 80.8 ;
    RECT 177.04 80.01 177.25 80.08 ;
    RECT 177.04 80.37 177.25 80.44 ;
    RECT 177.04 80.73 177.25 80.8 ;
    RECT 176.58 80.01 176.79 80.08 ;
    RECT 176.58 80.37 176.79 80.44 ;
    RECT 176.58 80.73 176.79 80.8 ;
    RECT 173.72 80.01 173.93 80.08 ;
    RECT 173.72 80.37 173.93 80.44 ;
    RECT 173.72 80.73 173.93 80.8 ;
    RECT 173.26 80.01 173.47 80.08 ;
    RECT 173.26 80.37 173.47 80.44 ;
    RECT 173.26 80.73 173.47 80.8 ;
    RECT 170.4 80.01 170.61 80.08 ;
    RECT 170.4 80.37 170.61 80.44 ;
    RECT 170.4 80.73 170.61 80.8 ;
    RECT 169.94 80.01 170.15 80.08 ;
    RECT 169.94 80.37 170.15 80.44 ;
    RECT 169.94 80.73 170.15 80.8 ;
    RECT 167.08 80.01 167.29 80.08 ;
    RECT 167.08 80.37 167.29 80.44 ;
    RECT 167.08 80.73 167.29 80.8 ;
    RECT 166.62 80.01 166.83 80.08 ;
    RECT 166.62 80.37 166.83 80.44 ;
    RECT 166.62 80.73 166.83 80.8 ;
    RECT 163.76 80.01 163.97 80.08 ;
    RECT 163.76 80.37 163.97 80.44 ;
    RECT 163.76 80.73 163.97 80.8 ;
    RECT 163.3 80.01 163.51 80.08 ;
    RECT 163.3 80.37 163.51 80.44 ;
    RECT 163.3 80.73 163.51 80.8 ;
    RECT 160.44 80.01 160.65 80.08 ;
    RECT 160.44 80.37 160.65 80.44 ;
    RECT 160.44 80.73 160.65 80.8 ;
    RECT 159.98 80.01 160.19 80.08 ;
    RECT 159.98 80.37 160.19 80.44 ;
    RECT 159.98 80.73 160.19 80.8 ;
    RECT 157.12 80.01 157.33 80.08 ;
    RECT 157.12 80.37 157.33 80.44 ;
    RECT 157.12 80.73 157.33 80.8 ;
    RECT 156.66 80.01 156.87 80.08 ;
    RECT 156.66 80.37 156.87 80.44 ;
    RECT 156.66 80.73 156.87 80.8 ;
    RECT 153.8 80.01 154.01 80.08 ;
    RECT 153.8 80.37 154.01 80.44 ;
    RECT 153.8 80.73 154.01 80.8 ;
    RECT 153.34 80.01 153.55 80.08 ;
    RECT 153.34 80.37 153.55 80.44 ;
    RECT 153.34 80.73 153.55 80.8 ;
    RECT 150.48 80.01 150.69 80.08 ;
    RECT 150.48 80.37 150.69 80.44 ;
    RECT 150.48 80.73 150.69 80.8 ;
    RECT 150.02 80.01 150.23 80.08 ;
    RECT 150.02 80.37 150.23 80.44 ;
    RECT 150.02 80.73 150.23 80.8 ;
    RECT 213.56 80.01 213.77 80.08 ;
    RECT 213.56 80.37 213.77 80.44 ;
    RECT 213.56 80.73 213.77 80.8 ;
    RECT 213.1 80.01 213.31 80.08 ;
    RECT 213.1 80.37 213.31 80.44 ;
    RECT 213.1 80.73 213.31 80.8 ;
    RECT 210.24 80.01 210.45 80.08 ;
    RECT 210.24 80.37 210.45 80.44 ;
    RECT 210.24 80.73 210.45 80.8 ;
    RECT 209.78 80.01 209.99 80.08 ;
    RECT 209.78 80.37 209.99 80.44 ;
    RECT 209.78 80.73 209.99 80.8 ;
    RECT 206.92 80.01 207.13 80.08 ;
    RECT 206.92 80.37 207.13 80.44 ;
    RECT 206.92 80.73 207.13 80.8 ;
    RECT 206.46 80.01 206.67 80.08 ;
    RECT 206.46 80.37 206.67 80.44 ;
    RECT 206.46 80.73 206.67 80.8 ;
    RECT 203.6 80.01 203.81 80.08 ;
    RECT 203.6 80.37 203.81 80.44 ;
    RECT 203.6 80.73 203.81 80.8 ;
    RECT 203.14 80.01 203.35 80.08 ;
    RECT 203.14 80.37 203.35 80.44 ;
    RECT 203.14 80.73 203.35 80.8 ;
    RECT 200.28 80.01 200.49 80.08 ;
    RECT 200.28 80.37 200.49 80.44 ;
    RECT 200.28 80.73 200.49 80.8 ;
    RECT 199.82 80.01 200.03 80.08 ;
    RECT 199.82 80.37 200.03 80.44 ;
    RECT 199.82 80.73 200.03 80.8 ;
    RECT 196.96 80.01 197.17 80.08 ;
    RECT 196.96 80.37 197.17 80.44 ;
    RECT 196.96 80.73 197.17 80.8 ;
    RECT 196.5 80.01 196.71 80.08 ;
    RECT 196.5 80.37 196.71 80.44 ;
    RECT 196.5 80.73 196.71 80.8 ;
    RECT 193.64 80.01 193.85 80.08 ;
    RECT 193.64 80.37 193.85 80.44 ;
    RECT 193.64 80.73 193.85 80.8 ;
    RECT 193.18 80.01 193.39 80.08 ;
    RECT 193.18 80.37 193.39 80.44 ;
    RECT 193.18 80.73 193.39 80.8 ;
    RECT 190.32 80.01 190.53 80.08 ;
    RECT 190.32 80.37 190.53 80.44 ;
    RECT 190.32 80.73 190.53 80.8 ;
    RECT 189.86 80.01 190.07 80.08 ;
    RECT 189.86 80.37 190.07 80.44 ;
    RECT 189.86 80.73 190.07 80.8 ;
    RECT 187.0 80.01 187.21 80.08 ;
    RECT 187.0 80.37 187.21 80.44 ;
    RECT 187.0 80.73 187.21 80.8 ;
    RECT 186.54 80.01 186.75 80.08 ;
    RECT 186.54 80.37 186.75 80.44 ;
    RECT 186.54 80.73 186.75 80.8 ;
    RECT 183.68 80.01 183.89 80.08 ;
    RECT 183.68 80.37 183.89 80.44 ;
    RECT 183.68 80.73 183.89 80.8 ;
    RECT 183.22 80.01 183.43 80.08 ;
    RECT 183.22 80.37 183.43 80.44 ;
    RECT 183.22 80.73 183.43 80.8 ;
    RECT 147.485 80.37 147.555 80.44 ;
    RECT 266.68 80.01 266.89 80.08 ;
    RECT 266.68 80.37 266.89 80.44 ;
    RECT 266.68 80.73 266.89 80.8 ;
    RECT 266.22 80.01 266.43 80.08 ;
    RECT 266.22 80.37 266.43 80.44 ;
    RECT 266.22 80.73 266.43 80.8 ;
    RECT 263.36 80.01 263.57 80.08 ;
    RECT 263.36 80.37 263.57 80.44 ;
    RECT 263.36 80.73 263.57 80.8 ;
    RECT 262.9 80.01 263.11 80.08 ;
    RECT 262.9 80.37 263.11 80.44 ;
    RECT 262.9 80.73 263.11 80.8 ;
    RECT 260.04 80.01 260.25 80.08 ;
    RECT 260.04 80.37 260.25 80.44 ;
    RECT 260.04 80.73 260.25 80.8 ;
    RECT 259.58 80.01 259.79 80.08 ;
    RECT 259.58 80.37 259.79 80.44 ;
    RECT 259.58 80.73 259.79 80.8 ;
    RECT 256.72 80.01 256.93 80.08 ;
    RECT 256.72 80.37 256.93 80.44 ;
    RECT 256.72 80.73 256.93 80.8 ;
    RECT 256.26 80.01 256.47 80.08 ;
    RECT 256.26 80.37 256.47 80.44 ;
    RECT 256.26 80.73 256.47 80.8 ;
    RECT 253.4 80.01 253.61 80.08 ;
    RECT 253.4 80.37 253.61 80.44 ;
    RECT 253.4 80.73 253.61 80.8 ;
    RECT 252.94 80.01 253.15 80.08 ;
    RECT 252.94 80.37 253.15 80.44 ;
    RECT 252.94 80.73 253.15 80.8 ;
    RECT 250.08 42.55 250.29 42.62 ;
    RECT 250.08 42.91 250.29 42.98 ;
    RECT 250.08 43.27 250.29 43.34 ;
    RECT 249.62 42.55 249.83 42.62 ;
    RECT 249.62 42.91 249.83 42.98 ;
    RECT 249.62 43.27 249.83 43.34 ;
    RECT 246.76 42.55 246.97 42.62 ;
    RECT 246.76 42.91 246.97 42.98 ;
    RECT 246.76 43.27 246.97 43.34 ;
    RECT 246.3 42.55 246.51 42.62 ;
    RECT 246.3 42.91 246.51 42.98 ;
    RECT 246.3 43.27 246.51 43.34 ;
    RECT 243.44 42.55 243.65 42.62 ;
    RECT 243.44 42.91 243.65 42.98 ;
    RECT 243.44 43.27 243.65 43.34 ;
    RECT 242.98 42.55 243.19 42.62 ;
    RECT 242.98 42.91 243.19 42.98 ;
    RECT 242.98 43.27 243.19 43.34 ;
    RECT 240.12 42.55 240.33 42.62 ;
    RECT 240.12 42.91 240.33 42.98 ;
    RECT 240.12 43.27 240.33 43.34 ;
    RECT 239.66 42.55 239.87 42.62 ;
    RECT 239.66 42.91 239.87 42.98 ;
    RECT 239.66 43.27 239.87 43.34 ;
    RECT 236.8 42.55 237.01 42.62 ;
    RECT 236.8 42.91 237.01 42.98 ;
    RECT 236.8 43.27 237.01 43.34 ;
    RECT 236.34 42.55 236.55 42.62 ;
    RECT 236.34 42.91 236.55 42.98 ;
    RECT 236.34 43.27 236.55 43.34 ;
    RECT 233.48 42.55 233.69 42.62 ;
    RECT 233.48 42.91 233.69 42.98 ;
    RECT 233.48 43.27 233.69 43.34 ;
    RECT 233.02 42.55 233.23 42.62 ;
    RECT 233.02 42.91 233.23 42.98 ;
    RECT 233.02 43.27 233.23 43.34 ;
    RECT 230.16 42.55 230.37 42.62 ;
    RECT 230.16 42.91 230.37 42.98 ;
    RECT 230.16 43.27 230.37 43.34 ;
    RECT 229.7 42.55 229.91 42.62 ;
    RECT 229.7 42.91 229.91 42.98 ;
    RECT 229.7 43.27 229.91 43.34 ;
    RECT 226.84 42.55 227.05 42.62 ;
    RECT 226.84 42.91 227.05 42.98 ;
    RECT 226.84 43.27 227.05 43.34 ;
    RECT 226.38 42.55 226.59 42.62 ;
    RECT 226.38 42.91 226.59 42.98 ;
    RECT 226.38 43.27 226.59 43.34 ;
    RECT 223.52 42.55 223.73 42.62 ;
    RECT 223.52 42.91 223.73 42.98 ;
    RECT 223.52 43.27 223.73 43.34 ;
    RECT 223.06 42.55 223.27 42.62 ;
    RECT 223.06 42.91 223.27 42.98 ;
    RECT 223.06 43.27 223.27 43.34 ;
    RECT 220.2 42.55 220.41 42.62 ;
    RECT 220.2 42.91 220.41 42.98 ;
    RECT 220.2 43.27 220.41 43.34 ;
    RECT 219.74 42.55 219.95 42.62 ;
    RECT 219.74 42.91 219.95 42.98 ;
    RECT 219.74 43.27 219.95 43.34 ;
    RECT 216.88 42.55 217.09 42.62 ;
    RECT 216.88 42.91 217.09 42.98 ;
    RECT 216.88 43.27 217.09 43.34 ;
    RECT 216.42 42.55 216.63 42.62 ;
    RECT 216.42 42.91 216.63 42.98 ;
    RECT 216.42 43.27 216.63 43.34 ;
    RECT 267.91 42.91 267.98 42.98 ;
    RECT 180.36 42.55 180.57 42.62 ;
    RECT 180.36 42.91 180.57 42.98 ;
    RECT 180.36 43.27 180.57 43.34 ;
    RECT 179.9 42.55 180.11 42.62 ;
    RECT 179.9 42.91 180.11 42.98 ;
    RECT 179.9 43.27 180.11 43.34 ;
    RECT 177.04 42.55 177.25 42.62 ;
    RECT 177.04 42.91 177.25 42.98 ;
    RECT 177.04 43.27 177.25 43.34 ;
    RECT 176.58 42.55 176.79 42.62 ;
    RECT 176.58 42.91 176.79 42.98 ;
    RECT 176.58 43.27 176.79 43.34 ;
    RECT 173.72 42.55 173.93 42.62 ;
    RECT 173.72 42.91 173.93 42.98 ;
    RECT 173.72 43.27 173.93 43.34 ;
    RECT 173.26 42.55 173.47 42.62 ;
    RECT 173.26 42.91 173.47 42.98 ;
    RECT 173.26 43.27 173.47 43.34 ;
    RECT 170.4 42.55 170.61 42.62 ;
    RECT 170.4 42.91 170.61 42.98 ;
    RECT 170.4 43.27 170.61 43.34 ;
    RECT 169.94 42.55 170.15 42.62 ;
    RECT 169.94 42.91 170.15 42.98 ;
    RECT 169.94 43.27 170.15 43.34 ;
    RECT 167.08 42.55 167.29 42.62 ;
    RECT 167.08 42.91 167.29 42.98 ;
    RECT 167.08 43.27 167.29 43.34 ;
    RECT 166.62 42.55 166.83 42.62 ;
    RECT 166.62 42.91 166.83 42.98 ;
    RECT 166.62 43.27 166.83 43.34 ;
    RECT 163.76 42.55 163.97 42.62 ;
    RECT 163.76 42.91 163.97 42.98 ;
    RECT 163.76 43.27 163.97 43.34 ;
    RECT 163.3 42.55 163.51 42.62 ;
    RECT 163.3 42.91 163.51 42.98 ;
    RECT 163.3 43.27 163.51 43.34 ;
    RECT 160.44 42.55 160.65 42.62 ;
    RECT 160.44 42.91 160.65 42.98 ;
    RECT 160.44 43.27 160.65 43.34 ;
    RECT 159.98 42.55 160.19 42.62 ;
    RECT 159.98 42.91 160.19 42.98 ;
    RECT 159.98 43.27 160.19 43.34 ;
    RECT 157.12 42.55 157.33 42.62 ;
    RECT 157.12 42.91 157.33 42.98 ;
    RECT 157.12 43.27 157.33 43.34 ;
    RECT 156.66 42.55 156.87 42.62 ;
    RECT 156.66 42.91 156.87 42.98 ;
    RECT 156.66 43.27 156.87 43.34 ;
    RECT 153.8 42.55 154.01 42.62 ;
    RECT 153.8 42.91 154.01 42.98 ;
    RECT 153.8 43.27 154.01 43.34 ;
    RECT 153.34 42.55 153.55 42.62 ;
    RECT 153.34 42.91 153.55 42.98 ;
    RECT 153.34 43.27 153.55 43.34 ;
    RECT 150.48 42.55 150.69 42.62 ;
    RECT 150.48 42.91 150.69 42.98 ;
    RECT 150.48 43.27 150.69 43.34 ;
    RECT 150.02 42.55 150.23 42.62 ;
    RECT 150.02 42.91 150.23 42.98 ;
    RECT 150.02 43.27 150.23 43.34 ;
    RECT 213.56 42.55 213.77 42.62 ;
    RECT 213.56 42.91 213.77 42.98 ;
    RECT 213.56 43.27 213.77 43.34 ;
    RECT 213.1 42.55 213.31 42.62 ;
    RECT 213.1 42.91 213.31 42.98 ;
    RECT 213.1 43.27 213.31 43.34 ;
    RECT 210.24 42.55 210.45 42.62 ;
    RECT 210.24 42.91 210.45 42.98 ;
    RECT 210.24 43.27 210.45 43.34 ;
    RECT 209.78 42.55 209.99 42.62 ;
    RECT 209.78 42.91 209.99 42.98 ;
    RECT 209.78 43.27 209.99 43.34 ;
    RECT 206.92 42.55 207.13 42.62 ;
    RECT 206.92 42.91 207.13 42.98 ;
    RECT 206.92 43.27 207.13 43.34 ;
    RECT 206.46 42.55 206.67 42.62 ;
    RECT 206.46 42.91 206.67 42.98 ;
    RECT 206.46 43.27 206.67 43.34 ;
    RECT 203.6 42.55 203.81 42.62 ;
    RECT 203.6 42.91 203.81 42.98 ;
    RECT 203.6 43.27 203.81 43.34 ;
    RECT 203.14 42.55 203.35 42.62 ;
    RECT 203.14 42.91 203.35 42.98 ;
    RECT 203.14 43.27 203.35 43.34 ;
    RECT 200.28 42.55 200.49 42.62 ;
    RECT 200.28 42.91 200.49 42.98 ;
    RECT 200.28 43.27 200.49 43.34 ;
    RECT 199.82 42.55 200.03 42.62 ;
    RECT 199.82 42.91 200.03 42.98 ;
    RECT 199.82 43.27 200.03 43.34 ;
    RECT 196.96 42.55 197.17 42.62 ;
    RECT 196.96 42.91 197.17 42.98 ;
    RECT 196.96 43.27 197.17 43.34 ;
    RECT 196.5 42.55 196.71 42.62 ;
    RECT 196.5 42.91 196.71 42.98 ;
    RECT 196.5 43.27 196.71 43.34 ;
    RECT 193.64 42.55 193.85 42.62 ;
    RECT 193.64 42.91 193.85 42.98 ;
    RECT 193.64 43.27 193.85 43.34 ;
    RECT 193.18 42.55 193.39 42.62 ;
    RECT 193.18 42.91 193.39 42.98 ;
    RECT 193.18 43.27 193.39 43.34 ;
    RECT 190.32 42.55 190.53 42.62 ;
    RECT 190.32 42.91 190.53 42.98 ;
    RECT 190.32 43.27 190.53 43.34 ;
    RECT 189.86 42.55 190.07 42.62 ;
    RECT 189.86 42.91 190.07 42.98 ;
    RECT 189.86 43.27 190.07 43.34 ;
    RECT 187.0 42.55 187.21 42.62 ;
    RECT 187.0 42.91 187.21 42.98 ;
    RECT 187.0 43.27 187.21 43.34 ;
    RECT 186.54 42.55 186.75 42.62 ;
    RECT 186.54 42.91 186.75 42.98 ;
    RECT 186.54 43.27 186.75 43.34 ;
    RECT 183.68 42.55 183.89 42.62 ;
    RECT 183.68 42.91 183.89 42.98 ;
    RECT 183.68 43.27 183.89 43.34 ;
    RECT 183.22 42.55 183.43 42.62 ;
    RECT 183.22 42.91 183.43 42.98 ;
    RECT 183.22 43.27 183.43 43.34 ;
    RECT 147.485 42.91 147.555 42.98 ;
    RECT 266.68 42.55 266.89 42.62 ;
    RECT 266.68 42.91 266.89 42.98 ;
    RECT 266.68 43.27 266.89 43.34 ;
    RECT 266.22 42.55 266.43 42.62 ;
    RECT 266.22 42.91 266.43 42.98 ;
    RECT 266.22 43.27 266.43 43.34 ;
    RECT 263.36 42.55 263.57 42.62 ;
    RECT 263.36 42.91 263.57 42.98 ;
    RECT 263.36 43.27 263.57 43.34 ;
    RECT 262.9 42.55 263.11 42.62 ;
    RECT 262.9 42.91 263.11 42.98 ;
    RECT 262.9 43.27 263.11 43.34 ;
    RECT 260.04 42.55 260.25 42.62 ;
    RECT 260.04 42.91 260.25 42.98 ;
    RECT 260.04 43.27 260.25 43.34 ;
    RECT 259.58 42.55 259.79 42.62 ;
    RECT 259.58 42.91 259.79 42.98 ;
    RECT 259.58 43.27 259.79 43.34 ;
    RECT 256.72 42.55 256.93 42.62 ;
    RECT 256.72 42.91 256.93 42.98 ;
    RECT 256.72 43.27 256.93 43.34 ;
    RECT 256.26 42.55 256.47 42.62 ;
    RECT 256.26 42.91 256.47 42.98 ;
    RECT 256.26 43.27 256.47 43.34 ;
    RECT 253.4 42.55 253.61 42.62 ;
    RECT 253.4 42.91 253.61 42.98 ;
    RECT 253.4 43.27 253.61 43.34 ;
    RECT 252.94 42.55 253.15 42.62 ;
    RECT 252.94 42.91 253.15 42.98 ;
    RECT 252.94 43.27 253.15 43.34 ;
    RECT 250.08 41.83 250.29 41.9 ;
    RECT 250.08 42.19 250.29 42.26 ;
    RECT 250.08 42.55 250.29 42.62 ;
    RECT 249.62 41.83 249.83 41.9 ;
    RECT 249.62 42.19 249.83 42.26 ;
    RECT 249.62 42.55 249.83 42.62 ;
    RECT 246.76 41.83 246.97 41.9 ;
    RECT 246.76 42.19 246.97 42.26 ;
    RECT 246.76 42.55 246.97 42.62 ;
    RECT 246.3 41.83 246.51 41.9 ;
    RECT 246.3 42.19 246.51 42.26 ;
    RECT 246.3 42.55 246.51 42.62 ;
    RECT 243.44 41.83 243.65 41.9 ;
    RECT 243.44 42.19 243.65 42.26 ;
    RECT 243.44 42.55 243.65 42.62 ;
    RECT 242.98 41.83 243.19 41.9 ;
    RECT 242.98 42.19 243.19 42.26 ;
    RECT 242.98 42.55 243.19 42.62 ;
    RECT 240.12 41.83 240.33 41.9 ;
    RECT 240.12 42.19 240.33 42.26 ;
    RECT 240.12 42.55 240.33 42.62 ;
    RECT 239.66 41.83 239.87 41.9 ;
    RECT 239.66 42.19 239.87 42.26 ;
    RECT 239.66 42.55 239.87 42.62 ;
    RECT 236.8 41.83 237.01 41.9 ;
    RECT 236.8 42.19 237.01 42.26 ;
    RECT 236.8 42.55 237.01 42.62 ;
    RECT 236.34 41.83 236.55 41.9 ;
    RECT 236.34 42.19 236.55 42.26 ;
    RECT 236.34 42.55 236.55 42.62 ;
    RECT 233.48 41.83 233.69 41.9 ;
    RECT 233.48 42.19 233.69 42.26 ;
    RECT 233.48 42.55 233.69 42.62 ;
    RECT 233.02 41.83 233.23 41.9 ;
    RECT 233.02 42.19 233.23 42.26 ;
    RECT 233.02 42.55 233.23 42.62 ;
    RECT 230.16 41.83 230.37 41.9 ;
    RECT 230.16 42.19 230.37 42.26 ;
    RECT 230.16 42.55 230.37 42.62 ;
    RECT 229.7 41.83 229.91 41.9 ;
    RECT 229.7 42.19 229.91 42.26 ;
    RECT 229.7 42.55 229.91 42.62 ;
    RECT 226.84 41.83 227.05 41.9 ;
    RECT 226.84 42.19 227.05 42.26 ;
    RECT 226.84 42.55 227.05 42.62 ;
    RECT 226.38 41.83 226.59 41.9 ;
    RECT 226.38 42.19 226.59 42.26 ;
    RECT 226.38 42.55 226.59 42.62 ;
    RECT 223.52 41.83 223.73 41.9 ;
    RECT 223.52 42.19 223.73 42.26 ;
    RECT 223.52 42.55 223.73 42.62 ;
    RECT 223.06 41.83 223.27 41.9 ;
    RECT 223.06 42.19 223.27 42.26 ;
    RECT 223.06 42.55 223.27 42.62 ;
    RECT 220.2 41.83 220.41 41.9 ;
    RECT 220.2 42.19 220.41 42.26 ;
    RECT 220.2 42.55 220.41 42.62 ;
    RECT 219.74 41.83 219.95 41.9 ;
    RECT 219.74 42.19 219.95 42.26 ;
    RECT 219.74 42.55 219.95 42.62 ;
    RECT 216.88 41.83 217.09 41.9 ;
    RECT 216.88 42.19 217.09 42.26 ;
    RECT 216.88 42.55 217.09 42.62 ;
    RECT 216.42 41.83 216.63 41.9 ;
    RECT 216.42 42.19 216.63 42.26 ;
    RECT 216.42 42.55 216.63 42.62 ;
    RECT 267.91 42.19 267.98 42.26 ;
    RECT 180.36 41.83 180.57 41.9 ;
    RECT 180.36 42.19 180.57 42.26 ;
    RECT 180.36 42.55 180.57 42.62 ;
    RECT 179.9 41.83 180.11 41.9 ;
    RECT 179.9 42.19 180.11 42.26 ;
    RECT 179.9 42.55 180.11 42.62 ;
    RECT 177.04 41.83 177.25 41.9 ;
    RECT 177.04 42.19 177.25 42.26 ;
    RECT 177.04 42.55 177.25 42.62 ;
    RECT 176.58 41.83 176.79 41.9 ;
    RECT 176.58 42.19 176.79 42.26 ;
    RECT 176.58 42.55 176.79 42.62 ;
    RECT 173.72 41.83 173.93 41.9 ;
    RECT 173.72 42.19 173.93 42.26 ;
    RECT 173.72 42.55 173.93 42.62 ;
    RECT 173.26 41.83 173.47 41.9 ;
    RECT 173.26 42.19 173.47 42.26 ;
    RECT 173.26 42.55 173.47 42.62 ;
    RECT 170.4 41.83 170.61 41.9 ;
    RECT 170.4 42.19 170.61 42.26 ;
    RECT 170.4 42.55 170.61 42.62 ;
    RECT 169.94 41.83 170.15 41.9 ;
    RECT 169.94 42.19 170.15 42.26 ;
    RECT 169.94 42.55 170.15 42.62 ;
    RECT 167.08 41.83 167.29 41.9 ;
    RECT 167.08 42.19 167.29 42.26 ;
    RECT 167.08 42.55 167.29 42.62 ;
    RECT 166.62 41.83 166.83 41.9 ;
    RECT 166.62 42.19 166.83 42.26 ;
    RECT 166.62 42.55 166.83 42.62 ;
    RECT 163.76 41.83 163.97 41.9 ;
    RECT 163.76 42.19 163.97 42.26 ;
    RECT 163.76 42.55 163.97 42.62 ;
    RECT 163.3 41.83 163.51 41.9 ;
    RECT 163.3 42.19 163.51 42.26 ;
    RECT 163.3 42.55 163.51 42.62 ;
    RECT 160.44 41.83 160.65 41.9 ;
    RECT 160.44 42.19 160.65 42.26 ;
    RECT 160.44 42.55 160.65 42.62 ;
    RECT 159.98 41.83 160.19 41.9 ;
    RECT 159.98 42.19 160.19 42.26 ;
    RECT 159.98 42.55 160.19 42.62 ;
    RECT 157.12 41.83 157.33 41.9 ;
    RECT 157.12 42.19 157.33 42.26 ;
    RECT 157.12 42.55 157.33 42.62 ;
    RECT 156.66 41.83 156.87 41.9 ;
    RECT 156.66 42.19 156.87 42.26 ;
    RECT 156.66 42.55 156.87 42.62 ;
    RECT 153.8 41.83 154.01 41.9 ;
    RECT 153.8 42.19 154.01 42.26 ;
    RECT 153.8 42.55 154.01 42.62 ;
    RECT 153.34 41.83 153.55 41.9 ;
    RECT 153.34 42.19 153.55 42.26 ;
    RECT 153.34 42.55 153.55 42.62 ;
    RECT 150.48 41.83 150.69 41.9 ;
    RECT 150.48 42.19 150.69 42.26 ;
    RECT 150.48 42.55 150.69 42.62 ;
    RECT 150.02 41.83 150.23 41.9 ;
    RECT 150.02 42.19 150.23 42.26 ;
    RECT 150.02 42.55 150.23 42.62 ;
    RECT 213.56 41.83 213.77 41.9 ;
    RECT 213.56 42.19 213.77 42.26 ;
    RECT 213.56 42.55 213.77 42.62 ;
    RECT 213.1 41.83 213.31 41.9 ;
    RECT 213.1 42.19 213.31 42.26 ;
    RECT 213.1 42.55 213.31 42.62 ;
    RECT 210.24 41.83 210.45 41.9 ;
    RECT 210.24 42.19 210.45 42.26 ;
    RECT 210.24 42.55 210.45 42.62 ;
    RECT 209.78 41.83 209.99 41.9 ;
    RECT 209.78 42.19 209.99 42.26 ;
    RECT 209.78 42.55 209.99 42.62 ;
    RECT 206.92 41.83 207.13 41.9 ;
    RECT 206.92 42.19 207.13 42.26 ;
    RECT 206.92 42.55 207.13 42.62 ;
    RECT 206.46 41.83 206.67 41.9 ;
    RECT 206.46 42.19 206.67 42.26 ;
    RECT 206.46 42.55 206.67 42.62 ;
    RECT 203.6 41.83 203.81 41.9 ;
    RECT 203.6 42.19 203.81 42.26 ;
    RECT 203.6 42.55 203.81 42.62 ;
    RECT 203.14 41.83 203.35 41.9 ;
    RECT 203.14 42.19 203.35 42.26 ;
    RECT 203.14 42.55 203.35 42.62 ;
    RECT 200.28 41.83 200.49 41.9 ;
    RECT 200.28 42.19 200.49 42.26 ;
    RECT 200.28 42.55 200.49 42.62 ;
    RECT 199.82 41.83 200.03 41.9 ;
    RECT 199.82 42.19 200.03 42.26 ;
    RECT 199.82 42.55 200.03 42.62 ;
    RECT 196.96 41.83 197.17 41.9 ;
    RECT 196.96 42.19 197.17 42.26 ;
    RECT 196.96 42.55 197.17 42.62 ;
    RECT 196.5 41.83 196.71 41.9 ;
    RECT 196.5 42.19 196.71 42.26 ;
    RECT 196.5 42.55 196.71 42.62 ;
    RECT 193.64 41.83 193.85 41.9 ;
    RECT 193.64 42.19 193.85 42.26 ;
    RECT 193.64 42.55 193.85 42.62 ;
    RECT 193.18 41.83 193.39 41.9 ;
    RECT 193.18 42.19 193.39 42.26 ;
    RECT 193.18 42.55 193.39 42.62 ;
    RECT 190.32 41.83 190.53 41.9 ;
    RECT 190.32 42.19 190.53 42.26 ;
    RECT 190.32 42.55 190.53 42.62 ;
    RECT 189.86 41.83 190.07 41.9 ;
    RECT 189.86 42.19 190.07 42.26 ;
    RECT 189.86 42.55 190.07 42.62 ;
    RECT 187.0 41.83 187.21 41.9 ;
    RECT 187.0 42.19 187.21 42.26 ;
    RECT 187.0 42.55 187.21 42.62 ;
    RECT 186.54 41.83 186.75 41.9 ;
    RECT 186.54 42.19 186.75 42.26 ;
    RECT 186.54 42.55 186.75 42.62 ;
    RECT 183.68 41.83 183.89 41.9 ;
    RECT 183.68 42.19 183.89 42.26 ;
    RECT 183.68 42.55 183.89 42.62 ;
    RECT 183.22 41.83 183.43 41.9 ;
    RECT 183.22 42.19 183.43 42.26 ;
    RECT 183.22 42.55 183.43 42.62 ;
    RECT 147.485 42.19 147.555 42.26 ;
    RECT 266.68 41.83 266.89 41.9 ;
    RECT 266.68 42.19 266.89 42.26 ;
    RECT 266.68 42.55 266.89 42.62 ;
    RECT 266.22 41.83 266.43 41.9 ;
    RECT 266.22 42.19 266.43 42.26 ;
    RECT 266.22 42.55 266.43 42.62 ;
    RECT 263.36 41.83 263.57 41.9 ;
    RECT 263.36 42.19 263.57 42.26 ;
    RECT 263.36 42.55 263.57 42.62 ;
    RECT 262.9 41.83 263.11 41.9 ;
    RECT 262.9 42.19 263.11 42.26 ;
    RECT 262.9 42.55 263.11 42.62 ;
    RECT 260.04 41.83 260.25 41.9 ;
    RECT 260.04 42.19 260.25 42.26 ;
    RECT 260.04 42.55 260.25 42.62 ;
    RECT 259.58 41.83 259.79 41.9 ;
    RECT 259.58 42.19 259.79 42.26 ;
    RECT 259.58 42.55 259.79 42.62 ;
    RECT 256.72 41.83 256.93 41.9 ;
    RECT 256.72 42.19 256.93 42.26 ;
    RECT 256.72 42.55 256.93 42.62 ;
    RECT 256.26 41.83 256.47 41.9 ;
    RECT 256.26 42.19 256.47 42.26 ;
    RECT 256.26 42.55 256.47 42.62 ;
    RECT 253.4 41.83 253.61 41.9 ;
    RECT 253.4 42.19 253.61 42.26 ;
    RECT 253.4 42.55 253.61 42.62 ;
    RECT 252.94 41.83 253.15 41.9 ;
    RECT 252.94 42.19 253.15 42.26 ;
    RECT 252.94 42.55 253.15 42.62 ;
    RECT 250.08 41.11 250.29 41.18 ;
    RECT 250.08 41.47 250.29 41.54 ;
    RECT 250.08 41.83 250.29 41.9 ;
    RECT 249.62 41.11 249.83 41.18 ;
    RECT 249.62 41.47 249.83 41.54 ;
    RECT 249.62 41.83 249.83 41.9 ;
    RECT 246.76 41.11 246.97 41.18 ;
    RECT 246.76 41.47 246.97 41.54 ;
    RECT 246.76 41.83 246.97 41.9 ;
    RECT 246.3 41.11 246.51 41.18 ;
    RECT 246.3 41.47 246.51 41.54 ;
    RECT 246.3 41.83 246.51 41.9 ;
    RECT 243.44 41.11 243.65 41.18 ;
    RECT 243.44 41.47 243.65 41.54 ;
    RECT 243.44 41.83 243.65 41.9 ;
    RECT 242.98 41.11 243.19 41.18 ;
    RECT 242.98 41.47 243.19 41.54 ;
    RECT 242.98 41.83 243.19 41.9 ;
    RECT 240.12 41.11 240.33 41.18 ;
    RECT 240.12 41.47 240.33 41.54 ;
    RECT 240.12 41.83 240.33 41.9 ;
    RECT 239.66 41.11 239.87 41.18 ;
    RECT 239.66 41.47 239.87 41.54 ;
    RECT 239.66 41.83 239.87 41.9 ;
    RECT 236.8 41.11 237.01 41.18 ;
    RECT 236.8 41.47 237.01 41.54 ;
    RECT 236.8 41.83 237.01 41.9 ;
    RECT 236.34 41.11 236.55 41.18 ;
    RECT 236.34 41.47 236.55 41.54 ;
    RECT 236.34 41.83 236.55 41.9 ;
    RECT 233.48 41.11 233.69 41.18 ;
    RECT 233.48 41.47 233.69 41.54 ;
    RECT 233.48 41.83 233.69 41.9 ;
    RECT 233.02 41.11 233.23 41.18 ;
    RECT 233.02 41.47 233.23 41.54 ;
    RECT 233.02 41.83 233.23 41.9 ;
    RECT 230.16 41.11 230.37 41.18 ;
    RECT 230.16 41.47 230.37 41.54 ;
    RECT 230.16 41.83 230.37 41.9 ;
    RECT 229.7 41.11 229.91 41.18 ;
    RECT 229.7 41.47 229.91 41.54 ;
    RECT 229.7 41.83 229.91 41.9 ;
    RECT 226.84 41.11 227.05 41.18 ;
    RECT 226.84 41.47 227.05 41.54 ;
    RECT 226.84 41.83 227.05 41.9 ;
    RECT 226.38 41.11 226.59 41.18 ;
    RECT 226.38 41.47 226.59 41.54 ;
    RECT 226.38 41.83 226.59 41.9 ;
    RECT 223.52 41.11 223.73 41.18 ;
    RECT 223.52 41.47 223.73 41.54 ;
    RECT 223.52 41.83 223.73 41.9 ;
    RECT 223.06 41.11 223.27 41.18 ;
    RECT 223.06 41.47 223.27 41.54 ;
    RECT 223.06 41.83 223.27 41.9 ;
    RECT 220.2 41.11 220.41 41.18 ;
    RECT 220.2 41.47 220.41 41.54 ;
    RECT 220.2 41.83 220.41 41.9 ;
    RECT 219.74 41.11 219.95 41.18 ;
    RECT 219.74 41.47 219.95 41.54 ;
    RECT 219.74 41.83 219.95 41.9 ;
    RECT 216.88 41.11 217.09 41.18 ;
    RECT 216.88 41.47 217.09 41.54 ;
    RECT 216.88 41.83 217.09 41.9 ;
    RECT 216.42 41.11 216.63 41.18 ;
    RECT 216.42 41.47 216.63 41.54 ;
    RECT 216.42 41.83 216.63 41.9 ;
    RECT 267.91 41.47 267.98 41.54 ;
    RECT 180.36 41.11 180.57 41.18 ;
    RECT 180.36 41.47 180.57 41.54 ;
    RECT 180.36 41.83 180.57 41.9 ;
    RECT 179.9 41.11 180.11 41.18 ;
    RECT 179.9 41.47 180.11 41.54 ;
    RECT 179.9 41.83 180.11 41.9 ;
    RECT 177.04 41.11 177.25 41.18 ;
    RECT 177.04 41.47 177.25 41.54 ;
    RECT 177.04 41.83 177.25 41.9 ;
    RECT 176.58 41.11 176.79 41.18 ;
    RECT 176.58 41.47 176.79 41.54 ;
    RECT 176.58 41.83 176.79 41.9 ;
    RECT 173.72 41.11 173.93 41.18 ;
    RECT 173.72 41.47 173.93 41.54 ;
    RECT 173.72 41.83 173.93 41.9 ;
    RECT 173.26 41.11 173.47 41.18 ;
    RECT 173.26 41.47 173.47 41.54 ;
    RECT 173.26 41.83 173.47 41.9 ;
    RECT 170.4 41.11 170.61 41.18 ;
    RECT 170.4 41.47 170.61 41.54 ;
    RECT 170.4 41.83 170.61 41.9 ;
    RECT 169.94 41.11 170.15 41.18 ;
    RECT 169.94 41.47 170.15 41.54 ;
    RECT 169.94 41.83 170.15 41.9 ;
    RECT 167.08 41.11 167.29 41.18 ;
    RECT 167.08 41.47 167.29 41.54 ;
    RECT 167.08 41.83 167.29 41.9 ;
    RECT 166.62 41.11 166.83 41.18 ;
    RECT 166.62 41.47 166.83 41.54 ;
    RECT 166.62 41.83 166.83 41.9 ;
    RECT 163.76 41.11 163.97 41.18 ;
    RECT 163.76 41.47 163.97 41.54 ;
    RECT 163.76 41.83 163.97 41.9 ;
    RECT 163.3 41.11 163.51 41.18 ;
    RECT 163.3 41.47 163.51 41.54 ;
    RECT 163.3 41.83 163.51 41.9 ;
    RECT 160.44 41.11 160.65 41.18 ;
    RECT 160.44 41.47 160.65 41.54 ;
    RECT 160.44 41.83 160.65 41.9 ;
    RECT 159.98 41.11 160.19 41.18 ;
    RECT 159.98 41.47 160.19 41.54 ;
    RECT 159.98 41.83 160.19 41.9 ;
    RECT 157.12 41.11 157.33 41.18 ;
    RECT 157.12 41.47 157.33 41.54 ;
    RECT 157.12 41.83 157.33 41.9 ;
    RECT 156.66 41.11 156.87 41.18 ;
    RECT 156.66 41.47 156.87 41.54 ;
    RECT 156.66 41.83 156.87 41.9 ;
    RECT 153.8 41.11 154.01 41.18 ;
    RECT 153.8 41.47 154.01 41.54 ;
    RECT 153.8 41.83 154.01 41.9 ;
    RECT 153.34 41.11 153.55 41.18 ;
    RECT 153.34 41.47 153.55 41.54 ;
    RECT 153.34 41.83 153.55 41.9 ;
    RECT 150.48 41.11 150.69 41.18 ;
    RECT 150.48 41.47 150.69 41.54 ;
    RECT 150.48 41.83 150.69 41.9 ;
    RECT 150.02 41.11 150.23 41.18 ;
    RECT 150.02 41.47 150.23 41.54 ;
    RECT 150.02 41.83 150.23 41.9 ;
    RECT 213.56 41.11 213.77 41.18 ;
    RECT 213.56 41.47 213.77 41.54 ;
    RECT 213.56 41.83 213.77 41.9 ;
    RECT 213.1 41.11 213.31 41.18 ;
    RECT 213.1 41.47 213.31 41.54 ;
    RECT 213.1 41.83 213.31 41.9 ;
    RECT 210.24 41.11 210.45 41.18 ;
    RECT 210.24 41.47 210.45 41.54 ;
    RECT 210.24 41.83 210.45 41.9 ;
    RECT 209.78 41.11 209.99 41.18 ;
    RECT 209.78 41.47 209.99 41.54 ;
    RECT 209.78 41.83 209.99 41.9 ;
    RECT 206.92 41.11 207.13 41.18 ;
    RECT 206.92 41.47 207.13 41.54 ;
    RECT 206.92 41.83 207.13 41.9 ;
    RECT 206.46 41.11 206.67 41.18 ;
    RECT 206.46 41.47 206.67 41.54 ;
    RECT 206.46 41.83 206.67 41.9 ;
    RECT 203.6 41.11 203.81 41.18 ;
    RECT 203.6 41.47 203.81 41.54 ;
    RECT 203.6 41.83 203.81 41.9 ;
    RECT 203.14 41.11 203.35 41.18 ;
    RECT 203.14 41.47 203.35 41.54 ;
    RECT 203.14 41.83 203.35 41.9 ;
    RECT 200.28 41.11 200.49 41.18 ;
    RECT 200.28 41.47 200.49 41.54 ;
    RECT 200.28 41.83 200.49 41.9 ;
    RECT 199.82 41.11 200.03 41.18 ;
    RECT 199.82 41.47 200.03 41.54 ;
    RECT 199.82 41.83 200.03 41.9 ;
    RECT 196.96 41.11 197.17 41.18 ;
    RECT 196.96 41.47 197.17 41.54 ;
    RECT 196.96 41.83 197.17 41.9 ;
    RECT 196.5 41.11 196.71 41.18 ;
    RECT 196.5 41.47 196.71 41.54 ;
    RECT 196.5 41.83 196.71 41.9 ;
    RECT 193.64 41.11 193.85 41.18 ;
    RECT 193.64 41.47 193.85 41.54 ;
    RECT 193.64 41.83 193.85 41.9 ;
    RECT 193.18 41.11 193.39 41.18 ;
    RECT 193.18 41.47 193.39 41.54 ;
    RECT 193.18 41.83 193.39 41.9 ;
    RECT 190.32 41.11 190.53 41.18 ;
    RECT 190.32 41.47 190.53 41.54 ;
    RECT 190.32 41.83 190.53 41.9 ;
    RECT 189.86 41.11 190.07 41.18 ;
    RECT 189.86 41.47 190.07 41.54 ;
    RECT 189.86 41.83 190.07 41.9 ;
    RECT 187.0 41.11 187.21 41.18 ;
    RECT 187.0 41.47 187.21 41.54 ;
    RECT 187.0 41.83 187.21 41.9 ;
    RECT 186.54 41.11 186.75 41.18 ;
    RECT 186.54 41.47 186.75 41.54 ;
    RECT 186.54 41.83 186.75 41.9 ;
    RECT 183.68 41.11 183.89 41.18 ;
    RECT 183.68 41.47 183.89 41.54 ;
    RECT 183.68 41.83 183.89 41.9 ;
    RECT 183.22 41.11 183.43 41.18 ;
    RECT 183.22 41.47 183.43 41.54 ;
    RECT 183.22 41.83 183.43 41.9 ;
    RECT 147.485 41.47 147.555 41.54 ;
    RECT 266.68 41.11 266.89 41.18 ;
    RECT 266.68 41.47 266.89 41.54 ;
    RECT 266.68 41.83 266.89 41.9 ;
    RECT 266.22 41.11 266.43 41.18 ;
    RECT 266.22 41.47 266.43 41.54 ;
    RECT 266.22 41.83 266.43 41.9 ;
    RECT 263.36 41.11 263.57 41.18 ;
    RECT 263.36 41.47 263.57 41.54 ;
    RECT 263.36 41.83 263.57 41.9 ;
    RECT 262.9 41.11 263.11 41.18 ;
    RECT 262.9 41.47 263.11 41.54 ;
    RECT 262.9 41.83 263.11 41.9 ;
    RECT 260.04 41.11 260.25 41.18 ;
    RECT 260.04 41.47 260.25 41.54 ;
    RECT 260.04 41.83 260.25 41.9 ;
    RECT 259.58 41.11 259.79 41.18 ;
    RECT 259.58 41.47 259.79 41.54 ;
    RECT 259.58 41.83 259.79 41.9 ;
    RECT 256.72 41.11 256.93 41.18 ;
    RECT 256.72 41.47 256.93 41.54 ;
    RECT 256.72 41.83 256.93 41.9 ;
    RECT 256.26 41.11 256.47 41.18 ;
    RECT 256.26 41.47 256.47 41.54 ;
    RECT 256.26 41.83 256.47 41.9 ;
    RECT 253.4 41.11 253.61 41.18 ;
    RECT 253.4 41.47 253.61 41.54 ;
    RECT 253.4 41.83 253.61 41.9 ;
    RECT 252.94 41.11 253.15 41.18 ;
    RECT 252.94 41.47 253.15 41.54 ;
    RECT 252.94 41.83 253.15 41.9 ;
    RECT 250.08 40.39 250.29 40.46 ;
    RECT 250.08 40.75 250.29 40.82 ;
    RECT 250.08 41.11 250.29 41.18 ;
    RECT 249.62 40.39 249.83 40.46 ;
    RECT 249.62 40.75 249.83 40.82 ;
    RECT 249.62 41.11 249.83 41.18 ;
    RECT 246.76 40.39 246.97 40.46 ;
    RECT 246.76 40.75 246.97 40.82 ;
    RECT 246.76 41.11 246.97 41.18 ;
    RECT 246.3 40.39 246.51 40.46 ;
    RECT 246.3 40.75 246.51 40.82 ;
    RECT 246.3 41.11 246.51 41.18 ;
    RECT 243.44 40.39 243.65 40.46 ;
    RECT 243.44 40.75 243.65 40.82 ;
    RECT 243.44 41.11 243.65 41.18 ;
    RECT 242.98 40.39 243.19 40.46 ;
    RECT 242.98 40.75 243.19 40.82 ;
    RECT 242.98 41.11 243.19 41.18 ;
    RECT 240.12 40.39 240.33 40.46 ;
    RECT 240.12 40.75 240.33 40.82 ;
    RECT 240.12 41.11 240.33 41.18 ;
    RECT 239.66 40.39 239.87 40.46 ;
    RECT 239.66 40.75 239.87 40.82 ;
    RECT 239.66 41.11 239.87 41.18 ;
    RECT 236.8 40.39 237.01 40.46 ;
    RECT 236.8 40.75 237.01 40.82 ;
    RECT 236.8 41.11 237.01 41.18 ;
    RECT 236.34 40.39 236.55 40.46 ;
    RECT 236.34 40.75 236.55 40.82 ;
    RECT 236.34 41.11 236.55 41.18 ;
    RECT 233.48 40.39 233.69 40.46 ;
    RECT 233.48 40.75 233.69 40.82 ;
    RECT 233.48 41.11 233.69 41.18 ;
    RECT 233.02 40.39 233.23 40.46 ;
    RECT 233.02 40.75 233.23 40.82 ;
    RECT 233.02 41.11 233.23 41.18 ;
    RECT 230.16 40.39 230.37 40.46 ;
    RECT 230.16 40.75 230.37 40.82 ;
    RECT 230.16 41.11 230.37 41.18 ;
    RECT 229.7 40.39 229.91 40.46 ;
    RECT 229.7 40.75 229.91 40.82 ;
    RECT 229.7 41.11 229.91 41.18 ;
    RECT 226.84 40.39 227.05 40.46 ;
    RECT 226.84 40.75 227.05 40.82 ;
    RECT 226.84 41.11 227.05 41.18 ;
    RECT 226.38 40.39 226.59 40.46 ;
    RECT 226.38 40.75 226.59 40.82 ;
    RECT 226.38 41.11 226.59 41.18 ;
    RECT 223.52 40.39 223.73 40.46 ;
    RECT 223.52 40.75 223.73 40.82 ;
    RECT 223.52 41.11 223.73 41.18 ;
    RECT 223.06 40.39 223.27 40.46 ;
    RECT 223.06 40.75 223.27 40.82 ;
    RECT 223.06 41.11 223.27 41.18 ;
    RECT 220.2 40.39 220.41 40.46 ;
    RECT 220.2 40.75 220.41 40.82 ;
    RECT 220.2 41.11 220.41 41.18 ;
    RECT 219.74 40.39 219.95 40.46 ;
    RECT 219.74 40.75 219.95 40.82 ;
    RECT 219.74 41.11 219.95 41.18 ;
    RECT 216.88 40.39 217.09 40.46 ;
    RECT 216.88 40.75 217.09 40.82 ;
    RECT 216.88 41.11 217.09 41.18 ;
    RECT 216.42 40.39 216.63 40.46 ;
    RECT 216.42 40.75 216.63 40.82 ;
    RECT 216.42 41.11 216.63 41.18 ;
    RECT 267.91 40.75 267.98 40.82 ;
    RECT 180.36 40.39 180.57 40.46 ;
    RECT 180.36 40.75 180.57 40.82 ;
    RECT 180.36 41.11 180.57 41.18 ;
    RECT 179.9 40.39 180.11 40.46 ;
    RECT 179.9 40.75 180.11 40.82 ;
    RECT 179.9 41.11 180.11 41.18 ;
    RECT 177.04 40.39 177.25 40.46 ;
    RECT 177.04 40.75 177.25 40.82 ;
    RECT 177.04 41.11 177.25 41.18 ;
    RECT 176.58 40.39 176.79 40.46 ;
    RECT 176.58 40.75 176.79 40.82 ;
    RECT 176.58 41.11 176.79 41.18 ;
    RECT 173.72 40.39 173.93 40.46 ;
    RECT 173.72 40.75 173.93 40.82 ;
    RECT 173.72 41.11 173.93 41.18 ;
    RECT 173.26 40.39 173.47 40.46 ;
    RECT 173.26 40.75 173.47 40.82 ;
    RECT 173.26 41.11 173.47 41.18 ;
    RECT 170.4 40.39 170.61 40.46 ;
    RECT 170.4 40.75 170.61 40.82 ;
    RECT 170.4 41.11 170.61 41.18 ;
    RECT 169.94 40.39 170.15 40.46 ;
    RECT 169.94 40.75 170.15 40.82 ;
    RECT 169.94 41.11 170.15 41.18 ;
    RECT 167.08 40.39 167.29 40.46 ;
    RECT 167.08 40.75 167.29 40.82 ;
    RECT 167.08 41.11 167.29 41.18 ;
    RECT 166.62 40.39 166.83 40.46 ;
    RECT 166.62 40.75 166.83 40.82 ;
    RECT 166.62 41.11 166.83 41.18 ;
    RECT 163.76 40.39 163.97 40.46 ;
    RECT 163.76 40.75 163.97 40.82 ;
    RECT 163.76 41.11 163.97 41.18 ;
    RECT 163.3 40.39 163.51 40.46 ;
    RECT 163.3 40.75 163.51 40.82 ;
    RECT 163.3 41.11 163.51 41.18 ;
    RECT 160.44 40.39 160.65 40.46 ;
    RECT 160.44 40.75 160.65 40.82 ;
    RECT 160.44 41.11 160.65 41.18 ;
    RECT 159.98 40.39 160.19 40.46 ;
    RECT 159.98 40.75 160.19 40.82 ;
    RECT 159.98 41.11 160.19 41.18 ;
    RECT 157.12 40.39 157.33 40.46 ;
    RECT 157.12 40.75 157.33 40.82 ;
    RECT 157.12 41.11 157.33 41.18 ;
    RECT 156.66 40.39 156.87 40.46 ;
    RECT 156.66 40.75 156.87 40.82 ;
    RECT 156.66 41.11 156.87 41.18 ;
    RECT 153.8 40.39 154.01 40.46 ;
    RECT 153.8 40.75 154.01 40.82 ;
    RECT 153.8 41.11 154.01 41.18 ;
    RECT 153.34 40.39 153.55 40.46 ;
    RECT 153.34 40.75 153.55 40.82 ;
    RECT 153.34 41.11 153.55 41.18 ;
    RECT 150.48 40.39 150.69 40.46 ;
    RECT 150.48 40.75 150.69 40.82 ;
    RECT 150.48 41.11 150.69 41.18 ;
    RECT 150.02 40.39 150.23 40.46 ;
    RECT 150.02 40.75 150.23 40.82 ;
    RECT 150.02 41.11 150.23 41.18 ;
    RECT 213.56 40.39 213.77 40.46 ;
    RECT 213.56 40.75 213.77 40.82 ;
    RECT 213.56 41.11 213.77 41.18 ;
    RECT 213.1 40.39 213.31 40.46 ;
    RECT 213.1 40.75 213.31 40.82 ;
    RECT 213.1 41.11 213.31 41.18 ;
    RECT 210.24 40.39 210.45 40.46 ;
    RECT 210.24 40.75 210.45 40.82 ;
    RECT 210.24 41.11 210.45 41.18 ;
    RECT 209.78 40.39 209.99 40.46 ;
    RECT 209.78 40.75 209.99 40.82 ;
    RECT 209.78 41.11 209.99 41.18 ;
    RECT 206.92 40.39 207.13 40.46 ;
    RECT 206.92 40.75 207.13 40.82 ;
    RECT 206.92 41.11 207.13 41.18 ;
    RECT 206.46 40.39 206.67 40.46 ;
    RECT 206.46 40.75 206.67 40.82 ;
    RECT 206.46 41.11 206.67 41.18 ;
    RECT 203.6 40.39 203.81 40.46 ;
    RECT 203.6 40.75 203.81 40.82 ;
    RECT 203.6 41.11 203.81 41.18 ;
    RECT 203.14 40.39 203.35 40.46 ;
    RECT 203.14 40.75 203.35 40.82 ;
    RECT 203.14 41.11 203.35 41.18 ;
    RECT 200.28 40.39 200.49 40.46 ;
    RECT 200.28 40.75 200.49 40.82 ;
    RECT 200.28 41.11 200.49 41.18 ;
    RECT 199.82 40.39 200.03 40.46 ;
    RECT 199.82 40.75 200.03 40.82 ;
    RECT 199.82 41.11 200.03 41.18 ;
    RECT 196.96 40.39 197.17 40.46 ;
    RECT 196.96 40.75 197.17 40.82 ;
    RECT 196.96 41.11 197.17 41.18 ;
    RECT 196.5 40.39 196.71 40.46 ;
    RECT 196.5 40.75 196.71 40.82 ;
    RECT 196.5 41.11 196.71 41.18 ;
    RECT 193.64 40.39 193.85 40.46 ;
    RECT 193.64 40.75 193.85 40.82 ;
    RECT 193.64 41.11 193.85 41.18 ;
    RECT 193.18 40.39 193.39 40.46 ;
    RECT 193.18 40.75 193.39 40.82 ;
    RECT 193.18 41.11 193.39 41.18 ;
    RECT 190.32 40.39 190.53 40.46 ;
    RECT 190.32 40.75 190.53 40.82 ;
    RECT 190.32 41.11 190.53 41.18 ;
    RECT 189.86 40.39 190.07 40.46 ;
    RECT 189.86 40.75 190.07 40.82 ;
    RECT 189.86 41.11 190.07 41.18 ;
    RECT 187.0 40.39 187.21 40.46 ;
    RECT 187.0 40.75 187.21 40.82 ;
    RECT 187.0 41.11 187.21 41.18 ;
    RECT 186.54 40.39 186.75 40.46 ;
    RECT 186.54 40.75 186.75 40.82 ;
    RECT 186.54 41.11 186.75 41.18 ;
    RECT 183.68 40.39 183.89 40.46 ;
    RECT 183.68 40.75 183.89 40.82 ;
    RECT 183.68 41.11 183.89 41.18 ;
    RECT 183.22 40.39 183.43 40.46 ;
    RECT 183.22 40.75 183.43 40.82 ;
    RECT 183.22 41.11 183.43 41.18 ;
    RECT 147.485 40.75 147.555 40.82 ;
    RECT 266.68 40.39 266.89 40.46 ;
    RECT 266.68 40.75 266.89 40.82 ;
    RECT 266.68 41.11 266.89 41.18 ;
    RECT 266.22 40.39 266.43 40.46 ;
    RECT 266.22 40.75 266.43 40.82 ;
    RECT 266.22 41.11 266.43 41.18 ;
    RECT 263.36 40.39 263.57 40.46 ;
    RECT 263.36 40.75 263.57 40.82 ;
    RECT 263.36 41.11 263.57 41.18 ;
    RECT 262.9 40.39 263.11 40.46 ;
    RECT 262.9 40.75 263.11 40.82 ;
    RECT 262.9 41.11 263.11 41.18 ;
    RECT 260.04 40.39 260.25 40.46 ;
    RECT 260.04 40.75 260.25 40.82 ;
    RECT 260.04 41.11 260.25 41.18 ;
    RECT 259.58 40.39 259.79 40.46 ;
    RECT 259.58 40.75 259.79 40.82 ;
    RECT 259.58 41.11 259.79 41.18 ;
    RECT 256.72 40.39 256.93 40.46 ;
    RECT 256.72 40.75 256.93 40.82 ;
    RECT 256.72 41.11 256.93 41.18 ;
    RECT 256.26 40.39 256.47 40.46 ;
    RECT 256.26 40.75 256.47 40.82 ;
    RECT 256.26 41.11 256.47 41.18 ;
    RECT 253.4 40.39 253.61 40.46 ;
    RECT 253.4 40.75 253.61 40.82 ;
    RECT 253.4 41.11 253.61 41.18 ;
    RECT 252.94 40.39 253.15 40.46 ;
    RECT 252.94 40.75 253.15 40.82 ;
    RECT 252.94 41.11 253.15 41.18 ;
    RECT 250.08 39.67 250.29 39.74 ;
    RECT 250.08 40.03 250.29 40.1 ;
    RECT 250.08 40.39 250.29 40.46 ;
    RECT 249.62 39.67 249.83 39.74 ;
    RECT 249.62 40.03 249.83 40.1 ;
    RECT 249.62 40.39 249.83 40.46 ;
    RECT 246.76 39.67 246.97 39.74 ;
    RECT 246.76 40.03 246.97 40.1 ;
    RECT 246.76 40.39 246.97 40.46 ;
    RECT 246.3 39.67 246.51 39.74 ;
    RECT 246.3 40.03 246.51 40.1 ;
    RECT 246.3 40.39 246.51 40.46 ;
    RECT 243.44 39.67 243.65 39.74 ;
    RECT 243.44 40.03 243.65 40.1 ;
    RECT 243.44 40.39 243.65 40.46 ;
    RECT 242.98 39.67 243.19 39.74 ;
    RECT 242.98 40.03 243.19 40.1 ;
    RECT 242.98 40.39 243.19 40.46 ;
    RECT 240.12 39.67 240.33 39.74 ;
    RECT 240.12 40.03 240.33 40.1 ;
    RECT 240.12 40.39 240.33 40.46 ;
    RECT 239.66 39.67 239.87 39.74 ;
    RECT 239.66 40.03 239.87 40.1 ;
    RECT 239.66 40.39 239.87 40.46 ;
    RECT 236.8 39.67 237.01 39.74 ;
    RECT 236.8 40.03 237.01 40.1 ;
    RECT 236.8 40.39 237.01 40.46 ;
    RECT 236.34 39.67 236.55 39.74 ;
    RECT 236.34 40.03 236.55 40.1 ;
    RECT 236.34 40.39 236.55 40.46 ;
    RECT 233.48 39.67 233.69 39.74 ;
    RECT 233.48 40.03 233.69 40.1 ;
    RECT 233.48 40.39 233.69 40.46 ;
    RECT 233.02 39.67 233.23 39.74 ;
    RECT 233.02 40.03 233.23 40.1 ;
    RECT 233.02 40.39 233.23 40.46 ;
    RECT 230.16 39.67 230.37 39.74 ;
    RECT 230.16 40.03 230.37 40.1 ;
    RECT 230.16 40.39 230.37 40.46 ;
    RECT 229.7 39.67 229.91 39.74 ;
    RECT 229.7 40.03 229.91 40.1 ;
    RECT 229.7 40.39 229.91 40.46 ;
    RECT 226.84 39.67 227.05 39.74 ;
    RECT 226.84 40.03 227.05 40.1 ;
    RECT 226.84 40.39 227.05 40.46 ;
    RECT 226.38 39.67 226.59 39.74 ;
    RECT 226.38 40.03 226.59 40.1 ;
    RECT 226.38 40.39 226.59 40.46 ;
    RECT 223.52 39.67 223.73 39.74 ;
    RECT 223.52 40.03 223.73 40.1 ;
    RECT 223.52 40.39 223.73 40.46 ;
    RECT 223.06 39.67 223.27 39.74 ;
    RECT 223.06 40.03 223.27 40.1 ;
    RECT 223.06 40.39 223.27 40.46 ;
    RECT 220.2 39.67 220.41 39.74 ;
    RECT 220.2 40.03 220.41 40.1 ;
    RECT 220.2 40.39 220.41 40.46 ;
    RECT 219.74 39.67 219.95 39.74 ;
    RECT 219.74 40.03 219.95 40.1 ;
    RECT 219.74 40.39 219.95 40.46 ;
    RECT 216.88 39.67 217.09 39.74 ;
    RECT 216.88 40.03 217.09 40.1 ;
    RECT 216.88 40.39 217.09 40.46 ;
    RECT 216.42 39.67 216.63 39.74 ;
    RECT 216.42 40.03 216.63 40.1 ;
    RECT 216.42 40.39 216.63 40.46 ;
    RECT 267.91 40.03 267.98 40.1 ;
    RECT 180.36 39.67 180.57 39.74 ;
    RECT 180.36 40.03 180.57 40.1 ;
    RECT 180.36 40.39 180.57 40.46 ;
    RECT 179.9 39.67 180.11 39.74 ;
    RECT 179.9 40.03 180.11 40.1 ;
    RECT 179.9 40.39 180.11 40.46 ;
    RECT 177.04 39.67 177.25 39.74 ;
    RECT 177.04 40.03 177.25 40.1 ;
    RECT 177.04 40.39 177.25 40.46 ;
    RECT 176.58 39.67 176.79 39.74 ;
    RECT 176.58 40.03 176.79 40.1 ;
    RECT 176.58 40.39 176.79 40.46 ;
    RECT 173.72 39.67 173.93 39.74 ;
    RECT 173.72 40.03 173.93 40.1 ;
    RECT 173.72 40.39 173.93 40.46 ;
    RECT 173.26 39.67 173.47 39.74 ;
    RECT 173.26 40.03 173.47 40.1 ;
    RECT 173.26 40.39 173.47 40.46 ;
    RECT 170.4 39.67 170.61 39.74 ;
    RECT 170.4 40.03 170.61 40.1 ;
    RECT 170.4 40.39 170.61 40.46 ;
    RECT 169.94 39.67 170.15 39.74 ;
    RECT 169.94 40.03 170.15 40.1 ;
    RECT 169.94 40.39 170.15 40.46 ;
    RECT 167.08 39.67 167.29 39.74 ;
    RECT 167.08 40.03 167.29 40.1 ;
    RECT 167.08 40.39 167.29 40.46 ;
    RECT 166.62 39.67 166.83 39.74 ;
    RECT 166.62 40.03 166.83 40.1 ;
    RECT 166.62 40.39 166.83 40.46 ;
    RECT 163.76 39.67 163.97 39.74 ;
    RECT 163.76 40.03 163.97 40.1 ;
    RECT 163.76 40.39 163.97 40.46 ;
    RECT 163.3 39.67 163.51 39.74 ;
    RECT 163.3 40.03 163.51 40.1 ;
    RECT 163.3 40.39 163.51 40.46 ;
    RECT 160.44 39.67 160.65 39.74 ;
    RECT 160.44 40.03 160.65 40.1 ;
    RECT 160.44 40.39 160.65 40.46 ;
    RECT 159.98 39.67 160.19 39.74 ;
    RECT 159.98 40.03 160.19 40.1 ;
    RECT 159.98 40.39 160.19 40.46 ;
    RECT 157.12 39.67 157.33 39.74 ;
    RECT 157.12 40.03 157.33 40.1 ;
    RECT 157.12 40.39 157.33 40.46 ;
    RECT 156.66 39.67 156.87 39.74 ;
    RECT 156.66 40.03 156.87 40.1 ;
    RECT 156.66 40.39 156.87 40.46 ;
    RECT 153.8 39.67 154.01 39.74 ;
    RECT 153.8 40.03 154.01 40.1 ;
    RECT 153.8 40.39 154.01 40.46 ;
    RECT 153.34 39.67 153.55 39.74 ;
    RECT 153.34 40.03 153.55 40.1 ;
    RECT 153.34 40.39 153.55 40.46 ;
    RECT 150.48 39.67 150.69 39.74 ;
    RECT 150.48 40.03 150.69 40.1 ;
    RECT 150.48 40.39 150.69 40.46 ;
    RECT 150.02 39.67 150.23 39.74 ;
    RECT 150.02 40.03 150.23 40.1 ;
    RECT 150.02 40.39 150.23 40.46 ;
    RECT 213.56 39.67 213.77 39.74 ;
    RECT 213.56 40.03 213.77 40.1 ;
    RECT 213.56 40.39 213.77 40.46 ;
    RECT 213.1 39.67 213.31 39.74 ;
    RECT 213.1 40.03 213.31 40.1 ;
    RECT 213.1 40.39 213.31 40.46 ;
    RECT 210.24 39.67 210.45 39.74 ;
    RECT 210.24 40.03 210.45 40.1 ;
    RECT 210.24 40.39 210.45 40.46 ;
    RECT 209.78 39.67 209.99 39.74 ;
    RECT 209.78 40.03 209.99 40.1 ;
    RECT 209.78 40.39 209.99 40.46 ;
    RECT 206.92 39.67 207.13 39.74 ;
    RECT 206.92 40.03 207.13 40.1 ;
    RECT 206.92 40.39 207.13 40.46 ;
    RECT 206.46 39.67 206.67 39.74 ;
    RECT 206.46 40.03 206.67 40.1 ;
    RECT 206.46 40.39 206.67 40.46 ;
    RECT 203.6 39.67 203.81 39.74 ;
    RECT 203.6 40.03 203.81 40.1 ;
    RECT 203.6 40.39 203.81 40.46 ;
    RECT 203.14 39.67 203.35 39.74 ;
    RECT 203.14 40.03 203.35 40.1 ;
    RECT 203.14 40.39 203.35 40.46 ;
    RECT 200.28 39.67 200.49 39.74 ;
    RECT 200.28 40.03 200.49 40.1 ;
    RECT 200.28 40.39 200.49 40.46 ;
    RECT 199.82 39.67 200.03 39.74 ;
    RECT 199.82 40.03 200.03 40.1 ;
    RECT 199.82 40.39 200.03 40.46 ;
    RECT 196.96 39.67 197.17 39.74 ;
    RECT 196.96 40.03 197.17 40.1 ;
    RECT 196.96 40.39 197.17 40.46 ;
    RECT 196.5 39.67 196.71 39.74 ;
    RECT 196.5 40.03 196.71 40.1 ;
    RECT 196.5 40.39 196.71 40.46 ;
    RECT 193.64 39.67 193.85 39.74 ;
    RECT 193.64 40.03 193.85 40.1 ;
    RECT 193.64 40.39 193.85 40.46 ;
    RECT 193.18 39.67 193.39 39.74 ;
    RECT 193.18 40.03 193.39 40.1 ;
    RECT 193.18 40.39 193.39 40.46 ;
    RECT 190.32 39.67 190.53 39.74 ;
    RECT 190.32 40.03 190.53 40.1 ;
    RECT 190.32 40.39 190.53 40.46 ;
    RECT 189.86 39.67 190.07 39.74 ;
    RECT 189.86 40.03 190.07 40.1 ;
    RECT 189.86 40.39 190.07 40.46 ;
    RECT 187.0 39.67 187.21 39.74 ;
    RECT 187.0 40.03 187.21 40.1 ;
    RECT 187.0 40.39 187.21 40.46 ;
    RECT 186.54 39.67 186.75 39.74 ;
    RECT 186.54 40.03 186.75 40.1 ;
    RECT 186.54 40.39 186.75 40.46 ;
    RECT 183.68 39.67 183.89 39.74 ;
    RECT 183.68 40.03 183.89 40.1 ;
    RECT 183.68 40.39 183.89 40.46 ;
    RECT 183.22 39.67 183.43 39.74 ;
    RECT 183.22 40.03 183.43 40.1 ;
    RECT 183.22 40.39 183.43 40.46 ;
    RECT 147.485 40.03 147.555 40.1 ;
    RECT 266.68 39.67 266.89 39.74 ;
    RECT 266.68 40.03 266.89 40.1 ;
    RECT 266.68 40.39 266.89 40.46 ;
    RECT 266.22 39.67 266.43 39.74 ;
    RECT 266.22 40.03 266.43 40.1 ;
    RECT 266.22 40.39 266.43 40.46 ;
    RECT 263.36 39.67 263.57 39.74 ;
    RECT 263.36 40.03 263.57 40.1 ;
    RECT 263.36 40.39 263.57 40.46 ;
    RECT 262.9 39.67 263.11 39.74 ;
    RECT 262.9 40.03 263.11 40.1 ;
    RECT 262.9 40.39 263.11 40.46 ;
    RECT 260.04 39.67 260.25 39.74 ;
    RECT 260.04 40.03 260.25 40.1 ;
    RECT 260.04 40.39 260.25 40.46 ;
    RECT 259.58 39.67 259.79 39.74 ;
    RECT 259.58 40.03 259.79 40.1 ;
    RECT 259.58 40.39 259.79 40.46 ;
    RECT 256.72 39.67 256.93 39.74 ;
    RECT 256.72 40.03 256.93 40.1 ;
    RECT 256.72 40.39 256.93 40.46 ;
    RECT 256.26 39.67 256.47 39.74 ;
    RECT 256.26 40.03 256.47 40.1 ;
    RECT 256.26 40.39 256.47 40.46 ;
    RECT 253.4 39.67 253.61 39.74 ;
    RECT 253.4 40.03 253.61 40.1 ;
    RECT 253.4 40.39 253.61 40.46 ;
    RECT 252.94 39.67 253.15 39.74 ;
    RECT 252.94 40.03 253.15 40.1 ;
    RECT 252.94 40.39 253.15 40.46 ;
    RECT 250.08 79.29 250.29 79.36 ;
    RECT 250.08 79.65 250.29 79.72 ;
    RECT 250.08 80.01 250.29 80.08 ;
    RECT 249.62 79.29 249.83 79.36 ;
    RECT 249.62 79.65 249.83 79.72 ;
    RECT 249.62 80.01 249.83 80.08 ;
    RECT 246.76 79.29 246.97 79.36 ;
    RECT 246.76 79.65 246.97 79.72 ;
    RECT 246.76 80.01 246.97 80.08 ;
    RECT 246.3 79.29 246.51 79.36 ;
    RECT 246.3 79.65 246.51 79.72 ;
    RECT 246.3 80.01 246.51 80.08 ;
    RECT 243.44 79.29 243.65 79.36 ;
    RECT 243.44 79.65 243.65 79.72 ;
    RECT 243.44 80.01 243.65 80.08 ;
    RECT 242.98 79.29 243.19 79.36 ;
    RECT 242.98 79.65 243.19 79.72 ;
    RECT 242.98 80.01 243.19 80.08 ;
    RECT 240.12 79.29 240.33 79.36 ;
    RECT 240.12 79.65 240.33 79.72 ;
    RECT 240.12 80.01 240.33 80.08 ;
    RECT 239.66 79.29 239.87 79.36 ;
    RECT 239.66 79.65 239.87 79.72 ;
    RECT 239.66 80.01 239.87 80.08 ;
    RECT 236.8 79.29 237.01 79.36 ;
    RECT 236.8 79.65 237.01 79.72 ;
    RECT 236.8 80.01 237.01 80.08 ;
    RECT 236.34 79.29 236.55 79.36 ;
    RECT 236.34 79.65 236.55 79.72 ;
    RECT 236.34 80.01 236.55 80.08 ;
    RECT 233.48 79.29 233.69 79.36 ;
    RECT 233.48 79.65 233.69 79.72 ;
    RECT 233.48 80.01 233.69 80.08 ;
    RECT 233.02 79.29 233.23 79.36 ;
    RECT 233.02 79.65 233.23 79.72 ;
    RECT 233.02 80.01 233.23 80.08 ;
    RECT 230.16 79.29 230.37 79.36 ;
    RECT 230.16 79.65 230.37 79.72 ;
    RECT 230.16 80.01 230.37 80.08 ;
    RECT 229.7 79.29 229.91 79.36 ;
    RECT 229.7 79.65 229.91 79.72 ;
    RECT 229.7 80.01 229.91 80.08 ;
    RECT 226.84 79.29 227.05 79.36 ;
    RECT 226.84 79.65 227.05 79.72 ;
    RECT 226.84 80.01 227.05 80.08 ;
    RECT 226.38 79.29 226.59 79.36 ;
    RECT 226.38 79.65 226.59 79.72 ;
    RECT 226.38 80.01 226.59 80.08 ;
    RECT 223.52 79.29 223.73 79.36 ;
    RECT 223.52 79.65 223.73 79.72 ;
    RECT 223.52 80.01 223.73 80.08 ;
    RECT 223.06 79.29 223.27 79.36 ;
    RECT 223.06 79.65 223.27 79.72 ;
    RECT 223.06 80.01 223.27 80.08 ;
    RECT 220.2 79.29 220.41 79.36 ;
    RECT 220.2 79.65 220.41 79.72 ;
    RECT 220.2 80.01 220.41 80.08 ;
    RECT 219.74 79.29 219.95 79.36 ;
    RECT 219.74 79.65 219.95 79.72 ;
    RECT 219.74 80.01 219.95 80.08 ;
    RECT 216.88 79.29 217.09 79.36 ;
    RECT 216.88 79.65 217.09 79.72 ;
    RECT 216.88 80.01 217.09 80.08 ;
    RECT 216.42 79.29 216.63 79.36 ;
    RECT 216.42 79.65 216.63 79.72 ;
    RECT 216.42 80.01 216.63 80.08 ;
    RECT 267.91 79.65 267.98 79.72 ;
    RECT 180.36 79.29 180.57 79.36 ;
    RECT 180.36 79.65 180.57 79.72 ;
    RECT 180.36 80.01 180.57 80.08 ;
    RECT 179.9 79.29 180.11 79.36 ;
    RECT 179.9 79.65 180.11 79.72 ;
    RECT 179.9 80.01 180.11 80.08 ;
    RECT 177.04 79.29 177.25 79.36 ;
    RECT 177.04 79.65 177.25 79.72 ;
    RECT 177.04 80.01 177.25 80.08 ;
    RECT 176.58 79.29 176.79 79.36 ;
    RECT 176.58 79.65 176.79 79.72 ;
    RECT 176.58 80.01 176.79 80.08 ;
    RECT 173.72 79.29 173.93 79.36 ;
    RECT 173.72 79.65 173.93 79.72 ;
    RECT 173.72 80.01 173.93 80.08 ;
    RECT 173.26 79.29 173.47 79.36 ;
    RECT 173.26 79.65 173.47 79.72 ;
    RECT 173.26 80.01 173.47 80.08 ;
    RECT 170.4 79.29 170.61 79.36 ;
    RECT 170.4 79.65 170.61 79.72 ;
    RECT 170.4 80.01 170.61 80.08 ;
    RECT 169.94 79.29 170.15 79.36 ;
    RECT 169.94 79.65 170.15 79.72 ;
    RECT 169.94 80.01 170.15 80.08 ;
    RECT 167.08 79.29 167.29 79.36 ;
    RECT 167.08 79.65 167.29 79.72 ;
    RECT 167.08 80.01 167.29 80.08 ;
    RECT 166.62 79.29 166.83 79.36 ;
    RECT 166.62 79.65 166.83 79.72 ;
    RECT 166.62 80.01 166.83 80.08 ;
    RECT 163.76 79.29 163.97 79.36 ;
    RECT 163.76 79.65 163.97 79.72 ;
    RECT 163.76 80.01 163.97 80.08 ;
    RECT 163.3 79.29 163.51 79.36 ;
    RECT 163.3 79.65 163.51 79.72 ;
    RECT 163.3 80.01 163.51 80.08 ;
    RECT 160.44 79.29 160.65 79.36 ;
    RECT 160.44 79.65 160.65 79.72 ;
    RECT 160.44 80.01 160.65 80.08 ;
    RECT 159.98 79.29 160.19 79.36 ;
    RECT 159.98 79.65 160.19 79.72 ;
    RECT 159.98 80.01 160.19 80.08 ;
    RECT 157.12 79.29 157.33 79.36 ;
    RECT 157.12 79.65 157.33 79.72 ;
    RECT 157.12 80.01 157.33 80.08 ;
    RECT 156.66 79.29 156.87 79.36 ;
    RECT 156.66 79.65 156.87 79.72 ;
    RECT 156.66 80.01 156.87 80.08 ;
    RECT 153.8 79.29 154.01 79.36 ;
    RECT 153.8 79.65 154.01 79.72 ;
    RECT 153.8 80.01 154.01 80.08 ;
    RECT 153.34 79.29 153.55 79.36 ;
    RECT 153.34 79.65 153.55 79.72 ;
    RECT 153.34 80.01 153.55 80.08 ;
    RECT 150.48 79.29 150.69 79.36 ;
    RECT 150.48 79.65 150.69 79.72 ;
    RECT 150.48 80.01 150.69 80.08 ;
    RECT 150.02 79.29 150.23 79.36 ;
    RECT 150.02 79.65 150.23 79.72 ;
    RECT 150.02 80.01 150.23 80.08 ;
    RECT 213.56 79.29 213.77 79.36 ;
    RECT 213.56 79.65 213.77 79.72 ;
    RECT 213.56 80.01 213.77 80.08 ;
    RECT 213.1 79.29 213.31 79.36 ;
    RECT 213.1 79.65 213.31 79.72 ;
    RECT 213.1 80.01 213.31 80.08 ;
    RECT 210.24 79.29 210.45 79.36 ;
    RECT 210.24 79.65 210.45 79.72 ;
    RECT 210.24 80.01 210.45 80.08 ;
    RECT 209.78 79.29 209.99 79.36 ;
    RECT 209.78 79.65 209.99 79.72 ;
    RECT 209.78 80.01 209.99 80.08 ;
    RECT 206.92 79.29 207.13 79.36 ;
    RECT 206.92 79.65 207.13 79.72 ;
    RECT 206.92 80.01 207.13 80.08 ;
    RECT 206.46 79.29 206.67 79.36 ;
    RECT 206.46 79.65 206.67 79.72 ;
    RECT 206.46 80.01 206.67 80.08 ;
    RECT 203.6 79.29 203.81 79.36 ;
    RECT 203.6 79.65 203.81 79.72 ;
    RECT 203.6 80.01 203.81 80.08 ;
    RECT 203.14 79.29 203.35 79.36 ;
    RECT 203.14 79.65 203.35 79.72 ;
    RECT 203.14 80.01 203.35 80.08 ;
    RECT 200.28 79.29 200.49 79.36 ;
    RECT 200.28 79.65 200.49 79.72 ;
    RECT 200.28 80.01 200.49 80.08 ;
    RECT 199.82 79.29 200.03 79.36 ;
    RECT 199.82 79.65 200.03 79.72 ;
    RECT 199.82 80.01 200.03 80.08 ;
    RECT 196.96 79.29 197.17 79.36 ;
    RECT 196.96 79.65 197.17 79.72 ;
    RECT 196.96 80.01 197.17 80.08 ;
    RECT 196.5 79.29 196.71 79.36 ;
    RECT 196.5 79.65 196.71 79.72 ;
    RECT 196.5 80.01 196.71 80.08 ;
    RECT 193.64 79.29 193.85 79.36 ;
    RECT 193.64 79.65 193.85 79.72 ;
    RECT 193.64 80.01 193.85 80.08 ;
    RECT 193.18 79.29 193.39 79.36 ;
    RECT 193.18 79.65 193.39 79.72 ;
    RECT 193.18 80.01 193.39 80.08 ;
    RECT 190.32 79.29 190.53 79.36 ;
    RECT 190.32 79.65 190.53 79.72 ;
    RECT 190.32 80.01 190.53 80.08 ;
    RECT 189.86 79.29 190.07 79.36 ;
    RECT 189.86 79.65 190.07 79.72 ;
    RECT 189.86 80.01 190.07 80.08 ;
    RECT 187.0 79.29 187.21 79.36 ;
    RECT 187.0 79.65 187.21 79.72 ;
    RECT 187.0 80.01 187.21 80.08 ;
    RECT 186.54 79.29 186.75 79.36 ;
    RECT 186.54 79.65 186.75 79.72 ;
    RECT 186.54 80.01 186.75 80.08 ;
    RECT 183.68 79.29 183.89 79.36 ;
    RECT 183.68 79.65 183.89 79.72 ;
    RECT 183.68 80.01 183.89 80.08 ;
    RECT 183.22 79.29 183.43 79.36 ;
    RECT 183.22 79.65 183.43 79.72 ;
    RECT 183.22 80.01 183.43 80.08 ;
    RECT 147.485 79.65 147.555 79.72 ;
    RECT 266.68 79.29 266.89 79.36 ;
    RECT 266.68 79.65 266.89 79.72 ;
    RECT 266.68 80.01 266.89 80.08 ;
    RECT 266.22 79.29 266.43 79.36 ;
    RECT 266.22 79.65 266.43 79.72 ;
    RECT 266.22 80.01 266.43 80.08 ;
    RECT 263.36 79.29 263.57 79.36 ;
    RECT 263.36 79.65 263.57 79.72 ;
    RECT 263.36 80.01 263.57 80.08 ;
    RECT 262.9 79.29 263.11 79.36 ;
    RECT 262.9 79.65 263.11 79.72 ;
    RECT 262.9 80.01 263.11 80.08 ;
    RECT 260.04 79.29 260.25 79.36 ;
    RECT 260.04 79.65 260.25 79.72 ;
    RECT 260.04 80.01 260.25 80.08 ;
    RECT 259.58 79.29 259.79 79.36 ;
    RECT 259.58 79.65 259.79 79.72 ;
    RECT 259.58 80.01 259.79 80.08 ;
    RECT 256.72 79.29 256.93 79.36 ;
    RECT 256.72 79.65 256.93 79.72 ;
    RECT 256.72 80.01 256.93 80.08 ;
    RECT 256.26 79.29 256.47 79.36 ;
    RECT 256.26 79.65 256.47 79.72 ;
    RECT 256.26 80.01 256.47 80.08 ;
    RECT 253.4 79.29 253.61 79.36 ;
    RECT 253.4 79.65 253.61 79.72 ;
    RECT 253.4 80.01 253.61 80.08 ;
    RECT 252.94 79.29 253.15 79.36 ;
    RECT 252.94 79.65 253.15 79.72 ;
    RECT 252.94 80.01 253.15 80.08 ;
    RECT 250.08 38.95 250.29 39.02 ;
    RECT 250.08 39.31 250.29 39.38 ;
    RECT 250.08 39.67 250.29 39.74 ;
    RECT 249.62 38.95 249.83 39.02 ;
    RECT 249.62 39.31 249.83 39.38 ;
    RECT 249.62 39.67 249.83 39.74 ;
    RECT 246.76 38.95 246.97 39.02 ;
    RECT 246.76 39.31 246.97 39.38 ;
    RECT 246.76 39.67 246.97 39.74 ;
    RECT 246.3 38.95 246.51 39.02 ;
    RECT 246.3 39.31 246.51 39.38 ;
    RECT 246.3 39.67 246.51 39.74 ;
    RECT 243.44 38.95 243.65 39.02 ;
    RECT 243.44 39.31 243.65 39.38 ;
    RECT 243.44 39.67 243.65 39.74 ;
    RECT 242.98 38.95 243.19 39.02 ;
    RECT 242.98 39.31 243.19 39.38 ;
    RECT 242.98 39.67 243.19 39.74 ;
    RECT 240.12 38.95 240.33 39.02 ;
    RECT 240.12 39.31 240.33 39.38 ;
    RECT 240.12 39.67 240.33 39.74 ;
    RECT 239.66 38.95 239.87 39.02 ;
    RECT 239.66 39.31 239.87 39.38 ;
    RECT 239.66 39.67 239.87 39.74 ;
    RECT 236.8 38.95 237.01 39.02 ;
    RECT 236.8 39.31 237.01 39.38 ;
    RECT 236.8 39.67 237.01 39.74 ;
    RECT 236.34 38.95 236.55 39.02 ;
    RECT 236.34 39.31 236.55 39.38 ;
    RECT 236.34 39.67 236.55 39.74 ;
    RECT 233.48 38.95 233.69 39.02 ;
    RECT 233.48 39.31 233.69 39.38 ;
    RECT 233.48 39.67 233.69 39.74 ;
    RECT 233.02 38.95 233.23 39.02 ;
    RECT 233.02 39.31 233.23 39.38 ;
    RECT 233.02 39.67 233.23 39.74 ;
    RECT 230.16 38.95 230.37 39.02 ;
    RECT 230.16 39.31 230.37 39.38 ;
    RECT 230.16 39.67 230.37 39.74 ;
    RECT 229.7 38.95 229.91 39.02 ;
    RECT 229.7 39.31 229.91 39.38 ;
    RECT 229.7 39.67 229.91 39.74 ;
    RECT 226.84 38.95 227.05 39.02 ;
    RECT 226.84 39.31 227.05 39.38 ;
    RECT 226.84 39.67 227.05 39.74 ;
    RECT 226.38 38.95 226.59 39.02 ;
    RECT 226.38 39.31 226.59 39.38 ;
    RECT 226.38 39.67 226.59 39.74 ;
    RECT 223.52 38.95 223.73 39.02 ;
    RECT 223.52 39.31 223.73 39.38 ;
    RECT 223.52 39.67 223.73 39.74 ;
    RECT 223.06 38.95 223.27 39.02 ;
    RECT 223.06 39.31 223.27 39.38 ;
    RECT 223.06 39.67 223.27 39.74 ;
    RECT 220.2 38.95 220.41 39.02 ;
    RECT 220.2 39.31 220.41 39.38 ;
    RECT 220.2 39.67 220.41 39.74 ;
    RECT 219.74 38.95 219.95 39.02 ;
    RECT 219.74 39.31 219.95 39.38 ;
    RECT 219.74 39.67 219.95 39.74 ;
    RECT 216.88 38.95 217.09 39.02 ;
    RECT 216.88 39.31 217.09 39.38 ;
    RECT 216.88 39.67 217.09 39.74 ;
    RECT 216.42 38.95 216.63 39.02 ;
    RECT 216.42 39.31 216.63 39.38 ;
    RECT 216.42 39.67 216.63 39.74 ;
    RECT 267.91 39.31 267.98 39.38 ;
    RECT 180.36 38.95 180.57 39.02 ;
    RECT 180.36 39.31 180.57 39.38 ;
    RECT 180.36 39.67 180.57 39.74 ;
    RECT 179.9 38.95 180.11 39.02 ;
    RECT 179.9 39.31 180.11 39.38 ;
    RECT 179.9 39.67 180.11 39.74 ;
    RECT 177.04 38.95 177.25 39.02 ;
    RECT 177.04 39.31 177.25 39.38 ;
    RECT 177.04 39.67 177.25 39.74 ;
    RECT 176.58 38.95 176.79 39.02 ;
    RECT 176.58 39.31 176.79 39.38 ;
    RECT 176.58 39.67 176.79 39.74 ;
    RECT 173.72 38.95 173.93 39.02 ;
    RECT 173.72 39.31 173.93 39.38 ;
    RECT 173.72 39.67 173.93 39.74 ;
    RECT 173.26 38.95 173.47 39.02 ;
    RECT 173.26 39.31 173.47 39.38 ;
    RECT 173.26 39.67 173.47 39.74 ;
    RECT 170.4 38.95 170.61 39.02 ;
    RECT 170.4 39.31 170.61 39.38 ;
    RECT 170.4 39.67 170.61 39.74 ;
    RECT 169.94 38.95 170.15 39.02 ;
    RECT 169.94 39.31 170.15 39.38 ;
    RECT 169.94 39.67 170.15 39.74 ;
    RECT 167.08 38.95 167.29 39.02 ;
    RECT 167.08 39.31 167.29 39.38 ;
    RECT 167.08 39.67 167.29 39.74 ;
    RECT 166.62 38.95 166.83 39.02 ;
    RECT 166.62 39.31 166.83 39.38 ;
    RECT 166.62 39.67 166.83 39.74 ;
    RECT 163.76 38.95 163.97 39.02 ;
    RECT 163.76 39.31 163.97 39.38 ;
    RECT 163.76 39.67 163.97 39.74 ;
    RECT 163.3 38.95 163.51 39.02 ;
    RECT 163.3 39.31 163.51 39.38 ;
    RECT 163.3 39.67 163.51 39.74 ;
    RECT 160.44 38.95 160.65 39.02 ;
    RECT 160.44 39.31 160.65 39.38 ;
    RECT 160.44 39.67 160.65 39.74 ;
    RECT 159.98 38.95 160.19 39.02 ;
    RECT 159.98 39.31 160.19 39.38 ;
    RECT 159.98 39.67 160.19 39.74 ;
    RECT 157.12 38.95 157.33 39.02 ;
    RECT 157.12 39.31 157.33 39.38 ;
    RECT 157.12 39.67 157.33 39.74 ;
    RECT 156.66 38.95 156.87 39.02 ;
    RECT 156.66 39.31 156.87 39.38 ;
    RECT 156.66 39.67 156.87 39.74 ;
    RECT 153.8 38.95 154.01 39.02 ;
    RECT 153.8 39.31 154.01 39.38 ;
    RECT 153.8 39.67 154.01 39.74 ;
    RECT 153.34 38.95 153.55 39.02 ;
    RECT 153.34 39.31 153.55 39.38 ;
    RECT 153.34 39.67 153.55 39.74 ;
    RECT 150.48 38.95 150.69 39.02 ;
    RECT 150.48 39.31 150.69 39.38 ;
    RECT 150.48 39.67 150.69 39.74 ;
    RECT 150.02 38.95 150.23 39.02 ;
    RECT 150.02 39.31 150.23 39.38 ;
    RECT 150.02 39.67 150.23 39.74 ;
    RECT 213.56 38.95 213.77 39.02 ;
    RECT 213.56 39.31 213.77 39.38 ;
    RECT 213.56 39.67 213.77 39.74 ;
    RECT 213.1 38.95 213.31 39.02 ;
    RECT 213.1 39.31 213.31 39.38 ;
    RECT 213.1 39.67 213.31 39.74 ;
    RECT 210.24 38.95 210.45 39.02 ;
    RECT 210.24 39.31 210.45 39.38 ;
    RECT 210.24 39.67 210.45 39.74 ;
    RECT 209.78 38.95 209.99 39.02 ;
    RECT 209.78 39.31 209.99 39.38 ;
    RECT 209.78 39.67 209.99 39.74 ;
    RECT 206.92 38.95 207.13 39.02 ;
    RECT 206.92 39.31 207.13 39.38 ;
    RECT 206.92 39.67 207.13 39.74 ;
    RECT 206.46 38.95 206.67 39.02 ;
    RECT 206.46 39.31 206.67 39.38 ;
    RECT 206.46 39.67 206.67 39.74 ;
    RECT 203.6 38.95 203.81 39.02 ;
    RECT 203.6 39.31 203.81 39.38 ;
    RECT 203.6 39.67 203.81 39.74 ;
    RECT 203.14 38.95 203.35 39.02 ;
    RECT 203.14 39.31 203.35 39.38 ;
    RECT 203.14 39.67 203.35 39.74 ;
    RECT 200.28 38.95 200.49 39.02 ;
    RECT 200.28 39.31 200.49 39.38 ;
    RECT 200.28 39.67 200.49 39.74 ;
    RECT 199.82 38.95 200.03 39.02 ;
    RECT 199.82 39.31 200.03 39.38 ;
    RECT 199.82 39.67 200.03 39.74 ;
    RECT 196.96 38.95 197.17 39.02 ;
    RECT 196.96 39.31 197.17 39.38 ;
    RECT 196.96 39.67 197.17 39.74 ;
    RECT 196.5 38.95 196.71 39.02 ;
    RECT 196.5 39.31 196.71 39.38 ;
    RECT 196.5 39.67 196.71 39.74 ;
    RECT 193.64 38.95 193.85 39.02 ;
    RECT 193.64 39.31 193.85 39.38 ;
    RECT 193.64 39.67 193.85 39.74 ;
    RECT 193.18 38.95 193.39 39.02 ;
    RECT 193.18 39.31 193.39 39.38 ;
    RECT 193.18 39.67 193.39 39.74 ;
    RECT 190.32 38.95 190.53 39.02 ;
    RECT 190.32 39.31 190.53 39.38 ;
    RECT 190.32 39.67 190.53 39.74 ;
    RECT 189.86 38.95 190.07 39.02 ;
    RECT 189.86 39.31 190.07 39.38 ;
    RECT 189.86 39.67 190.07 39.74 ;
    RECT 187.0 38.95 187.21 39.02 ;
    RECT 187.0 39.31 187.21 39.38 ;
    RECT 187.0 39.67 187.21 39.74 ;
    RECT 186.54 38.95 186.75 39.02 ;
    RECT 186.54 39.31 186.75 39.38 ;
    RECT 186.54 39.67 186.75 39.74 ;
    RECT 183.68 38.95 183.89 39.02 ;
    RECT 183.68 39.31 183.89 39.38 ;
    RECT 183.68 39.67 183.89 39.74 ;
    RECT 183.22 38.95 183.43 39.02 ;
    RECT 183.22 39.31 183.43 39.38 ;
    RECT 183.22 39.67 183.43 39.74 ;
    RECT 147.485 39.31 147.555 39.38 ;
    RECT 266.68 38.95 266.89 39.02 ;
    RECT 266.68 39.31 266.89 39.38 ;
    RECT 266.68 39.67 266.89 39.74 ;
    RECT 266.22 38.95 266.43 39.02 ;
    RECT 266.22 39.31 266.43 39.38 ;
    RECT 266.22 39.67 266.43 39.74 ;
    RECT 263.36 38.95 263.57 39.02 ;
    RECT 263.36 39.31 263.57 39.38 ;
    RECT 263.36 39.67 263.57 39.74 ;
    RECT 262.9 38.95 263.11 39.02 ;
    RECT 262.9 39.31 263.11 39.38 ;
    RECT 262.9 39.67 263.11 39.74 ;
    RECT 260.04 38.95 260.25 39.02 ;
    RECT 260.04 39.31 260.25 39.38 ;
    RECT 260.04 39.67 260.25 39.74 ;
    RECT 259.58 38.95 259.79 39.02 ;
    RECT 259.58 39.31 259.79 39.38 ;
    RECT 259.58 39.67 259.79 39.74 ;
    RECT 256.72 38.95 256.93 39.02 ;
    RECT 256.72 39.31 256.93 39.38 ;
    RECT 256.72 39.67 256.93 39.74 ;
    RECT 256.26 38.95 256.47 39.02 ;
    RECT 256.26 39.31 256.47 39.38 ;
    RECT 256.26 39.67 256.47 39.74 ;
    RECT 253.4 38.95 253.61 39.02 ;
    RECT 253.4 39.31 253.61 39.38 ;
    RECT 253.4 39.67 253.61 39.74 ;
    RECT 252.94 38.95 253.15 39.02 ;
    RECT 252.94 39.31 253.15 39.38 ;
    RECT 252.94 39.67 253.15 39.74 ;
    RECT 250.08 78.57 250.29 78.64 ;
    RECT 250.08 78.93 250.29 79.0 ;
    RECT 250.08 79.29 250.29 79.36 ;
    RECT 249.62 78.57 249.83 78.64 ;
    RECT 249.62 78.93 249.83 79.0 ;
    RECT 249.62 79.29 249.83 79.36 ;
    RECT 246.76 78.57 246.97 78.64 ;
    RECT 246.76 78.93 246.97 79.0 ;
    RECT 246.76 79.29 246.97 79.36 ;
    RECT 246.3 78.57 246.51 78.64 ;
    RECT 246.3 78.93 246.51 79.0 ;
    RECT 246.3 79.29 246.51 79.36 ;
    RECT 243.44 78.57 243.65 78.64 ;
    RECT 243.44 78.93 243.65 79.0 ;
    RECT 243.44 79.29 243.65 79.36 ;
    RECT 242.98 78.57 243.19 78.64 ;
    RECT 242.98 78.93 243.19 79.0 ;
    RECT 242.98 79.29 243.19 79.36 ;
    RECT 240.12 78.57 240.33 78.64 ;
    RECT 240.12 78.93 240.33 79.0 ;
    RECT 240.12 79.29 240.33 79.36 ;
    RECT 239.66 78.57 239.87 78.64 ;
    RECT 239.66 78.93 239.87 79.0 ;
    RECT 239.66 79.29 239.87 79.36 ;
    RECT 236.8 78.57 237.01 78.64 ;
    RECT 236.8 78.93 237.01 79.0 ;
    RECT 236.8 79.29 237.01 79.36 ;
    RECT 236.34 78.57 236.55 78.64 ;
    RECT 236.34 78.93 236.55 79.0 ;
    RECT 236.34 79.29 236.55 79.36 ;
    RECT 233.48 78.57 233.69 78.64 ;
    RECT 233.48 78.93 233.69 79.0 ;
    RECT 233.48 79.29 233.69 79.36 ;
    RECT 233.02 78.57 233.23 78.64 ;
    RECT 233.02 78.93 233.23 79.0 ;
    RECT 233.02 79.29 233.23 79.36 ;
    RECT 230.16 78.57 230.37 78.64 ;
    RECT 230.16 78.93 230.37 79.0 ;
    RECT 230.16 79.29 230.37 79.36 ;
    RECT 229.7 78.57 229.91 78.64 ;
    RECT 229.7 78.93 229.91 79.0 ;
    RECT 229.7 79.29 229.91 79.36 ;
    RECT 226.84 78.57 227.05 78.64 ;
    RECT 226.84 78.93 227.05 79.0 ;
    RECT 226.84 79.29 227.05 79.36 ;
    RECT 226.38 78.57 226.59 78.64 ;
    RECT 226.38 78.93 226.59 79.0 ;
    RECT 226.38 79.29 226.59 79.36 ;
    RECT 223.52 78.57 223.73 78.64 ;
    RECT 223.52 78.93 223.73 79.0 ;
    RECT 223.52 79.29 223.73 79.36 ;
    RECT 223.06 78.57 223.27 78.64 ;
    RECT 223.06 78.93 223.27 79.0 ;
    RECT 223.06 79.29 223.27 79.36 ;
    RECT 220.2 78.57 220.41 78.64 ;
    RECT 220.2 78.93 220.41 79.0 ;
    RECT 220.2 79.29 220.41 79.36 ;
    RECT 219.74 78.57 219.95 78.64 ;
    RECT 219.74 78.93 219.95 79.0 ;
    RECT 219.74 79.29 219.95 79.36 ;
    RECT 216.88 78.57 217.09 78.64 ;
    RECT 216.88 78.93 217.09 79.0 ;
    RECT 216.88 79.29 217.09 79.36 ;
    RECT 216.42 78.57 216.63 78.64 ;
    RECT 216.42 78.93 216.63 79.0 ;
    RECT 216.42 79.29 216.63 79.36 ;
    RECT 267.91 78.93 267.98 79.0 ;
    RECT 180.36 78.57 180.57 78.64 ;
    RECT 180.36 78.93 180.57 79.0 ;
    RECT 180.36 79.29 180.57 79.36 ;
    RECT 179.9 78.57 180.11 78.64 ;
    RECT 179.9 78.93 180.11 79.0 ;
    RECT 179.9 79.29 180.11 79.36 ;
    RECT 177.04 78.57 177.25 78.64 ;
    RECT 177.04 78.93 177.25 79.0 ;
    RECT 177.04 79.29 177.25 79.36 ;
    RECT 176.58 78.57 176.79 78.64 ;
    RECT 176.58 78.93 176.79 79.0 ;
    RECT 176.58 79.29 176.79 79.36 ;
    RECT 173.72 78.57 173.93 78.64 ;
    RECT 173.72 78.93 173.93 79.0 ;
    RECT 173.72 79.29 173.93 79.36 ;
    RECT 173.26 78.57 173.47 78.64 ;
    RECT 173.26 78.93 173.47 79.0 ;
    RECT 173.26 79.29 173.47 79.36 ;
    RECT 170.4 78.57 170.61 78.64 ;
    RECT 170.4 78.93 170.61 79.0 ;
    RECT 170.4 79.29 170.61 79.36 ;
    RECT 169.94 78.57 170.15 78.64 ;
    RECT 169.94 78.93 170.15 79.0 ;
    RECT 169.94 79.29 170.15 79.36 ;
    RECT 167.08 78.57 167.29 78.64 ;
    RECT 167.08 78.93 167.29 79.0 ;
    RECT 167.08 79.29 167.29 79.36 ;
    RECT 166.62 78.57 166.83 78.64 ;
    RECT 166.62 78.93 166.83 79.0 ;
    RECT 166.62 79.29 166.83 79.36 ;
    RECT 163.76 78.57 163.97 78.64 ;
    RECT 163.76 78.93 163.97 79.0 ;
    RECT 163.76 79.29 163.97 79.36 ;
    RECT 163.3 78.57 163.51 78.64 ;
    RECT 163.3 78.93 163.51 79.0 ;
    RECT 163.3 79.29 163.51 79.36 ;
    RECT 160.44 78.57 160.65 78.64 ;
    RECT 160.44 78.93 160.65 79.0 ;
    RECT 160.44 79.29 160.65 79.36 ;
    RECT 159.98 78.57 160.19 78.64 ;
    RECT 159.98 78.93 160.19 79.0 ;
    RECT 159.98 79.29 160.19 79.36 ;
    RECT 157.12 78.57 157.33 78.64 ;
    RECT 157.12 78.93 157.33 79.0 ;
    RECT 157.12 79.29 157.33 79.36 ;
    RECT 156.66 78.57 156.87 78.64 ;
    RECT 156.66 78.93 156.87 79.0 ;
    RECT 156.66 79.29 156.87 79.36 ;
    RECT 153.8 78.57 154.01 78.64 ;
    RECT 153.8 78.93 154.01 79.0 ;
    RECT 153.8 79.29 154.01 79.36 ;
    RECT 153.34 78.57 153.55 78.64 ;
    RECT 153.34 78.93 153.55 79.0 ;
    RECT 153.34 79.29 153.55 79.36 ;
    RECT 150.48 78.57 150.69 78.64 ;
    RECT 150.48 78.93 150.69 79.0 ;
    RECT 150.48 79.29 150.69 79.36 ;
    RECT 150.02 78.57 150.23 78.64 ;
    RECT 150.02 78.93 150.23 79.0 ;
    RECT 150.02 79.29 150.23 79.36 ;
    RECT 213.56 78.57 213.77 78.64 ;
    RECT 213.56 78.93 213.77 79.0 ;
    RECT 213.56 79.29 213.77 79.36 ;
    RECT 213.1 78.57 213.31 78.64 ;
    RECT 213.1 78.93 213.31 79.0 ;
    RECT 213.1 79.29 213.31 79.36 ;
    RECT 210.24 78.57 210.45 78.64 ;
    RECT 210.24 78.93 210.45 79.0 ;
    RECT 210.24 79.29 210.45 79.36 ;
    RECT 209.78 78.57 209.99 78.64 ;
    RECT 209.78 78.93 209.99 79.0 ;
    RECT 209.78 79.29 209.99 79.36 ;
    RECT 206.92 78.57 207.13 78.64 ;
    RECT 206.92 78.93 207.13 79.0 ;
    RECT 206.92 79.29 207.13 79.36 ;
    RECT 206.46 78.57 206.67 78.64 ;
    RECT 206.46 78.93 206.67 79.0 ;
    RECT 206.46 79.29 206.67 79.36 ;
    RECT 203.6 78.57 203.81 78.64 ;
    RECT 203.6 78.93 203.81 79.0 ;
    RECT 203.6 79.29 203.81 79.36 ;
    RECT 203.14 78.57 203.35 78.64 ;
    RECT 203.14 78.93 203.35 79.0 ;
    RECT 203.14 79.29 203.35 79.36 ;
    RECT 200.28 78.57 200.49 78.64 ;
    RECT 200.28 78.93 200.49 79.0 ;
    RECT 200.28 79.29 200.49 79.36 ;
    RECT 199.82 78.57 200.03 78.64 ;
    RECT 199.82 78.93 200.03 79.0 ;
    RECT 199.82 79.29 200.03 79.36 ;
    RECT 196.96 78.57 197.17 78.64 ;
    RECT 196.96 78.93 197.17 79.0 ;
    RECT 196.96 79.29 197.17 79.36 ;
    RECT 196.5 78.57 196.71 78.64 ;
    RECT 196.5 78.93 196.71 79.0 ;
    RECT 196.5 79.29 196.71 79.36 ;
    RECT 193.64 78.57 193.85 78.64 ;
    RECT 193.64 78.93 193.85 79.0 ;
    RECT 193.64 79.29 193.85 79.36 ;
    RECT 193.18 78.57 193.39 78.64 ;
    RECT 193.18 78.93 193.39 79.0 ;
    RECT 193.18 79.29 193.39 79.36 ;
    RECT 190.32 78.57 190.53 78.64 ;
    RECT 190.32 78.93 190.53 79.0 ;
    RECT 190.32 79.29 190.53 79.36 ;
    RECT 189.86 78.57 190.07 78.64 ;
    RECT 189.86 78.93 190.07 79.0 ;
    RECT 189.86 79.29 190.07 79.36 ;
    RECT 187.0 78.57 187.21 78.64 ;
    RECT 187.0 78.93 187.21 79.0 ;
    RECT 187.0 79.29 187.21 79.36 ;
    RECT 186.54 78.57 186.75 78.64 ;
    RECT 186.54 78.93 186.75 79.0 ;
    RECT 186.54 79.29 186.75 79.36 ;
    RECT 183.68 78.57 183.89 78.64 ;
    RECT 183.68 78.93 183.89 79.0 ;
    RECT 183.68 79.29 183.89 79.36 ;
    RECT 183.22 78.57 183.43 78.64 ;
    RECT 183.22 78.93 183.43 79.0 ;
    RECT 183.22 79.29 183.43 79.36 ;
    RECT 147.485 78.93 147.555 79.0 ;
    RECT 266.68 78.57 266.89 78.64 ;
    RECT 266.68 78.93 266.89 79.0 ;
    RECT 266.68 79.29 266.89 79.36 ;
    RECT 266.22 78.57 266.43 78.64 ;
    RECT 266.22 78.93 266.43 79.0 ;
    RECT 266.22 79.29 266.43 79.36 ;
    RECT 263.36 78.57 263.57 78.64 ;
    RECT 263.36 78.93 263.57 79.0 ;
    RECT 263.36 79.29 263.57 79.36 ;
    RECT 262.9 78.57 263.11 78.64 ;
    RECT 262.9 78.93 263.11 79.0 ;
    RECT 262.9 79.29 263.11 79.36 ;
    RECT 260.04 78.57 260.25 78.64 ;
    RECT 260.04 78.93 260.25 79.0 ;
    RECT 260.04 79.29 260.25 79.36 ;
    RECT 259.58 78.57 259.79 78.64 ;
    RECT 259.58 78.93 259.79 79.0 ;
    RECT 259.58 79.29 259.79 79.36 ;
    RECT 256.72 78.57 256.93 78.64 ;
    RECT 256.72 78.93 256.93 79.0 ;
    RECT 256.72 79.29 256.93 79.36 ;
    RECT 256.26 78.57 256.47 78.64 ;
    RECT 256.26 78.93 256.47 79.0 ;
    RECT 256.26 79.29 256.47 79.36 ;
    RECT 253.4 78.57 253.61 78.64 ;
    RECT 253.4 78.93 253.61 79.0 ;
    RECT 253.4 79.29 253.61 79.36 ;
    RECT 252.94 78.57 253.15 78.64 ;
    RECT 252.94 78.93 253.15 79.0 ;
    RECT 252.94 79.29 253.15 79.36 ;
    RECT 250.08 38.23 250.29 38.3 ;
    RECT 250.08 38.59 250.29 38.66 ;
    RECT 250.08 38.95 250.29 39.02 ;
    RECT 249.62 38.23 249.83 38.3 ;
    RECT 249.62 38.59 249.83 38.66 ;
    RECT 249.62 38.95 249.83 39.02 ;
    RECT 246.76 38.23 246.97 38.3 ;
    RECT 246.76 38.59 246.97 38.66 ;
    RECT 246.76 38.95 246.97 39.02 ;
    RECT 246.3 38.23 246.51 38.3 ;
    RECT 246.3 38.59 246.51 38.66 ;
    RECT 246.3 38.95 246.51 39.02 ;
    RECT 243.44 38.23 243.65 38.3 ;
    RECT 243.44 38.59 243.65 38.66 ;
    RECT 243.44 38.95 243.65 39.02 ;
    RECT 242.98 38.23 243.19 38.3 ;
    RECT 242.98 38.59 243.19 38.66 ;
    RECT 242.98 38.95 243.19 39.02 ;
    RECT 240.12 38.23 240.33 38.3 ;
    RECT 240.12 38.59 240.33 38.66 ;
    RECT 240.12 38.95 240.33 39.02 ;
    RECT 239.66 38.23 239.87 38.3 ;
    RECT 239.66 38.59 239.87 38.66 ;
    RECT 239.66 38.95 239.87 39.02 ;
    RECT 236.8 38.23 237.01 38.3 ;
    RECT 236.8 38.59 237.01 38.66 ;
    RECT 236.8 38.95 237.01 39.02 ;
    RECT 236.34 38.23 236.55 38.3 ;
    RECT 236.34 38.59 236.55 38.66 ;
    RECT 236.34 38.95 236.55 39.02 ;
    RECT 233.48 38.23 233.69 38.3 ;
    RECT 233.48 38.59 233.69 38.66 ;
    RECT 233.48 38.95 233.69 39.02 ;
    RECT 233.02 38.23 233.23 38.3 ;
    RECT 233.02 38.59 233.23 38.66 ;
    RECT 233.02 38.95 233.23 39.02 ;
    RECT 230.16 38.23 230.37 38.3 ;
    RECT 230.16 38.59 230.37 38.66 ;
    RECT 230.16 38.95 230.37 39.02 ;
    RECT 229.7 38.23 229.91 38.3 ;
    RECT 229.7 38.59 229.91 38.66 ;
    RECT 229.7 38.95 229.91 39.02 ;
    RECT 226.84 38.23 227.05 38.3 ;
    RECT 226.84 38.59 227.05 38.66 ;
    RECT 226.84 38.95 227.05 39.02 ;
    RECT 226.38 38.23 226.59 38.3 ;
    RECT 226.38 38.59 226.59 38.66 ;
    RECT 226.38 38.95 226.59 39.02 ;
    RECT 223.52 38.23 223.73 38.3 ;
    RECT 223.52 38.59 223.73 38.66 ;
    RECT 223.52 38.95 223.73 39.02 ;
    RECT 223.06 38.23 223.27 38.3 ;
    RECT 223.06 38.59 223.27 38.66 ;
    RECT 223.06 38.95 223.27 39.02 ;
    RECT 220.2 38.23 220.41 38.3 ;
    RECT 220.2 38.59 220.41 38.66 ;
    RECT 220.2 38.95 220.41 39.02 ;
    RECT 219.74 38.23 219.95 38.3 ;
    RECT 219.74 38.59 219.95 38.66 ;
    RECT 219.74 38.95 219.95 39.02 ;
    RECT 216.88 38.23 217.09 38.3 ;
    RECT 216.88 38.59 217.09 38.66 ;
    RECT 216.88 38.95 217.09 39.02 ;
    RECT 216.42 38.23 216.63 38.3 ;
    RECT 216.42 38.59 216.63 38.66 ;
    RECT 216.42 38.95 216.63 39.02 ;
    RECT 267.91 38.59 267.98 38.66 ;
    RECT 180.36 38.23 180.57 38.3 ;
    RECT 180.36 38.59 180.57 38.66 ;
    RECT 180.36 38.95 180.57 39.02 ;
    RECT 179.9 38.23 180.11 38.3 ;
    RECT 179.9 38.59 180.11 38.66 ;
    RECT 179.9 38.95 180.11 39.02 ;
    RECT 177.04 38.23 177.25 38.3 ;
    RECT 177.04 38.59 177.25 38.66 ;
    RECT 177.04 38.95 177.25 39.02 ;
    RECT 176.58 38.23 176.79 38.3 ;
    RECT 176.58 38.59 176.79 38.66 ;
    RECT 176.58 38.95 176.79 39.02 ;
    RECT 173.72 38.23 173.93 38.3 ;
    RECT 173.72 38.59 173.93 38.66 ;
    RECT 173.72 38.95 173.93 39.02 ;
    RECT 173.26 38.23 173.47 38.3 ;
    RECT 173.26 38.59 173.47 38.66 ;
    RECT 173.26 38.95 173.47 39.02 ;
    RECT 170.4 38.23 170.61 38.3 ;
    RECT 170.4 38.59 170.61 38.66 ;
    RECT 170.4 38.95 170.61 39.02 ;
    RECT 169.94 38.23 170.15 38.3 ;
    RECT 169.94 38.59 170.15 38.66 ;
    RECT 169.94 38.95 170.15 39.02 ;
    RECT 167.08 38.23 167.29 38.3 ;
    RECT 167.08 38.59 167.29 38.66 ;
    RECT 167.08 38.95 167.29 39.02 ;
    RECT 166.62 38.23 166.83 38.3 ;
    RECT 166.62 38.59 166.83 38.66 ;
    RECT 166.62 38.95 166.83 39.02 ;
    RECT 163.76 38.23 163.97 38.3 ;
    RECT 163.76 38.59 163.97 38.66 ;
    RECT 163.76 38.95 163.97 39.02 ;
    RECT 163.3 38.23 163.51 38.3 ;
    RECT 163.3 38.59 163.51 38.66 ;
    RECT 163.3 38.95 163.51 39.02 ;
    RECT 160.44 38.23 160.65 38.3 ;
    RECT 160.44 38.59 160.65 38.66 ;
    RECT 160.44 38.95 160.65 39.02 ;
    RECT 159.98 38.23 160.19 38.3 ;
    RECT 159.98 38.59 160.19 38.66 ;
    RECT 159.98 38.95 160.19 39.02 ;
    RECT 157.12 38.23 157.33 38.3 ;
    RECT 157.12 38.59 157.33 38.66 ;
    RECT 157.12 38.95 157.33 39.02 ;
    RECT 156.66 38.23 156.87 38.3 ;
    RECT 156.66 38.59 156.87 38.66 ;
    RECT 156.66 38.95 156.87 39.02 ;
    RECT 153.8 38.23 154.01 38.3 ;
    RECT 153.8 38.59 154.01 38.66 ;
    RECT 153.8 38.95 154.01 39.02 ;
    RECT 153.34 38.23 153.55 38.3 ;
    RECT 153.34 38.59 153.55 38.66 ;
    RECT 153.34 38.95 153.55 39.02 ;
    RECT 150.48 38.23 150.69 38.3 ;
    RECT 150.48 38.59 150.69 38.66 ;
    RECT 150.48 38.95 150.69 39.02 ;
    RECT 150.02 38.23 150.23 38.3 ;
    RECT 150.02 38.59 150.23 38.66 ;
    RECT 150.02 38.95 150.23 39.02 ;
    RECT 213.56 38.23 213.77 38.3 ;
    RECT 213.56 38.59 213.77 38.66 ;
    RECT 213.56 38.95 213.77 39.02 ;
    RECT 213.1 38.23 213.31 38.3 ;
    RECT 213.1 38.59 213.31 38.66 ;
    RECT 213.1 38.95 213.31 39.02 ;
    RECT 210.24 38.23 210.45 38.3 ;
    RECT 210.24 38.59 210.45 38.66 ;
    RECT 210.24 38.95 210.45 39.02 ;
    RECT 209.78 38.23 209.99 38.3 ;
    RECT 209.78 38.59 209.99 38.66 ;
    RECT 209.78 38.95 209.99 39.02 ;
    RECT 206.92 38.23 207.13 38.3 ;
    RECT 206.92 38.59 207.13 38.66 ;
    RECT 206.92 38.95 207.13 39.02 ;
    RECT 206.46 38.23 206.67 38.3 ;
    RECT 206.46 38.59 206.67 38.66 ;
    RECT 206.46 38.95 206.67 39.02 ;
    RECT 203.6 38.23 203.81 38.3 ;
    RECT 203.6 38.59 203.81 38.66 ;
    RECT 203.6 38.95 203.81 39.02 ;
    RECT 203.14 38.23 203.35 38.3 ;
    RECT 203.14 38.59 203.35 38.66 ;
    RECT 203.14 38.95 203.35 39.02 ;
    RECT 200.28 38.23 200.49 38.3 ;
    RECT 200.28 38.59 200.49 38.66 ;
    RECT 200.28 38.95 200.49 39.02 ;
    RECT 199.82 38.23 200.03 38.3 ;
    RECT 199.82 38.59 200.03 38.66 ;
    RECT 199.82 38.95 200.03 39.02 ;
    RECT 196.96 38.23 197.17 38.3 ;
    RECT 196.96 38.59 197.17 38.66 ;
    RECT 196.96 38.95 197.17 39.02 ;
    RECT 196.5 38.23 196.71 38.3 ;
    RECT 196.5 38.59 196.71 38.66 ;
    RECT 196.5 38.95 196.71 39.02 ;
    RECT 193.64 38.23 193.85 38.3 ;
    RECT 193.64 38.59 193.85 38.66 ;
    RECT 193.64 38.95 193.85 39.02 ;
    RECT 193.18 38.23 193.39 38.3 ;
    RECT 193.18 38.59 193.39 38.66 ;
    RECT 193.18 38.95 193.39 39.02 ;
    RECT 190.32 38.23 190.53 38.3 ;
    RECT 190.32 38.59 190.53 38.66 ;
    RECT 190.32 38.95 190.53 39.02 ;
    RECT 189.86 38.23 190.07 38.3 ;
    RECT 189.86 38.59 190.07 38.66 ;
    RECT 189.86 38.95 190.07 39.02 ;
    RECT 187.0 38.23 187.21 38.3 ;
    RECT 187.0 38.59 187.21 38.66 ;
    RECT 187.0 38.95 187.21 39.02 ;
    RECT 186.54 38.23 186.75 38.3 ;
    RECT 186.54 38.59 186.75 38.66 ;
    RECT 186.54 38.95 186.75 39.02 ;
    RECT 183.68 38.23 183.89 38.3 ;
    RECT 183.68 38.59 183.89 38.66 ;
    RECT 183.68 38.95 183.89 39.02 ;
    RECT 183.22 38.23 183.43 38.3 ;
    RECT 183.22 38.59 183.43 38.66 ;
    RECT 183.22 38.95 183.43 39.02 ;
    RECT 147.485 38.59 147.555 38.66 ;
    RECT 266.68 38.23 266.89 38.3 ;
    RECT 266.68 38.59 266.89 38.66 ;
    RECT 266.68 38.95 266.89 39.02 ;
    RECT 266.22 38.23 266.43 38.3 ;
    RECT 266.22 38.59 266.43 38.66 ;
    RECT 266.22 38.95 266.43 39.02 ;
    RECT 263.36 38.23 263.57 38.3 ;
    RECT 263.36 38.59 263.57 38.66 ;
    RECT 263.36 38.95 263.57 39.02 ;
    RECT 262.9 38.23 263.11 38.3 ;
    RECT 262.9 38.59 263.11 38.66 ;
    RECT 262.9 38.95 263.11 39.02 ;
    RECT 260.04 38.23 260.25 38.3 ;
    RECT 260.04 38.59 260.25 38.66 ;
    RECT 260.04 38.95 260.25 39.02 ;
    RECT 259.58 38.23 259.79 38.3 ;
    RECT 259.58 38.59 259.79 38.66 ;
    RECT 259.58 38.95 259.79 39.02 ;
    RECT 256.72 38.23 256.93 38.3 ;
    RECT 256.72 38.59 256.93 38.66 ;
    RECT 256.72 38.95 256.93 39.02 ;
    RECT 256.26 38.23 256.47 38.3 ;
    RECT 256.26 38.59 256.47 38.66 ;
    RECT 256.26 38.95 256.47 39.02 ;
    RECT 253.4 38.23 253.61 38.3 ;
    RECT 253.4 38.59 253.61 38.66 ;
    RECT 253.4 38.95 253.61 39.02 ;
    RECT 252.94 38.23 253.15 38.3 ;
    RECT 252.94 38.59 253.15 38.66 ;
    RECT 252.94 38.95 253.15 39.02 ;
    RECT 250.08 77.85 250.29 77.92 ;
    RECT 250.08 78.21 250.29 78.28 ;
    RECT 250.08 78.57 250.29 78.64 ;
    RECT 249.62 77.85 249.83 77.92 ;
    RECT 249.62 78.21 249.83 78.28 ;
    RECT 249.62 78.57 249.83 78.64 ;
    RECT 246.76 77.85 246.97 77.92 ;
    RECT 246.76 78.21 246.97 78.28 ;
    RECT 246.76 78.57 246.97 78.64 ;
    RECT 246.3 77.85 246.51 77.92 ;
    RECT 246.3 78.21 246.51 78.28 ;
    RECT 246.3 78.57 246.51 78.64 ;
    RECT 243.44 77.85 243.65 77.92 ;
    RECT 243.44 78.21 243.65 78.28 ;
    RECT 243.44 78.57 243.65 78.64 ;
    RECT 242.98 77.85 243.19 77.92 ;
    RECT 242.98 78.21 243.19 78.28 ;
    RECT 242.98 78.57 243.19 78.64 ;
    RECT 240.12 77.85 240.33 77.92 ;
    RECT 240.12 78.21 240.33 78.28 ;
    RECT 240.12 78.57 240.33 78.64 ;
    RECT 239.66 77.85 239.87 77.92 ;
    RECT 239.66 78.21 239.87 78.28 ;
    RECT 239.66 78.57 239.87 78.64 ;
    RECT 236.8 77.85 237.01 77.92 ;
    RECT 236.8 78.21 237.01 78.28 ;
    RECT 236.8 78.57 237.01 78.64 ;
    RECT 236.34 77.85 236.55 77.92 ;
    RECT 236.34 78.21 236.55 78.28 ;
    RECT 236.34 78.57 236.55 78.64 ;
    RECT 233.48 77.85 233.69 77.92 ;
    RECT 233.48 78.21 233.69 78.28 ;
    RECT 233.48 78.57 233.69 78.64 ;
    RECT 233.02 77.85 233.23 77.92 ;
    RECT 233.02 78.21 233.23 78.28 ;
    RECT 233.02 78.57 233.23 78.64 ;
    RECT 230.16 77.85 230.37 77.92 ;
    RECT 230.16 78.21 230.37 78.28 ;
    RECT 230.16 78.57 230.37 78.64 ;
    RECT 229.7 77.85 229.91 77.92 ;
    RECT 229.7 78.21 229.91 78.28 ;
    RECT 229.7 78.57 229.91 78.64 ;
    RECT 226.84 77.85 227.05 77.92 ;
    RECT 226.84 78.21 227.05 78.28 ;
    RECT 226.84 78.57 227.05 78.64 ;
    RECT 226.38 77.85 226.59 77.92 ;
    RECT 226.38 78.21 226.59 78.28 ;
    RECT 226.38 78.57 226.59 78.64 ;
    RECT 223.52 77.85 223.73 77.92 ;
    RECT 223.52 78.21 223.73 78.28 ;
    RECT 223.52 78.57 223.73 78.64 ;
    RECT 223.06 77.85 223.27 77.92 ;
    RECT 223.06 78.21 223.27 78.28 ;
    RECT 223.06 78.57 223.27 78.64 ;
    RECT 220.2 77.85 220.41 77.92 ;
    RECT 220.2 78.21 220.41 78.28 ;
    RECT 220.2 78.57 220.41 78.64 ;
    RECT 219.74 77.85 219.95 77.92 ;
    RECT 219.74 78.21 219.95 78.28 ;
    RECT 219.74 78.57 219.95 78.64 ;
    RECT 216.88 77.85 217.09 77.92 ;
    RECT 216.88 78.21 217.09 78.28 ;
    RECT 216.88 78.57 217.09 78.64 ;
    RECT 216.42 77.85 216.63 77.92 ;
    RECT 216.42 78.21 216.63 78.28 ;
    RECT 216.42 78.57 216.63 78.64 ;
    RECT 267.91 78.21 267.98 78.28 ;
    RECT 180.36 77.85 180.57 77.92 ;
    RECT 180.36 78.21 180.57 78.28 ;
    RECT 180.36 78.57 180.57 78.64 ;
    RECT 179.9 77.85 180.11 77.92 ;
    RECT 179.9 78.21 180.11 78.28 ;
    RECT 179.9 78.57 180.11 78.64 ;
    RECT 177.04 77.85 177.25 77.92 ;
    RECT 177.04 78.21 177.25 78.28 ;
    RECT 177.04 78.57 177.25 78.64 ;
    RECT 176.58 77.85 176.79 77.92 ;
    RECT 176.58 78.21 176.79 78.28 ;
    RECT 176.58 78.57 176.79 78.64 ;
    RECT 173.72 77.85 173.93 77.92 ;
    RECT 173.72 78.21 173.93 78.28 ;
    RECT 173.72 78.57 173.93 78.64 ;
    RECT 173.26 77.85 173.47 77.92 ;
    RECT 173.26 78.21 173.47 78.28 ;
    RECT 173.26 78.57 173.47 78.64 ;
    RECT 170.4 77.85 170.61 77.92 ;
    RECT 170.4 78.21 170.61 78.28 ;
    RECT 170.4 78.57 170.61 78.64 ;
    RECT 169.94 77.85 170.15 77.92 ;
    RECT 169.94 78.21 170.15 78.28 ;
    RECT 169.94 78.57 170.15 78.64 ;
    RECT 167.08 77.85 167.29 77.92 ;
    RECT 167.08 78.21 167.29 78.28 ;
    RECT 167.08 78.57 167.29 78.64 ;
    RECT 166.62 77.85 166.83 77.92 ;
    RECT 166.62 78.21 166.83 78.28 ;
    RECT 166.62 78.57 166.83 78.64 ;
    RECT 163.76 77.85 163.97 77.92 ;
    RECT 163.76 78.21 163.97 78.28 ;
    RECT 163.76 78.57 163.97 78.64 ;
    RECT 163.3 77.85 163.51 77.92 ;
    RECT 163.3 78.21 163.51 78.28 ;
    RECT 163.3 78.57 163.51 78.64 ;
    RECT 160.44 77.85 160.65 77.92 ;
    RECT 160.44 78.21 160.65 78.28 ;
    RECT 160.44 78.57 160.65 78.64 ;
    RECT 159.98 77.85 160.19 77.92 ;
    RECT 159.98 78.21 160.19 78.28 ;
    RECT 159.98 78.57 160.19 78.64 ;
    RECT 157.12 77.85 157.33 77.92 ;
    RECT 157.12 78.21 157.33 78.28 ;
    RECT 157.12 78.57 157.33 78.64 ;
    RECT 156.66 77.85 156.87 77.92 ;
    RECT 156.66 78.21 156.87 78.28 ;
    RECT 156.66 78.57 156.87 78.64 ;
    RECT 153.8 77.85 154.01 77.92 ;
    RECT 153.8 78.21 154.01 78.28 ;
    RECT 153.8 78.57 154.01 78.64 ;
    RECT 153.34 77.85 153.55 77.92 ;
    RECT 153.34 78.21 153.55 78.28 ;
    RECT 153.34 78.57 153.55 78.64 ;
    RECT 150.48 77.85 150.69 77.92 ;
    RECT 150.48 78.21 150.69 78.28 ;
    RECT 150.48 78.57 150.69 78.64 ;
    RECT 150.02 77.85 150.23 77.92 ;
    RECT 150.02 78.21 150.23 78.28 ;
    RECT 150.02 78.57 150.23 78.64 ;
    RECT 213.56 77.85 213.77 77.92 ;
    RECT 213.56 78.21 213.77 78.28 ;
    RECT 213.56 78.57 213.77 78.64 ;
    RECT 213.1 77.85 213.31 77.92 ;
    RECT 213.1 78.21 213.31 78.28 ;
    RECT 213.1 78.57 213.31 78.64 ;
    RECT 210.24 77.85 210.45 77.92 ;
    RECT 210.24 78.21 210.45 78.28 ;
    RECT 210.24 78.57 210.45 78.64 ;
    RECT 209.78 77.85 209.99 77.92 ;
    RECT 209.78 78.21 209.99 78.28 ;
    RECT 209.78 78.57 209.99 78.64 ;
    RECT 206.92 77.85 207.13 77.92 ;
    RECT 206.92 78.21 207.13 78.28 ;
    RECT 206.92 78.57 207.13 78.64 ;
    RECT 206.46 77.85 206.67 77.92 ;
    RECT 206.46 78.21 206.67 78.28 ;
    RECT 206.46 78.57 206.67 78.64 ;
    RECT 203.6 77.85 203.81 77.92 ;
    RECT 203.6 78.21 203.81 78.28 ;
    RECT 203.6 78.57 203.81 78.64 ;
    RECT 203.14 77.85 203.35 77.92 ;
    RECT 203.14 78.21 203.35 78.28 ;
    RECT 203.14 78.57 203.35 78.64 ;
    RECT 200.28 77.85 200.49 77.92 ;
    RECT 200.28 78.21 200.49 78.28 ;
    RECT 200.28 78.57 200.49 78.64 ;
    RECT 199.82 77.85 200.03 77.92 ;
    RECT 199.82 78.21 200.03 78.28 ;
    RECT 199.82 78.57 200.03 78.64 ;
    RECT 196.96 77.85 197.17 77.92 ;
    RECT 196.96 78.21 197.17 78.28 ;
    RECT 196.96 78.57 197.17 78.64 ;
    RECT 196.5 77.85 196.71 77.92 ;
    RECT 196.5 78.21 196.71 78.28 ;
    RECT 196.5 78.57 196.71 78.64 ;
    RECT 193.64 77.85 193.85 77.92 ;
    RECT 193.64 78.21 193.85 78.28 ;
    RECT 193.64 78.57 193.85 78.64 ;
    RECT 193.18 77.85 193.39 77.92 ;
    RECT 193.18 78.21 193.39 78.28 ;
    RECT 193.18 78.57 193.39 78.64 ;
    RECT 190.32 77.85 190.53 77.92 ;
    RECT 190.32 78.21 190.53 78.28 ;
    RECT 190.32 78.57 190.53 78.64 ;
    RECT 189.86 77.85 190.07 77.92 ;
    RECT 189.86 78.21 190.07 78.28 ;
    RECT 189.86 78.57 190.07 78.64 ;
    RECT 187.0 77.85 187.21 77.92 ;
    RECT 187.0 78.21 187.21 78.28 ;
    RECT 187.0 78.57 187.21 78.64 ;
    RECT 186.54 77.85 186.75 77.92 ;
    RECT 186.54 78.21 186.75 78.28 ;
    RECT 186.54 78.57 186.75 78.64 ;
    RECT 183.68 77.85 183.89 77.92 ;
    RECT 183.68 78.21 183.89 78.28 ;
    RECT 183.68 78.57 183.89 78.64 ;
    RECT 183.22 77.85 183.43 77.92 ;
    RECT 183.22 78.21 183.43 78.28 ;
    RECT 183.22 78.57 183.43 78.64 ;
    RECT 147.485 78.21 147.555 78.28 ;
    RECT 266.68 77.85 266.89 77.92 ;
    RECT 266.68 78.21 266.89 78.28 ;
    RECT 266.68 78.57 266.89 78.64 ;
    RECT 266.22 77.85 266.43 77.92 ;
    RECT 266.22 78.21 266.43 78.28 ;
    RECT 266.22 78.57 266.43 78.64 ;
    RECT 263.36 77.85 263.57 77.92 ;
    RECT 263.36 78.21 263.57 78.28 ;
    RECT 263.36 78.57 263.57 78.64 ;
    RECT 262.9 77.85 263.11 77.92 ;
    RECT 262.9 78.21 263.11 78.28 ;
    RECT 262.9 78.57 263.11 78.64 ;
    RECT 260.04 77.85 260.25 77.92 ;
    RECT 260.04 78.21 260.25 78.28 ;
    RECT 260.04 78.57 260.25 78.64 ;
    RECT 259.58 77.85 259.79 77.92 ;
    RECT 259.58 78.21 259.79 78.28 ;
    RECT 259.58 78.57 259.79 78.64 ;
    RECT 256.72 77.85 256.93 77.92 ;
    RECT 256.72 78.21 256.93 78.28 ;
    RECT 256.72 78.57 256.93 78.64 ;
    RECT 256.26 77.85 256.47 77.92 ;
    RECT 256.26 78.21 256.47 78.28 ;
    RECT 256.26 78.57 256.47 78.64 ;
    RECT 253.4 77.85 253.61 77.92 ;
    RECT 253.4 78.21 253.61 78.28 ;
    RECT 253.4 78.57 253.61 78.64 ;
    RECT 252.94 77.85 253.15 77.92 ;
    RECT 252.94 78.21 253.15 78.28 ;
    RECT 252.94 78.57 253.15 78.64 ;
    RECT 250.08 37.51 250.29 37.58 ;
    RECT 250.08 37.87 250.29 37.94 ;
    RECT 250.08 38.23 250.29 38.3 ;
    RECT 249.62 37.51 249.83 37.58 ;
    RECT 249.62 37.87 249.83 37.94 ;
    RECT 249.62 38.23 249.83 38.3 ;
    RECT 246.76 37.51 246.97 37.58 ;
    RECT 246.76 37.87 246.97 37.94 ;
    RECT 246.76 38.23 246.97 38.3 ;
    RECT 246.3 37.51 246.51 37.58 ;
    RECT 246.3 37.87 246.51 37.94 ;
    RECT 246.3 38.23 246.51 38.3 ;
    RECT 243.44 37.51 243.65 37.58 ;
    RECT 243.44 37.87 243.65 37.94 ;
    RECT 243.44 38.23 243.65 38.3 ;
    RECT 242.98 37.51 243.19 37.58 ;
    RECT 242.98 37.87 243.19 37.94 ;
    RECT 242.98 38.23 243.19 38.3 ;
    RECT 240.12 37.51 240.33 37.58 ;
    RECT 240.12 37.87 240.33 37.94 ;
    RECT 240.12 38.23 240.33 38.3 ;
    RECT 239.66 37.51 239.87 37.58 ;
    RECT 239.66 37.87 239.87 37.94 ;
    RECT 239.66 38.23 239.87 38.3 ;
    RECT 236.8 37.51 237.01 37.58 ;
    RECT 236.8 37.87 237.01 37.94 ;
    RECT 236.8 38.23 237.01 38.3 ;
    RECT 236.34 37.51 236.55 37.58 ;
    RECT 236.34 37.87 236.55 37.94 ;
    RECT 236.34 38.23 236.55 38.3 ;
    RECT 233.48 37.51 233.69 37.58 ;
    RECT 233.48 37.87 233.69 37.94 ;
    RECT 233.48 38.23 233.69 38.3 ;
    RECT 233.02 37.51 233.23 37.58 ;
    RECT 233.02 37.87 233.23 37.94 ;
    RECT 233.02 38.23 233.23 38.3 ;
    RECT 230.16 37.51 230.37 37.58 ;
    RECT 230.16 37.87 230.37 37.94 ;
    RECT 230.16 38.23 230.37 38.3 ;
    RECT 229.7 37.51 229.91 37.58 ;
    RECT 229.7 37.87 229.91 37.94 ;
    RECT 229.7 38.23 229.91 38.3 ;
    RECT 226.84 37.51 227.05 37.58 ;
    RECT 226.84 37.87 227.05 37.94 ;
    RECT 226.84 38.23 227.05 38.3 ;
    RECT 226.38 37.51 226.59 37.58 ;
    RECT 226.38 37.87 226.59 37.94 ;
    RECT 226.38 38.23 226.59 38.3 ;
    RECT 223.52 37.51 223.73 37.58 ;
    RECT 223.52 37.87 223.73 37.94 ;
    RECT 223.52 38.23 223.73 38.3 ;
    RECT 223.06 37.51 223.27 37.58 ;
    RECT 223.06 37.87 223.27 37.94 ;
    RECT 223.06 38.23 223.27 38.3 ;
    RECT 220.2 37.51 220.41 37.58 ;
    RECT 220.2 37.87 220.41 37.94 ;
    RECT 220.2 38.23 220.41 38.3 ;
    RECT 219.74 37.51 219.95 37.58 ;
    RECT 219.74 37.87 219.95 37.94 ;
    RECT 219.74 38.23 219.95 38.3 ;
    RECT 216.88 37.51 217.09 37.58 ;
    RECT 216.88 37.87 217.09 37.94 ;
    RECT 216.88 38.23 217.09 38.3 ;
    RECT 216.42 37.51 216.63 37.58 ;
    RECT 216.42 37.87 216.63 37.94 ;
    RECT 216.42 38.23 216.63 38.3 ;
    RECT 267.91 37.87 267.98 37.94 ;
    RECT 180.36 37.51 180.57 37.58 ;
    RECT 180.36 37.87 180.57 37.94 ;
    RECT 180.36 38.23 180.57 38.3 ;
    RECT 179.9 37.51 180.11 37.58 ;
    RECT 179.9 37.87 180.11 37.94 ;
    RECT 179.9 38.23 180.11 38.3 ;
    RECT 177.04 37.51 177.25 37.58 ;
    RECT 177.04 37.87 177.25 37.94 ;
    RECT 177.04 38.23 177.25 38.3 ;
    RECT 176.58 37.51 176.79 37.58 ;
    RECT 176.58 37.87 176.79 37.94 ;
    RECT 176.58 38.23 176.79 38.3 ;
    RECT 173.72 37.51 173.93 37.58 ;
    RECT 173.72 37.87 173.93 37.94 ;
    RECT 173.72 38.23 173.93 38.3 ;
    RECT 173.26 37.51 173.47 37.58 ;
    RECT 173.26 37.87 173.47 37.94 ;
    RECT 173.26 38.23 173.47 38.3 ;
    RECT 170.4 37.51 170.61 37.58 ;
    RECT 170.4 37.87 170.61 37.94 ;
    RECT 170.4 38.23 170.61 38.3 ;
    RECT 169.94 37.51 170.15 37.58 ;
    RECT 169.94 37.87 170.15 37.94 ;
    RECT 169.94 38.23 170.15 38.3 ;
    RECT 167.08 37.51 167.29 37.58 ;
    RECT 167.08 37.87 167.29 37.94 ;
    RECT 167.08 38.23 167.29 38.3 ;
    RECT 166.62 37.51 166.83 37.58 ;
    RECT 166.62 37.87 166.83 37.94 ;
    RECT 166.62 38.23 166.83 38.3 ;
    RECT 163.76 37.51 163.97 37.58 ;
    RECT 163.76 37.87 163.97 37.94 ;
    RECT 163.76 38.23 163.97 38.3 ;
    RECT 163.3 37.51 163.51 37.58 ;
    RECT 163.3 37.87 163.51 37.94 ;
    RECT 163.3 38.23 163.51 38.3 ;
    RECT 160.44 37.51 160.65 37.58 ;
    RECT 160.44 37.87 160.65 37.94 ;
    RECT 160.44 38.23 160.65 38.3 ;
    RECT 159.98 37.51 160.19 37.58 ;
    RECT 159.98 37.87 160.19 37.94 ;
    RECT 159.98 38.23 160.19 38.3 ;
    RECT 157.12 37.51 157.33 37.58 ;
    RECT 157.12 37.87 157.33 37.94 ;
    RECT 157.12 38.23 157.33 38.3 ;
    RECT 156.66 37.51 156.87 37.58 ;
    RECT 156.66 37.87 156.87 37.94 ;
    RECT 156.66 38.23 156.87 38.3 ;
    RECT 153.8 37.51 154.01 37.58 ;
    RECT 153.8 37.87 154.01 37.94 ;
    RECT 153.8 38.23 154.01 38.3 ;
    RECT 153.34 37.51 153.55 37.58 ;
    RECT 153.34 37.87 153.55 37.94 ;
    RECT 153.34 38.23 153.55 38.3 ;
    RECT 150.48 37.51 150.69 37.58 ;
    RECT 150.48 37.87 150.69 37.94 ;
    RECT 150.48 38.23 150.69 38.3 ;
    RECT 150.02 37.51 150.23 37.58 ;
    RECT 150.02 37.87 150.23 37.94 ;
    RECT 150.02 38.23 150.23 38.3 ;
    RECT 213.56 37.51 213.77 37.58 ;
    RECT 213.56 37.87 213.77 37.94 ;
    RECT 213.56 38.23 213.77 38.3 ;
    RECT 213.1 37.51 213.31 37.58 ;
    RECT 213.1 37.87 213.31 37.94 ;
    RECT 213.1 38.23 213.31 38.3 ;
    RECT 210.24 37.51 210.45 37.58 ;
    RECT 210.24 37.87 210.45 37.94 ;
    RECT 210.24 38.23 210.45 38.3 ;
    RECT 209.78 37.51 209.99 37.58 ;
    RECT 209.78 37.87 209.99 37.94 ;
    RECT 209.78 38.23 209.99 38.3 ;
    RECT 206.92 37.51 207.13 37.58 ;
    RECT 206.92 37.87 207.13 37.94 ;
    RECT 206.92 38.23 207.13 38.3 ;
    RECT 206.46 37.51 206.67 37.58 ;
    RECT 206.46 37.87 206.67 37.94 ;
    RECT 206.46 38.23 206.67 38.3 ;
    RECT 203.6 37.51 203.81 37.58 ;
    RECT 203.6 37.87 203.81 37.94 ;
    RECT 203.6 38.23 203.81 38.3 ;
    RECT 203.14 37.51 203.35 37.58 ;
    RECT 203.14 37.87 203.35 37.94 ;
    RECT 203.14 38.23 203.35 38.3 ;
    RECT 200.28 37.51 200.49 37.58 ;
    RECT 200.28 37.87 200.49 37.94 ;
    RECT 200.28 38.23 200.49 38.3 ;
    RECT 199.82 37.51 200.03 37.58 ;
    RECT 199.82 37.87 200.03 37.94 ;
    RECT 199.82 38.23 200.03 38.3 ;
    RECT 196.96 37.51 197.17 37.58 ;
    RECT 196.96 37.87 197.17 37.94 ;
    RECT 196.96 38.23 197.17 38.3 ;
    RECT 196.5 37.51 196.71 37.58 ;
    RECT 196.5 37.87 196.71 37.94 ;
    RECT 196.5 38.23 196.71 38.3 ;
    RECT 193.64 37.51 193.85 37.58 ;
    RECT 193.64 37.87 193.85 37.94 ;
    RECT 193.64 38.23 193.85 38.3 ;
    RECT 193.18 37.51 193.39 37.58 ;
    RECT 193.18 37.87 193.39 37.94 ;
    RECT 193.18 38.23 193.39 38.3 ;
    RECT 190.32 37.51 190.53 37.58 ;
    RECT 190.32 37.87 190.53 37.94 ;
    RECT 190.32 38.23 190.53 38.3 ;
    RECT 189.86 37.51 190.07 37.58 ;
    RECT 189.86 37.87 190.07 37.94 ;
    RECT 189.86 38.23 190.07 38.3 ;
    RECT 187.0 37.51 187.21 37.58 ;
    RECT 187.0 37.87 187.21 37.94 ;
    RECT 187.0 38.23 187.21 38.3 ;
    RECT 186.54 37.51 186.75 37.58 ;
    RECT 186.54 37.87 186.75 37.94 ;
    RECT 186.54 38.23 186.75 38.3 ;
    RECT 183.68 37.51 183.89 37.58 ;
    RECT 183.68 37.87 183.89 37.94 ;
    RECT 183.68 38.23 183.89 38.3 ;
    RECT 183.22 37.51 183.43 37.58 ;
    RECT 183.22 37.87 183.43 37.94 ;
    RECT 183.22 38.23 183.43 38.3 ;
    RECT 147.485 37.87 147.555 37.94 ;
    RECT 266.68 37.51 266.89 37.58 ;
    RECT 266.68 37.87 266.89 37.94 ;
    RECT 266.68 38.23 266.89 38.3 ;
    RECT 266.22 37.51 266.43 37.58 ;
    RECT 266.22 37.87 266.43 37.94 ;
    RECT 266.22 38.23 266.43 38.3 ;
    RECT 263.36 37.51 263.57 37.58 ;
    RECT 263.36 37.87 263.57 37.94 ;
    RECT 263.36 38.23 263.57 38.3 ;
    RECT 262.9 37.51 263.11 37.58 ;
    RECT 262.9 37.87 263.11 37.94 ;
    RECT 262.9 38.23 263.11 38.3 ;
    RECT 260.04 37.51 260.25 37.58 ;
    RECT 260.04 37.87 260.25 37.94 ;
    RECT 260.04 38.23 260.25 38.3 ;
    RECT 259.58 37.51 259.79 37.58 ;
    RECT 259.58 37.87 259.79 37.94 ;
    RECT 259.58 38.23 259.79 38.3 ;
    RECT 256.72 37.51 256.93 37.58 ;
    RECT 256.72 37.87 256.93 37.94 ;
    RECT 256.72 38.23 256.93 38.3 ;
    RECT 256.26 37.51 256.47 37.58 ;
    RECT 256.26 37.87 256.47 37.94 ;
    RECT 256.26 38.23 256.47 38.3 ;
    RECT 253.4 37.51 253.61 37.58 ;
    RECT 253.4 37.87 253.61 37.94 ;
    RECT 253.4 38.23 253.61 38.3 ;
    RECT 252.94 37.51 253.15 37.58 ;
    RECT 252.94 37.87 253.15 37.94 ;
    RECT 252.94 38.23 253.15 38.3 ;
    RECT 250.08 77.13 250.29 77.2 ;
    RECT 250.08 77.49 250.29 77.56 ;
    RECT 250.08 77.85 250.29 77.92 ;
    RECT 249.62 77.13 249.83 77.2 ;
    RECT 249.62 77.49 249.83 77.56 ;
    RECT 249.62 77.85 249.83 77.92 ;
    RECT 246.76 77.13 246.97 77.2 ;
    RECT 246.76 77.49 246.97 77.56 ;
    RECT 246.76 77.85 246.97 77.92 ;
    RECT 246.3 77.13 246.51 77.2 ;
    RECT 246.3 77.49 246.51 77.56 ;
    RECT 246.3 77.85 246.51 77.92 ;
    RECT 243.44 77.13 243.65 77.2 ;
    RECT 243.44 77.49 243.65 77.56 ;
    RECT 243.44 77.85 243.65 77.92 ;
    RECT 242.98 77.13 243.19 77.2 ;
    RECT 242.98 77.49 243.19 77.56 ;
    RECT 242.98 77.85 243.19 77.92 ;
    RECT 240.12 77.13 240.33 77.2 ;
    RECT 240.12 77.49 240.33 77.56 ;
    RECT 240.12 77.85 240.33 77.92 ;
    RECT 239.66 77.13 239.87 77.2 ;
    RECT 239.66 77.49 239.87 77.56 ;
    RECT 239.66 77.85 239.87 77.92 ;
    RECT 236.8 77.13 237.01 77.2 ;
    RECT 236.8 77.49 237.01 77.56 ;
    RECT 236.8 77.85 237.01 77.92 ;
    RECT 236.34 77.13 236.55 77.2 ;
    RECT 236.34 77.49 236.55 77.56 ;
    RECT 236.34 77.85 236.55 77.92 ;
    RECT 233.48 77.13 233.69 77.2 ;
    RECT 233.48 77.49 233.69 77.56 ;
    RECT 233.48 77.85 233.69 77.92 ;
    RECT 233.02 77.13 233.23 77.2 ;
    RECT 233.02 77.49 233.23 77.56 ;
    RECT 233.02 77.85 233.23 77.92 ;
    RECT 230.16 77.13 230.37 77.2 ;
    RECT 230.16 77.49 230.37 77.56 ;
    RECT 230.16 77.85 230.37 77.92 ;
    RECT 229.7 77.13 229.91 77.2 ;
    RECT 229.7 77.49 229.91 77.56 ;
    RECT 229.7 77.85 229.91 77.92 ;
    RECT 226.84 77.13 227.05 77.2 ;
    RECT 226.84 77.49 227.05 77.56 ;
    RECT 226.84 77.85 227.05 77.92 ;
    RECT 226.38 77.13 226.59 77.2 ;
    RECT 226.38 77.49 226.59 77.56 ;
    RECT 226.38 77.85 226.59 77.92 ;
    RECT 223.52 77.13 223.73 77.2 ;
    RECT 223.52 77.49 223.73 77.56 ;
    RECT 223.52 77.85 223.73 77.92 ;
    RECT 223.06 77.13 223.27 77.2 ;
    RECT 223.06 77.49 223.27 77.56 ;
    RECT 223.06 77.85 223.27 77.92 ;
    RECT 220.2 77.13 220.41 77.2 ;
    RECT 220.2 77.49 220.41 77.56 ;
    RECT 220.2 77.85 220.41 77.92 ;
    RECT 219.74 77.13 219.95 77.2 ;
    RECT 219.74 77.49 219.95 77.56 ;
    RECT 219.74 77.85 219.95 77.92 ;
    RECT 216.88 77.13 217.09 77.2 ;
    RECT 216.88 77.49 217.09 77.56 ;
    RECT 216.88 77.85 217.09 77.92 ;
    RECT 216.42 77.13 216.63 77.2 ;
    RECT 216.42 77.49 216.63 77.56 ;
    RECT 216.42 77.85 216.63 77.92 ;
    RECT 267.91 77.49 267.98 77.56 ;
    RECT 180.36 77.13 180.57 77.2 ;
    RECT 180.36 77.49 180.57 77.56 ;
    RECT 180.36 77.85 180.57 77.92 ;
    RECT 179.9 77.13 180.11 77.2 ;
    RECT 179.9 77.49 180.11 77.56 ;
    RECT 179.9 77.85 180.11 77.92 ;
    RECT 177.04 77.13 177.25 77.2 ;
    RECT 177.04 77.49 177.25 77.56 ;
    RECT 177.04 77.85 177.25 77.92 ;
    RECT 176.58 77.13 176.79 77.2 ;
    RECT 176.58 77.49 176.79 77.56 ;
    RECT 176.58 77.85 176.79 77.92 ;
    RECT 173.72 77.13 173.93 77.2 ;
    RECT 173.72 77.49 173.93 77.56 ;
    RECT 173.72 77.85 173.93 77.92 ;
    RECT 173.26 77.13 173.47 77.2 ;
    RECT 173.26 77.49 173.47 77.56 ;
    RECT 173.26 77.85 173.47 77.92 ;
    RECT 170.4 77.13 170.61 77.2 ;
    RECT 170.4 77.49 170.61 77.56 ;
    RECT 170.4 77.85 170.61 77.92 ;
    RECT 169.94 77.13 170.15 77.2 ;
    RECT 169.94 77.49 170.15 77.56 ;
    RECT 169.94 77.85 170.15 77.92 ;
    RECT 167.08 77.13 167.29 77.2 ;
    RECT 167.08 77.49 167.29 77.56 ;
    RECT 167.08 77.85 167.29 77.92 ;
    RECT 166.62 77.13 166.83 77.2 ;
    RECT 166.62 77.49 166.83 77.56 ;
    RECT 166.62 77.85 166.83 77.92 ;
    RECT 163.76 77.13 163.97 77.2 ;
    RECT 163.76 77.49 163.97 77.56 ;
    RECT 163.76 77.85 163.97 77.92 ;
    RECT 163.3 77.13 163.51 77.2 ;
    RECT 163.3 77.49 163.51 77.56 ;
    RECT 163.3 77.85 163.51 77.92 ;
    RECT 160.44 77.13 160.65 77.2 ;
    RECT 160.44 77.49 160.65 77.56 ;
    RECT 160.44 77.85 160.65 77.92 ;
    RECT 159.98 77.13 160.19 77.2 ;
    RECT 159.98 77.49 160.19 77.56 ;
    RECT 159.98 77.85 160.19 77.92 ;
    RECT 157.12 77.13 157.33 77.2 ;
    RECT 157.12 77.49 157.33 77.56 ;
    RECT 157.12 77.85 157.33 77.92 ;
    RECT 156.66 77.13 156.87 77.2 ;
    RECT 156.66 77.49 156.87 77.56 ;
    RECT 156.66 77.85 156.87 77.92 ;
    RECT 153.8 77.13 154.01 77.2 ;
    RECT 153.8 77.49 154.01 77.56 ;
    RECT 153.8 77.85 154.01 77.92 ;
    RECT 153.34 77.13 153.55 77.2 ;
    RECT 153.34 77.49 153.55 77.56 ;
    RECT 153.34 77.85 153.55 77.92 ;
    RECT 150.48 77.13 150.69 77.2 ;
    RECT 150.48 77.49 150.69 77.56 ;
    RECT 150.48 77.85 150.69 77.92 ;
    RECT 150.02 77.13 150.23 77.2 ;
    RECT 150.02 77.49 150.23 77.56 ;
    RECT 150.02 77.85 150.23 77.92 ;
    RECT 213.56 77.13 213.77 77.2 ;
    RECT 213.56 77.49 213.77 77.56 ;
    RECT 213.56 77.85 213.77 77.92 ;
    RECT 213.1 77.13 213.31 77.2 ;
    RECT 213.1 77.49 213.31 77.56 ;
    RECT 213.1 77.85 213.31 77.92 ;
    RECT 210.24 77.13 210.45 77.2 ;
    RECT 210.24 77.49 210.45 77.56 ;
    RECT 210.24 77.85 210.45 77.92 ;
    RECT 209.78 77.13 209.99 77.2 ;
    RECT 209.78 77.49 209.99 77.56 ;
    RECT 209.78 77.85 209.99 77.92 ;
    RECT 206.92 77.13 207.13 77.2 ;
    RECT 206.92 77.49 207.13 77.56 ;
    RECT 206.92 77.85 207.13 77.92 ;
    RECT 206.46 77.13 206.67 77.2 ;
    RECT 206.46 77.49 206.67 77.56 ;
    RECT 206.46 77.85 206.67 77.92 ;
    RECT 203.6 77.13 203.81 77.2 ;
    RECT 203.6 77.49 203.81 77.56 ;
    RECT 203.6 77.85 203.81 77.92 ;
    RECT 203.14 77.13 203.35 77.2 ;
    RECT 203.14 77.49 203.35 77.56 ;
    RECT 203.14 77.85 203.35 77.92 ;
    RECT 200.28 77.13 200.49 77.2 ;
    RECT 200.28 77.49 200.49 77.56 ;
    RECT 200.28 77.85 200.49 77.92 ;
    RECT 199.82 77.13 200.03 77.2 ;
    RECT 199.82 77.49 200.03 77.56 ;
    RECT 199.82 77.85 200.03 77.92 ;
    RECT 196.96 77.13 197.17 77.2 ;
    RECT 196.96 77.49 197.17 77.56 ;
    RECT 196.96 77.85 197.17 77.92 ;
    RECT 196.5 77.13 196.71 77.2 ;
    RECT 196.5 77.49 196.71 77.56 ;
    RECT 196.5 77.85 196.71 77.92 ;
    RECT 193.64 77.13 193.85 77.2 ;
    RECT 193.64 77.49 193.85 77.56 ;
    RECT 193.64 77.85 193.85 77.92 ;
    RECT 193.18 77.13 193.39 77.2 ;
    RECT 193.18 77.49 193.39 77.56 ;
    RECT 193.18 77.85 193.39 77.92 ;
    RECT 190.32 77.13 190.53 77.2 ;
    RECT 190.32 77.49 190.53 77.56 ;
    RECT 190.32 77.85 190.53 77.92 ;
    RECT 189.86 77.13 190.07 77.2 ;
    RECT 189.86 77.49 190.07 77.56 ;
    RECT 189.86 77.85 190.07 77.92 ;
    RECT 187.0 77.13 187.21 77.2 ;
    RECT 187.0 77.49 187.21 77.56 ;
    RECT 187.0 77.85 187.21 77.92 ;
    RECT 186.54 77.13 186.75 77.2 ;
    RECT 186.54 77.49 186.75 77.56 ;
    RECT 186.54 77.85 186.75 77.92 ;
    RECT 183.68 77.13 183.89 77.2 ;
    RECT 183.68 77.49 183.89 77.56 ;
    RECT 183.68 77.85 183.89 77.92 ;
    RECT 183.22 77.13 183.43 77.2 ;
    RECT 183.22 77.49 183.43 77.56 ;
    RECT 183.22 77.85 183.43 77.92 ;
    RECT 147.485 77.49 147.555 77.56 ;
    RECT 266.68 77.13 266.89 77.2 ;
    RECT 266.68 77.49 266.89 77.56 ;
    RECT 266.68 77.85 266.89 77.92 ;
    RECT 266.22 77.13 266.43 77.2 ;
    RECT 266.22 77.49 266.43 77.56 ;
    RECT 266.22 77.85 266.43 77.92 ;
    RECT 263.36 77.13 263.57 77.2 ;
    RECT 263.36 77.49 263.57 77.56 ;
    RECT 263.36 77.85 263.57 77.92 ;
    RECT 262.9 77.13 263.11 77.2 ;
    RECT 262.9 77.49 263.11 77.56 ;
    RECT 262.9 77.85 263.11 77.92 ;
    RECT 260.04 77.13 260.25 77.2 ;
    RECT 260.04 77.49 260.25 77.56 ;
    RECT 260.04 77.85 260.25 77.92 ;
    RECT 259.58 77.13 259.79 77.2 ;
    RECT 259.58 77.49 259.79 77.56 ;
    RECT 259.58 77.85 259.79 77.92 ;
    RECT 256.72 77.13 256.93 77.2 ;
    RECT 256.72 77.49 256.93 77.56 ;
    RECT 256.72 77.85 256.93 77.92 ;
    RECT 256.26 77.13 256.47 77.2 ;
    RECT 256.26 77.49 256.47 77.56 ;
    RECT 256.26 77.85 256.47 77.92 ;
    RECT 253.4 77.13 253.61 77.2 ;
    RECT 253.4 77.49 253.61 77.56 ;
    RECT 253.4 77.85 253.61 77.92 ;
    RECT 252.94 77.13 253.15 77.2 ;
    RECT 252.94 77.49 253.15 77.56 ;
    RECT 252.94 77.85 253.15 77.92 ;
    RECT 250.08 36.79 250.29 36.86 ;
    RECT 250.08 37.15 250.29 37.22 ;
    RECT 250.08 37.51 250.29 37.58 ;
    RECT 249.62 36.79 249.83 36.86 ;
    RECT 249.62 37.15 249.83 37.22 ;
    RECT 249.62 37.51 249.83 37.58 ;
    RECT 246.76 36.79 246.97 36.86 ;
    RECT 246.76 37.15 246.97 37.22 ;
    RECT 246.76 37.51 246.97 37.58 ;
    RECT 246.3 36.79 246.51 36.86 ;
    RECT 246.3 37.15 246.51 37.22 ;
    RECT 246.3 37.51 246.51 37.58 ;
    RECT 243.44 36.79 243.65 36.86 ;
    RECT 243.44 37.15 243.65 37.22 ;
    RECT 243.44 37.51 243.65 37.58 ;
    RECT 242.98 36.79 243.19 36.86 ;
    RECT 242.98 37.15 243.19 37.22 ;
    RECT 242.98 37.51 243.19 37.58 ;
    RECT 240.12 36.79 240.33 36.86 ;
    RECT 240.12 37.15 240.33 37.22 ;
    RECT 240.12 37.51 240.33 37.58 ;
    RECT 239.66 36.79 239.87 36.86 ;
    RECT 239.66 37.15 239.87 37.22 ;
    RECT 239.66 37.51 239.87 37.58 ;
    RECT 236.8 36.79 237.01 36.86 ;
    RECT 236.8 37.15 237.01 37.22 ;
    RECT 236.8 37.51 237.01 37.58 ;
    RECT 236.34 36.79 236.55 36.86 ;
    RECT 236.34 37.15 236.55 37.22 ;
    RECT 236.34 37.51 236.55 37.58 ;
    RECT 233.48 36.79 233.69 36.86 ;
    RECT 233.48 37.15 233.69 37.22 ;
    RECT 233.48 37.51 233.69 37.58 ;
    RECT 233.02 36.79 233.23 36.86 ;
    RECT 233.02 37.15 233.23 37.22 ;
    RECT 233.02 37.51 233.23 37.58 ;
    RECT 230.16 36.79 230.37 36.86 ;
    RECT 230.16 37.15 230.37 37.22 ;
    RECT 230.16 37.51 230.37 37.58 ;
    RECT 229.7 36.79 229.91 36.86 ;
    RECT 229.7 37.15 229.91 37.22 ;
    RECT 229.7 37.51 229.91 37.58 ;
    RECT 226.84 36.79 227.05 36.86 ;
    RECT 226.84 37.15 227.05 37.22 ;
    RECT 226.84 37.51 227.05 37.58 ;
    RECT 226.38 36.79 226.59 36.86 ;
    RECT 226.38 37.15 226.59 37.22 ;
    RECT 226.38 37.51 226.59 37.58 ;
    RECT 223.52 36.79 223.73 36.86 ;
    RECT 223.52 37.15 223.73 37.22 ;
    RECT 223.52 37.51 223.73 37.58 ;
    RECT 223.06 36.79 223.27 36.86 ;
    RECT 223.06 37.15 223.27 37.22 ;
    RECT 223.06 37.51 223.27 37.58 ;
    RECT 220.2 36.79 220.41 36.86 ;
    RECT 220.2 37.15 220.41 37.22 ;
    RECT 220.2 37.51 220.41 37.58 ;
    RECT 219.74 36.79 219.95 36.86 ;
    RECT 219.74 37.15 219.95 37.22 ;
    RECT 219.74 37.51 219.95 37.58 ;
    RECT 216.88 36.79 217.09 36.86 ;
    RECT 216.88 37.15 217.09 37.22 ;
    RECT 216.88 37.51 217.09 37.58 ;
    RECT 216.42 36.79 216.63 36.86 ;
    RECT 216.42 37.15 216.63 37.22 ;
    RECT 216.42 37.51 216.63 37.58 ;
    RECT 267.91 37.15 267.98 37.22 ;
    RECT 180.36 36.79 180.57 36.86 ;
    RECT 180.36 37.15 180.57 37.22 ;
    RECT 180.36 37.51 180.57 37.58 ;
    RECT 179.9 36.79 180.11 36.86 ;
    RECT 179.9 37.15 180.11 37.22 ;
    RECT 179.9 37.51 180.11 37.58 ;
    RECT 177.04 36.79 177.25 36.86 ;
    RECT 177.04 37.15 177.25 37.22 ;
    RECT 177.04 37.51 177.25 37.58 ;
    RECT 176.58 36.79 176.79 36.86 ;
    RECT 176.58 37.15 176.79 37.22 ;
    RECT 176.58 37.51 176.79 37.58 ;
    RECT 173.72 36.79 173.93 36.86 ;
    RECT 173.72 37.15 173.93 37.22 ;
    RECT 173.72 37.51 173.93 37.58 ;
    RECT 173.26 36.79 173.47 36.86 ;
    RECT 173.26 37.15 173.47 37.22 ;
    RECT 173.26 37.51 173.47 37.58 ;
    RECT 170.4 36.79 170.61 36.86 ;
    RECT 170.4 37.15 170.61 37.22 ;
    RECT 170.4 37.51 170.61 37.58 ;
    RECT 169.94 36.79 170.15 36.86 ;
    RECT 169.94 37.15 170.15 37.22 ;
    RECT 169.94 37.51 170.15 37.58 ;
    RECT 167.08 36.79 167.29 36.86 ;
    RECT 167.08 37.15 167.29 37.22 ;
    RECT 167.08 37.51 167.29 37.58 ;
    RECT 166.62 36.79 166.83 36.86 ;
    RECT 166.62 37.15 166.83 37.22 ;
    RECT 166.62 37.51 166.83 37.58 ;
    RECT 163.76 36.79 163.97 36.86 ;
    RECT 163.76 37.15 163.97 37.22 ;
    RECT 163.76 37.51 163.97 37.58 ;
    RECT 163.3 36.79 163.51 36.86 ;
    RECT 163.3 37.15 163.51 37.22 ;
    RECT 163.3 37.51 163.51 37.58 ;
    RECT 160.44 36.79 160.65 36.86 ;
    RECT 160.44 37.15 160.65 37.22 ;
    RECT 160.44 37.51 160.65 37.58 ;
    RECT 159.98 36.79 160.19 36.86 ;
    RECT 159.98 37.15 160.19 37.22 ;
    RECT 159.98 37.51 160.19 37.58 ;
    RECT 157.12 36.79 157.33 36.86 ;
    RECT 157.12 37.15 157.33 37.22 ;
    RECT 157.12 37.51 157.33 37.58 ;
    RECT 156.66 36.79 156.87 36.86 ;
    RECT 156.66 37.15 156.87 37.22 ;
    RECT 156.66 37.51 156.87 37.58 ;
    RECT 153.8 36.79 154.01 36.86 ;
    RECT 153.8 37.15 154.01 37.22 ;
    RECT 153.8 37.51 154.01 37.58 ;
    RECT 153.34 36.79 153.55 36.86 ;
    RECT 153.34 37.15 153.55 37.22 ;
    RECT 153.34 37.51 153.55 37.58 ;
    RECT 150.48 36.79 150.69 36.86 ;
    RECT 150.48 37.15 150.69 37.22 ;
    RECT 150.48 37.51 150.69 37.58 ;
    RECT 150.02 36.79 150.23 36.86 ;
    RECT 150.02 37.15 150.23 37.22 ;
    RECT 150.02 37.51 150.23 37.58 ;
    RECT 213.56 36.79 213.77 36.86 ;
    RECT 213.56 37.15 213.77 37.22 ;
    RECT 213.56 37.51 213.77 37.58 ;
    RECT 213.1 36.79 213.31 36.86 ;
    RECT 213.1 37.15 213.31 37.22 ;
    RECT 213.1 37.51 213.31 37.58 ;
    RECT 210.24 36.79 210.45 36.86 ;
    RECT 210.24 37.15 210.45 37.22 ;
    RECT 210.24 37.51 210.45 37.58 ;
    RECT 209.78 36.79 209.99 36.86 ;
    RECT 209.78 37.15 209.99 37.22 ;
    RECT 209.78 37.51 209.99 37.58 ;
    RECT 206.92 36.79 207.13 36.86 ;
    RECT 206.92 37.15 207.13 37.22 ;
    RECT 206.92 37.51 207.13 37.58 ;
    RECT 206.46 36.79 206.67 36.86 ;
    RECT 206.46 37.15 206.67 37.22 ;
    RECT 206.46 37.51 206.67 37.58 ;
    RECT 203.6 36.79 203.81 36.86 ;
    RECT 203.6 37.15 203.81 37.22 ;
    RECT 203.6 37.51 203.81 37.58 ;
    RECT 203.14 36.79 203.35 36.86 ;
    RECT 203.14 37.15 203.35 37.22 ;
    RECT 203.14 37.51 203.35 37.58 ;
    RECT 200.28 36.79 200.49 36.86 ;
    RECT 200.28 37.15 200.49 37.22 ;
    RECT 200.28 37.51 200.49 37.58 ;
    RECT 199.82 36.79 200.03 36.86 ;
    RECT 199.82 37.15 200.03 37.22 ;
    RECT 199.82 37.51 200.03 37.58 ;
    RECT 196.96 36.79 197.17 36.86 ;
    RECT 196.96 37.15 197.17 37.22 ;
    RECT 196.96 37.51 197.17 37.58 ;
    RECT 196.5 36.79 196.71 36.86 ;
    RECT 196.5 37.15 196.71 37.22 ;
    RECT 196.5 37.51 196.71 37.58 ;
    RECT 193.64 36.79 193.85 36.86 ;
    RECT 193.64 37.15 193.85 37.22 ;
    RECT 193.64 37.51 193.85 37.58 ;
    RECT 193.18 36.79 193.39 36.86 ;
    RECT 193.18 37.15 193.39 37.22 ;
    RECT 193.18 37.51 193.39 37.58 ;
    RECT 190.32 36.79 190.53 36.86 ;
    RECT 190.32 37.15 190.53 37.22 ;
    RECT 190.32 37.51 190.53 37.58 ;
    RECT 189.86 36.79 190.07 36.86 ;
    RECT 189.86 37.15 190.07 37.22 ;
    RECT 189.86 37.51 190.07 37.58 ;
    RECT 187.0 36.79 187.21 36.86 ;
    RECT 187.0 37.15 187.21 37.22 ;
    RECT 187.0 37.51 187.21 37.58 ;
    RECT 186.54 36.79 186.75 36.86 ;
    RECT 186.54 37.15 186.75 37.22 ;
    RECT 186.54 37.51 186.75 37.58 ;
    RECT 183.68 36.79 183.89 36.86 ;
    RECT 183.68 37.15 183.89 37.22 ;
    RECT 183.68 37.51 183.89 37.58 ;
    RECT 183.22 36.79 183.43 36.86 ;
    RECT 183.22 37.15 183.43 37.22 ;
    RECT 183.22 37.51 183.43 37.58 ;
    RECT 147.485 37.15 147.555 37.22 ;
    RECT 266.68 36.79 266.89 36.86 ;
    RECT 266.68 37.15 266.89 37.22 ;
    RECT 266.68 37.51 266.89 37.58 ;
    RECT 266.22 36.79 266.43 36.86 ;
    RECT 266.22 37.15 266.43 37.22 ;
    RECT 266.22 37.51 266.43 37.58 ;
    RECT 263.36 36.79 263.57 36.86 ;
    RECT 263.36 37.15 263.57 37.22 ;
    RECT 263.36 37.51 263.57 37.58 ;
    RECT 262.9 36.79 263.11 36.86 ;
    RECT 262.9 37.15 263.11 37.22 ;
    RECT 262.9 37.51 263.11 37.58 ;
    RECT 260.04 36.79 260.25 36.86 ;
    RECT 260.04 37.15 260.25 37.22 ;
    RECT 260.04 37.51 260.25 37.58 ;
    RECT 259.58 36.79 259.79 36.86 ;
    RECT 259.58 37.15 259.79 37.22 ;
    RECT 259.58 37.51 259.79 37.58 ;
    RECT 256.72 36.79 256.93 36.86 ;
    RECT 256.72 37.15 256.93 37.22 ;
    RECT 256.72 37.51 256.93 37.58 ;
    RECT 256.26 36.79 256.47 36.86 ;
    RECT 256.26 37.15 256.47 37.22 ;
    RECT 256.26 37.51 256.47 37.58 ;
    RECT 253.4 36.79 253.61 36.86 ;
    RECT 253.4 37.15 253.61 37.22 ;
    RECT 253.4 37.51 253.61 37.58 ;
    RECT 252.94 36.79 253.15 36.86 ;
    RECT 252.94 37.15 253.15 37.22 ;
    RECT 252.94 37.51 253.15 37.58 ;
    RECT 250.08 76.41 250.29 76.48 ;
    RECT 250.08 76.77 250.29 76.84 ;
    RECT 250.08 77.13 250.29 77.2 ;
    RECT 249.62 76.41 249.83 76.48 ;
    RECT 249.62 76.77 249.83 76.84 ;
    RECT 249.62 77.13 249.83 77.2 ;
    RECT 246.76 76.41 246.97 76.48 ;
    RECT 246.76 76.77 246.97 76.84 ;
    RECT 246.76 77.13 246.97 77.2 ;
    RECT 246.3 76.41 246.51 76.48 ;
    RECT 246.3 76.77 246.51 76.84 ;
    RECT 246.3 77.13 246.51 77.2 ;
    RECT 243.44 76.41 243.65 76.48 ;
    RECT 243.44 76.77 243.65 76.84 ;
    RECT 243.44 77.13 243.65 77.2 ;
    RECT 242.98 76.41 243.19 76.48 ;
    RECT 242.98 76.77 243.19 76.84 ;
    RECT 242.98 77.13 243.19 77.2 ;
    RECT 240.12 76.41 240.33 76.48 ;
    RECT 240.12 76.77 240.33 76.84 ;
    RECT 240.12 77.13 240.33 77.2 ;
    RECT 239.66 76.41 239.87 76.48 ;
    RECT 239.66 76.77 239.87 76.84 ;
    RECT 239.66 77.13 239.87 77.2 ;
    RECT 236.8 76.41 237.01 76.48 ;
    RECT 236.8 76.77 237.01 76.84 ;
    RECT 236.8 77.13 237.01 77.2 ;
    RECT 236.34 76.41 236.55 76.48 ;
    RECT 236.34 76.77 236.55 76.84 ;
    RECT 236.34 77.13 236.55 77.2 ;
    RECT 233.48 76.41 233.69 76.48 ;
    RECT 233.48 76.77 233.69 76.84 ;
    RECT 233.48 77.13 233.69 77.2 ;
    RECT 233.02 76.41 233.23 76.48 ;
    RECT 233.02 76.77 233.23 76.84 ;
    RECT 233.02 77.13 233.23 77.2 ;
    RECT 230.16 76.41 230.37 76.48 ;
    RECT 230.16 76.77 230.37 76.84 ;
    RECT 230.16 77.13 230.37 77.2 ;
    RECT 229.7 76.41 229.91 76.48 ;
    RECT 229.7 76.77 229.91 76.84 ;
    RECT 229.7 77.13 229.91 77.2 ;
    RECT 226.84 76.41 227.05 76.48 ;
    RECT 226.84 76.77 227.05 76.84 ;
    RECT 226.84 77.13 227.05 77.2 ;
    RECT 226.38 76.41 226.59 76.48 ;
    RECT 226.38 76.77 226.59 76.84 ;
    RECT 226.38 77.13 226.59 77.2 ;
    RECT 223.52 76.41 223.73 76.48 ;
    RECT 223.52 76.77 223.73 76.84 ;
    RECT 223.52 77.13 223.73 77.2 ;
    RECT 223.06 76.41 223.27 76.48 ;
    RECT 223.06 76.77 223.27 76.84 ;
    RECT 223.06 77.13 223.27 77.2 ;
    RECT 220.2 76.41 220.41 76.48 ;
    RECT 220.2 76.77 220.41 76.84 ;
    RECT 220.2 77.13 220.41 77.2 ;
    RECT 219.74 76.41 219.95 76.48 ;
    RECT 219.74 76.77 219.95 76.84 ;
    RECT 219.74 77.13 219.95 77.2 ;
    RECT 216.88 76.41 217.09 76.48 ;
    RECT 216.88 76.77 217.09 76.84 ;
    RECT 216.88 77.13 217.09 77.2 ;
    RECT 216.42 76.41 216.63 76.48 ;
    RECT 216.42 76.77 216.63 76.84 ;
    RECT 216.42 77.13 216.63 77.2 ;
    RECT 267.91 76.77 267.98 76.84 ;
    RECT 180.36 76.41 180.57 76.48 ;
    RECT 180.36 76.77 180.57 76.84 ;
    RECT 180.36 77.13 180.57 77.2 ;
    RECT 179.9 76.41 180.11 76.48 ;
    RECT 179.9 76.77 180.11 76.84 ;
    RECT 179.9 77.13 180.11 77.2 ;
    RECT 177.04 76.41 177.25 76.48 ;
    RECT 177.04 76.77 177.25 76.84 ;
    RECT 177.04 77.13 177.25 77.2 ;
    RECT 176.58 76.41 176.79 76.48 ;
    RECT 176.58 76.77 176.79 76.84 ;
    RECT 176.58 77.13 176.79 77.2 ;
    RECT 173.72 76.41 173.93 76.48 ;
    RECT 173.72 76.77 173.93 76.84 ;
    RECT 173.72 77.13 173.93 77.2 ;
    RECT 173.26 76.41 173.47 76.48 ;
    RECT 173.26 76.77 173.47 76.84 ;
    RECT 173.26 77.13 173.47 77.2 ;
    RECT 170.4 76.41 170.61 76.48 ;
    RECT 170.4 76.77 170.61 76.84 ;
    RECT 170.4 77.13 170.61 77.2 ;
    RECT 169.94 76.41 170.15 76.48 ;
    RECT 169.94 76.77 170.15 76.84 ;
    RECT 169.94 77.13 170.15 77.2 ;
    RECT 167.08 76.41 167.29 76.48 ;
    RECT 167.08 76.77 167.29 76.84 ;
    RECT 167.08 77.13 167.29 77.2 ;
    RECT 166.62 76.41 166.83 76.48 ;
    RECT 166.62 76.77 166.83 76.84 ;
    RECT 166.62 77.13 166.83 77.2 ;
    RECT 163.76 76.41 163.97 76.48 ;
    RECT 163.76 76.77 163.97 76.84 ;
    RECT 163.76 77.13 163.97 77.2 ;
    RECT 163.3 76.41 163.51 76.48 ;
    RECT 163.3 76.77 163.51 76.84 ;
    RECT 163.3 77.13 163.51 77.2 ;
    RECT 160.44 76.41 160.65 76.48 ;
    RECT 160.44 76.77 160.65 76.84 ;
    RECT 160.44 77.13 160.65 77.2 ;
    RECT 159.98 76.41 160.19 76.48 ;
    RECT 159.98 76.77 160.19 76.84 ;
    RECT 159.98 77.13 160.19 77.2 ;
    RECT 157.12 76.41 157.33 76.48 ;
    RECT 157.12 76.77 157.33 76.84 ;
    RECT 157.12 77.13 157.33 77.2 ;
    RECT 156.66 76.41 156.87 76.48 ;
    RECT 156.66 76.77 156.87 76.84 ;
    RECT 156.66 77.13 156.87 77.2 ;
    RECT 153.8 76.41 154.01 76.48 ;
    RECT 153.8 76.77 154.01 76.84 ;
    RECT 153.8 77.13 154.01 77.2 ;
    RECT 153.34 76.41 153.55 76.48 ;
    RECT 153.34 76.77 153.55 76.84 ;
    RECT 153.34 77.13 153.55 77.2 ;
    RECT 150.48 76.41 150.69 76.48 ;
    RECT 150.48 76.77 150.69 76.84 ;
    RECT 150.48 77.13 150.69 77.2 ;
    RECT 150.02 76.41 150.23 76.48 ;
    RECT 150.02 76.77 150.23 76.84 ;
    RECT 150.02 77.13 150.23 77.2 ;
    RECT 213.56 76.41 213.77 76.48 ;
    RECT 213.56 76.77 213.77 76.84 ;
    RECT 213.56 77.13 213.77 77.2 ;
    RECT 213.1 76.41 213.31 76.48 ;
    RECT 213.1 76.77 213.31 76.84 ;
    RECT 213.1 77.13 213.31 77.2 ;
    RECT 210.24 76.41 210.45 76.48 ;
    RECT 210.24 76.77 210.45 76.84 ;
    RECT 210.24 77.13 210.45 77.2 ;
    RECT 209.78 76.41 209.99 76.48 ;
    RECT 209.78 76.77 209.99 76.84 ;
    RECT 209.78 77.13 209.99 77.2 ;
    RECT 206.92 76.41 207.13 76.48 ;
    RECT 206.92 76.77 207.13 76.84 ;
    RECT 206.92 77.13 207.13 77.2 ;
    RECT 206.46 76.41 206.67 76.48 ;
    RECT 206.46 76.77 206.67 76.84 ;
    RECT 206.46 77.13 206.67 77.2 ;
    RECT 203.6 76.41 203.81 76.48 ;
    RECT 203.6 76.77 203.81 76.84 ;
    RECT 203.6 77.13 203.81 77.2 ;
    RECT 203.14 76.41 203.35 76.48 ;
    RECT 203.14 76.77 203.35 76.84 ;
    RECT 203.14 77.13 203.35 77.2 ;
    RECT 200.28 76.41 200.49 76.48 ;
    RECT 200.28 76.77 200.49 76.84 ;
    RECT 200.28 77.13 200.49 77.2 ;
    RECT 199.82 76.41 200.03 76.48 ;
    RECT 199.82 76.77 200.03 76.84 ;
    RECT 199.82 77.13 200.03 77.2 ;
    RECT 196.96 76.41 197.17 76.48 ;
    RECT 196.96 76.77 197.17 76.84 ;
    RECT 196.96 77.13 197.17 77.2 ;
    RECT 196.5 76.41 196.71 76.48 ;
    RECT 196.5 76.77 196.71 76.84 ;
    RECT 196.5 77.13 196.71 77.2 ;
    RECT 193.64 76.41 193.85 76.48 ;
    RECT 193.64 76.77 193.85 76.84 ;
    RECT 193.64 77.13 193.85 77.2 ;
    RECT 193.18 76.41 193.39 76.48 ;
    RECT 193.18 76.77 193.39 76.84 ;
    RECT 193.18 77.13 193.39 77.2 ;
    RECT 190.32 76.41 190.53 76.48 ;
    RECT 190.32 76.77 190.53 76.84 ;
    RECT 190.32 77.13 190.53 77.2 ;
    RECT 189.86 76.41 190.07 76.48 ;
    RECT 189.86 76.77 190.07 76.84 ;
    RECT 189.86 77.13 190.07 77.2 ;
    RECT 187.0 76.41 187.21 76.48 ;
    RECT 187.0 76.77 187.21 76.84 ;
    RECT 187.0 77.13 187.21 77.2 ;
    RECT 186.54 76.41 186.75 76.48 ;
    RECT 186.54 76.77 186.75 76.84 ;
    RECT 186.54 77.13 186.75 77.2 ;
    RECT 183.68 76.41 183.89 76.48 ;
    RECT 183.68 76.77 183.89 76.84 ;
    RECT 183.68 77.13 183.89 77.2 ;
    RECT 183.22 76.41 183.43 76.48 ;
    RECT 183.22 76.77 183.43 76.84 ;
    RECT 183.22 77.13 183.43 77.2 ;
    RECT 147.485 76.77 147.555 76.84 ;
    RECT 266.68 76.41 266.89 76.48 ;
    RECT 266.68 76.77 266.89 76.84 ;
    RECT 266.68 77.13 266.89 77.2 ;
    RECT 266.22 76.41 266.43 76.48 ;
    RECT 266.22 76.77 266.43 76.84 ;
    RECT 266.22 77.13 266.43 77.2 ;
    RECT 263.36 76.41 263.57 76.48 ;
    RECT 263.36 76.77 263.57 76.84 ;
    RECT 263.36 77.13 263.57 77.2 ;
    RECT 262.9 76.41 263.11 76.48 ;
    RECT 262.9 76.77 263.11 76.84 ;
    RECT 262.9 77.13 263.11 77.2 ;
    RECT 260.04 76.41 260.25 76.48 ;
    RECT 260.04 76.77 260.25 76.84 ;
    RECT 260.04 77.13 260.25 77.2 ;
    RECT 259.58 76.41 259.79 76.48 ;
    RECT 259.58 76.77 259.79 76.84 ;
    RECT 259.58 77.13 259.79 77.2 ;
    RECT 256.72 76.41 256.93 76.48 ;
    RECT 256.72 76.77 256.93 76.84 ;
    RECT 256.72 77.13 256.93 77.2 ;
    RECT 256.26 76.41 256.47 76.48 ;
    RECT 256.26 76.77 256.47 76.84 ;
    RECT 256.26 77.13 256.47 77.2 ;
    RECT 253.4 76.41 253.61 76.48 ;
    RECT 253.4 76.77 253.61 76.84 ;
    RECT 253.4 77.13 253.61 77.2 ;
    RECT 252.94 76.41 253.15 76.48 ;
    RECT 252.94 76.77 253.15 76.84 ;
    RECT 252.94 77.13 253.15 77.2 ;
    RECT 61.25 52.63 61.46 52.7 ;
    RECT 61.25 52.99 61.46 53.06 ;
    RECT 61.25 53.35 61.46 53.42 ;
    RECT 61.71 52.63 61.92 52.7 ;
    RECT 61.71 52.99 61.92 53.06 ;
    RECT 61.71 53.35 61.92 53.42 ;
    RECT 57.93 52.63 58.14 52.7 ;
    RECT 57.93 52.99 58.14 53.06 ;
    RECT 57.93 53.35 58.14 53.42 ;
    RECT 58.39 52.63 58.6 52.7 ;
    RECT 58.39 52.99 58.6 53.06 ;
    RECT 58.39 53.35 58.6 53.42 ;
    RECT 54.61 52.63 54.82 52.7 ;
    RECT 54.61 52.99 54.82 53.06 ;
    RECT 54.61 53.35 54.82 53.42 ;
    RECT 55.07 52.63 55.28 52.7 ;
    RECT 55.07 52.99 55.28 53.06 ;
    RECT 55.07 53.35 55.28 53.42 ;
    RECT 51.29 52.63 51.5 52.7 ;
    RECT 51.29 52.99 51.5 53.06 ;
    RECT 51.29 53.35 51.5 53.42 ;
    RECT 51.75 52.63 51.96 52.7 ;
    RECT 51.75 52.99 51.96 53.06 ;
    RECT 51.75 53.35 51.96 53.42 ;
    RECT 47.97 52.63 48.18 52.7 ;
    RECT 47.97 52.99 48.18 53.06 ;
    RECT 47.97 53.35 48.18 53.42 ;
    RECT 48.43 52.63 48.64 52.7 ;
    RECT 48.43 52.99 48.64 53.06 ;
    RECT 48.43 53.35 48.64 53.42 ;
    RECT 44.65 52.63 44.86 52.7 ;
    RECT 44.65 52.99 44.86 53.06 ;
    RECT 44.65 53.35 44.86 53.42 ;
    RECT 45.11 52.63 45.32 52.7 ;
    RECT 45.11 52.99 45.32 53.06 ;
    RECT 45.11 53.35 45.32 53.42 ;
    RECT 41.33 52.63 41.54 52.7 ;
    RECT 41.33 52.99 41.54 53.06 ;
    RECT 41.33 53.35 41.54 53.42 ;
    RECT 41.79 52.63 42.0 52.7 ;
    RECT 41.79 52.99 42.0 53.06 ;
    RECT 41.79 53.35 42.0 53.42 ;
    RECT 38.01 52.63 38.22 52.7 ;
    RECT 38.01 52.99 38.22 53.06 ;
    RECT 38.01 53.35 38.22 53.42 ;
    RECT 38.47 52.63 38.68 52.7 ;
    RECT 38.47 52.99 38.68 53.06 ;
    RECT 38.47 53.35 38.68 53.42 ;
    RECT 0.4 52.99 0.47 53.06 ;
    RECT 34.69 52.63 34.9 52.7 ;
    RECT 34.69 52.99 34.9 53.06 ;
    RECT 34.69 53.35 34.9 53.42 ;
    RECT 35.15 52.63 35.36 52.7 ;
    RECT 35.15 52.99 35.36 53.06 ;
    RECT 35.15 53.35 35.36 53.42 ;
    RECT 117.69 52.63 117.9 52.7 ;
    RECT 117.69 52.99 117.9 53.06 ;
    RECT 117.69 53.35 117.9 53.42 ;
    RECT 118.15 52.63 118.36 52.7 ;
    RECT 118.15 52.99 118.36 53.06 ;
    RECT 118.15 53.35 118.36 53.42 ;
    RECT 114.37 52.63 114.58 52.7 ;
    RECT 114.37 52.99 114.58 53.06 ;
    RECT 114.37 53.35 114.58 53.42 ;
    RECT 114.83 52.63 115.04 52.7 ;
    RECT 114.83 52.99 115.04 53.06 ;
    RECT 114.83 53.35 115.04 53.42 ;
    RECT 111.05 52.63 111.26 52.7 ;
    RECT 111.05 52.99 111.26 53.06 ;
    RECT 111.05 53.35 111.26 53.42 ;
    RECT 111.51 52.63 111.72 52.7 ;
    RECT 111.51 52.99 111.72 53.06 ;
    RECT 111.51 53.35 111.72 53.42 ;
    RECT 107.73 52.63 107.94 52.7 ;
    RECT 107.73 52.99 107.94 53.06 ;
    RECT 107.73 53.35 107.94 53.42 ;
    RECT 108.19 52.63 108.4 52.7 ;
    RECT 108.19 52.99 108.4 53.06 ;
    RECT 108.19 53.35 108.4 53.42 ;
    RECT 104.41 52.63 104.62 52.7 ;
    RECT 104.41 52.99 104.62 53.06 ;
    RECT 104.41 53.35 104.62 53.42 ;
    RECT 104.87 52.63 105.08 52.7 ;
    RECT 104.87 52.99 105.08 53.06 ;
    RECT 104.87 53.35 105.08 53.42 ;
    RECT 101.09 52.63 101.3 52.7 ;
    RECT 101.09 52.99 101.3 53.06 ;
    RECT 101.09 53.35 101.3 53.42 ;
    RECT 101.55 52.63 101.76 52.7 ;
    RECT 101.55 52.99 101.76 53.06 ;
    RECT 101.55 53.35 101.76 53.42 ;
    RECT 97.77 52.63 97.98 52.7 ;
    RECT 97.77 52.99 97.98 53.06 ;
    RECT 97.77 53.35 97.98 53.42 ;
    RECT 98.23 52.63 98.44 52.7 ;
    RECT 98.23 52.99 98.44 53.06 ;
    RECT 98.23 53.35 98.44 53.42 ;
    RECT 94.45 52.63 94.66 52.7 ;
    RECT 94.45 52.99 94.66 53.06 ;
    RECT 94.45 53.35 94.66 53.42 ;
    RECT 94.91 52.63 95.12 52.7 ;
    RECT 94.91 52.99 95.12 53.06 ;
    RECT 94.91 53.35 95.12 53.42 ;
    RECT 91.13 52.63 91.34 52.7 ;
    RECT 91.13 52.99 91.34 53.06 ;
    RECT 91.13 53.35 91.34 53.42 ;
    RECT 91.59 52.63 91.8 52.7 ;
    RECT 91.59 52.99 91.8 53.06 ;
    RECT 91.59 53.35 91.8 53.42 ;
    RECT 87.81 52.63 88.02 52.7 ;
    RECT 87.81 52.99 88.02 53.06 ;
    RECT 87.81 53.35 88.02 53.42 ;
    RECT 88.27 52.63 88.48 52.7 ;
    RECT 88.27 52.99 88.48 53.06 ;
    RECT 88.27 53.35 88.48 53.42 ;
    RECT 84.49 52.63 84.7 52.7 ;
    RECT 84.49 52.99 84.7 53.06 ;
    RECT 84.49 53.35 84.7 53.42 ;
    RECT 84.95 52.63 85.16 52.7 ;
    RECT 84.95 52.99 85.16 53.06 ;
    RECT 84.95 53.35 85.16 53.42 ;
    RECT 81.17 52.63 81.38 52.7 ;
    RECT 81.17 52.99 81.38 53.06 ;
    RECT 81.17 53.35 81.38 53.42 ;
    RECT 81.63 52.63 81.84 52.7 ;
    RECT 81.63 52.99 81.84 53.06 ;
    RECT 81.63 53.35 81.84 53.42 ;
    RECT 77.85 52.63 78.06 52.7 ;
    RECT 77.85 52.99 78.06 53.06 ;
    RECT 77.85 53.35 78.06 53.42 ;
    RECT 78.31 52.63 78.52 52.7 ;
    RECT 78.31 52.99 78.52 53.06 ;
    RECT 78.31 53.35 78.52 53.42 ;
    RECT 74.53 52.63 74.74 52.7 ;
    RECT 74.53 52.99 74.74 53.06 ;
    RECT 74.53 53.35 74.74 53.42 ;
    RECT 74.99 52.63 75.2 52.7 ;
    RECT 74.99 52.99 75.2 53.06 ;
    RECT 74.99 53.35 75.2 53.42 ;
    RECT 71.21 52.63 71.42 52.7 ;
    RECT 71.21 52.99 71.42 53.06 ;
    RECT 71.21 53.35 71.42 53.42 ;
    RECT 71.67 52.63 71.88 52.7 ;
    RECT 71.67 52.99 71.88 53.06 ;
    RECT 71.67 53.35 71.88 53.42 ;
    RECT 31.37 52.63 31.58 52.7 ;
    RECT 31.37 52.99 31.58 53.06 ;
    RECT 31.37 53.35 31.58 53.42 ;
    RECT 31.83 52.63 32.04 52.7 ;
    RECT 31.83 52.99 32.04 53.06 ;
    RECT 31.83 53.35 32.04 53.42 ;
    RECT 67.89 52.63 68.1 52.7 ;
    RECT 67.89 52.99 68.1 53.06 ;
    RECT 67.89 53.35 68.1 53.42 ;
    RECT 68.35 52.63 68.56 52.7 ;
    RECT 68.35 52.99 68.56 53.06 ;
    RECT 68.35 53.35 68.56 53.42 ;
    RECT 28.05 52.63 28.26 52.7 ;
    RECT 28.05 52.99 28.26 53.06 ;
    RECT 28.05 53.35 28.26 53.42 ;
    RECT 28.51 52.63 28.72 52.7 ;
    RECT 28.51 52.99 28.72 53.06 ;
    RECT 28.51 53.35 28.72 53.42 ;
    RECT 24.73 52.63 24.94 52.7 ;
    RECT 24.73 52.99 24.94 53.06 ;
    RECT 24.73 53.35 24.94 53.42 ;
    RECT 25.19 52.63 25.4 52.7 ;
    RECT 25.19 52.99 25.4 53.06 ;
    RECT 25.19 53.35 25.4 53.42 ;
    RECT 21.41 52.63 21.62 52.7 ;
    RECT 21.41 52.99 21.62 53.06 ;
    RECT 21.41 53.35 21.62 53.42 ;
    RECT 21.87 52.63 22.08 52.7 ;
    RECT 21.87 52.99 22.08 53.06 ;
    RECT 21.87 53.35 22.08 53.42 ;
    RECT 18.09 52.63 18.3 52.7 ;
    RECT 18.09 52.99 18.3 53.06 ;
    RECT 18.09 53.35 18.3 53.42 ;
    RECT 18.55 52.63 18.76 52.7 ;
    RECT 18.55 52.99 18.76 53.06 ;
    RECT 18.55 53.35 18.76 53.42 ;
    RECT 120.825 52.99 120.895 53.06 ;
    RECT 14.77 52.63 14.98 52.7 ;
    RECT 14.77 52.99 14.98 53.06 ;
    RECT 14.77 53.35 14.98 53.42 ;
    RECT 15.23 52.63 15.44 52.7 ;
    RECT 15.23 52.99 15.44 53.06 ;
    RECT 15.23 53.35 15.44 53.42 ;
    RECT 11.45 52.63 11.66 52.7 ;
    RECT 11.45 52.99 11.66 53.06 ;
    RECT 11.45 53.35 11.66 53.42 ;
    RECT 11.91 52.63 12.12 52.7 ;
    RECT 11.91 52.99 12.12 53.06 ;
    RECT 11.91 53.35 12.12 53.42 ;
    RECT 8.13 52.63 8.34 52.7 ;
    RECT 8.13 52.99 8.34 53.06 ;
    RECT 8.13 53.35 8.34 53.42 ;
    RECT 8.59 52.63 8.8 52.7 ;
    RECT 8.59 52.99 8.8 53.06 ;
    RECT 8.59 53.35 8.8 53.42 ;
    RECT 4.81 52.63 5.02 52.7 ;
    RECT 4.81 52.99 5.02 53.06 ;
    RECT 4.81 53.35 5.02 53.42 ;
    RECT 5.27 52.63 5.48 52.7 ;
    RECT 5.27 52.99 5.48 53.06 ;
    RECT 5.27 53.35 5.48 53.42 ;
    RECT 1.49 52.63 1.7 52.7 ;
    RECT 1.49 52.99 1.7 53.06 ;
    RECT 1.49 53.35 1.7 53.42 ;
    RECT 1.95 52.63 2.16 52.7 ;
    RECT 1.95 52.99 2.16 53.06 ;
    RECT 1.95 53.35 2.16 53.42 ;
    RECT 64.57 52.63 64.78 52.7 ;
    RECT 64.57 52.99 64.78 53.06 ;
    RECT 64.57 53.35 64.78 53.42 ;
    RECT 65.03 52.63 65.24 52.7 ;
    RECT 65.03 52.99 65.24 53.06 ;
    RECT 65.03 53.35 65.24 53.42 ;
    RECT 61.25 51.91 61.46 51.98 ;
    RECT 61.25 52.27 61.46 52.34 ;
    RECT 61.25 52.63 61.46 52.7 ;
    RECT 61.71 51.91 61.92 51.98 ;
    RECT 61.71 52.27 61.92 52.34 ;
    RECT 61.71 52.63 61.92 52.7 ;
    RECT 57.93 51.91 58.14 51.98 ;
    RECT 57.93 52.27 58.14 52.34 ;
    RECT 57.93 52.63 58.14 52.7 ;
    RECT 58.39 51.91 58.6 51.98 ;
    RECT 58.39 52.27 58.6 52.34 ;
    RECT 58.39 52.63 58.6 52.7 ;
    RECT 54.61 51.91 54.82 51.98 ;
    RECT 54.61 52.27 54.82 52.34 ;
    RECT 54.61 52.63 54.82 52.7 ;
    RECT 55.07 51.91 55.28 51.98 ;
    RECT 55.07 52.27 55.28 52.34 ;
    RECT 55.07 52.63 55.28 52.7 ;
    RECT 51.29 51.91 51.5 51.98 ;
    RECT 51.29 52.27 51.5 52.34 ;
    RECT 51.29 52.63 51.5 52.7 ;
    RECT 51.75 51.91 51.96 51.98 ;
    RECT 51.75 52.27 51.96 52.34 ;
    RECT 51.75 52.63 51.96 52.7 ;
    RECT 47.97 51.91 48.18 51.98 ;
    RECT 47.97 52.27 48.18 52.34 ;
    RECT 47.97 52.63 48.18 52.7 ;
    RECT 48.43 51.91 48.64 51.98 ;
    RECT 48.43 52.27 48.64 52.34 ;
    RECT 48.43 52.63 48.64 52.7 ;
    RECT 44.65 51.91 44.86 51.98 ;
    RECT 44.65 52.27 44.86 52.34 ;
    RECT 44.65 52.63 44.86 52.7 ;
    RECT 45.11 51.91 45.32 51.98 ;
    RECT 45.11 52.27 45.32 52.34 ;
    RECT 45.11 52.63 45.32 52.7 ;
    RECT 41.33 51.91 41.54 51.98 ;
    RECT 41.33 52.27 41.54 52.34 ;
    RECT 41.33 52.63 41.54 52.7 ;
    RECT 41.79 51.91 42.0 51.98 ;
    RECT 41.79 52.27 42.0 52.34 ;
    RECT 41.79 52.63 42.0 52.7 ;
    RECT 38.01 51.91 38.22 51.98 ;
    RECT 38.01 52.27 38.22 52.34 ;
    RECT 38.01 52.63 38.22 52.7 ;
    RECT 38.47 51.91 38.68 51.98 ;
    RECT 38.47 52.27 38.68 52.34 ;
    RECT 38.47 52.63 38.68 52.7 ;
    RECT 0.4 52.27 0.47 52.34 ;
    RECT 34.69 51.91 34.9 51.98 ;
    RECT 34.69 52.27 34.9 52.34 ;
    RECT 34.69 52.63 34.9 52.7 ;
    RECT 35.15 51.91 35.36 51.98 ;
    RECT 35.15 52.27 35.36 52.34 ;
    RECT 35.15 52.63 35.36 52.7 ;
    RECT 117.69 51.91 117.9 51.98 ;
    RECT 117.69 52.27 117.9 52.34 ;
    RECT 117.69 52.63 117.9 52.7 ;
    RECT 118.15 51.91 118.36 51.98 ;
    RECT 118.15 52.27 118.36 52.34 ;
    RECT 118.15 52.63 118.36 52.7 ;
    RECT 114.37 51.91 114.58 51.98 ;
    RECT 114.37 52.27 114.58 52.34 ;
    RECT 114.37 52.63 114.58 52.7 ;
    RECT 114.83 51.91 115.04 51.98 ;
    RECT 114.83 52.27 115.04 52.34 ;
    RECT 114.83 52.63 115.04 52.7 ;
    RECT 111.05 51.91 111.26 51.98 ;
    RECT 111.05 52.27 111.26 52.34 ;
    RECT 111.05 52.63 111.26 52.7 ;
    RECT 111.51 51.91 111.72 51.98 ;
    RECT 111.51 52.27 111.72 52.34 ;
    RECT 111.51 52.63 111.72 52.7 ;
    RECT 107.73 51.91 107.94 51.98 ;
    RECT 107.73 52.27 107.94 52.34 ;
    RECT 107.73 52.63 107.94 52.7 ;
    RECT 108.19 51.91 108.4 51.98 ;
    RECT 108.19 52.27 108.4 52.34 ;
    RECT 108.19 52.63 108.4 52.7 ;
    RECT 104.41 51.91 104.62 51.98 ;
    RECT 104.41 52.27 104.62 52.34 ;
    RECT 104.41 52.63 104.62 52.7 ;
    RECT 104.87 51.91 105.08 51.98 ;
    RECT 104.87 52.27 105.08 52.34 ;
    RECT 104.87 52.63 105.08 52.7 ;
    RECT 101.09 51.91 101.3 51.98 ;
    RECT 101.09 52.27 101.3 52.34 ;
    RECT 101.09 52.63 101.3 52.7 ;
    RECT 101.55 51.91 101.76 51.98 ;
    RECT 101.55 52.27 101.76 52.34 ;
    RECT 101.55 52.63 101.76 52.7 ;
    RECT 97.77 51.91 97.98 51.98 ;
    RECT 97.77 52.27 97.98 52.34 ;
    RECT 97.77 52.63 97.98 52.7 ;
    RECT 98.23 51.91 98.44 51.98 ;
    RECT 98.23 52.27 98.44 52.34 ;
    RECT 98.23 52.63 98.44 52.7 ;
    RECT 94.45 51.91 94.66 51.98 ;
    RECT 94.45 52.27 94.66 52.34 ;
    RECT 94.45 52.63 94.66 52.7 ;
    RECT 94.91 51.91 95.12 51.98 ;
    RECT 94.91 52.27 95.12 52.34 ;
    RECT 94.91 52.63 95.12 52.7 ;
    RECT 91.13 51.91 91.34 51.98 ;
    RECT 91.13 52.27 91.34 52.34 ;
    RECT 91.13 52.63 91.34 52.7 ;
    RECT 91.59 51.91 91.8 51.98 ;
    RECT 91.59 52.27 91.8 52.34 ;
    RECT 91.59 52.63 91.8 52.7 ;
    RECT 87.81 51.91 88.02 51.98 ;
    RECT 87.81 52.27 88.02 52.34 ;
    RECT 87.81 52.63 88.02 52.7 ;
    RECT 88.27 51.91 88.48 51.98 ;
    RECT 88.27 52.27 88.48 52.34 ;
    RECT 88.27 52.63 88.48 52.7 ;
    RECT 84.49 51.91 84.7 51.98 ;
    RECT 84.49 52.27 84.7 52.34 ;
    RECT 84.49 52.63 84.7 52.7 ;
    RECT 84.95 51.91 85.16 51.98 ;
    RECT 84.95 52.27 85.16 52.34 ;
    RECT 84.95 52.63 85.16 52.7 ;
    RECT 81.17 51.91 81.38 51.98 ;
    RECT 81.17 52.27 81.38 52.34 ;
    RECT 81.17 52.63 81.38 52.7 ;
    RECT 81.63 51.91 81.84 51.98 ;
    RECT 81.63 52.27 81.84 52.34 ;
    RECT 81.63 52.63 81.84 52.7 ;
    RECT 77.85 51.91 78.06 51.98 ;
    RECT 77.85 52.27 78.06 52.34 ;
    RECT 77.85 52.63 78.06 52.7 ;
    RECT 78.31 51.91 78.52 51.98 ;
    RECT 78.31 52.27 78.52 52.34 ;
    RECT 78.31 52.63 78.52 52.7 ;
    RECT 74.53 51.91 74.74 51.98 ;
    RECT 74.53 52.27 74.74 52.34 ;
    RECT 74.53 52.63 74.74 52.7 ;
    RECT 74.99 51.91 75.2 51.98 ;
    RECT 74.99 52.27 75.2 52.34 ;
    RECT 74.99 52.63 75.2 52.7 ;
    RECT 71.21 51.91 71.42 51.98 ;
    RECT 71.21 52.27 71.42 52.34 ;
    RECT 71.21 52.63 71.42 52.7 ;
    RECT 71.67 51.91 71.88 51.98 ;
    RECT 71.67 52.27 71.88 52.34 ;
    RECT 71.67 52.63 71.88 52.7 ;
    RECT 31.37 51.91 31.58 51.98 ;
    RECT 31.37 52.27 31.58 52.34 ;
    RECT 31.37 52.63 31.58 52.7 ;
    RECT 31.83 51.91 32.04 51.98 ;
    RECT 31.83 52.27 32.04 52.34 ;
    RECT 31.83 52.63 32.04 52.7 ;
    RECT 67.89 51.91 68.1 51.98 ;
    RECT 67.89 52.27 68.1 52.34 ;
    RECT 67.89 52.63 68.1 52.7 ;
    RECT 68.35 51.91 68.56 51.98 ;
    RECT 68.35 52.27 68.56 52.34 ;
    RECT 68.35 52.63 68.56 52.7 ;
    RECT 28.05 51.91 28.26 51.98 ;
    RECT 28.05 52.27 28.26 52.34 ;
    RECT 28.05 52.63 28.26 52.7 ;
    RECT 28.51 51.91 28.72 51.98 ;
    RECT 28.51 52.27 28.72 52.34 ;
    RECT 28.51 52.63 28.72 52.7 ;
    RECT 24.73 51.91 24.94 51.98 ;
    RECT 24.73 52.27 24.94 52.34 ;
    RECT 24.73 52.63 24.94 52.7 ;
    RECT 25.19 51.91 25.4 51.98 ;
    RECT 25.19 52.27 25.4 52.34 ;
    RECT 25.19 52.63 25.4 52.7 ;
    RECT 21.41 51.91 21.62 51.98 ;
    RECT 21.41 52.27 21.62 52.34 ;
    RECT 21.41 52.63 21.62 52.7 ;
    RECT 21.87 51.91 22.08 51.98 ;
    RECT 21.87 52.27 22.08 52.34 ;
    RECT 21.87 52.63 22.08 52.7 ;
    RECT 18.09 51.91 18.3 51.98 ;
    RECT 18.09 52.27 18.3 52.34 ;
    RECT 18.09 52.63 18.3 52.7 ;
    RECT 18.55 51.91 18.76 51.98 ;
    RECT 18.55 52.27 18.76 52.34 ;
    RECT 18.55 52.63 18.76 52.7 ;
    RECT 120.825 52.27 120.895 52.34 ;
    RECT 14.77 51.91 14.98 51.98 ;
    RECT 14.77 52.27 14.98 52.34 ;
    RECT 14.77 52.63 14.98 52.7 ;
    RECT 15.23 51.91 15.44 51.98 ;
    RECT 15.23 52.27 15.44 52.34 ;
    RECT 15.23 52.63 15.44 52.7 ;
    RECT 11.45 51.91 11.66 51.98 ;
    RECT 11.45 52.27 11.66 52.34 ;
    RECT 11.45 52.63 11.66 52.7 ;
    RECT 11.91 51.91 12.12 51.98 ;
    RECT 11.91 52.27 12.12 52.34 ;
    RECT 11.91 52.63 12.12 52.7 ;
    RECT 8.13 51.91 8.34 51.98 ;
    RECT 8.13 52.27 8.34 52.34 ;
    RECT 8.13 52.63 8.34 52.7 ;
    RECT 8.59 51.91 8.8 51.98 ;
    RECT 8.59 52.27 8.8 52.34 ;
    RECT 8.59 52.63 8.8 52.7 ;
    RECT 4.81 51.91 5.02 51.98 ;
    RECT 4.81 52.27 5.02 52.34 ;
    RECT 4.81 52.63 5.02 52.7 ;
    RECT 5.27 51.91 5.48 51.98 ;
    RECT 5.27 52.27 5.48 52.34 ;
    RECT 5.27 52.63 5.48 52.7 ;
    RECT 1.49 51.91 1.7 51.98 ;
    RECT 1.49 52.27 1.7 52.34 ;
    RECT 1.49 52.63 1.7 52.7 ;
    RECT 1.95 51.91 2.16 51.98 ;
    RECT 1.95 52.27 2.16 52.34 ;
    RECT 1.95 52.63 2.16 52.7 ;
    RECT 64.57 51.91 64.78 51.98 ;
    RECT 64.57 52.27 64.78 52.34 ;
    RECT 64.57 52.63 64.78 52.7 ;
    RECT 65.03 51.91 65.24 51.98 ;
    RECT 65.03 52.27 65.24 52.34 ;
    RECT 65.03 52.63 65.24 52.7 ;
    RECT 61.25 51.19 61.46 51.26 ;
    RECT 61.25 51.55 61.46 51.62 ;
    RECT 61.25 51.91 61.46 51.98 ;
    RECT 61.71 51.19 61.92 51.26 ;
    RECT 61.71 51.55 61.92 51.62 ;
    RECT 61.71 51.91 61.92 51.98 ;
    RECT 57.93 51.19 58.14 51.26 ;
    RECT 57.93 51.55 58.14 51.62 ;
    RECT 57.93 51.91 58.14 51.98 ;
    RECT 58.39 51.19 58.6 51.26 ;
    RECT 58.39 51.55 58.6 51.62 ;
    RECT 58.39 51.91 58.6 51.98 ;
    RECT 54.61 51.19 54.82 51.26 ;
    RECT 54.61 51.55 54.82 51.62 ;
    RECT 54.61 51.91 54.82 51.98 ;
    RECT 55.07 51.19 55.28 51.26 ;
    RECT 55.07 51.55 55.28 51.62 ;
    RECT 55.07 51.91 55.28 51.98 ;
    RECT 51.29 51.19 51.5 51.26 ;
    RECT 51.29 51.55 51.5 51.62 ;
    RECT 51.29 51.91 51.5 51.98 ;
    RECT 51.75 51.19 51.96 51.26 ;
    RECT 51.75 51.55 51.96 51.62 ;
    RECT 51.75 51.91 51.96 51.98 ;
    RECT 47.97 51.19 48.18 51.26 ;
    RECT 47.97 51.55 48.18 51.62 ;
    RECT 47.97 51.91 48.18 51.98 ;
    RECT 48.43 51.19 48.64 51.26 ;
    RECT 48.43 51.55 48.64 51.62 ;
    RECT 48.43 51.91 48.64 51.98 ;
    RECT 44.65 51.19 44.86 51.26 ;
    RECT 44.65 51.55 44.86 51.62 ;
    RECT 44.65 51.91 44.86 51.98 ;
    RECT 45.11 51.19 45.32 51.26 ;
    RECT 45.11 51.55 45.32 51.62 ;
    RECT 45.11 51.91 45.32 51.98 ;
    RECT 41.33 51.19 41.54 51.26 ;
    RECT 41.33 51.55 41.54 51.62 ;
    RECT 41.33 51.91 41.54 51.98 ;
    RECT 41.79 51.19 42.0 51.26 ;
    RECT 41.79 51.55 42.0 51.62 ;
    RECT 41.79 51.91 42.0 51.98 ;
    RECT 38.01 51.19 38.22 51.26 ;
    RECT 38.01 51.55 38.22 51.62 ;
    RECT 38.01 51.91 38.22 51.98 ;
    RECT 38.47 51.19 38.68 51.26 ;
    RECT 38.47 51.55 38.68 51.62 ;
    RECT 38.47 51.91 38.68 51.98 ;
    RECT 0.4 51.55 0.47 51.62 ;
    RECT 34.69 51.19 34.9 51.26 ;
    RECT 34.69 51.55 34.9 51.62 ;
    RECT 34.69 51.91 34.9 51.98 ;
    RECT 35.15 51.19 35.36 51.26 ;
    RECT 35.15 51.55 35.36 51.62 ;
    RECT 35.15 51.91 35.36 51.98 ;
    RECT 117.69 51.19 117.9 51.26 ;
    RECT 117.69 51.55 117.9 51.62 ;
    RECT 117.69 51.91 117.9 51.98 ;
    RECT 118.15 51.19 118.36 51.26 ;
    RECT 118.15 51.55 118.36 51.62 ;
    RECT 118.15 51.91 118.36 51.98 ;
    RECT 114.37 51.19 114.58 51.26 ;
    RECT 114.37 51.55 114.58 51.62 ;
    RECT 114.37 51.91 114.58 51.98 ;
    RECT 114.83 51.19 115.04 51.26 ;
    RECT 114.83 51.55 115.04 51.62 ;
    RECT 114.83 51.91 115.04 51.98 ;
    RECT 111.05 51.19 111.26 51.26 ;
    RECT 111.05 51.55 111.26 51.62 ;
    RECT 111.05 51.91 111.26 51.98 ;
    RECT 111.51 51.19 111.72 51.26 ;
    RECT 111.51 51.55 111.72 51.62 ;
    RECT 111.51 51.91 111.72 51.98 ;
    RECT 107.73 51.19 107.94 51.26 ;
    RECT 107.73 51.55 107.94 51.62 ;
    RECT 107.73 51.91 107.94 51.98 ;
    RECT 108.19 51.19 108.4 51.26 ;
    RECT 108.19 51.55 108.4 51.62 ;
    RECT 108.19 51.91 108.4 51.98 ;
    RECT 104.41 51.19 104.62 51.26 ;
    RECT 104.41 51.55 104.62 51.62 ;
    RECT 104.41 51.91 104.62 51.98 ;
    RECT 104.87 51.19 105.08 51.26 ;
    RECT 104.87 51.55 105.08 51.62 ;
    RECT 104.87 51.91 105.08 51.98 ;
    RECT 101.09 51.19 101.3 51.26 ;
    RECT 101.09 51.55 101.3 51.62 ;
    RECT 101.09 51.91 101.3 51.98 ;
    RECT 101.55 51.19 101.76 51.26 ;
    RECT 101.55 51.55 101.76 51.62 ;
    RECT 101.55 51.91 101.76 51.98 ;
    RECT 97.77 51.19 97.98 51.26 ;
    RECT 97.77 51.55 97.98 51.62 ;
    RECT 97.77 51.91 97.98 51.98 ;
    RECT 98.23 51.19 98.44 51.26 ;
    RECT 98.23 51.55 98.44 51.62 ;
    RECT 98.23 51.91 98.44 51.98 ;
    RECT 94.45 51.19 94.66 51.26 ;
    RECT 94.45 51.55 94.66 51.62 ;
    RECT 94.45 51.91 94.66 51.98 ;
    RECT 94.91 51.19 95.12 51.26 ;
    RECT 94.91 51.55 95.12 51.62 ;
    RECT 94.91 51.91 95.12 51.98 ;
    RECT 91.13 51.19 91.34 51.26 ;
    RECT 91.13 51.55 91.34 51.62 ;
    RECT 91.13 51.91 91.34 51.98 ;
    RECT 91.59 51.19 91.8 51.26 ;
    RECT 91.59 51.55 91.8 51.62 ;
    RECT 91.59 51.91 91.8 51.98 ;
    RECT 87.81 51.19 88.02 51.26 ;
    RECT 87.81 51.55 88.02 51.62 ;
    RECT 87.81 51.91 88.02 51.98 ;
    RECT 88.27 51.19 88.48 51.26 ;
    RECT 88.27 51.55 88.48 51.62 ;
    RECT 88.27 51.91 88.48 51.98 ;
    RECT 84.49 51.19 84.7 51.26 ;
    RECT 84.49 51.55 84.7 51.62 ;
    RECT 84.49 51.91 84.7 51.98 ;
    RECT 84.95 51.19 85.16 51.26 ;
    RECT 84.95 51.55 85.16 51.62 ;
    RECT 84.95 51.91 85.16 51.98 ;
    RECT 81.17 51.19 81.38 51.26 ;
    RECT 81.17 51.55 81.38 51.62 ;
    RECT 81.17 51.91 81.38 51.98 ;
    RECT 81.63 51.19 81.84 51.26 ;
    RECT 81.63 51.55 81.84 51.62 ;
    RECT 81.63 51.91 81.84 51.98 ;
    RECT 77.85 51.19 78.06 51.26 ;
    RECT 77.85 51.55 78.06 51.62 ;
    RECT 77.85 51.91 78.06 51.98 ;
    RECT 78.31 51.19 78.52 51.26 ;
    RECT 78.31 51.55 78.52 51.62 ;
    RECT 78.31 51.91 78.52 51.98 ;
    RECT 74.53 51.19 74.74 51.26 ;
    RECT 74.53 51.55 74.74 51.62 ;
    RECT 74.53 51.91 74.74 51.98 ;
    RECT 74.99 51.19 75.2 51.26 ;
    RECT 74.99 51.55 75.2 51.62 ;
    RECT 74.99 51.91 75.2 51.98 ;
    RECT 71.21 51.19 71.42 51.26 ;
    RECT 71.21 51.55 71.42 51.62 ;
    RECT 71.21 51.91 71.42 51.98 ;
    RECT 71.67 51.19 71.88 51.26 ;
    RECT 71.67 51.55 71.88 51.62 ;
    RECT 71.67 51.91 71.88 51.98 ;
    RECT 31.37 51.19 31.58 51.26 ;
    RECT 31.37 51.55 31.58 51.62 ;
    RECT 31.37 51.91 31.58 51.98 ;
    RECT 31.83 51.19 32.04 51.26 ;
    RECT 31.83 51.55 32.04 51.62 ;
    RECT 31.83 51.91 32.04 51.98 ;
    RECT 67.89 51.19 68.1 51.26 ;
    RECT 67.89 51.55 68.1 51.62 ;
    RECT 67.89 51.91 68.1 51.98 ;
    RECT 68.35 51.19 68.56 51.26 ;
    RECT 68.35 51.55 68.56 51.62 ;
    RECT 68.35 51.91 68.56 51.98 ;
    RECT 28.05 51.19 28.26 51.26 ;
    RECT 28.05 51.55 28.26 51.62 ;
    RECT 28.05 51.91 28.26 51.98 ;
    RECT 28.51 51.19 28.72 51.26 ;
    RECT 28.51 51.55 28.72 51.62 ;
    RECT 28.51 51.91 28.72 51.98 ;
    RECT 24.73 51.19 24.94 51.26 ;
    RECT 24.73 51.55 24.94 51.62 ;
    RECT 24.73 51.91 24.94 51.98 ;
    RECT 25.19 51.19 25.4 51.26 ;
    RECT 25.19 51.55 25.4 51.62 ;
    RECT 25.19 51.91 25.4 51.98 ;
    RECT 21.41 51.19 21.62 51.26 ;
    RECT 21.41 51.55 21.62 51.62 ;
    RECT 21.41 51.91 21.62 51.98 ;
    RECT 21.87 51.19 22.08 51.26 ;
    RECT 21.87 51.55 22.08 51.62 ;
    RECT 21.87 51.91 22.08 51.98 ;
    RECT 18.09 51.19 18.3 51.26 ;
    RECT 18.09 51.55 18.3 51.62 ;
    RECT 18.09 51.91 18.3 51.98 ;
    RECT 18.55 51.19 18.76 51.26 ;
    RECT 18.55 51.55 18.76 51.62 ;
    RECT 18.55 51.91 18.76 51.98 ;
    RECT 120.825 51.55 120.895 51.62 ;
    RECT 14.77 51.19 14.98 51.26 ;
    RECT 14.77 51.55 14.98 51.62 ;
    RECT 14.77 51.91 14.98 51.98 ;
    RECT 15.23 51.19 15.44 51.26 ;
    RECT 15.23 51.55 15.44 51.62 ;
    RECT 15.23 51.91 15.44 51.98 ;
    RECT 11.45 51.19 11.66 51.26 ;
    RECT 11.45 51.55 11.66 51.62 ;
    RECT 11.45 51.91 11.66 51.98 ;
    RECT 11.91 51.19 12.12 51.26 ;
    RECT 11.91 51.55 12.12 51.62 ;
    RECT 11.91 51.91 12.12 51.98 ;
    RECT 8.13 51.19 8.34 51.26 ;
    RECT 8.13 51.55 8.34 51.62 ;
    RECT 8.13 51.91 8.34 51.98 ;
    RECT 8.59 51.19 8.8 51.26 ;
    RECT 8.59 51.55 8.8 51.62 ;
    RECT 8.59 51.91 8.8 51.98 ;
    RECT 4.81 51.19 5.02 51.26 ;
    RECT 4.81 51.55 5.02 51.62 ;
    RECT 4.81 51.91 5.02 51.98 ;
    RECT 5.27 51.19 5.48 51.26 ;
    RECT 5.27 51.55 5.48 51.62 ;
    RECT 5.27 51.91 5.48 51.98 ;
    RECT 1.49 51.19 1.7 51.26 ;
    RECT 1.49 51.55 1.7 51.62 ;
    RECT 1.49 51.91 1.7 51.98 ;
    RECT 1.95 51.19 2.16 51.26 ;
    RECT 1.95 51.55 2.16 51.62 ;
    RECT 1.95 51.91 2.16 51.98 ;
    RECT 64.57 51.19 64.78 51.26 ;
    RECT 64.57 51.55 64.78 51.62 ;
    RECT 64.57 51.91 64.78 51.98 ;
    RECT 65.03 51.19 65.24 51.26 ;
    RECT 65.03 51.55 65.24 51.62 ;
    RECT 65.03 51.91 65.24 51.98 ;
    RECT 61.25 50.47 61.46 50.54 ;
    RECT 61.25 50.83 61.46 50.9 ;
    RECT 61.25 51.19 61.46 51.26 ;
    RECT 61.71 50.47 61.92 50.54 ;
    RECT 61.71 50.83 61.92 50.9 ;
    RECT 61.71 51.19 61.92 51.26 ;
    RECT 57.93 50.47 58.14 50.54 ;
    RECT 57.93 50.83 58.14 50.9 ;
    RECT 57.93 51.19 58.14 51.26 ;
    RECT 58.39 50.47 58.6 50.54 ;
    RECT 58.39 50.83 58.6 50.9 ;
    RECT 58.39 51.19 58.6 51.26 ;
    RECT 54.61 50.47 54.82 50.54 ;
    RECT 54.61 50.83 54.82 50.9 ;
    RECT 54.61 51.19 54.82 51.26 ;
    RECT 55.07 50.47 55.28 50.54 ;
    RECT 55.07 50.83 55.28 50.9 ;
    RECT 55.07 51.19 55.28 51.26 ;
    RECT 51.29 50.47 51.5 50.54 ;
    RECT 51.29 50.83 51.5 50.9 ;
    RECT 51.29 51.19 51.5 51.26 ;
    RECT 51.75 50.47 51.96 50.54 ;
    RECT 51.75 50.83 51.96 50.9 ;
    RECT 51.75 51.19 51.96 51.26 ;
    RECT 47.97 50.47 48.18 50.54 ;
    RECT 47.97 50.83 48.18 50.9 ;
    RECT 47.97 51.19 48.18 51.26 ;
    RECT 48.43 50.47 48.64 50.54 ;
    RECT 48.43 50.83 48.64 50.9 ;
    RECT 48.43 51.19 48.64 51.26 ;
    RECT 44.65 50.47 44.86 50.54 ;
    RECT 44.65 50.83 44.86 50.9 ;
    RECT 44.65 51.19 44.86 51.26 ;
    RECT 45.11 50.47 45.32 50.54 ;
    RECT 45.11 50.83 45.32 50.9 ;
    RECT 45.11 51.19 45.32 51.26 ;
    RECT 41.33 50.47 41.54 50.54 ;
    RECT 41.33 50.83 41.54 50.9 ;
    RECT 41.33 51.19 41.54 51.26 ;
    RECT 41.79 50.47 42.0 50.54 ;
    RECT 41.79 50.83 42.0 50.9 ;
    RECT 41.79 51.19 42.0 51.26 ;
    RECT 38.01 50.47 38.22 50.54 ;
    RECT 38.01 50.83 38.22 50.9 ;
    RECT 38.01 51.19 38.22 51.26 ;
    RECT 38.47 50.47 38.68 50.54 ;
    RECT 38.47 50.83 38.68 50.9 ;
    RECT 38.47 51.19 38.68 51.26 ;
    RECT 0.4 50.83 0.47 50.9 ;
    RECT 34.69 50.47 34.9 50.54 ;
    RECT 34.69 50.83 34.9 50.9 ;
    RECT 34.69 51.19 34.9 51.26 ;
    RECT 35.15 50.47 35.36 50.54 ;
    RECT 35.15 50.83 35.36 50.9 ;
    RECT 35.15 51.19 35.36 51.26 ;
    RECT 117.69 50.47 117.9 50.54 ;
    RECT 117.69 50.83 117.9 50.9 ;
    RECT 117.69 51.19 117.9 51.26 ;
    RECT 118.15 50.47 118.36 50.54 ;
    RECT 118.15 50.83 118.36 50.9 ;
    RECT 118.15 51.19 118.36 51.26 ;
    RECT 114.37 50.47 114.58 50.54 ;
    RECT 114.37 50.83 114.58 50.9 ;
    RECT 114.37 51.19 114.58 51.26 ;
    RECT 114.83 50.47 115.04 50.54 ;
    RECT 114.83 50.83 115.04 50.9 ;
    RECT 114.83 51.19 115.04 51.26 ;
    RECT 111.05 50.47 111.26 50.54 ;
    RECT 111.05 50.83 111.26 50.9 ;
    RECT 111.05 51.19 111.26 51.26 ;
    RECT 111.51 50.47 111.72 50.54 ;
    RECT 111.51 50.83 111.72 50.9 ;
    RECT 111.51 51.19 111.72 51.26 ;
    RECT 107.73 50.47 107.94 50.54 ;
    RECT 107.73 50.83 107.94 50.9 ;
    RECT 107.73 51.19 107.94 51.26 ;
    RECT 108.19 50.47 108.4 50.54 ;
    RECT 108.19 50.83 108.4 50.9 ;
    RECT 108.19 51.19 108.4 51.26 ;
    RECT 104.41 50.47 104.62 50.54 ;
    RECT 104.41 50.83 104.62 50.9 ;
    RECT 104.41 51.19 104.62 51.26 ;
    RECT 104.87 50.47 105.08 50.54 ;
    RECT 104.87 50.83 105.08 50.9 ;
    RECT 104.87 51.19 105.08 51.26 ;
    RECT 101.09 50.47 101.3 50.54 ;
    RECT 101.09 50.83 101.3 50.9 ;
    RECT 101.09 51.19 101.3 51.26 ;
    RECT 101.55 50.47 101.76 50.54 ;
    RECT 101.55 50.83 101.76 50.9 ;
    RECT 101.55 51.19 101.76 51.26 ;
    RECT 97.77 50.47 97.98 50.54 ;
    RECT 97.77 50.83 97.98 50.9 ;
    RECT 97.77 51.19 97.98 51.26 ;
    RECT 98.23 50.47 98.44 50.54 ;
    RECT 98.23 50.83 98.44 50.9 ;
    RECT 98.23 51.19 98.44 51.26 ;
    RECT 94.45 50.47 94.66 50.54 ;
    RECT 94.45 50.83 94.66 50.9 ;
    RECT 94.45 51.19 94.66 51.26 ;
    RECT 94.91 50.47 95.12 50.54 ;
    RECT 94.91 50.83 95.12 50.9 ;
    RECT 94.91 51.19 95.12 51.26 ;
    RECT 91.13 50.47 91.34 50.54 ;
    RECT 91.13 50.83 91.34 50.9 ;
    RECT 91.13 51.19 91.34 51.26 ;
    RECT 91.59 50.47 91.8 50.54 ;
    RECT 91.59 50.83 91.8 50.9 ;
    RECT 91.59 51.19 91.8 51.26 ;
    RECT 87.81 50.47 88.02 50.54 ;
    RECT 87.81 50.83 88.02 50.9 ;
    RECT 87.81 51.19 88.02 51.26 ;
    RECT 88.27 50.47 88.48 50.54 ;
    RECT 88.27 50.83 88.48 50.9 ;
    RECT 88.27 51.19 88.48 51.26 ;
    RECT 84.49 50.47 84.7 50.54 ;
    RECT 84.49 50.83 84.7 50.9 ;
    RECT 84.49 51.19 84.7 51.26 ;
    RECT 84.95 50.47 85.16 50.54 ;
    RECT 84.95 50.83 85.16 50.9 ;
    RECT 84.95 51.19 85.16 51.26 ;
    RECT 81.17 50.47 81.38 50.54 ;
    RECT 81.17 50.83 81.38 50.9 ;
    RECT 81.17 51.19 81.38 51.26 ;
    RECT 81.63 50.47 81.84 50.54 ;
    RECT 81.63 50.83 81.84 50.9 ;
    RECT 81.63 51.19 81.84 51.26 ;
    RECT 77.85 50.47 78.06 50.54 ;
    RECT 77.85 50.83 78.06 50.9 ;
    RECT 77.85 51.19 78.06 51.26 ;
    RECT 78.31 50.47 78.52 50.54 ;
    RECT 78.31 50.83 78.52 50.9 ;
    RECT 78.31 51.19 78.52 51.26 ;
    RECT 74.53 50.47 74.74 50.54 ;
    RECT 74.53 50.83 74.74 50.9 ;
    RECT 74.53 51.19 74.74 51.26 ;
    RECT 74.99 50.47 75.2 50.54 ;
    RECT 74.99 50.83 75.2 50.9 ;
    RECT 74.99 51.19 75.2 51.26 ;
    RECT 71.21 50.47 71.42 50.54 ;
    RECT 71.21 50.83 71.42 50.9 ;
    RECT 71.21 51.19 71.42 51.26 ;
    RECT 71.67 50.47 71.88 50.54 ;
    RECT 71.67 50.83 71.88 50.9 ;
    RECT 71.67 51.19 71.88 51.26 ;
    RECT 31.37 50.47 31.58 50.54 ;
    RECT 31.37 50.83 31.58 50.9 ;
    RECT 31.37 51.19 31.58 51.26 ;
    RECT 31.83 50.47 32.04 50.54 ;
    RECT 31.83 50.83 32.04 50.9 ;
    RECT 31.83 51.19 32.04 51.26 ;
    RECT 67.89 50.47 68.1 50.54 ;
    RECT 67.89 50.83 68.1 50.9 ;
    RECT 67.89 51.19 68.1 51.26 ;
    RECT 68.35 50.47 68.56 50.54 ;
    RECT 68.35 50.83 68.56 50.9 ;
    RECT 68.35 51.19 68.56 51.26 ;
    RECT 28.05 50.47 28.26 50.54 ;
    RECT 28.05 50.83 28.26 50.9 ;
    RECT 28.05 51.19 28.26 51.26 ;
    RECT 28.51 50.47 28.72 50.54 ;
    RECT 28.51 50.83 28.72 50.9 ;
    RECT 28.51 51.19 28.72 51.26 ;
    RECT 24.73 50.47 24.94 50.54 ;
    RECT 24.73 50.83 24.94 50.9 ;
    RECT 24.73 51.19 24.94 51.26 ;
    RECT 25.19 50.47 25.4 50.54 ;
    RECT 25.19 50.83 25.4 50.9 ;
    RECT 25.19 51.19 25.4 51.26 ;
    RECT 21.41 50.47 21.62 50.54 ;
    RECT 21.41 50.83 21.62 50.9 ;
    RECT 21.41 51.19 21.62 51.26 ;
    RECT 21.87 50.47 22.08 50.54 ;
    RECT 21.87 50.83 22.08 50.9 ;
    RECT 21.87 51.19 22.08 51.26 ;
    RECT 18.09 50.47 18.3 50.54 ;
    RECT 18.09 50.83 18.3 50.9 ;
    RECT 18.09 51.19 18.3 51.26 ;
    RECT 18.55 50.47 18.76 50.54 ;
    RECT 18.55 50.83 18.76 50.9 ;
    RECT 18.55 51.19 18.76 51.26 ;
    RECT 120.825 50.83 120.895 50.9 ;
    RECT 14.77 50.47 14.98 50.54 ;
    RECT 14.77 50.83 14.98 50.9 ;
    RECT 14.77 51.19 14.98 51.26 ;
    RECT 15.23 50.47 15.44 50.54 ;
    RECT 15.23 50.83 15.44 50.9 ;
    RECT 15.23 51.19 15.44 51.26 ;
    RECT 11.45 50.47 11.66 50.54 ;
    RECT 11.45 50.83 11.66 50.9 ;
    RECT 11.45 51.19 11.66 51.26 ;
    RECT 11.91 50.47 12.12 50.54 ;
    RECT 11.91 50.83 12.12 50.9 ;
    RECT 11.91 51.19 12.12 51.26 ;
    RECT 8.13 50.47 8.34 50.54 ;
    RECT 8.13 50.83 8.34 50.9 ;
    RECT 8.13 51.19 8.34 51.26 ;
    RECT 8.59 50.47 8.8 50.54 ;
    RECT 8.59 50.83 8.8 50.9 ;
    RECT 8.59 51.19 8.8 51.26 ;
    RECT 4.81 50.47 5.02 50.54 ;
    RECT 4.81 50.83 5.02 50.9 ;
    RECT 4.81 51.19 5.02 51.26 ;
    RECT 5.27 50.47 5.48 50.54 ;
    RECT 5.27 50.83 5.48 50.9 ;
    RECT 5.27 51.19 5.48 51.26 ;
    RECT 1.49 50.47 1.7 50.54 ;
    RECT 1.49 50.83 1.7 50.9 ;
    RECT 1.49 51.19 1.7 51.26 ;
    RECT 1.95 50.47 2.16 50.54 ;
    RECT 1.95 50.83 2.16 50.9 ;
    RECT 1.95 51.19 2.16 51.26 ;
    RECT 64.57 50.47 64.78 50.54 ;
    RECT 64.57 50.83 64.78 50.9 ;
    RECT 64.57 51.19 64.78 51.26 ;
    RECT 65.03 50.47 65.24 50.54 ;
    RECT 65.03 50.83 65.24 50.9 ;
    RECT 65.03 51.19 65.24 51.26 ;
    RECT 61.25 93.69 61.46 93.76 ;
    RECT 61.25 94.05 61.46 94.12 ;
    RECT 61.25 94.41 61.46 94.48 ;
    RECT 61.71 93.69 61.92 93.76 ;
    RECT 61.71 94.05 61.92 94.12 ;
    RECT 61.71 94.41 61.92 94.48 ;
    RECT 57.93 93.69 58.14 93.76 ;
    RECT 57.93 94.05 58.14 94.12 ;
    RECT 57.93 94.41 58.14 94.48 ;
    RECT 58.39 93.69 58.6 93.76 ;
    RECT 58.39 94.05 58.6 94.12 ;
    RECT 58.39 94.41 58.6 94.48 ;
    RECT 54.61 93.69 54.82 93.76 ;
    RECT 54.61 94.05 54.82 94.12 ;
    RECT 54.61 94.41 54.82 94.48 ;
    RECT 55.07 93.69 55.28 93.76 ;
    RECT 55.07 94.05 55.28 94.12 ;
    RECT 55.07 94.41 55.28 94.48 ;
    RECT 51.29 93.69 51.5 93.76 ;
    RECT 51.29 94.05 51.5 94.12 ;
    RECT 51.29 94.41 51.5 94.48 ;
    RECT 51.75 93.69 51.96 93.76 ;
    RECT 51.75 94.05 51.96 94.12 ;
    RECT 51.75 94.41 51.96 94.48 ;
    RECT 47.97 93.69 48.18 93.76 ;
    RECT 47.97 94.05 48.18 94.12 ;
    RECT 47.97 94.41 48.18 94.48 ;
    RECT 48.43 93.69 48.64 93.76 ;
    RECT 48.43 94.05 48.64 94.12 ;
    RECT 48.43 94.41 48.64 94.48 ;
    RECT 44.65 93.69 44.86 93.76 ;
    RECT 44.65 94.05 44.86 94.12 ;
    RECT 44.65 94.41 44.86 94.48 ;
    RECT 45.11 93.69 45.32 93.76 ;
    RECT 45.11 94.05 45.32 94.12 ;
    RECT 45.11 94.41 45.32 94.48 ;
    RECT 41.33 93.69 41.54 93.76 ;
    RECT 41.33 94.05 41.54 94.12 ;
    RECT 41.33 94.41 41.54 94.48 ;
    RECT 41.79 93.69 42.0 93.76 ;
    RECT 41.79 94.05 42.0 94.12 ;
    RECT 41.79 94.41 42.0 94.48 ;
    RECT 38.01 93.69 38.22 93.76 ;
    RECT 38.01 94.05 38.22 94.12 ;
    RECT 38.01 94.41 38.22 94.48 ;
    RECT 38.47 93.69 38.68 93.76 ;
    RECT 38.47 94.05 38.68 94.12 ;
    RECT 38.47 94.41 38.68 94.48 ;
    RECT 0.4 94.05 0.47 94.12 ;
    RECT 34.69 93.69 34.9 93.76 ;
    RECT 34.69 94.05 34.9 94.12 ;
    RECT 34.69 94.41 34.9 94.48 ;
    RECT 35.15 93.69 35.36 93.76 ;
    RECT 35.15 94.05 35.36 94.12 ;
    RECT 35.15 94.41 35.36 94.48 ;
    RECT 117.69 93.69 117.9 93.76 ;
    RECT 117.69 94.05 117.9 94.12 ;
    RECT 117.69 94.41 117.9 94.48 ;
    RECT 118.15 93.69 118.36 93.76 ;
    RECT 118.15 94.05 118.36 94.12 ;
    RECT 118.15 94.41 118.36 94.48 ;
    RECT 114.37 93.69 114.58 93.76 ;
    RECT 114.37 94.05 114.58 94.12 ;
    RECT 114.37 94.41 114.58 94.48 ;
    RECT 114.83 93.69 115.04 93.76 ;
    RECT 114.83 94.05 115.04 94.12 ;
    RECT 114.83 94.41 115.04 94.48 ;
    RECT 111.05 93.69 111.26 93.76 ;
    RECT 111.05 94.05 111.26 94.12 ;
    RECT 111.05 94.41 111.26 94.48 ;
    RECT 111.51 93.69 111.72 93.76 ;
    RECT 111.51 94.05 111.72 94.12 ;
    RECT 111.51 94.41 111.72 94.48 ;
    RECT 107.73 93.69 107.94 93.76 ;
    RECT 107.73 94.05 107.94 94.12 ;
    RECT 107.73 94.41 107.94 94.48 ;
    RECT 108.19 93.69 108.4 93.76 ;
    RECT 108.19 94.05 108.4 94.12 ;
    RECT 108.19 94.41 108.4 94.48 ;
    RECT 104.41 93.69 104.62 93.76 ;
    RECT 104.41 94.05 104.62 94.12 ;
    RECT 104.41 94.41 104.62 94.48 ;
    RECT 104.87 93.69 105.08 93.76 ;
    RECT 104.87 94.05 105.08 94.12 ;
    RECT 104.87 94.41 105.08 94.48 ;
    RECT 101.09 93.69 101.3 93.76 ;
    RECT 101.09 94.05 101.3 94.12 ;
    RECT 101.09 94.41 101.3 94.48 ;
    RECT 101.55 93.69 101.76 93.76 ;
    RECT 101.55 94.05 101.76 94.12 ;
    RECT 101.55 94.41 101.76 94.48 ;
    RECT 97.77 93.69 97.98 93.76 ;
    RECT 97.77 94.05 97.98 94.12 ;
    RECT 97.77 94.41 97.98 94.48 ;
    RECT 98.23 93.69 98.44 93.76 ;
    RECT 98.23 94.05 98.44 94.12 ;
    RECT 98.23 94.41 98.44 94.48 ;
    RECT 94.45 93.69 94.66 93.76 ;
    RECT 94.45 94.05 94.66 94.12 ;
    RECT 94.45 94.41 94.66 94.48 ;
    RECT 94.91 93.69 95.12 93.76 ;
    RECT 94.91 94.05 95.12 94.12 ;
    RECT 94.91 94.41 95.12 94.48 ;
    RECT 91.13 93.69 91.34 93.76 ;
    RECT 91.13 94.05 91.34 94.12 ;
    RECT 91.13 94.41 91.34 94.48 ;
    RECT 91.59 93.69 91.8 93.76 ;
    RECT 91.59 94.05 91.8 94.12 ;
    RECT 91.59 94.41 91.8 94.48 ;
    RECT 87.81 93.69 88.02 93.76 ;
    RECT 87.81 94.05 88.02 94.12 ;
    RECT 87.81 94.41 88.02 94.48 ;
    RECT 88.27 93.69 88.48 93.76 ;
    RECT 88.27 94.05 88.48 94.12 ;
    RECT 88.27 94.41 88.48 94.48 ;
    RECT 84.49 93.69 84.7 93.76 ;
    RECT 84.49 94.05 84.7 94.12 ;
    RECT 84.49 94.41 84.7 94.48 ;
    RECT 84.95 93.69 85.16 93.76 ;
    RECT 84.95 94.05 85.16 94.12 ;
    RECT 84.95 94.41 85.16 94.48 ;
    RECT 81.17 93.69 81.38 93.76 ;
    RECT 81.17 94.05 81.38 94.12 ;
    RECT 81.17 94.41 81.38 94.48 ;
    RECT 81.63 93.69 81.84 93.76 ;
    RECT 81.63 94.05 81.84 94.12 ;
    RECT 81.63 94.41 81.84 94.48 ;
    RECT 77.85 93.69 78.06 93.76 ;
    RECT 77.85 94.05 78.06 94.12 ;
    RECT 77.85 94.41 78.06 94.48 ;
    RECT 78.31 93.69 78.52 93.76 ;
    RECT 78.31 94.05 78.52 94.12 ;
    RECT 78.31 94.41 78.52 94.48 ;
    RECT 74.53 93.69 74.74 93.76 ;
    RECT 74.53 94.05 74.74 94.12 ;
    RECT 74.53 94.41 74.74 94.48 ;
    RECT 74.99 93.69 75.2 93.76 ;
    RECT 74.99 94.05 75.2 94.12 ;
    RECT 74.99 94.41 75.2 94.48 ;
    RECT 71.21 93.69 71.42 93.76 ;
    RECT 71.21 94.05 71.42 94.12 ;
    RECT 71.21 94.41 71.42 94.48 ;
    RECT 71.67 93.69 71.88 93.76 ;
    RECT 71.67 94.05 71.88 94.12 ;
    RECT 71.67 94.41 71.88 94.48 ;
    RECT 31.37 93.69 31.58 93.76 ;
    RECT 31.37 94.05 31.58 94.12 ;
    RECT 31.37 94.41 31.58 94.48 ;
    RECT 31.83 93.69 32.04 93.76 ;
    RECT 31.83 94.05 32.04 94.12 ;
    RECT 31.83 94.41 32.04 94.48 ;
    RECT 67.89 93.69 68.1 93.76 ;
    RECT 67.89 94.05 68.1 94.12 ;
    RECT 67.89 94.41 68.1 94.48 ;
    RECT 68.35 93.69 68.56 93.76 ;
    RECT 68.35 94.05 68.56 94.12 ;
    RECT 68.35 94.41 68.56 94.48 ;
    RECT 28.05 93.69 28.26 93.76 ;
    RECT 28.05 94.05 28.26 94.12 ;
    RECT 28.05 94.41 28.26 94.48 ;
    RECT 28.51 93.69 28.72 93.76 ;
    RECT 28.51 94.05 28.72 94.12 ;
    RECT 28.51 94.41 28.72 94.48 ;
    RECT 24.73 93.69 24.94 93.76 ;
    RECT 24.73 94.05 24.94 94.12 ;
    RECT 24.73 94.41 24.94 94.48 ;
    RECT 25.19 93.69 25.4 93.76 ;
    RECT 25.19 94.05 25.4 94.12 ;
    RECT 25.19 94.41 25.4 94.48 ;
    RECT 21.41 93.69 21.62 93.76 ;
    RECT 21.41 94.05 21.62 94.12 ;
    RECT 21.41 94.41 21.62 94.48 ;
    RECT 21.87 93.69 22.08 93.76 ;
    RECT 21.87 94.05 22.08 94.12 ;
    RECT 21.87 94.41 22.08 94.48 ;
    RECT 18.09 93.69 18.3 93.76 ;
    RECT 18.09 94.05 18.3 94.12 ;
    RECT 18.09 94.41 18.3 94.48 ;
    RECT 18.55 93.69 18.76 93.76 ;
    RECT 18.55 94.05 18.76 94.12 ;
    RECT 18.55 94.41 18.76 94.48 ;
    RECT 120.825 94.05 120.895 94.12 ;
    RECT 14.77 93.69 14.98 93.76 ;
    RECT 14.77 94.05 14.98 94.12 ;
    RECT 14.77 94.41 14.98 94.48 ;
    RECT 15.23 93.69 15.44 93.76 ;
    RECT 15.23 94.05 15.44 94.12 ;
    RECT 15.23 94.41 15.44 94.48 ;
    RECT 11.45 93.69 11.66 93.76 ;
    RECT 11.45 94.05 11.66 94.12 ;
    RECT 11.45 94.41 11.66 94.48 ;
    RECT 11.91 93.69 12.12 93.76 ;
    RECT 11.91 94.05 12.12 94.12 ;
    RECT 11.91 94.41 12.12 94.48 ;
    RECT 8.13 93.69 8.34 93.76 ;
    RECT 8.13 94.05 8.34 94.12 ;
    RECT 8.13 94.41 8.34 94.48 ;
    RECT 8.59 93.69 8.8 93.76 ;
    RECT 8.59 94.05 8.8 94.12 ;
    RECT 8.59 94.41 8.8 94.48 ;
    RECT 4.81 93.69 5.02 93.76 ;
    RECT 4.81 94.05 5.02 94.12 ;
    RECT 4.81 94.41 5.02 94.48 ;
    RECT 5.27 93.69 5.48 93.76 ;
    RECT 5.27 94.05 5.48 94.12 ;
    RECT 5.27 94.41 5.48 94.48 ;
    RECT 1.49 93.69 1.7 93.76 ;
    RECT 1.49 94.05 1.7 94.12 ;
    RECT 1.49 94.41 1.7 94.48 ;
    RECT 1.95 93.69 2.16 93.76 ;
    RECT 1.95 94.05 2.16 94.12 ;
    RECT 1.95 94.41 2.16 94.48 ;
    RECT 64.57 93.69 64.78 93.76 ;
    RECT 64.57 94.05 64.78 94.12 ;
    RECT 64.57 94.41 64.78 94.48 ;
    RECT 65.03 93.69 65.24 93.76 ;
    RECT 65.03 94.05 65.24 94.12 ;
    RECT 65.03 94.41 65.24 94.48 ;
    RECT 61.25 92.97 61.46 93.04 ;
    RECT 61.25 93.33 61.46 93.4 ;
    RECT 61.25 93.69 61.46 93.76 ;
    RECT 61.71 92.97 61.92 93.04 ;
    RECT 61.71 93.33 61.92 93.4 ;
    RECT 61.71 93.69 61.92 93.76 ;
    RECT 57.93 92.97 58.14 93.04 ;
    RECT 57.93 93.33 58.14 93.4 ;
    RECT 57.93 93.69 58.14 93.76 ;
    RECT 58.39 92.97 58.6 93.04 ;
    RECT 58.39 93.33 58.6 93.4 ;
    RECT 58.39 93.69 58.6 93.76 ;
    RECT 54.61 92.97 54.82 93.04 ;
    RECT 54.61 93.33 54.82 93.4 ;
    RECT 54.61 93.69 54.82 93.76 ;
    RECT 55.07 92.97 55.28 93.04 ;
    RECT 55.07 93.33 55.28 93.4 ;
    RECT 55.07 93.69 55.28 93.76 ;
    RECT 51.29 92.97 51.5 93.04 ;
    RECT 51.29 93.33 51.5 93.4 ;
    RECT 51.29 93.69 51.5 93.76 ;
    RECT 51.75 92.97 51.96 93.04 ;
    RECT 51.75 93.33 51.96 93.4 ;
    RECT 51.75 93.69 51.96 93.76 ;
    RECT 47.97 92.97 48.18 93.04 ;
    RECT 47.97 93.33 48.18 93.4 ;
    RECT 47.97 93.69 48.18 93.76 ;
    RECT 48.43 92.97 48.64 93.04 ;
    RECT 48.43 93.33 48.64 93.4 ;
    RECT 48.43 93.69 48.64 93.76 ;
    RECT 44.65 92.97 44.86 93.04 ;
    RECT 44.65 93.33 44.86 93.4 ;
    RECT 44.65 93.69 44.86 93.76 ;
    RECT 45.11 92.97 45.32 93.04 ;
    RECT 45.11 93.33 45.32 93.4 ;
    RECT 45.11 93.69 45.32 93.76 ;
    RECT 41.33 92.97 41.54 93.04 ;
    RECT 41.33 93.33 41.54 93.4 ;
    RECT 41.33 93.69 41.54 93.76 ;
    RECT 41.79 92.97 42.0 93.04 ;
    RECT 41.79 93.33 42.0 93.4 ;
    RECT 41.79 93.69 42.0 93.76 ;
    RECT 38.01 92.97 38.22 93.04 ;
    RECT 38.01 93.33 38.22 93.4 ;
    RECT 38.01 93.69 38.22 93.76 ;
    RECT 38.47 92.97 38.68 93.04 ;
    RECT 38.47 93.33 38.68 93.4 ;
    RECT 38.47 93.69 38.68 93.76 ;
    RECT 0.4 93.33 0.47 93.4 ;
    RECT 34.69 92.97 34.9 93.04 ;
    RECT 34.69 93.33 34.9 93.4 ;
    RECT 34.69 93.69 34.9 93.76 ;
    RECT 35.15 92.97 35.36 93.04 ;
    RECT 35.15 93.33 35.36 93.4 ;
    RECT 35.15 93.69 35.36 93.76 ;
    RECT 117.69 92.97 117.9 93.04 ;
    RECT 117.69 93.33 117.9 93.4 ;
    RECT 117.69 93.69 117.9 93.76 ;
    RECT 118.15 92.97 118.36 93.04 ;
    RECT 118.15 93.33 118.36 93.4 ;
    RECT 118.15 93.69 118.36 93.76 ;
    RECT 114.37 92.97 114.58 93.04 ;
    RECT 114.37 93.33 114.58 93.4 ;
    RECT 114.37 93.69 114.58 93.76 ;
    RECT 114.83 92.97 115.04 93.04 ;
    RECT 114.83 93.33 115.04 93.4 ;
    RECT 114.83 93.69 115.04 93.76 ;
    RECT 111.05 92.97 111.26 93.04 ;
    RECT 111.05 93.33 111.26 93.4 ;
    RECT 111.05 93.69 111.26 93.76 ;
    RECT 111.51 92.97 111.72 93.04 ;
    RECT 111.51 93.33 111.72 93.4 ;
    RECT 111.51 93.69 111.72 93.76 ;
    RECT 107.73 92.97 107.94 93.04 ;
    RECT 107.73 93.33 107.94 93.4 ;
    RECT 107.73 93.69 107.94 93.76 ;
    RECT 108.19 92.97 108.4 93.04 ;
    RECT 108.19 93.33 108.4 93.4 ;
    RECT 108.19 93.69 108.4 93.76 ;
    RECT 104.41 92.97 104.62 93.04 ;
    RECT 104.41 93.33 104.62 93.4 ;
    RECT 104.41 93.69 104.62 93.76 ;
    RECT 104.87 92.97 105.08 93.04 ;
    RECT 104.87 93.33 105.08 93.4 ;
    RECT 104.87 93.69 105.08 93.76 ;
    RECT 101.09 92.97 101.3 93.04 ;
    RECT 101.09 93.33 101.3 93.4 ;
    RECT 101.09 93.69 101.3 93.76 ;
    RECT 101.55 92.97 101.76 93.04 ;
    RECT 101.55 93.33 101.76 93.4 ;
    RECT 101.55 93.69 101.76 93.76 ;
    RECT 97.77 92.97 97.98 93.04 ;
    RECT 97.77 93.33 97.98 93.4 ;
    RECT 97.77 93.69 97.98 93.76 ;
    RECT 98.23 92.97 98.44 93.04 ;
    RECT 98.23 93.33 98.44 93.4 ;
    RECT 98.23 93.69 98.44 93.76 ;
    RECT 94.45 92.97 94.66 93.04 ;
    RECT 94.45 93.33 94.66 93.4 ;
    RECT 94.45 93.69 94.66 93.76 ;
    RECT 94.91 92.97 95.12 93.04 ;
    RECT 94.91 93.33 95.12 93.4 ;
    RECT 94.91 93.69 95.12 93.76 ;
    RECT 91.13 92.97 91.34 93.04 ;
    RECT 91.13 93.33 91.34 93.4 ;
    RECT 91.13 93.69 91.34 93.76 ;
    RECT 91.59 92.97 91.8 93.04 ;
    RECT 91.59 93.33 91.8 93.4 ;
    RECT 91.59 93.69 91.8 93.76 ;
    RECT 87.81 92.97 88.02 93.04 ;
    RECT 87.81 93.33 88.02 93.4 ;
    RECT 87.81 93.69 88.02 93.76 ;
    RECT 88.27 92.97 88.48 93.04 ;
    RECT 88.27 93.33 88.48 93.4 ;
    RECT 88.27 93.69 88.48 93.76 ;
    RECT 84.49 92.97 84.7 93.04 ;
    RECT 84.49 93.33 84.7 93.4 ;
    RECT 84.49 93.69 84.7 93.76 ;
    RECT 84.95 92.97 85.16 93.04 ;
    RECT 84.95 93.33 85.16 93.4 ;
    RECT 84.95 93.69 85.16 93.76 ;
    RECT 81.17 92.97 81.38 93.04 ;
    RECT 81.17 93.33 81.38 93.4 ;
    RECT 81.17 93.69 81.38 93.76 ;
    RECT 81.63 92.97 81.84 93.04 ;
    RECT 81.63 93.33 81.84 93.4 ;
    RECT 81.63 93.69 81.84 93.76 ;
    RECT 77.85 92.97 78.06 93.04 ;
    RECT 77.85 93.33 78.06 93.4 ;
    RECT 77.85 93.69 78.06 93.76 ;
    RECT 78.31 92.97 78.52 93.04 ;
    RECT 78.31 93.33 78.52 93.4 ;
    RECT 78.31 93.69 78.52 93.76 ;
    RECT 74.53 92.97 74.74 93.04 ;
    RECT 74.53 93.33 74.74 93.4 ;
    RECT 74.53 93.69 74.74 93.76 ;
    RECT 74.99 92.97 75.2 93.04 ;
    RECT 74.99 93.33 75.2 93.4 ;
    RECT 74.99 93.69 75.2 93.76 ;
    RECT 71.21 92.97 71.42 93.04 ;
    RECT 71.21 93.33 71.42 93.4 ;
    RECT 71.21 93.69 71.42 93.76 ;
    RECT 71.67 92.97 71.88 93.04 ;
    RECT 71.67 93.33 71.88 93.4 ;
    RECT 71.67 93.69 71.88 93.76 ;
    RECT 31.37 92.97 31.58 93.04 ;
    RECT 31.37 93.33 31.58 93.4 ;
    RECT 31.37 93.69 31.58 93.76 ;
    RECT 31.83 92.97 32.04 93.04 ;
    RECT 31.83 93.33 32.04 93.4 ;
    RECT 31.83 93.69 32.04 93.76 ;
    RECT 67.89 92.97 68.1 93.04 ;
    RECT 67.89 93.33 68.1 93.4 ;
    RECT 67.89 93.69 68.1 93.76 ;
    RECT 68.35 92.97 68.56 93.04 ;
    RECT 68.35 93.33 68.56 93.4 ;
    RECT 68.35 93.69 68.56 93.76 ;
    RECT 28.05 92.97 28.26 93.04 ;
    RECT 28.05 93.33 28.26 93.4 ;
    RECT 28.05 93.69 28.26 93.76 ;
    RECT 28.51 92.97 28.72 93.04 ;
    RECT 28.51 93.33 28.72 93.4 ;
    RECT 28.51 93.69 28.72 93.76 ;
    RECT 24.73 92.97 24.94 93.04 ;
    RECT 24.73 93.33 24.94 93.4 ;
    RECT 24.73 93.69 24.94 93.76 ;
    RECT 25.19 92.97 25.4 93.04 ;
    RECT 25.19 93.33 25.4 93.4 ;
    RECT 25.19 93.69 25.4 93.76 ;
    RECT 21.41 92.97 21.62 93.04 ;
    RECT 21.41 93.33 21.62 93.4 ;
    RECT 21.41 93.69 21.62 93.76 ;
    RECT 21.87 92.97 22.08 93.04 ;
    RECT 21.87 93.33 22.08 93.4 ;
    RECT 21.87 93.69 22.08 93.76 ;
    RECT 18.09 92.97 18.3 93.04 ;
    RECT 18.09 93.33 18.3 93.4 ;
    RECT 18.09 93.69 18.3 93.76 ;
    RECT 18.55 92.97 18.76 93.04 ;
    RECT 18.55 93.33 18.76 93.4 ;
    RECT 18.55 93.69 18.76 93.76 ;
    RECT 120.825 93.33 120.895 93.4 ;
    RECT 14.77 92.97 14.98 93.04 ;
    RECT 14.77 93.33 14.98 93.4 ;
    RECT 14.77 93.69 14.98 93.76 ;
    RECT 15.23 92.97 15.44 93.04 ;
    RECT 15.23 93.33 15.44 93.4 ;
    RECT 15.23 93.69 15.44 93.76 ;
    RECT 11.45 92.97 11.66 93.04 ;
    RECT 11.45 93.33 11.66 93.4 ;
    RECT 11.45 93.69 11.66 93.76 ;
    RECT 11.91 92.97 12.12 93.04 ;
    RECT 11.91 93.33 12.12 93.4 ;
    RECT 11.91 93.69 12.12 93.76 ;
    RECT 8.13 92.97 8.34 93.04 ;
    RECT 8.13 93.33 8.34 93.4 ;
    RECT 8.13 93.69 8.34 93.76 ;
    RECT 8.59 92.97 8.8 93.04 ;
    RECT 8.59 93.33 8.8 93.4 ;
    RECT 8.59 93.69 8.8 93.76 ;
    RECT 4.81 92.97 5.02 93.04 ;
    RECT 4.81 93.33 5.02 93.4 ;
    RECT 4.81 93.69 5.02 93.76 ;
    RECT 5.27 92.97 5.48 93.04 ;
    RECT 5.27 93.33 5.48 93.4 ;
    RECT 5.27 93.69 5.48 93.76 ;
    RECT 1.49 92.97 1.7 93.04 ;
    RECT 1.49 93.33 1.7 93.4 ;
    RECT 1.49 93.69 1.7 93.76 ;
    RECT 1.95 92.97 2.16 93.04 ;
    RECT 1.95 93.33 2.16 93.4 ;
    RECT 1.95 93.69 2.16 93.76 ;
    RECT 64.57 92.97 64.78 93.04 ;
    RECT 64.57 93.33 64.78 93.4 ;
    RECT 64.57 93.69 64.78 93.76 ;
    RECT 65.03 92.97 65.24 93.04 ;
    RECT 65.03 93.33 65.24 93.4 ;
    RECT 65.03 93.69 65.24 93.76 ;
    RECT 61.25 92.25 61.46 92.32 ;
    RECT 61.25 92.61 61.46 92.68 ;
    RECT 61.25 92.97 61.46 93.04 ;
    RECT 61.71 92.25 61.92 92.32 ;
    RECT 61.71 92.61 61.92 92.68 ;
    RECT 61.71 92.97 61.92 93.04 ;
    RECT 57.93 92.25 58.14 92.32 ;
    RECT 57.93 92.61 58.14 92.68 ;
    RECT 57.93 92.97 58.14 93.04 ;
    RECT 58.39 92.25 58.6 92.32 ;
    RECT 58.39 92.61 58.6 92.68 ;
    RECT 58.39 92.97 58.6 93.04 ;
    RECT 54.61 92.25 54.82 92.32 ;
    RECT 54.61 92.61 54.82 92.68 ;
    RECT 54.61 92.97 54.82 93.04 ;
    RECT 55.07 92.25 55.28 92.32 ;
    RECT 55.07 92.61 55.28 92.68 ;
    RECT 55.07 92.97 55.28 93.04 ;
    RECT 51.29 92.25 51.5 92.32 ;
    RECT 51.29 92.61 51.5 92.68 ;
    RECT 51.29 92.97 51.5 93.04 ;
    RECT 51.75 92.25 51.96 92.32 ;
    RECT 51.75 92.61 51.96 92.68 ;
    RECT 51.75 92.97 51.96 93.04 ;
    RECT 47.97 92.25 48.18 92.32 ;
    RECT 47.97 92.61 48.18 92.68 ;
    RECT 47.97 92.97 48.18 93.04 ;
    RECT 48.43 92.25 48.64 92.32 ;
    RECT 48.43 92.61 48.64 92.68 ;
    RECT 48.43 92.97 48.64 93.04 ;
    RECT 44.65 92.25 44.86 92.32 ;
    RECT 44.65 92.61 44.86 92.68 ;
    RECT 44.65 92.97 44.86 93.04 ;
    RECT 45.11 92.25 45.32 92.32 ;
    RECT 45.11 92.61 45.32 92.68 ;
    RECT 45.11 92.97 45.32 93.04 ;
    RECT 41.33 92.25 41.54 92.32 ;
    RECT 41.33 92.61 41.54 92.68 ;
    RECT 41.33 92.97 41.54 93.04 ;
    RECT 41.79 92.25 42.0 92.32 ;
    RECT 41.79 92.61 42.0 92.68 ;
    RECT 41.79 92.97 42.0 93.04 ;
    RECT 38.01 92.25 38.22 92.32 ;
    RECT 38.01 92.61 38.22 92.68 ;
    RECT 38.01 92.97 38.22 93.04 ;
    RECT 38.47 92.25 38.68 92.32 ;
    RECT 38.47 92.61 38.68 92.68 ;
    RECT 38.47 92.97 38.68 93.04 ;
    RECT 0.4 92.61 0.47 92.68 ;
    RECT 34.69 92.25 34.9 92.32 ;
    RECT 34.69 92.61 34.9 92.68 ;
    RECT 34.69 92.97 34.9 93.04 ;
    RECT 35.15 92.25 35.36 92.32 ;
    RECT 35.15 92.61 35.36 92.68 ;
    RECT 35.15 92.97 35.36 93.04 ;
    RECT 117.69 92.25 117.9 92.32 ;
    RECT 117.69 92.61 117.9 92.68 ;
    RECT 117.69 92.97 117.9 93.04 ;
    RECT 118.15 92.25 118.36 92.32 ;
    RECT 118.15 92.61 118.36 92.68 ;
    RECT 118.15 92.97 118.36 93.04 ;
    RECT 114.37 92.25 114.58 92.32 ;
    RECT 114.37 92.61 114.58 92.68 ;
    RECT 114.37 92.97 114.58 93.04 ;
    RECT 114.83 92.25 115.04 92.32 ;
    RECT 114.83 92.61 115.04 92.68 ;
    RECT 114.83 92.97 115.04 93.04 ;
    RECT 111.05 92.25 111.26 92.32 ;
    RECT 111.05 92.61 111.26 92.68 ;
    RECT 111.05 92.97 111.26 93.04 ;
    RECT 111.51 92.25 111.72 92.32 ;
    RECT 111.51 92.61 111.72 92.68 ;
    RECT 111.51 92.97 111.72 93.04 ;
    RECT 107.73 92.25 107.94 92.32 ;
    RECT 107.73 92.61 107.94 92.68 ;
    RECT 107.73 92.97 107.94 93.04 ;
    RECT 108.19 92.25 108.4 92.32 ;
    RECT 108.19 92.61 108.4 92.68 ;
    RECT 108.19 92.97 108.4 93.04 ;
    RECT 104.41 92.25 104.62 92.32 ;
    RECT 104.41 92.61 104.62 92.68 ;
    RECT 104.41 92.97 104.62 93.04 ;
    RECT 104.87 92.25 105.08 92.32 ;
    RECT 104.87 92.61 105.08 92.68 ;
    RECT 104.87 92.97 105.08 93.04 ;
    RECT 101.09 92.25 101.3 92.32 ;
    RECT 101.09 92.61 101.3 92.68 ;
    RECT 101.09 92.97 101.3 93.04 ;
    RECT 101.55 92.25 101.76 92.32 ;
    RECT 101.55 92.61 101.76 92.68 ;
    RECT 101.55 92.97 101.76 93.04 ;
    RECT 97.77 92.25 97.98 92.32 ;
    RECT 97.77 92.61 97.98 92.68 ;
    RECT 97.77 92.97 97.98 93.04 ;
    RECT 98.23 92.25 98.44 92.32 ;
    RECT 98.23 92.61 98.44 92.68 ;
    RECT 98.23 92.97 98.44 93.04 ;
    RECT 94.45 92.25 94.66 92.32 ;
    RECT 94.45 92.61 94.66 92.68 ;
    RECT 94.45 92.97 94.66 93.04 ;
    RECT 94.91 92.25 95.12 92.32 ;
    RECT 94.91 92.61 95.12 92.68 ;
    RECT 94.91 92.97 95.12 93.04 ;
    RECT 91.13 92.25 91.34 92.32 ;
    RECT 91.13 92.61 91.34 92.68 ;
    RECT 91.13 92.97 91.34 93.04 ;
    RECT 91.59 92.25 91.8 92.32 ;
    RECT 91.59 92.61 91.8 92.68 ;
    RECT 91.59 92.97 91.8 93.04 ;
    RECT 87.81 92.25 88.02 92.32 ;
    RECT 87.81 92.61 88.02 92.68 ;
    RECT 87.81 92.97 88.02 93.04 ;
    RECT 88.27 92.25 88.48 92.32 ;
    RECT 88.27 92.61 88.48 92.68 ;
    RECT 88.27 92.97 88.48 93.04 ;
    RECT 84.49 92.25 84.7 92.32 ;
    RECT 84.49 92.61 84.7 92.68 ;
    RECT 84.49 92.97 84.7 93.04 ;
    RECT 84.95 92.25 85.16 92.32 ;
    RECT 84.95 92.61 85.16 92.68 ;
    RECT 84.95 92.97 85.16 93.04 ;
    RECT 81.17 92.25 81.38 92.32 ;
    RECT 81.17 92.61 81.38 92.68 ;
    RECT 81.17 92.97 81.38 93.04 ;
    RECT 81.63 92.25 81.84 92.32 ;
    RECT 81.63 92.61 81.84 92.68 ;
    RECT 81.63 92.97 81.84 93.04 ;
    RECT 77.85 92.25 78.06 92.32 ;
    RECT 77.85 92.61 78.06 92.68 ;
    RECT 77.85 92.97 78.06 93.04 ;
    RECT 78.31 92.25 78.52 92.32 ;
    RECT 78.31 92.61 78.52 92.68 ;
    RECT 78.31 92.97 78.52 93.04 ;
    RECT 74.53 92.25 74.74 92.32 ;
    RECT 74.53 92.61 74.74 92.68 ;
    RECT 74.53 92.97 74.74 93.04 ;
    RECT 74.99 92.25 75.2 92.32 ;
    RECT 74.99 92.61 75.2 92.68 ;
    RECT 74.99 92.97 75.2 93.04 ;
    RECT 71.21 92.25 71.42 92.32 ;
    RECT 71.21 92.61 71.42 92.68 ;
    RECT 71.21 92.97 71.42 93.04 ;
    RECT 71.67 92.25 71.88 92.32 ;
    RECT 71.67 92.61 71.88 92.68 ;
    RECT 71.67 92.97 71.88 93.04 ;
    RECT 31.37 92.25 31.58 92.32 ;
    RECT 31.37 92.61 31.58 92.68 ;
    RECT 31.37 92.97 31.58 93.04 ;
    RECT 31.83 92.25 32.04 92.32 ;
    RECT 31.83 92.61 32.04 92.68 ;
    RECT 31.83 92.97 32.04 93.04 ;
    RECT 67.89 92.25 68.1 92.32 ;
    RECT 67.89 92.61 68.1 92.68 ;
    RECT 67.89 92.97 68.1 93.04 ;
    RECT 68.35 92.25 68.56 92.32 ;
    RECT 68.35 92.61 68.56 92.68 ;
    RECT 68.35 92.97 68.56 93.04 ;
    RECT 28.05 92.25 28.26 92.32 ;
    RECT 28.05 92.61 28.26 92.68 ;
    RECT 28.05 92.97 28.26 93.04 ;
    RECT 28.51 92.25 28.72 92.32 ;
    RECT 28.51 92.61 28.72 92.68 ;
    RECT 28.51 92.97 28.72 93.04 ;
    RECT 24.73 92.25 24.94 92.32 ;
    RECT 24.73 92.61 24.94 92.68 ;
    RECT 24.73 92.97 24.94 93.04 ;
    RECT 25.19 92.25 25.4 92.32 ;
    RECT 25.19 92.61 25.4 92.68 ;
    RECT 25.19 92.97 25.4 93.04 ;
    RECT 21.41 92.25 21.62 92.32 ;
    RECT 21.41 92.61 21.62 92.68 ;
    RECT 21.41 92.97 21.62 93.04 ;
    RECT 21.87 92.25 22.08 92.32 ;
    RECT 21.87 92.61 22.08 92.68 ;
    RECT 21.87 92.97 22.08 93.04 ;
    RECT 18.09 92.25 18.3 92.32 ;
    RECT 18.09 92.61 18.3 92.68 ;
    RECT 18.09 92.97 18.3 93.04 ;
    RECT 18.55 92.25 18.76 92.32 ;
    RECT 18.55 92.61 18.76 92.68 ;
    RECT 18.55 92.97 18.76 93.04 ;
    RECT 120.825 92.61 120.895 92.68 ;
    RECT 14.77 92.25 14.98 92.32 ;
    RECT 14.77 92.61 14.98 92.68 ;
    RECT 14.77 92.97 14.98 93.04 ;
    RECT 15.23 92.25 15.44 92.32 ;
    RECT 15.23 92.61 15.44 92.68 ;
    RECT 15.23 92.97 15.44 93.04 ;
    RECT 11.45 92.25 11.66 92.32 ;
    RECT 11.45 92.61 11.66 92.68 ;
    RECT 11.45 92.97 11.66 93.04 ;
    RECT 11.91 92.25 12.12 92.32 ;
    RECT 11.91 92.61 12.12 92.68 ;
    RECT 11.91 92.97 12.12 93.04 ;
    RECT 8.13 92.25 8.34 92.32 ;
    RECT 8.13 92.61 8.34 92.68 ;
    RECT 8.13 92.97 8.34 93.04 ;
    RECT 8.59 92.25 8.8 92.32 ;
    RECT 8.59 92.61 8.8 92.68 ;
    RECT 8.59 92.97 8.8 93.04 ;
    RECT 4.81 92.25 5.02 92.32 ;
    RECT 4.81 92.61 5.02 92.68 ;
    RECT 4.81 92.97 5.02 93.04 ;
    RECT 5.27 92.25 5.48 92.32 ;
    RECT 5.27 92.61 5.48 92.68 ;
    RECT 5.27 92.97 5.48 93.04 ;
    RECT 1.49 92.25 1.7 92.32 ;
    RECT 1.49 92.61 1.7 92.68 ;
    RECT 1.49 92.97 1.7 93.04 ;
    RECT 1.95 92.25 2.16 92.32 ;
    RECT 1.95 92.61 2.16 92.68 ;
    RECT 1.95 92.97 2.16 93.04 ;
    RECT 64.57 92.25 64.78 92.32 ;
    RECT 64.57 92.61 64.78 92.68 ;
    RECT 64.57 92.97 64.78 93.04 ;
    RECT 65.03 92.25 65.24 92.32 ;
    RECT 65.03 92.61 65.24 92.68 ;
    RECT 65.03 92.97 65.24 93.04 ;
    RECT 61.25 91.53 61.46 91.6 ;
    RECT 61.25 91.89 61.46 91.96 ;
    RECT 61.25 92.25 61.46 92.32 ;
    RECT 61.71 91.53 61.92 91.6 ;
    RECT 61.71 91.89 61.92 91.96 ;
    RECT 61.71 92.25 61.92 92.32 ;
    RECT 57.93 91.53 58.14 91.6 ;
    RECT 57.93 91.89 58.14 91.96 ;
    RECT 57.93 92.25 58.14 92.32 ;
    RECT 58.39 91.53 58.6 91.6 ;
    RECT 58.39 91.89 58.6 91.96 ;
    RECT 58.39 92.25 58.6 92.32 ;
    RECT 54.61 91.53 54.82 91.6 ;
    RECT 54.61 91.89 54.82 91.96 ;
    RECT 54.61 92.25 54.82 92.32 ;
    RECT 55.07 91.53 55.28 91.6 ;
    RECT 55.07 91.89 55.28 91.96 ;
    RECT 55.07 92.25 55.28 92.32 ;
    RECT 51.29 91.53 51.5 91.6 ;
    RECT 51.29 91.89 51.5 91.96 ;
    RECT 51.29 92.25 51.5 92.32 ;
    RECT 51.75 91.53 51.96 91.6 ;
    RECT 51.75 91.89 51.96 91.96 ;
    RECT 51.75 92.25 51.96 92.32 ;
    RECT 47.97 91.53 48.18 91.6 ;
    RECT 47.97 91.89 48.18 91.96 ;
    RECT 47.97 92.25 48.18 92.32 ;
    RECT 48.43 91.53 48.64 91.6 ;
    RECT 48.43 91.89 48.64 91.96 ;
    RECT 48.43 92.25 48.64 92.32 ;
    RECT 44.65 91.53 44.86 91.6 ;
    RECT 44.65 91.89 44.86 91.96 ;
    RECT 44.65 92.25 44.86 92.32 ;
    RECT 45.11 91.53 45.32 91.6 ;
    RECT 45.11 91.89 45.32 91.96 ;
    RECT 45.11 92.25 45.32 92.32 ;
    RECT 41.33 91.53 41.54 91.6 ;
    RECT 41.33 91.89 41.54 91.96 ;
    RECT 41.33 92.25 41.54 92.32 ;
    RECT 41.79 91.53 42.0 91.6 ;
    RECT 41.79 91.89 42.0 91.96 ;
    RECT 41.79 92.25 42.0 92.32 ;
    RECT 38.01 91.53 38.22 91.6 ;
    RECT 38.01 91.89 38.22 91.96 ;
    RECT 38.01 92.25 38.22 92.32 ;
    RECT 38.47 91.53 38.68 91.6 ;
    RECT 38.47 91.89 38.68 91.96 ;
    RECT 38.47 92.25 38.68 92.32 ;
    RECT 0.4 91.89 0.47 91.96 ;
    RECT 34.69 91.53 34.9 91.6 ;
    RECT 34.69 91.89 34.9 91.96 ;
    RECT 34.69 92.25 34.9 92.32 ;
    RECT 35.15 91.53 35.36 91.6 ;
    RECT 35.15 91.89 35.36 91.96 ;
    RECT 35.15 92.25 35.36 92.32 ;
    RECT 117.69 91.53 117.9 91.6 ;
    RECT 117.69 91.89 117.9 91.96 ;
    RECT 117.69 92.25 117.9 92.32 ;
    RECT 118.15 91.53 118.36 91.6 ;
    RECT 118.15 91.89 118.36 91.96 ;
    RECT 118.15 92.25 118.36 92.32 ;
    RECT 114.37 91.53 114.58 91.6 ;
    RECT 114.37 91.89 114.58 91.96 ;
    RECT 114.37 92.25 114.58 92.32 ;
    RECT 114.83 91.53 115.04 91.6 ;
    RECT 114.83 91.89 115.04 91.96 ;
    RECT 114.83 92.25 115.04 92.32 ;
    RECT 111.05 91.53 111.26 91.6 ;
    RECT 111.05 91.89 111.26 91.96 ;
    RECT 111.05 92.25 111.26 92.32 ;
    RECT 111.51 91.53 111.72 91.6 ;
    RECT 111.51 91.89 111.72 91.96 ;
    RECT 111.51 92.25 111.72 92.32 ;
    RECT 107.73 91.53 107.94 91.6 ;
    RECT 107.73 91.89 107.94 91.96 ;
    RECT 107.73 92.25 107.94 92.32 ;
    RECT 108.19 91.53 108.4 91.6 ;
    RECT 108.19 91.89 108.4 91.96 ;
    RECT 108.19 92.25 108.4 92.32 ;
    RECT 104.41 91.53 104.62 91.6 ;
    RECT 104.41 91.89 104.62 91.96 ;
    RECT 104.41 92.25 104.62 92.32 ;
    RECT 104.87 91.53 105.08 91.6 ;
    RECT 104.87 91.89 105.08 91.96 ;
    RECT 104.87 92.25 105.08 92.32 ;
    RECT 101.09 91.53 101.3 91.6 ;
    RECT 101.09 91.89 101.3 91.96 ;
    RECT 101.09 92.25 101.3 92.32 ;
    RECT 101.55 91.53 101.76 91.6 ;
    RECT 101.55 91.89 101.76 91.96 ;
    RECT 101.55 92.25 101.76 92.32 ;
    RECT 97.77 91.53 97.98 91.6 ;
    RECT 97.77 91.89 97.98 91.96 ;
    RECT 97.77 92.25 97.98 92.32 ;
    RECT 98.23 91.53 98.44 91.6 ;
    RECT 98.23 91.89 98.44 91.96 ;
    RECT 98.23 92.25 98.44 92.32 ;
    RECT 94.45 91.53 94.66 91.6 ;
    RECT 94.45 91.89 94.66 91.96 ;
    RECT 94.45 92.25 94.66 92.32 ;
    RECT 94.91 91.53 95.12 91.6 ;
    RECT 94.91 91.89 95.12 91.96 ;
    RECT 94.91 92.25 95.12 92.32 ;
    RECT 91.13 91.53 91.34 91.6 ;
    RECT 91.13 91.89 91.34 91.96 ;
    RECT 91.13 92.25 91.34 92.32 ;
    RECT 91.59 91.53 91.8 91.6 ;
    RECT 91.59 91.89 91.8 91.96 ;
    RECT 91.59 92.25 91.8 92.32 ;
    RECT 87.81 91.53 88.02 91.6 ;
    RECT 87.81 91.89 88.02 91.96 ;
    RECT 87.81 92.25 88.02 92.32 ;
    RECT 88.27 91.53 88.48 91.6 ;
    RECT 88.27 91.89 88.48 91.96 ;
    RECT 88.27 92.25 88.48 92.32 ;
    RECT 84.49 91.53 84.7 91.6 ;
    RECT 84.49 91.89 84.7 91.96 ;
    RECT 84.49 92.25 84.7 92.32 ;
    RECT 84.95 91.53 85.16 91.6 ;
    RECT 84.95 91.89 85.16 91.96 ;
    RECT 84.95 92.25 85.16 92.32 ;
    RECT 81.17 91.53 81.38 91.6 ;
    RECT 81.17 91.89 81.38 91.96 ;
    RECT 81.17 92.25 81.38 92.32 ;
    RECT 81.63 91.53 81.84 91.6 ;
    RECT 81.63 91.89 81.84 91.96 ;
    RECT 81.63 92.25 81.84 92.32 ;
    RECT 77.85 91.53 78.06 91.6 ;
    RECT 77.85 91.89 78.06 91.96 ;
    RECT 77.85 92.25 78.06 92.32 ;
    RECT 78.31 91.53 78.52 91.6 ;
    RECT 78.31 91.89 78.52 91.96 ;
    RECT 78.31 92.25 78.52 92.32 ;
    RECT 74.53 91.53 74.74 91.6 ;
    RECT 74.53 91.89 74.74 91.96 ;
    RECT 74.53 92.25 74.74 92.32 ;
    RECT 74.99 91.53 75.2 91.6 ;
    RECT 74.99 91.89 75.2 91.96 ;
    RECT 74.99 92.25 75.2 92.32 ;
    RECT 71.21 91.53 71.42 91.6 ;
    RECT 71.21 91.89 71.42 91.96 ;
    RECT 71.21 92.25 71.42 92.32 ;
    RECT 71.67 91.53 71.88 91.6 ;
    RECT 71.67 91.89 71.88 91.96 ;
    RECT 71.67 92.25 71.88 92.32 ;
    RECT 31.37 91.53 31.58 91.6 ;
    RECT 31.37 91.89 31.58 91.96 ;
    RECT 31.37 92.25 31.58 92.32 ;
    RECT 31.83 91.53 32.04 91.6 ;
    RECT 31.83 91.89 32.04 91.96 ;
    RECT 31.83 92.25 32.04 92.32 ;
    RECT 67.89 91.53 68.1 91.6 ;
    RECT 67.89 91.89 68.1 91.96 ;
    RECT 67.89 92.25 68.1 92.32 ;
    RECT 68.35 91.53 68.56 91.6 ;
    RECT 68.35 91.89 68.56 91.96 ;
    RECT 68.35 92.25 68.56 92.32 ;
    RECT 28.05 91.53 28.26 91.6 ;
    RECT 28.05 91.89 28.26 91.96 ;
    RECT 28.05 92.25 28.26 92.32 ;
    RECT 28.51 91.53 28.72 91.6 ;
    RECT 28.51 91.89 28.72 91.96 ;
    RECT 28.51 92.25 28.72 92.32 ;
    RECT 24.73 91.53 24.94 91.6 ;
    RECT 24.73 91.89 24.94 91.96 ;
    RECT 24.73 92.25 24.94 92.32 ;
    RECT 25.19 91.53 25.4 91.6 ;
    RECT 25.19 91.89 25.4 91.96 ;
    RECT 25.19 92.25 25.4 92.32 ;
    RECT 21.41 91.53 21.62 91.6 ;
    RECT 21.41 91.89 21.62 91.96 ;
    RECT 21.41 92.25 21.62 92.32 ;
    RECT 21.87 91.53 22.08 91.6 ;
    RECT 21.87 91.89 22.08 91.96 ;
    RECT 21.87 92.25 22.08 92.32 ;
    RECT 18.09 91.53 18.3 91.6 ;
    RECT 18.09 91.89 18.3 91.96 ;
    RECT 18.09 92.25 18.3 92.32 ;
    RECT 18.55 91.53 18.76 91.6 ;
    RECT 18.55 91.89 18.76 91.96 ;
    RECT 18.55 92.25 18.76 92.32 ;
    RECT 120.825 91.89 120.895 91.96 ;
    RECT 14.77 91.53 14.98 91.6 ;
    RECT 14.77 91.89 14.98 91.96 ;
    RECT 14.77 92.25 14.98 92.32 ;
    RECT 15.23 91.53 15.44 91.6 ;
    RECT 15.23 91.89 15.44 91.96 ;
    RECT 15.23 92.25 15.44 92.32 ;
    RECT 11.45 91.53 11.66 91.6 ;
    RECT 11.45 91.89 11.66 91.96 ;
    RECT 11.45 92.25 11.66 92.32 ;
    RECT 11.91 91.53 12.12 91.6 ;
    RECT 11.91 91.89 12.12 91.96 ;
    RECT 11.91 92.25 12.12 92.32 ;
    RECT 8.13 91.53 8.34 91.6 ;
    RECT 8.13 91.89 8.34 91.96 ;
    RECT 8.13 92.25 8.34 92.32 ;
    RECT 8.59 91.53 8.8 91.6 ;
    RECT 8.59 91.89 8.8 91.96 ;
    RECT 8.59 92.25 8.8 92.32 ;
    RECT 4.81 91.53 5.02 91.6 ;
    RECT 4.81 91.89 5.02 91.96 ;
    RECT 4.81 92.25 5.02 92.32 ;
    RECT 5.27 91.53 5.48 91.6 ;
    RECT 5.27 91.89 5.48 91.96 ;
    RECT 5.27 92.25 5.48 92.32 ;
    RECT 1.49 91.53 1.7 91.6 ;
    RECT 1.49 91.89 1.7 91.96 ;
    RECT 1.49 92.25 1.7 92.32 ;
    RECT 1.95 91.53 2.16 91.6 ;
    RECT 1.95 91.89 2.16 91.96 ;
    RECT 1.95 92.25 2.16 92.32 ;
    RECT 64.57 91.53 64.78 91.6 ;
    RECT 64.57 91.89 64.78 91.96 ;
    RECT 64.57 92.25 64.78 92.32 ;
    RECT 65.03 91.53 65.24 91.6 ;
    RECT 65.03 91.89 65.24 91.96 ;
    RECT 65.03 92.25 65.24 92.32 ;
    RECT 61.25 90.81 61.46 90.88 ;
    RECT 61.25 91.17 61.46 91.24 ;
    RECT 61.25 91.53 61.46 91.6 ;
    RECT 61.71 90.81 61.92 90.88 ;
    RECT 61.71 91.17 61.92 91.24 ;
    RECT 61.71 91.53 61.92 91.6 ;
    RECT 57.93 90.81 58.14 90.88 ;
    RECT 57.93 91.17 58.14 91.24 ;
    RECT 57.93 91.53 58.14 91.6 ;
    RECT 58.39 90.81 58.6 90.88 ;
    RECT 58.39 91.17 58.6 91.24 ;
    RECT 58.39 91.53 58.6 91.6 ;
    RECT 54.61 90.81 54.82 90.88 ;
    RECT 54.61 91.17 54.82 91.24 ;
    RECT 54.61 91.53 54.82 91.6 ;
    RECT 55.07 90.81 55.28 90.88 ;
    RECT 55.07 91.17 55.28 91.24 ;
    RECT 55.07 91.53 55.28 91.6 ;
    RECT 51.29 90.81 51.5 90.88 ;
    RECT 51.29 91.17 51.5 91.24 ;
    RECT 51.29 91.53 51.5 91.6 ;
    RECT 51.75 90.81 51.96 90.88 ;
    RECT 51.75 91.17 51.96 91.24 ;
    RECT 51.75 91.53 51.96 91.6 ;
    RECT 47.97 90.81 48.18 90.88 ;
    RECT 47.97 91.17 48.18 91.24 ;
    RECT 47.97 91.53 48.18 91.6 ;
    RECT 48.43 90.81 48.64 90.88 ;
    RECT 48.43 91.17 48.64 91.24 ;
    RECT 48.43 91.53 48.64 91.6 ;
    RECT 44.65 90.81 44.86 90.88 ;
    RECT 44.65 91.17 44.86 91.24 ;
    RECT 44.65 91.53 44.86 91.6 ;
    RECT 45.11 90.81 45.32 90.88 ;
    RECT 45.11 91.17 45.32 91.24 ;
    RECT 45.11 91.53 45.32 91.6 ;
    RECT 41.33 90.81 41.54 90.88 ;
    RECT 41.33 91.17 41.54 91.24 ;
    RECT 41.33 91.53 41.54 91.6 ;
    RECT 41.79 90.81 42.0 90.88 ;
    RECT 41.79 91.17 42.0 91.24 ;
    RECT 41.79 91.53 42.0 91.6 ;
    RECT 38.01 90.81 38.22 90.88 ;
    RECT 38.01 91.17 38.22 91.24 ;
    RECT 38.01 91.53 38.22 91.6 ;
    RECT 38.47 90.81 38.68 90.88 ;
    RECT 38.47 91.17 38.68 91.24 ;
    RECT 38.47 91.53 38.68 91.6 ;
    RECT 0.4 91.17 0.47 91.24 ;
    RECT 34.69 90.81 34.9 90.88 ;
    RECT 34.69 91.17 34.9 91.24 ;
    RECT 34.69 91.53 34.9 91.6 ;
    RECT 35.15 90.81 35.36 90.88 ;
    RECT 35.15 91.17 35.36 91.24 ;
    RECT 35.15 91.53 35.36 91.6 ;
    RECT 117.69 90.81 117.9 90.88 ;
    RECT 117.69 91.17 117.9 91.24 ;
    RECT 117.69 91.53 117.9 91.6 ;
    RECT 118.15 90.81 118.36 90.88 ;
    RECT 118.15 91.17 118.36 91.24 ;
    RECT 118.15 91.53 118.36 91.6 ;
    RECT 114.37 90.81 114.58 90.88 ;
    RECT 114.37 91.17 114.58 91.24 ;
    RECT 114.37 91.53 114.58 91.6 ;
    RECT 114.83 90.81 115.04 90.88 ;
    RECT 114.83 91.17 115.04 91.24 ;
    RECT 114.83 91.53 115.04 91.6 ;
    RECT 111.05 90.81 111.26 90.88 ;
    RECT 111.05 91.17 111.26 91.24 ;
    RECT 111.05 91.53 111.26 91.6 ;
    RECT 111.51 90.81 111.72 90.88 ;
    RECT 111.51 91.17 111.72 91.24 ;
    RECT 111.51 91.53 111.72 91.6 ;
    RECT 107.73 90.81 107.94 90.88 ;
    RECT 107.73 91.17 107.94 91.24 ;
    RECT 107.73 91.53 107.94 91.6 ;
    RECT 108.19 90.81 108.4 90.88 ;
    RECT 108.19 91.17 108.4 91.24 ;
    RECT 108.19 91.53 108.4 91.6 ;
    RECT 104.41 90.81 104.62 90.88 ;
    RECT 104.41 91.17 104.62 91.24 ;
    RECT 104.41 91.53 104.62 91.6 ;
    RECT 104.87 90.81 105.08 90.88 ;
    RECT 104.87 91.17 105.08 91.24 ;
    RECT 104.87 91.53 105.08 91.6 ;
    RECT 101.09 90.81 101.3 90.88 ;
    RECT 101.09 91.17 101.3 91.24 ;
    RECT 101.09 91.53 101.3 91.6 ;
    RECT 101.55 90.81 101.76 90.88 ;
    RECT 101.55 91.17 101.76 91.24 ;
    RECT 101.55 91.53 101.76 91.6 ;
    RECT 97.77 90.81 97.98 90.88 ;
    RECT 97.77 91.17 97.98 91.24 ;
    RECT 97.77 91.53 97.98 91.6 ;
    RECT 98.23 90.81 98.44 90.88 ;
    RECT 98.23 91.17 98.44 91.24 ;
    RECT 98.23 91.53 98.44 91.6 ;
    RECT 94.45 90.81 94.66 90.88 ;
    RECT 94.45 91.17 94.66 91.24 ;
    RECT 94.45 91.53 94.66 91.6 ;
    RECT 94.91 90.81 95.12 90.88 ;
    RECT 94.91 91.17 95.12 91.24 ;
    RECT 94.91 91.53 95.12 91.6 ;
    RECT 91.13 90.81 91.34 90.88 ;
    RECT 91.13 91.17 91.34 91.24 ;
    RECT 91.13 91.53 91.34 91.6 ;
    RECT 91.59 90.81 91.8 90.88 ;
    RECT 91.59 91.17 91.8 91.24 ;
    RECT 91.59 91.53 91.8 91.6 ;
    RECT 87.81 90.81 88.02 90.88 ;
    RECT 87.81 91.17 88.02 91.24 ;
    RECT 87.81 91.53 88.02 91.6 ;
    RECT 88.27 90.81 88.48 90.88 ;
    RECT 88.27 91.17 88.48 91.24 ;
    RECT 88.27 91.53 88.48 91.6 ;
    RECT 84.49 90.81 84.7 90.88 ;
    RECT 84.49 91.17 84.7 91.24 ;
    RECT 84.49 91.53 84.7 91.6 ;
    RECT 84.95 90.81 85.16 90.88 ;
    RECT 84.95 91.17 85.16 91.24 ;
    RECT 84.95 91.53 85.16 91.6 ;
    RECT 81.17 90.81 81.38 90.88 ;
    RECT 81.17 91.17 81.38 91.24 ;
    RECT 81.17 91.53 81.38 91.6 ;
    RECT 81.63 90.81 81.84 90.88 ;
    RECT 81.63 91.17 81.84 91.24 ;
    RECT 81.63 91.53 81.84 91.6 ;
    RECT 77.85 90.81 78.06 90.88 ;
    RECT 77.85 91.17 78.06 91.24 ;
    RECT 77.85 91.53 78.06 91.6 ;
    RECT 78.31 90.81 78.52 90.88 ;
    RECT 78.31 91.17 78.52 91.24 ;
    RECT 78.31 91.53 78.52 91.6 ;
    RECT 74.53 90.81 74.74 90.88 ;
    RECT 74.53 91.17 74.74 91.24 ;
    RECT 74.53 91.53 74.74 91.6 ;
    RECT 74.99 90.81 75.2 90.88 ;
    RECT 74.99 91.17 75.2 91.24 ;
    RECT 74.99 91.53 75.2 91.6 ;
    RECT 71.21 90.81 71.42 90.88 ;
    RECT 71.21 91.17 71.42 91.24 ;
    RECT 71.21 91.53 71.42 91.6 ;
    RECT 71.67 90.81 71.88 90.88 ;
    RECT 71.67 91.17 71.88 91.24 ;
    RECT 71.67 91.53 71.88 91.6 ;
    RECT 31.37 90.81 31.58 90.88 ;
    RECT 31.37 91.17 31.58 91.24 ;
    RECT 31.37 91.53 31.58 91.6 ;
    RECT 31.83 90.81 32.04 90.88 ;
    RECT 31.83 91.17 32.04 91.24 ;
    RECT 31.83 91.53 32.04 91.6 ;
    RECT 67.89 90.81 68.1 90.88 ;
    RECT 67.89 91.17 68.1 91.24 ;
    RECT 67.89 91.53 68.1 91.6 ;
    RECT 68.35 90.81 68.56 90.88 ;
    RECT 68.35 91.17 68.56 91.24 ;
    RECT 68.35 91.53 68.56 91.6 ;
    RECT 28.05 90.81 28.26 90.88 ;
    RECT 28.05 91.17 28.26 91.24 ;
    RECT 28.05 91.53 28.26 91.6 ;
    RECT 28.51 90.81 28.72 90.88 ;
    RECT 28.51 91.17 28.72 91.24 ;
    RECT 28.51 91.53 28.72 91.6 ;
    RECT 24.73 90.81 24.94 90.88 ;
    RECT 24.73 91.17 24.94 91.24 ;
    RECT 24.73 91.53 24.94 91.6 ;
    RECT 25.19 90.81 25.4 90.88 ;
    RECT 25.19 91.17 25.4 91.24 ;
    RECT 25.19 91.53 25.4 91.6 ;
    RECT 21.41 90.81 21.62 90.88 ;
    RECT 21.41 91.17 21.62 91.24 ;
    RECT 21.41 91.53 21.62 91.6 ;
    RECT 21.87 90.81 22.08 90.88 ;
    RECT 21.87 91.17 22.08 91.24 ;
    RECT 21.87 91.53 22.08 91.6 ;
    RECT 18.09 90.81 18.3 90.88 ;
    RECT 18.09 91.17 18.3 91.24 ;
    RECT 18.09 91.53 18.3 91.6 ;
    RECT 18.55 90.81 18.76 90.88 ;
    RECT 18.55 91.17 18.76 91.24 ;
    RECT 18.55 91.53 18.76 91.6 ;
    RECT 120.825 91.17 120.895 91.24 ;
    RECT 14.77 90.81 14.98 90.88 ;
    RECT 14.77 91.17 14.98 91.24 ;
    RECT 14.77 91.53 14.98 91.6 ;
    RECT 15.23 90.81 15.44 90.88 ;
    RECT 15.23 91.17 15.44 91.24 ;
    RECT 15.23 91.53 15.44 91.6 ;
    RECT 11.45 90.81 11.66 90.88 ;
    RECT 11.45 91.17 11.66 91.24 ;
    RECT 11.45 91.53 11.66 91.6 ;
    RECT 11.91 90.81 12.12 90.88 ;
    RECT 11.91 91.17 12.12 91.24 ;
    RECT 11.91 91.53 12.12 91.6 ;
    RECT 8.13 90.81 8.34 90.88 ;
    RECT 8.13 91.17 8.34 91.24 ;
    RECT 8.13 91.53 8.34 91.6 ;
    RECT 8.59 90.81 8.8 90.88 ;
    RECT 8.59 91.17 8.8 91.24 ;
    RECT 8.59 91.53 8.8 91.6 ;
    RECT 4.81 90.81 5.02 90.88 ;
    RECT 4.81 91.17 5.02 91.24 ;
    RECT 4.81 91.53 5.02 91.6 ;
    RECT 5.27 90.81 5.48 90.88 ;
    RECT 5.27 91.17 5.48 91.24 ;
    RECT 5.27 91.53 5.48 91.6 ;
    RECT 1.49 90.81 1.7 90.88 ;
    RECT 1.49 91.17 1.7 91.24 ;
    RECT 1.49 91.53 1.7 91.6 ;
    RECT 1.95 90.81 2.16 90.88 ;
    RECT 1.95 91.17 2.16 91.24 ;
    RECT 1.95 91.53 2.16 91.6 ;
    RECT 64.57 90.81 64.78 90.88 ;
    RECT 64.57 91.17 64.78 91.24 ;
    RECT 64.57 91.53 64.78 91.6 ;
    RECT 65.03 90.81 65.24 90.88 ;
    RECT 65.03 91.17 65.24 91.24 ;
    RECT 65.03 91.53 65.24 91.6 ;
    RECT 61.25 90.09 61.46 90.16 ;
    RECT 61.25 90.45 61.46 90.52 ;
    RECT 61.25 90.81 61.46 90.88 ;
    RECT 61.71 90.09 61.92 90.16 ;
    RECT 61.71 90.45 61.92 90.52 ;
    RECT 61.71 90.81 61.92 90.88 ;
    RECT 57.93 90.09 58.14 90.16 ;
    RECT 57.93 90.45 58.14 90.52 ;
    RECT 57.93 90.81 58.14 90.88 ;
    RECT 58.39 90.09 58.6 90.16 ;
    RECT 58.39 90.45 58.6 90.52 ;
    RECT 58.39 90.81 58.6 90.88 ;
    RECT 54.61 90.09 54.82 90.16 ;
    RECT 54.61 90.45 54.82 90.52 ;
    RECT 54.61 90.81 54.82 90.88 ;
    RECT 55.07 90.09 55.28 90.16 ;
    RECT 55.07 90.45 55.28 90.52 ;
    RECT 55.07 90.81 55.28 90.88 ;
    RECT 51.29 90.09 51.5 90.16 ;
    RECT 51.29 90.45 51.5 90.52 ;
    RECT 51.29 90.81 51.5 90.88 ;
    RECT 51.75 90.09 51.96 90.16 ;
    RECT 51.75 90.45 51.96 90.52 ;
    RECT 51.75 90.81 51.96 90.88 ;
    RECT 47.97 90.09 48.18 90.16 ;
    RECT 47.97 90.45 48.18 90.52 ;
    RECT 47.97 90.81 48.18 90.88 ;
    RECT 48.43 90.09 48.64 90.16 ;
    RECT 48.43 90.45 48.64 90.52 ;
    RECT 48.43 90.81 48.64 90.88 ;
    RECT 44.65 90.09 44.86 90.16 ;
    RECT 44.65 90.45 44.86 90.52 ;
    RECT 44.65 90.81 44.86 90.88 ;
    RECT 45.11 90.09 45.32 90.16 ;
    RECT 45.11 90.45 45.32 90.52 ;
    RECT 45.11 90.81 45.32 90.88 ;
    RECT 41.33 90.09 41.54 90.16 ;
    RECT 41.33 90.45 41.54 90.52 ;
    RECT 41.33 90.81 41.54 90.88 ;
    RECT 41.79 90.09 42.0 90.16 ;
    RECT 41.79 90.45 42.0 90.52 ;
    RECT 41.79 90.81 42.0 90.88 ;
    RECT 38.01 90.09 38.22 90.16 ;
    RECT 38.01 90.45 38.22 90.52 ;
    RECT 38.01 90.81 38.22 90.88 ;
    RECT 38.47 90.09 38.68 90.16 ;
    RECT 38.47 90.45 38.68 90.52 ;
    RECT 38.47 90.81 38.68 90.88 ;
    RECT 0.4 90.45 0.47 90.52 ;
    RECT 34.69 90.09 34.9 90.16 ;
    RECT 34.69 90.45 34.9 90.52 ;
    RECT 34.69 90.81 34.9 90.88 ;
    RECT 35.15 90.09 35.36 90.16 ;
    RECT 35.15 90.45 35.36 90.52 ;
    RECT 35.15 90.81 35.36 90.88 ;
    RECT 117.69 90.09 117.9 90.16 ;
    RECT 117.69 90.45 117.9 90.52 ;
    RECT 117.69 90.81 117.9 90.88 ;
    RECT 118.15 90.09 118.36 90.16 ;
    RECT 118.15 90.45 118.36 90.52 ;
    RECT 118.15 90.81 118.36 90.88 ;
    RECT 114.37 90.09 114.58 90.16 ;
    RECT 114.37 90.45 114.58 90.52 ;
    RECT 114.37 90.81 114.58 90.88 ;
    RECT 114.83 90.09 115.04 90.16 ;
    RECT 114.83 90.45 115.04 90.52 ;
    RECT 114.83 90.81 115.04 90.88 ;
    RECT 111.05 90.09 111.26 90.16 ;
    RECT 111.05 90.45 111.26 90.52 ;
    RECT 111.05 90.81 111.26 90.88 ;
    RECT 111.51 90.09 111.72 90.16 ;
    RECT 111.51 90.45 111.72 90.52 ;
    RECT 111.51 90.81 111.72 90.88 ;
    RECT 107.73 90.09 107.94 90.16 ;
    RECT 107.73 90.45 107.94 90.52 ;
    RECT 107.73 90.81 107.94 90.88 ;
    RECT 108.19 90.09 108.4 90.16 ;
    RECT 108.19 90.45 108.4 90.52 ;
    RECT 108.19 90.81 108.4 90.88 ;
    RECT 104.41 90.09 104.62 90.16 ;
    RECT 104.41 90.45 104.62 90.52 ;
    RECT 104.41 90.81 104.62 90.88 ;
    RECT 104.87 90.09 105.08 90.16 ;
    RECT 104.87 90.45 105.08 90.52 ;
    RECT 104.87 90.81 105.08 90.88 ;
    RECT 101.09 90.09 101.3 90.16 ;
    RECT 101.09 90.45 101.3 90.52 ;
    RECT 101.09 90.81 101.3 90.88 ;
    RECT 101.55 90.09 101.76 90.16 ;
    RECT 101.55 90.45 101.76 90.52 ;
    RECT 101.55 90.81 101.76 90.88 ;
    RECT 97.77 90.09 97.98 90.16 ;
    RECT 97.77 90.45 97.98 90.52 ;
    RECT 97.77 90.81 97.98 90.88 ;
    RECT 98.23 90.09 98.44 90.16 ;
    RECT 98.23 90.45 98.44 90.52 ;
    RECT 98.23 90.81 98.44 90.88 ;
    RECT 94.45 90.09 94.66 90.16 ;
    RECT 94.45 90.45 94.66 90.52 ;
    RECT 94.45 90.81 94.66 90.88 ;
    RECT 94.91 90.09 95.12 90.16 ;
    RECT 94.91 90.45 95.12 90.52 ;
    RECT 94.91 90.81 95.12 90.88 ;
    RECT 91.13 90.09 91.34 90.16 ;
    RECT 91.13 90.45 91.34 90.52 ;
    RECT 91.13 90.81 91.34 90.88 ;
    RECT 91.59 90.09 91.8 90.16 ;
    RECT 91.59 90.45 91.8 90.52 ;
    RECT 91.59 90.81 91.8 90.88 ;
    RECT 87.81 90.09 88.02 90.16 ;
    RECT 87.81 90.45 88.02 90.52 ;
    RECT 87.81 90.81 88.02 90.88 ;
    RECT 88.27 90.09 88.48 90.16 ;
    RECT 88.27 90.45 88.48 90.52 ;
    RECT 88.27 90.81 88.48 90.88 ;
    RECT 84.49 90.09 84.7 90.16 ;
    RECT 84.49 90.45 84.7 90.52 ;
    RECT 84.49 90.81 84.7 90.88 ;
    RECT 84.95 90.09 85.16 90.16 ;
    RECT 84.95 90.45 85.16 90.52 ;
    RECT 84.95 90.81 85.16 90.88 ;
    RECT 81.17 90.09 81.38 90.16 ;
    RECT 81.17 90.45 81.38 90.52 ;
    RECT 81.17 90.81 81.38 90.88 ;
    RECT 81.63 90.09 81.84 90.16 ;
    RECT 81.63 90.45 81.84 90.52 ;
    RECT 81.63 90.81 81.84 90.88 ;
    RECT 77.85 90.09 78.06 90.16 ;
    RECT 77.85 90.45 78.06 90.52 ;
    RECT 77.85 90.81 78.06 90.88 ;
    RECT 78.31 90.09 78.52 90.16 ;
    RECT 78.31 90.45 78.52 90.52 ;
    RECT 78.31 90.81 78.52 90.88 ;
    RECT 74.53 90.09 74.74 90.16 ;
    RECT 74.53 90.45 74.74 90.52 ;
    RECT 74.53 90.81 74.74 90.88 ;
    RECT 74.99 90.09 75.2 90.16 ;
    RECT 74.99 90.45 75.2 90.52 ;
    RECT 74.99 90.81 75.2 90.88 ;
    RECT 71.21 90.09 71.42 90.16 ;
    RECT 71.21 90.45 71.42 90.52 ;
    RECT 71.21 90.81 71.42 90.88 ;
    RECT 71.67 90.09 71.88 90.16 ;
    RECT 71.67 90.45 71.88 90.52 ;
    RECT 71.67 90.81 71.88 90.88 ;
    RECT 31.37 90.09 31.58 90.16 ;
    RECT 31.37 90.45 31.58 90.52 ;
    RECT 31.37 90.81 31.58 90.88 ;
    RECT 31.83 90.09 32.04 90.16 ;
    RECT 31.83 90.45 32.04 90.52 ;
    RECT 31.83 90.81 32.04 90.88 ;
    RECT 67.89 90.09 68.1 90.16 ;
    RECT 67.89 90.45 68.1 90.52 ;
    RECT 67.89 90.81 68.1 90.88 ;
    RECT 68.35 90.09 68.56 90.16 ;
    RECT 68.35 90.45 68.56 90.52 ;
    RECT 68.35 90.81 68.56 90.88 ;
    RECT 28.05 90.09 28.26 90.16 ;
    RECT 28.05 90.45 28.26 90.52 ;
    RECT 28.05 90.81 28.26 90.88 ;
    RECT 28.51 90.09 28.72 90.16 ;
    RECT 28.51 90.45 28.72 90.52 ;
    RECT 28.51 90.81 28.72 90.88 ;
    RECT 24.73 90.09 24.94 90.16 ;
    RECT 24.73 90.45 24.94 90.52 ;
    RECT 24.73 90.81 24.94 90.88 ;
    RECT 25.19 90.09 25.4 90.16 ;
    RECT 25.19 90.45 25.4 90.52 ;
    RECT 25.19 90.81 25.4 90.88 ;
    RECT 21.41 90.09 21.62 90.16 ;
    RECT 21.41 90.45 21.62 90.52 ;
    RECT 21.41 90.81 21.62 90.88 ;
    RECT 21.87 90.09 22.08 90.16 ;
    RECT 21.87 90.45 22.08 90.52 ;
    RECT 21.87 90.81 22.08 90.88 ;
    RECT 18.09 90.09 18.3 90.16 ;
    RECT 18.09 90.45 18.3 90.52 ;
    RECT 18.09 90.81 18.3 90.88 ;
    RECT 18.55 90.09 18.76 90.16 ;
    RECT 18.55 90.45 18.76 90.52 ;
    RECT 18.55 90.81 18.76 90.88 ;
    RECT 120.825 90.45 120.895 90.52 ;
    RECT 14.77 90.09 14.98 90.16 ;
    RECT 14.77 90.45 14.98 90.52 ;
    RECT 14.77 90.81 14.98 90.88 ;
    RECT 15.23 90.09 15.44 90.16 ;
    RECT 15.23 90.45 15.44 90.52 ;
    RECT 15.23 90.81 15.44 90.88 ;
    RECT 11.45 90.09 11.66 90.16 ;
    RECT 11.45 90.45 11.66 90.52 ;
    RECT 11.45 90.81 11.66 90.88 ;
    RECT 11.91 90.09 12.12 90.16 ;
    RECT 11.91 90.45 12.12 90.52 ;
    RECT 11.91 90.81 12.12 90.88 ;
    RECT 8.13 90.09 8.34 90.16 ;
    RECT 8.13 90.45 8.34 90.52 ;
    RECT 8.13 90.81 8.34 90.88 ;
    RECT 8.59 90.09 8.8 90.16 ;
    RECT 8.59 90.45 8.8 90.52 ;
    RECT 8.59 90.81 8.8 90.88 ;
    RECT 4.81 90.09 5.02 90.16 ;
    RECT 4.81 90.45 5.02 90.52 ;
    RECT 4.81 90.81 5.02 90.88 ;
    RECT 5.27 90.09 5.48 90.16 ;
    RECT 5.27 90.45 5.48 90.52 ;
    RECT 5.27 90.81 5.48 90.88 ;
    RECT 1.49 90.09 1.7 90.16 ;
    RECT 1.49 90.45 1.7 90.52 ;
    RECT 1.49 90.81 1.7 90.88 ;
    RECT 1.95 90.09 2.16 90.16 ;
    RECT 1.95 90.45 2.16 90.52 ;
    RECT 1.95 90.81 2.16 90.88 ;
    RECT 64.57 90.09 64.78 90.16 ;
    RECT 64.57 90.45 64.78 90.52 ;
    RECT 64.57 90.81 64.78 90.88 ;
    RECT 65.03 90.09 65.24 90.16 ;
    RECT 65.03 90.45 65.24 90.52 ;
    RECT 65.03 90.81 65.24 90.88 ;
    RECT 61.25 89.37 61.46 89.44 ;
    RECT 61.25 89.73 61.46 89.8 ;
    RECT 61.25 90.09 61.46 90.16 ;
    RECT 61.71 89.37 61.92 89.44 ;
    RECT 61.71 89.73 61.92 89.8 ;
    RECT 61.71 90.09 61.92 90.16 ;
    RECT 57.93 89.37 58.14 89.44 ;
    RECT 57.93 89.73 58.14 89.8 ;
    RECT 57.93 90.09 58.14 90.16 ;
    RECT 58.39 89.37 58.6 89.44 ;
    RECT 58.39 89.73 58.6 89.8 ;
    RECT 58.39 90.09 58.6 90.16 ;
    RECT 54.61 89.37 54.82 89.44 ;
    RECT 54.61 89.73 54.82 89.8 ;
    RECT 54.61 90.09 54.82 90.16 ;
    RECT 55.07 89.37 55.28 89.44 ;
    RECT 55.07 89.73 55.28 89.8 ;
    RECT 55.07 90.09 55.28 90.16 ;
    RECT 51.29 89.37 51.5 89.44 ;
    RECT 51.29 89.73 51.5 89.8 ;
    RECT 51.29 90.09 51.5 90.16 ;
    RECT 51.75 89.37 51.96 89.44 ;
    RECT 51.75 89.73 51.96 89.8 ;
    RECT 51.75 90.09 51.96 90.16 ;
    RECT 47.97 89.37 48.18 89.44 ;
    RECT 47.97 89.73 48.18 89.8 ;
    RECT 47.97 90.09 48.18 90.16 ;
    RECT 48.43 89.37 48.64 89.44 ;
    RECT 48.43 89.73 48.64 89.8 ;
    RECT 48.43 90.09 48.64 90.16 ;
    RECT 44.65 89.37 44.86 89.44 ;
    RECT 44.65 89.73 44.86 89.8 ;
    RECT 44.65 90.09 44.86 90.16 ;
    RECT 45.11 89.37 45.32 89.44 ;
    RECT 45.11 89.73 45.32 89.8 ;
    RECT 45.11 90.09 45.32 90.16 ;
    RECT 41.33 89.37 41.54 89.44 ;
    RECT 41.33 89.73 41.54 89.8 ;
    RECT 41.33 90.09 41.54 90.16 ;
    RECT 41.79 89.37 42.0 89.44 ;
    RECT 41.79 89.73 42.0 89.8 ;
    RECT 41.79 90.09 42.0 90.16 ;
    RECT 38.01 89.37 38.22 89.44 ;
    RECT 38.01 89.73 38.22 89.8 ;
    RECT 38.01 90.09 38.22 90.16 ;
    RECT 38.47 89.37 38.68 89.44 ;
    RECT 38.47 89.73 38.68 89.8 ;
    RECT 38.47 90.09 38.68 90.16 ;
    RECT 0.4 89.73 0.47 89.8 ;
    RECT 34.69 89.37 34.9 89.44 ;
    RECT 34.69 89.73 34.9 89.8 ;
    RECT 34.69 90.09 34.9 90.16 ;
    RECT 35.15 89.37 35.36 89.44 ;
    RECT 35.15 89.73 35.36 89.8 ;
    RECT 35.15 90.09 35.36 90.16 ;
    RECT 117.69 89.37 117.9 89.44 ;
    RECT 117.69 89.73 117.9 89.8 ;
    RECT 117.69 90.09 117.9 90.16 ;
    RECT 118.15 89.37 118.36 89.44 ;
    RECT 118.15 89.73 118.36 89.8 ;
    RECT 118.15 90.09 118.36 90.16 ;
    RECT 114.37 89.37 114.58 89.44 ;
    RECT 114.37 89.73 114.58 89.8 ;
    RECT 114.37 90.09 114.58 90.16 ;
    RECT 114.83 89.37 115.04 89.44 ;
    RECT 114.83 89.73 115.04 89.8 ;
    RECT 114.83 90.09 115.04 90.16 ;
    RECT 111.05 89.37 111.26 89.44 ;
    RECT 111.05 89.73 111.26 89.8 ;
    RECT 111.05 90.09 111.26 90.16 ;
    RECT 111.51 89.37 111.72 89.44 ;
    RECT 111.51 89.73 111.72 89.8 ;
    RECT 111.51 90.09 111.72 90.16 ;
    RECT 107.73 89.37 107.94 89.44 ;
    RECT 107.73 89.73 107.94 89.8 ;
    RECT 107.73 90.09 107.94 90.16 ;
    RECT 108.19 89.37 108.4 89.44 ;
    RECT 108.19 89.73 108.4 89.8 ;
    RECT 108.19 90.09 108.4 90.16 ;
    RECT 104.41 89.37 104.62 89.44 ;
    RECT 104.41 89.73 104.62 89.8 ;
    RECT 104.41 90.09 104.62 90.16 ;
    RECT 104.87 89.37 105.08 89.44 ;
    RECT 104.87 89.73 105.08 89.8 ;
    RECT 104.87 90.09 105.08 90.16 ;
    RECT 101.09 89.37 101.3 89.44 ;
    RECT 101.09 89.73 101.3 89.8 ;
    RECT 101.09 90.09 101.3 90.16 ;
    RECT 101.55 89.37 101.76 89.44 ;
    RECT 101.55 89.73 101.76 89.8 ;
    RECT 101.55 90.09 101.76 90.16 ;
    RECT 97.77 89.37 97.98 89.44 ;
    RECT 97.77 89.73 97.98 89.8 ;
    RECT 97.77 90.09 97.98 90.16 ;
    RECT 98.23 89.37 98.44 89.44 ;
    RECT 98.23 89.73 98.44 89.8 ;
    RECT 98.23 90.09 98.44 90.16 ;
    RECT 94.45 89.37 94.66 89.44 ;
    RECT 94.45 89.73 94.66 89.8 ;
    RECT 94.45 90.09 94.66 90.16 ;
    RECT 94.91 89.37 95.12 89.44 ;
    RECT 94.91 89.73 95.12 89.8 ;
    RECT 94.91 90.09 95.12 90.16 ;
    RECT 91.13 89.37 91.34 89.44 ;
    RECT 91.13 89.73 91.34 89.8 ;
    RECT 91.13 90.09 91.34 90.16 ;
    RECT 91.59 89.37 91.8 89.44 ;
    RECT 91.59 89.73 91.8 89.8 ;
    RECT 91.59 90.09 91.8 90.16 ;
    RECT 87.81 89.37 88.02 89.44 ;
    RECT 87.81 89.73 88.02 89.8 ;
    RECT 87.81 90.09 88.02 90.16 ;
    RECT 88.27 89.37 88.48 89.44 ;
    RECT 88.27 89.73 88.48 89.8 ;
    RECT 88.27 90.09 88.48 90.16 ;
    RECT 84.49 89.37 84.7 89.44 ;
    RECT 84.49 89.73 84.7 89.8 ;
    RECT 84.49 90.09 84.7 90.16 ;
    RECT 84.95 89.37 85.16 89.44 ;
    RECT 84.95 89.73 85.16 89.8 ;
    RECT 84.95 90.09 85.16 90.16 ;
    RECT 81.17 89.37 81.38 89.44 ;
    RECT 81.17 89.73 81.38 89.8 ;
    RECT 81.17 90.09 81.38 90.16 ;
    RECT 81.63 89.37 81.84 89.44 ;
    RECT 81.63 89.73 81.84 89.8 ;
    RECT 81.63 90.09 81.84 90.16 ;
    RECT 77.85 89.37 78.06 89.44 ;
    RECT 77.85 89.73 78.06 89.8 ;
    RECT 77.85 90.09 78.06 90.16 ;
    RECT 78.31 89.37 78.52 89.44 ;
    RECT 78.31 89.73 78.52 89.8 ;
    RECT 78.31 90.09 78.52 90.16 ;
    RECT 74.53 89.37 74.74 89.44 ;
    RECT 74.53 89.73 74.74 89.8 ;
    RECT 74.53 90.09 74.74 90.16 ;
    RECT 74.99 89.37 75.2 89.44 ;
    RECT 74.99 89.73 75.2 89.8 ;
    RECT 74.99 90.09 75.2 90.16 ;
    RECT 71.21 89.37 71.42 89.44 ;
    RECT 71.21 89.73 71.42 89.8 ;
    RECT 71.21 90.09 71.42 90.16 ;
    RECT 71.67 89.37 71.88 89.44 ;
    RECT 71.67 89.73 71.88 89.8 ;
    RECT 71.67 90.09 71.88 90.16 ;
    RECT 31.37 89.37 31.58 89.44 ;
    RECT 31.37 89.73 31.58 89.8 ;
    RECT 31.37 90.09 31.58 90.16 ;
    RECT 31.83 89.37 32.04 89.44 ;
    RECT 31.83 89.73 32.04 89.8 ;
    RECT 31.83 90.09 32.04 90.16 ;
    RECT 67.89 89.37 68.1 89.44 ;
    RECT 67.89 89.73 68.1 89.8 ;
    RECT 67.89 90.09 68.1 90.16 ;
    RECT 68.35 89.37 68.56 89.44 ;
    RECT 68.35 89.73 68.56 89.8 ;
    RECT 68.35 90.09 68.56 90.16 ;
    RECT 28.05 89.37 28.26 89.44 ;
    RECT 28.05 89.73 28.26 89.8 ;
    RECT 28.05 90.09 28.26 90.16 ;
    RECT 28.51 89.37 28.72 89.44 ;
    RECT 28.51 89.73 28.72 89.8 ;
    RECT 28.51 90.09 28.72 90.16 ;
    RECT 24.73 89.37 24.94 89.44 ;
    RECT 24.73 89.73 24.94 89.8 ;
    RECT 24.73 90.09 24.94 90.16 ;
    RECT 25.19 89.37 25.4 89.44 ;
    RECT 25.19 89.73 25.4 89.8 ;
    RECT 25.19 90.09 25.4 90.16 ;
    RECT 21.41 89.37 21.62 89.44 ;
    RECT 21.41 89.73 21.62 89.8 ;
    RECT 21.41 90.09 21.62 90.16 ;
    RECT 21.87 89.37 22.08 89.44 ;
    RECT 21.87 89.73 22.08 89.8 ;
    RECT 21.87 90.09 22.08 90.16 ;
    RECT 18.09 89.37 18.3 89.44 ;
    RECT 18.09 89.73 18.3 89.8 ;
    RECT 18.09 90.09 18.3 90.16 ;
    RECT 18.55 89.37 18.76 89.44 ;
    RECT 18.55 89.73 18.76 89.8 ;
    RECT 18.55 90.09 18.76 90.16 ;
    RECT 120.825 89.73 120.895 89.8 ;
    RECT 14.77 89.37 14.98 89.44 ;
    RECT 14.77 89.73 14.98 89.8 ;
    RECT 14.77 90.09 14.98 90.16 ;
    RECT 15.23 89.37 15.44 89.44 ;
    RECT 15.23 89.73 15.44 89.8 ;
    RECT 15.23 90.09 15.44 90.16 ;
    RECT 11.45 89.37 11.66 89.44 ;
    RECT 11.45 89.73 11.66 89.8 ;
    RECT 11.45 90.09 11.66 90.16 ;
    RECT 11.91 89.37 12.12 89.44 ;
    RECT 11.91 89.73 12.12 89.8 ;
    RECT 11.91 90.09 12.12 90.16 ;
    RECT 8.13 89.37 8.34 89.44 ;
    RECT 8.13 89.73 8.34 89.8 ;
    RECT 8.13 90.09 8.34 90.16 ;
    RECT 8.59 89.37 8.8 89.44 ;
    RECT 8.59 89.73 8.8 89.8 ;
    RECT 8.59 90.09 8.8 90.16 ;
    RECT 4.81 89.37 5.02 89.44 ;
    RECT 4.81 89.73 5.02 89.8 ;
    RECT 4.81 90.09 5.02 90.16 ;
    RECT 5.27 89.37 5.48 89.44 ;
    RECT 5.27 89.73 5.48 89.8 ;
    RECT 5.27 90.09 5.48 90.16 ;
    RECT 1.49 89.37 1.7 89.44 ;
    RECT 1.49 89.73 1.7 89.8 ;
    RECT 1.49 90.09 1.7 90.16 ;
    RECT 1.95 89.37 2.16 89.44 ;
    RECT 1.95 89.73 2.16 89.8 ;
    RECT 1.95 90.09 2.16 90.16 ;
    RECT 64.57 89.37 64.78 89.44 ;
    RECT 64.57 89.73 64.78 89.8 ;
    RECT 64.57 90.09 64.78 90.16 ;
    RECT 65.03 89.37 65.24 89.44 ;
    RECT 65.03 89.73 65.24 89.8 ;
    RECT 65.03 90.09 65.24 90.16 ;
    RECT 61.25 14.47 61.46 14.54 ;
    RECT 61.25 14.83 61.46 14.9 ;
    RECT 61.25 15.19 61.46 15.26 ;
    RECT 61.71 14.47 61.92 14.54 ;
    RECT 61.71 14.83 61.92 14.9 ;
    RECT 61.71 15.19 61.92 15.26 ;
    RECT 57.93 14.47 58.14 14.54 ;
    RECT 57.93 14.83 58.14 14.9 ;
    RECT 57.93 15.19 58.14 15.26 ;
    RECT 58.39 14.47 58.6 14.54 ;
    RECT 58.39 14.83 58.6 14.9 ;
    RECT 58.39 15.19 58.6 15.26 ;
    RECT 54.61 14.47 54.82 14.54 ;
    RECT 54.61 14.83 54.82 14.9 ;
    RECT 54.61 15.19 54.82 15.26 ;
    RECT 55.07 14.47 55.28 14.54 ;
    RECT 55.07 14.83 55.28 14.9 ;
    RECT 55.07 15.19 55.28 15.26 ;
    RECT 51.29 14.47 51.5 14.54 ;
    RECT 51.29 14.83 51.5 14.9 ;
    RECT 51.29 15.19 51.5 15.26 ;
    RECT 51.75 14.47 51.96 14.54 ;
    RECT 51.75 14.83 51.96 14.9 ;
    RECT 51.75 15.19 51.96 15.26 ;
    RECT 47.97 14.47 48.18 14.54 ;
    RECT 47.97 14.83 48.18 14.9 ;
    RECT 47.97 15.19 48.18 15.26 ;
    RECT 48.43 14.47 48.64 14.54 ;
    RECT 48.43 14.83 48.64 14.9 ;
    RECT 48.43 15.19 48.64 15.26 ;
    RECT 44.65 14.47 44.86 14.54 ;
    RECT 44.65 14.83 44.86 14.9 ;
    RECT 44.65 15.19 44.86 15.26 ;
    RECT 45.11 14.47 45.32 14.54 ;
    RECT 45.11 14.83 45.32 14.9 ;
    RECT 45.11 15.19 45.32 15.26 ;
    RECT 41.33 14.47 41.54 14.54 ;
    RECT 41.33 14.83 41.54 14.9 ;
    RECT 41.33 15.19 41.54 15.26 ;
    RECT 41.79 14.47 42.0 14.54 ;
    RECT 41.79 14.83 42.0 14.9 ;
    RECT 41.79 15.19 42.0 15.26 ;
    RECT 38.01 14.47 38.22 14.54 ;
    RECT 38.01 14.83 38.22 14.9 ;
    RECT 38.01 15.19 38.22 15.26 ;
    RECT 38.47 14.47 38.68 14.54 ;
    RECT 38.47 14.83 38.68 14.9 ;
    RECT 38.47 15.19 38.68 15.26 ;
    RECT 34.69 14.47 34.9 14.54 ;
    RECT 34.69 14.83 34.9 14.9 ;
    RECT 34.69 15.19 34.9 15.26 ;
    RECT 35.15 14.47 35.36 14.54 ;
    RECT 35.15 14.83 35.36 14.9 ;
    RECT 35.15 15.19 35.36 15.26 ;
    RECT 0.4 14.83 0.47 14.9 ;
    RECT 114.37 14.47 114.58 14.54 ;
    RECT 114.37 14.83 114.58 14.9 ;
    RECT 114.37 15.19 114.58 15.26 ;
    RECT 114.83 14.47 115.04 14.54 ;
    RECT 114.83 14.83 115.04 14.9 ;
    RECT 114.83 15.19 115.04 15.26 ;
    RECT 111.05 14.47 111.26 14.54 ;
    RECT 111.05 14.83 111.26 14.9 ;
    RECT 111.05 15.19 111.26 15.26 ;
    RECT 111.51 14.47 111.72 14.54 ;
    RECT 111.51 14.83 111.72 14.9 ;
    RECT 111.51 15.19 111.72 15.26 ;
    RECT 107.73 14.47 107.94 14.54 ;
    RECT 107.73 14.83 107.94 14.9 ;
    RECT 107.73 15.19 107.94 15.26 ;
    RECT 108.19 14.47 108.4 14.54 ;
    RECT 108.19 14.83 108.4 14.9 ;
    RECT 108.19 15.19 108.4 15.26 ;
    RECT 104.41 14.47 104.62 14.54 ;
    RECT 104.41 14.83 104.62 14.9 ;
    RECT 104.41 15.19 104.62 15.26 ;
    RECT 104.87 14.47 105.08 14.54 ;
    RECT 104.87 14.83 105.08 14.9 ;
    RECT 104.87 15.19 105.08 15.26 ;
    RECT 101.09 14.47 101.3 14.54 ;
    RECT 101.09 14.83 101.3 14.9 ;
    RECT 101.09 15.19 101.3 15.26 ;
    RECT 101.55 14.47 101.76 14.54 ;
    RECT 101.55 14.83 101.76 14.9 ;
    RECT 101.55 15.19 101.76 15.26 ;
    RECT 97.77 14.47 97.98 14.54 ;
    RECT 97.77 14.83 97.98 14.9 ;
    RECT 97.77 15.19 97.98 15.26 ;
    RECT 98.23 14.47 98.44 14.54 ;
    RECT 98.23 14.83 98.44 14.9 ;
    RECT 98.23 15.19 98.44 15.26 ;
    RECT 94.45 14.47 94.66 14.54 ;
    RECT 94.45 14.83 94.66 14.9 ;
    RECT 94.45 15.19 94.66 15.26 ;
    RECT 94.91 14.47 95.12 14.54 ;
    RECT 94.91 14.83 95.12 14.9 ;
    RECT 94.91 15.19 95.12 15.26 ;
    RECT 91.13 14.47 91.34 14.54 ;
    RECT 91.13 14.83 91.34 14.9 ;
    RECT 91.13 15.19 91.34 15.26 ;
    RECT 91.59 14.47 91.8 14.54 ;
    RECT 91.59 14.83 91.8 14.9 ;
    RECT 91.59 15.19 91.8 15.26 ;
    RECT 87.81 14.47 88.02 14.54 ;
    RECT 87.81 14.83 88.02 14.9 ;
    RECT 87.81 15.19 88.02 15.26 ;
    RECT 88.27 14.47 88.48 14.54 ;
    RECT 88.27 14.83 88.48 14.9 ;
    RECT 88.27 15.19 88.48 15.26 ;
    RECT 84.49 14.47 84.7 14.54 ;
    RECT 84.49 14.83 84.7 14.9 ;
    RECT 84.49 15.19 84.7 15.26 ;
    RECT 84.95 14.47 85.16 14.54 ;
    RECT 84.95 14.83 85.16 14.9 ;
    RECT 84.95 15.19 85.16 15.26 ;
    RECT 81.17 14.47 81.38 14.54 ;
    RECT 81.17 14.83 81.38 14.9 ;
    RECT 81.17 15.19 81.38 15.26 ;
    RECT 81.63 14.47 81.84 14.54 ;
    RECT 81.63 14.83 81.84 14.9 ;
    RECT 81.63 15.19 81.84 15.26 ;
    RECT 77.85 14.47 78.06 14.54 ;
    RECT 77.85 14.83 78.06 14.9 ;
    RECT 77.85 15.19 78.06 15.26 ;
    RECT 78.31 14.47 78.52 14.54 ;
    RECT 78.31 14.83 78.52 14.9 ;
    RECT 78.31 15.19 78.52 15.26 ;
    RECT 74.53 14.47 74.74 14.54 ;
    RECT 74.53 14.83 74.74 14.9 ;
    RECT 74.53 15.19 74.74 15.26 ;
    RECT 74.99 14.47 75.2 14.54 ;
    RECT 74.99 14.83 75.2 14.9 ;
    RECT 74.99 15.19 75.2 15.26 ;
    RECT 71.21 14.47 71.42 14.54 ;
    RECT 71.21 14.83 71.42 14.9 ;
    RECT 71.21 15.19 71.42 15.26 ;
    RECT 71.67 14.47 71.88 14.54 ;
    RECT 71.67 14.83 71.88 14.9 ;
    RECT 71.67 15.19 71.88 15.26 ;
    RECT 31.37 14.47 31.58 14.54 ;
    RECT 31.37 14.83 31.58 14.9 ;
    RECT 31.37 15.19 31.58 15.26 ;
    RECT 31.83 14.47 32.04 14.54 ;
    RECT 31.83 14.83 32.04 14.9 ;
    RECT 31.83 15.19 32.04 15.26 ;
    RECT 67.89 14.47 68.1 14.54 ;
    RECT 67.89 14.83 68.1 14.9 ;
    RECT 67.89 15.19 68.1 15.26 ;
    RECT 68.35 14.47 68.56 14.54 ;
    RECT 68.35 14.83 68.56 14.9 ;
    RECT 68.35 15.19 68.56 15.26 ;
    RECT 28.05 14.47 28.26 14.54 ;
    RECT 28.05 14.83 28.26 14.9 ;
    RECT 28.05 15.19 28.26 15.26 ;
    RECT 28.51 14.47 28.72 14.54 ;
    RECT 28.51 14.83 28.72 14.9 ;
    RECT 28.51 15.19 28.72 15.26 ;
    RECT 24.73 14.47 24.94 14.54 ;
    RECT 24.73 14.83 24.94 14.9 ;
    RECT 24.73 15.19 24.94 15.26 ;
    RECT 25.19 14.47 25.4 14.54 ;
    RECT 25.19 14.83 25.4 14.9 ;
    RECT 25.19 15.19 25.4 15.26 ;
    RECT 21.41 14.47 21.62 14.54 ;
    RECT 21.41 14.83 21.62 14.9 ;
    RECT 21.41 15.19 21.62 15.26 ;
    RECT 21.87 14.47 22.08 14.54 ;
    RECT 21.87 14.83 22.08 14.9 ;
    RECT 21.87 15.19 22.08 15.26 ;
    RECT 18.09 14.47 18.3 14.54 ;
    RECT 18.09 14.83 18.3 14.9 ;
    RECT 18.09 15.19 18.3 15.26 ;
    RECT 18.55 14.47 18.76 14.54 ;
    RECT 18.55 14.83 18.76 14.9 ;
    RECT 18.55 15.19 18.76 15.26 ;
    RECT 14.77 14.47 14.98 14.54 ;
    RECT 14.77 14.83 14.98 14.9 ;
    RECT 14.77 15.19 14.98 15.26 ;
    RECT 15.23 14.47 15.44 14.54 ;
    RECT 15.23 14.83 15.44 14.9 ;
    RECT 15.23 15.19 15.44 15.26 ;
    RECT 11.45 14.47 11.66 14.54 ;
    RECT 11.45 14.83 11.66 14.9 ;
    RECT 11.45 15.19 11.66 15.26 ;
    RECT 11.91 14.47 12.12 14.54 ;
    RECT 11.91 14.83 12.12 14.9 ;
    RECT 11.91 15.19 12.12 15.26 ;
    RECT 8.13 14.47 8.34 14.54 ;
    RECT 8.13 14.83 8.34 14.9 ;
    RECT 8.13 15.19 8.34 15.26 ;
    RECT 8.59 14.47 8.8 14.54 ;
    RECT 8.59 14.83 8.8 14.9 ;
    RECT 8.59 15.19 8.8 15.26 ;
    RECT 120.825 14.83 120.895 14.9 ;
    RECT 4.81 14.47 5.02 14.54 ;
    RECT 4.81 14.83 5.02 14.9 ;
    RECT 4.81 15.19 5.02 15.26 ;
    RECT 5.27 14.47 5.48 14.54 ;
    RECT 5.27 14.83 5.48 14.9 ;
    RECT 5.27 15.19 5.48 15.26 ;
    RECT 117.69 14.47 117.9 14.54 ;
    RECT 117.69 14.83 117.9 14.9 ;
    RECT 117.69 15.19 117.9 15.26 ;
    RECT 118.15 14.47 118.36 14.54 ;
    RECT 118.15 14.83 118.36 14.9 ;
    RECT 118.15 15.19 118.36 15.26 ;
    RECT 1.49 14.47 1.7 14.54 ;
    RECT 1.49 14.83 1.7 14.9 ;
    RECT 1.49 15.19 1.7 15.26 ;
    RECT 1.95 14.47 2.16 14.54 ;
    RECT 1.95 14.83 2.16 14.9 ;
    RECT 1.95 15.19 2.16 15.26 ;
    RECT 64.57 14.47 64.78 14.54 ;
    RECT 64.57 14.83 64.78 14.9 ;
    RECT 64.57 15.19 64.78 15.26 ;
    RECT 65.03 14.47 65.24 14.54 ;
    RECT 65.03 14.83 65.24 14.9 ;
    RECT 65.03 15.19 65.24 15.26 ;
    RECT 61.25 88.65 61.46 88.72 ;
    RECT 61.25 89.01 61.46 89.08 ;
    RECT 61.25 89.37 61.46 89.44 ;
    RECT 61.71 88.65 61.92 88.72 ;
    RECT 61.71 89.01 61.92 89.08 ;
    RECT 61.71 89.37 61.92 89.44 ;
    RECT 57.93 88.65 58.14 88.72 ;
    RECT 57.93 89.01 58.14 89.08 ;
    RECT 57.93 89.37 58.14 89.44 ;
    RECT 58.39 88.65 58.6 88.72 ;
    RECT 58.39 89.01 58.6 89.08 ;
    RECT 58.39 89.37 58.6 89.44 ;
    RECT 54.61 88.65 54.82 88.72 ;
    RECT 54.61 89.01 54.82 89.08 ;
    RECT 54.61 89.37 54.82 89.44 ;
    RECT 55.07 88.65 55.28 88.72 ;
    RECT 55.07 89.01 55.28 89.08 ;
    RECT 55.07 89.37 55.28 89.44 ;
    RECT 51.29 88.65 51.5 88.72 ;
    RECT 51.29 89.01 51.5 89.08 ;
    RECT 51.29 89.37 51.5 89.44 ;
    RECT 51.75 88.65 51.96 88.72 ;
    RECT 51.75 89.01 51.96 89.08 ;
    RECT 51.75 89.37 51.96 89.44 ;
    RECT 47.97 88.65 48.18 88.72 ;
    RECT 47.97 89.01 48.18 89.08 ;
    RECT 47.97 89.37 48.18 89.44 ;
    RECT 48.43 88.65 48.64 88.72 ;
    RECT 48.43 89.01 48.64 89.08 ;
    RECT 48.43 89.37 48.64 89.44 ;
    RECT 44.65 88.65 44.86 88.72 ;
    RECT 44.65 89.01 44.86 89.08 ;
    RECT 44.65 89.37 44.86 89.44 ;
    RECT 45.11 88.65 45.32 88.72 ;
    RECT 45.11 89.01 45.32 89.08 ;
    RECT 45.11 89.37 45.32 89.44 ;
    RECT 41.33 88.65 41.54 88.72 ;
    RECT 41.33 89.01 41.54 89.08 ;
    RECT 41.33 89.37 41.54 89.44 ;
    RECT 41.79 88.65 42.0 88.72 ;
    RECT 41.79 89.01 42.0 89.08 ;
    RECT 41.79 89.37 42.0 89.44 ;
    RECT 38.01 88.65 38.22 88.72 ;
    RECT 38.01 89.01 38.22 89.08 ;
    RECT 38.01 89.37 38.22 89.44 ;
    RECT 38.47 88.65 38.68 88.72 ;
    RECT 38.47 89.01 38.68 89.08 ;
    RECT 38.47 89.37 38.68 89.44 ;
    RECT 0.4 89.01 0.47 89.08 ;
    RECT 34.69 88.65 34.9 88.72 ;
    RECT 34.69 89.01 34.9 89.08 ;
    RECT 34.69 89.37 34.9 89.44 ;
    RECT 35.15 88.65 35.36 88.72 ;
    RECT 35.15 89.01 35.36 89.08 ;
    RECT 35.15 89.37 35.36 89.44 ;
    RECT 117.69 88.65 117.9 88.72 ;
    RECT 117.69 89.01 117.9 89.08 ;
    RECT 117.69 89.37 117.9 89.44 ;
    RECT 118.15 88.65 118.36 88.72 ;
    RECT 118.15 89.01 118.36 89.08 ;
    RECT 118.15 89.37 118.36 89.44 ;
    RECT 114.37 88.65 114.58 88.72 ;
    RECT 114.37 89.01 114.58 89.08 ;
    RECT 114.37 89.37 114.58 89.44 ;
    RECT 114.83 88.65 115.04 88.72 ;
    RECT 114.83 89.01 115.04 89.08 ;
    RECT 114.83 89.37 115.04 89.44 ;
    RECT 111.05 88.65 111.26 88.72 ;
    RECT 111.05 89.01 111.26 89.08 ;
    RECT 111.05 89.37 111.26 89.44 ;
    RECT 111.51 88.65 111.72 88.72 ;
    RECT 111.51 89.01 111.72 89.08 ;
    RECT 111.51 89.37 111.72 89.44 ;
    RECT 107.73 88.65 107.94 88.72 ;
    RECT 107.73 89.01 107.94 89.08 ;
    RECT 107.73 89.37 107.94 89.44 ;
    RECT 108.19 88.65 108.4 88.72 ;
    RECT 108.19 89.01 108.4 89.08 ;
    RECT 108.19 89.37 108.4 89.44 ;
    RECT 104.41 88.65 104.62 88.72 ;
    RECT 104.41 89.01 104.62 89.08 ;
    RECT 104.41 89.37 104.62 89.44 ;
    RECT 104.87 88.65 105.08 88.72 ;
    RECT 104.87 89.01 105.08 89.08 ;
    RECT 104.87 89.37 105.08 89.44 ;
    RECT 101.09 88.65 101.3 88.72 ;
    RECT 101.09 89.01 101.3 89.08 ;
    RECT 101.09 89.37 101.3 89.44 ;
    RECT 101.55 88.65 101.76 88.72 ;
    RECT 101.55 89.01 101.76 89.08 ;
    RECT 101.55 89.37 101.76 89.44 ;
    RECT 97.77 88.65 97.98 88.72 ;
    RECT 97.77 89.01 97.98 89.08 ;
    RECT 97.77 89.37 97.98 89.44 ;
    RECT 98.23 88.65 98.44 88.72 ;
    RECT 98.23 89.01 98.44 89.08 ;
    RECT 98.23 89.37 98.44 89.44 ;
    RECT 94.45 88.65 94.66 88.72 ;
    RECT 94.45 89.01 94.66 89.08 ;
    RECT 94.45 89.37 94.66 89.44 ;
    RECT 94.91 88.65 95.12 88.72 ;
    RECT 94.91 89.01 95.12 89.08 ;
    RECT 94.91 89.37 95.12 89.44 ;
    RECT 91.13 88.65 91.34 88.72 ;
    RECT 91.13 89.01 91.34 89.08 ;
    RECT 91.13 89.37 91.34 89.44 ;
    RECT 91.59 88.65 91.8 88.72 ;
    RECT 91.59 89.01 91.8 89.08 ;
    RECT 91.59 89.37 91.8 89.44 ;
    RECT 87.81 88.65 88.02 88.72 ;
    RECT 87.81 89.01 88.02 89.08 ;
    RECT 87.81 89.37 88.02 89.44 ;
    RECT 88.27 88.65 88.48 88.72 ;
    RECT 88.27 89.01 88.48 89.08 ;
    RECT 88.27 89.37 88.48 89.44 ;
    RECT 84.49 88.65 84.7 88.72 ;
    RECT 84.49 89.01 84.7 89.08 ;
    RECT 84.49 89.37 84.7 89.44 ;
    RECT 84.95 88.65 85.16 88.72 ;
    RECT 84.95 89.01 85.16 89.08 ;
    RECT 84.95 89.37 85.16 89.44 ;
    RECT 81.17 88.65 81.38 88.72 ;
    RECT 81.17 89.01 81.38 89.08 ;
    RECT 81.17 89.37 81.38 89.44 ;
    RECT 81.63 88.65 81.84 88.72 ;
    RECT 81.63 89.01 81.84 89.08 ;
    RECT 81.63 89.37 81.84 89.44 ;
    RECT 77.85 88.65 78.06 88.72 ;
    RECT 77.85 89.01 78.06 89.08 ;
    RECT 77.85 89.37 78.06 89.44 ;
    RECT 78.31 88.65 78.52 88.72 ;
    RECT 78.31 89.01 78.52 89.08 ;
    RECT 78.31 89.37 78.52 89.44 ;
    RECT 74.53 88.65 74.74 88.72 ;
    RECT 74.53 89.01 74.74 89.08 ;
    RECT 74.53 89.37 74.74 89.44 ;
    RECT 74.99 88.65 75.2 88.72 ;
    RECT 74.99 89.01 75.2 89.08 ;
    RECT 74.99 89.37 75.2 89.44 ;
    RECT 71.21 88.65 71.42 88.72 ;
    RECT 71.21 89.01 71.42 89.08 ;
    RECT 71.21 89.37 71.42 89.44 ;
    RECT 71.67 88.65 71.88 88.72 ;
    RECT 71.67 89.01 71.88 89.08 ;
    RECT 71.67 89.37 71.88 89.44 ;
    RECT 31.37 88.65 31.58 88.72 ;
    RECT 31.37 89.01 31.58 89.08 ;
    RECT 31.37 89.37 31.58 89.44 ;
    RECT 31.83 88.65 32.04 88.72 ;
    RECT 31.83 89.01 32.04 89.08 ;
    RECT 31.83 89.37 32.04 89.44 ;
    RECT 67.89 88.65 68.1 88.72 ;
    RECT 67.89 89.01 68.1 89.08 ;
    RECT 67.89 89.37 68.1 89.44 ;
    RECT 68.35 88.65 68.56 88.72 ;
    RECT 68.35 89.01 68.56 89.08 ;
    RECT 68.35 89.37 68.56 89.44 ;
    RECT 28.05 88.65 28.26 88.72 ;
    RECT 28.05 89.01 28.26 89.08 ;
    RECT 28.05 89.37 28.26 89.44 ;
    RECT 28.51 88.65 28.72 88.72 ;
    RECT 28.51 89.01 28.72 89.08 ;
    RECT 28.51 89.37 28.72 89.44 ;
    RECT 24.73 88.65 24.94 88.72 ;
    RECT 24.73 89.01 24.94 89.08 ;
    RECT 24.73 89.37 24.94 89.44 ;
    RECT 25.19 88.65 25.4 88.72 ;
    RECT 25.19 89.01 25.4 89.08 ;
    RECT 25.19 89.37 25.4 89.44 ;
    RECT 21.41 88.65 21.62 88.72 ;
    RECT 21.41 89.01 21.62 89.08 ;
    RECT 21.41 89.37 21.62 89.44 ;
    RECT 21.87 88.65 22.08 88.72 ;
    RECT 21.87 89.01 22.08 89.08 ;
    RECT 21.87 89.37 22.08 89.44 ;
    RECT 18.09 88.65 18.3 88.72 ;
    RECT 18.09 89.01 18.3 89.08 ;
    RECT 18.09 89.37 18.3 89.44 ;
    RECT 18.55 88.65 18.76 88.72 ;
    RECT 18.55 89.01 18.76 89.08 ;
    RECT 18.55 89.37 18.76 89.44 ;
    RECT 120.825 89.01 120.895 89.08 ;
    RECT 14.77 88.65 14.98 88.72 ;
    RECT 14.77 89.01 14.98 89.08 ;
    RECT 14.77 89.37 14.98 89.44 ;
    RECT 15.23 88.65 15.44 88.72 ;
    RECT 15.23 89.01 15.44 89.08 ;
    RECT 15.23 89.37 15.44 89.44 ;
    RECT 11.45 88.65 11.66 88.72 ;
    RECT 11.45 89.01 11.66 89.08 ;
    RECT 11.45 89.37 11.66 89.44 ;
    RECT 11.91 88.65 12.12 88.72 ;
    RECT 11.91 89.01 12.12 89.08 ;
    RECT 11.91 89.37 12.12 89.44 ;
    RECT 8.13 88.65 8.34 88.72 ;
    RECT 8.13 89.01 8.34 89.08 ;
    RECT 8.13 89.37 8.34 89.44 ;
    RECT 8.59 88.65 8.8 88.72 ;
    RECT 8.59 89.01 8.8 89.08 ;
    RECT 8.59 89.37 8.8 89.44 ;
    RECT 4.81 88.65 5.02 88.72 ;
    RECT 4.81 89.01 5.02 89.08 ;
    RECT 4.81 89.37 5.02 89.44 ;
    RECT 5.27 88.65 5.48 88.72 ;
    RECT 5.27 89.01 5.48 89.08 ;
    RECT 5.27 89.37 5.48 89.44 ;
    RECT 1.49 88.65 1.7 88.72 ;
    RECT 1.49 89.01 1.7 89.08 ;
    RECT 1.49 89.37 1.7 89.44 ;
    RECT 1.95 88.65 2.16 88.72 ;
    RECT 1.95 89.01 2.16 89.08 ;
    RECT 1.95 89.37 2.16 89.44 ;
    RECT 64.57 88.65 64.78 88.72 ;
    RECT 64.57 89.01 64.78 89.08 ;
    RECT 64.57 89.37 64.78 89.44 ;
    RECT 65.03 88.65 65.24 88.72 ;
    RECT 65.03 89.01 65.24 89.08 ;
    RECT 65.03 89.37 65.24 89.44 ;
    RECT 61.25 20.95 61.46 21.02 ;
    RECT 61.25 21.31 61.46 21.38 ;
    RECT 61.25 21.67 61.46 21.74 ;
    RECT 61.71 20.95 61.92 21.02 ;
    RECT 61.71 21.31 61.92 21.38 ;
    RECT 61.71 21.67 61.92 21.74 ;
    RECT 57.93 20.95 58.14 21.02 ;
    RECT 57.93 21.31 58.14 21.38 ;
    RECT 57.93 21.67 58.14 21.74 ;
    RECT 58.39 20.95 58.6 21.02 ;
    RECT 58.39 21.31 58.6 21.38 ;
    RECT 58.39 21.67 58.6 21.74 ;
    RECT 54.61 20.95 54.82 21.02 ;
    RECT 54.61 21.31 54.82 21.38 ;
    RECT 54.61 21.67 54.82 21.74 ;
    RECT 55.07 20.95 55.28 21.02 ;
    RECT 55.07 21.31 55.28 21.38 ;
    RECT 55.07 21.67 55.28 21.74 ;
    RECT 51.29 20.95 51.5 21.02 ;
    RECT 51.29 21.31 51.5 21.38 ;
    RECT 51.29 21.67 51.5 21.74 ;
    RECT 51.75 20.95 51.96 21.02 ;
    RECT 51.75 21.31 51.96 21.38 ;
    RECT 51.75 21.67 51.96 21.74 ;
    RECT 47.97 20.95 48.18 21.02 ;
    RECT 47.97 21.31 48.18 21.38 ;
    RECT 47.97 21.67 48.18 21.74 ;
    RECT 48.43 20.95 48.64 21.02 ;
    RECT 48.43 21.31 48.64 21.38 ;
    RECT 48.43 21.67 48.64 21.74 ;
    RECT 44.65 20.95 44.86 21.02 ;
    RECT 44.65 21.31 44.86 21.38 ;
    RECT 44.65 21.67 44.86 21.74 ;
    RECT 45.11 20.95 45.32 21.02 ;
    RECT 45.11 21.31 45.32 21.38 ;
    RECT 45.11 21.67 45.32 21.74 ;
    RECT 41.33 20.95 41.54 21.02 ;
    RECT 41.33 21.31 41.54 21.38 ;
    RECT 41.33 21.67 41.54 21.74 ;
    RECT 41.79 20.95 42.0 21.02 ;
    RECT 41.79 21.31 42.0 21.38 ;
    RECT 41.79 21.67 42.0 21.74 ;
    RECT 38.01 20.95 38.22 21.02 ;
    RECT 38.01 21.31 38.22 21.38 ;
    RECT 38.01 21.67 38.22 21.74 ;
    RECT 38.47 20.95 38.68 21.02 ;
    RECT 38.47 21.31 38.68 21.38 ;
    RECT 38.47 21.67 38.68 21.74 ;
    RECT 0.4 21.31 0.47 21.38 ;
    RECT 34.69 20.95 34.9 21.02 ;
    RECT 34.69 21.31 34.9 21.38 ;
    RECT 34.69 21.67 34.9 21.74 ;
    RECT 35.15 20.95 35.36 21.02 ;
    RECT 35.15 21.31 35.36 21.38 ;
    RECT 35.15 21.67 35.36 21.74 ;
    RECT 117.69 20.95 117.9 21.02 ;
    RECT 117.69 21.31 117.9 21.38 ;
    RECT 117.69 21.67 117.9 21.74 ;
    RECT 118.15 20.95 118.36 21.02 ;
    RECT 118.15 21.31 118.36 21.38 ;
    RECT 118.15 21.67 118.36 21.74 ;
    RECT 114.37 20.95 114.58 21.02 ;
    RECT 114.37 21.31 114.58 21.38 ;
    RECT 114.37 21.67 114.58 21.74 ;
    RECT 114.83 20.95 115.04 21.02 ;
    RECT 114.83 21.31 115.04 21.38 ;
    RECT 114.83 21.67 115.04 21.74 ;
    RECT 111.05 20.95 111.26 21.02 ;
    RECT 111.05 21.31 111.26 21.38 ;
    RECT 111.05 21.67 111.26 21.74 ;
    RECT 111.51 20.95 111.72 21.02 ;
    RECT 111.51 21.31 111.72 21.38 ;
    RECT 111.51 21.67 111.72 21.74 ;
    RECT 107.73 20.95 107.94 21.02 ;
    RECT 107.73 21.31 107.94 21.38 ;
    RECT 107.73 21.67 107.94 21.74 ;
    RECT 108.19 20.95 108.4 21.02 ;
    RECT 108.19 21.31 108.4 21.38 ;
    RECT 108.19 21.67 108.4 21.74 ;
    RECT 104.41 20.95 104.62 21.02 ;
    RECT 104.41 21.31 104.62 21.38 ;
    RECT 104.41 21.67 104.62 21.74 ;
    RECT 104.87 20.95 105.08 21.02 ;
    RECT 104.87 21.31 105.08 21.38 ;
    RECT 104.87 21.67 105.08 21.74 ;
    RECT 101.09 20.95 101.3 21.02 ;
    RECT 101.09 21.31 101.3 21.38 ;
    RECT 101.09 21.67 101.3 21.74 ;
    RECT 101.55 20.95 101.76 21.02 ;
    RECT 101.55 21.31 101.76 21.38 ;
    RECT 101.55 21.67 101.76 21.74 ;
    RECT 97.77 20.95 97.98 21.02 ;
    RECT 97.77 21.31 97.98 21.38 ;
    RECT 97.77 21.67 97.98 21.74 ;
    RECT 98.23 20.95 98.44 21.02 ;
    RECT 98.23 21.31 98.44 21.38 ;
    RECT 98.23 21.67 98.44 21.74 ;
    RECT 94.45 20.95 94.66 21.02 ;
    RECT 94.45 21.31 94.66 21.38 ;
    RECT 94.45 21.67 94.66 21.74 ;
    RECT 94.91 20.95 95.12 21.02 ;
    RECT 94.91 21.31 95.12 21.38 ;
    RECT 94.91 21.67 95.12 21.74 ;
    RECT 91.13 20.95 91.34 21.02 ;
    RECT 91.13 21.31 91.34 21.38 ;
    RECT 91.13 21.67 91.34 21.74 ;
    RECT 91.59 20.95 91.8 21.02 ;
    RECT 91.59 21.31 91.8 21.38 ;
    RECT 91.59 21.67 91.8 21.74 ;
    RECT 87.81 20.95 88.02 21.02 ;
    RECT 87.81 21.31 88.02 21.38 ;
    RECT 87.81 21.67 88.02 21.74 ;
    RECT 88.27 20.95 88.48 21.02 ;
    RECT 88.27 21.31 88.48 21.38 ;
    RECT 88.27 21.67 88.48 21.74 ;
    RECT 84.49 20.95 84.7 21.02 ;
    RECT 84.49 21.31 84.7 21.38 ;
    RECT 84.49 21.67 84.7 21.74 ;
    RECT 84.95 20.95 85.16 21.02 ;
    RECT 84.95 21.31 85.16 21.38 ;
    RECT 84.95 21.67 85.16 21.74 ;
    RECT 81.17 20.95 81.38 21.02 ;
    RECT 81.17 21.31 81.38 21.38 ;
    RECT 81.17 21.67 81.38 21.74 ;
    RECT 81.63 20.95 81.84 21.02 ;
    RECT 81.63 21.31 81.84 21.38 ;
    RECT 81.63 21.67 81.84 21.74 ;
    RECT 77.85 20.95 78.06 21.02 ;
    RECT 77.85 21.31 78.06 21.38 ;
    RECT 77.85 21.67 78.06 21.74 ;
    RECT 78.31 20.95 78.52 21.02 ;
    RECT 78.31 21.31 78.52 21.38 ;
    RECT 78.31 21.67 78.52 21.74 ;
    RECT 74.53 20.95 74.74 21.02 ;
    RECT 74.53 21.31 74.74 21.38 ;
    RECT 74.53 21.67 74.74 21.74 ;
    RECT 74.99 20.95 75.2 21.02 ;
    RECT 74.99 21.31 75.2 21.38 ;
    RECT 74.99 21.67 75.2 21.74 ;
    RECT 71.21 20.95 71.42 21.02 ;
    RECT 71.21 21.31 71.42 21.38 ;
    RECT 71.21 21.67 71.42 21.74 ;
    RECT 71.67 20.95 71.88 21.02 ;
    RECT 71.67 21.31 71.88 21.38 ;
    RECT 71.67 21.67 71.88 21.74 ;
    RECT 31.37 20.95 31.58 21.02 ;
    RECT 31.37 21.31 31.58 21.38 ;
    RECT 31.37 21.67 31.58 21.74 ;
    RECT 31.83 20.95 32.04 21.02 ;
    RECT 31.83 21.31 32.04 21.38 ;
    RECT 31.83 21.67 32.04 21.74 ;
    RECT 67.89 20.95 68.1 21.02 ;
    RECT 67.89 21.31 68.1 21.38 ;
    RECT 67.89 21.67 68.1 21.74 ;
    RECT 68.35 20.95 68.56 21.02 ;
    RECT 68.35 21.31 68.56 21.38 ;
    RECT 68.35 21.67 68.56 21.74 ;
    RECT 28.05 20.95 28.26 21.02 ;
    RECT 28.05 21.31 28.26 21.38 ;
    RECT 28.05 21.67 28.26 21.74 ;
    RECT 28.51 20.95 28.72 21.02 ;
    RECT 28.51 21.31 28.72 21.38 ;
    RECT 28.51 21.67 28.72 21.74 ;
    RECT 24.73 20.95 24.94 21.02 ;
    RECT 24.73 21.31 24.94 21.38 ;
    RECT 24.73 21.67 24.94 21.74 ;
    RECT 25.19 20.95 25.4 21.02 ;
    RECT 25.19 21.31 25.4 21.38 ;
    RECT 25.19 21.67 25.4 21.74 ;
    RECT 21.41 20.95 21.62 21.02 ;
    RECT 21.41 21.31 21.62 21.38 ;
    RECT 21.41 21.67 21.62 21.74 ;
    RECT 21.87 20.95 22.08 21.02 ;
    RECT 21.87 21.31 22.08 21.38 ;
    RECT 21.87 21.67 22.08 21.74 ;
    RECT 18.09 20.95 18.3 21.02 ;
    RECT 18.09 21.31 18.3 21.38 ;
    RECT 18.09 21.67 18.3 21.74 ;
    RECT 18.55 20.95 18.76 21.02 ;
    RECT 18.55 21.31 18.76 21.38 ;
    RECT 18.55 21.67 18.76 21.74 ;
    RECT 120.825 21.31 120.895 21.38 ;
    RECT 14.77 20.95 14.98 21.02 ;
    RECT 14.77 21.31 14.98 21.38 ;
    RECT 14.77 21.67 14.98 21.74 ;
    RECT 15.23 20.95 15.44 21.02 ;
    RECT 15.23 21.31 15.44 21.38 ;
    RECT 15.23 21.67 15.44 21.74 ;
    RECT 11.45 20.95 11.66 21.02 ;
    RECT 11.45 21.31 11.66 21.38 ;
    RECT 11.45 21.67 11.66 21.74 ;
    RECT 11.91 20.95 12.12 21.02 ;
    RECT 11.91 21.31 12.12 21.38 ;
    RECT 11.91 21.67 12.12 21.74 ;
    RECT 8.13 20.95 8.34 21.02 ;
    RECT 8.13 21.31 8.34 21.38 ;
    RECT 8.13 21.67 8.34 21.74 ;
    RECT 8.59 20.95 8.8 21.02 ;
    RECT 8.59 21.31 8.8 21.38 ;
    RECT 8.59 21.67 8.8 21.74 ;
    RECT 4.81 20.95 5.02 21.02 ;
    RECT 4.81 21.31 5.02 21.38 ;
    RECT 4.81 21.67 5.02 21.74 ;
    RECT 5.27 20.95 5.48 21.02 ;
    RECT 5.27 21.31 5.48 21.38 ;
    RECT 5.27 21.67 5.48 21.74 ;
    RECT 1.49 20.95 1.7 21.02 ;
    RECT 1.49 21.31 1.7 21.38 ;
    RECT 1.49 21.67 1.7 21.74 ;
    RECT 1.95 20.95 2.16 21.02 ;
    RECT 1.95 21.31 2.16 21.38 ;
    RECT 1.95 21.67 2.16 21.74 ;
    RECT 64.57 20.95 64.78 21.02 ;
    RECT 64.57 21.31 64.78 21.38 ;
    RECT 64.57 21.67 64.78 21.74 ;
    RECT 65.03 20.95 65.24 21.02 ;
    RECT 65.03 21.31 65.24 21.38 ;
    RECT 65.03 21.67 65.24 21.74 ;
    RECT 61.25 87.93 61.46 88.0 ;
    RECT 61.25 88.29 61.46 88.36 ;
    RECT 61.25 88.65 61.46 88.72 ;
    RECT 61.71 87.93 61.92 88.0 ;
    RECT 61.71 88.29 61.92 88.36 ;
    RECT 61.71 88.65 61.92 88.72 ;
    RECT 57.93 87.93 58.14 88.0 ;
    RECT 57.93 88.29 58.14 88.36 ;
    RECT 57.93 88.65 58.14 88.72 ;
    RECT 58.39 87.93 58.6 88.0 ;
    RECT 58.39 88.29 58.6 88.36 ;
    RECT 58.39 88.65 58.6 88.72 ;
    RECT 54.61 87.93 54.82 88.0 ;
    RECT 54.61 88.29 54.82 88.36 ;
    RECT 54.61 88.65 54.82 88.72 ;
    RECT 55.07 87.93 55.28 88.0 ;
    RECT 55.07 88.29 55.28 88.36 ;
    RECT 55.07 88.65 55.28 88.72 ;
    RECT 51.29 87.93 51.5 88.0 ;
    RECT 51.29 88.29 51.5 88.36 ;
    RECT 51.29 88.65 51.5 88.72 ;
    RECT 51.75 87.93 51.96 88.0 ;
    RECT 51.75 88.29 51.96 88.36 ;
    RECT 51.75 88.65 51.96 88.72 ;
    RECT 47.97 87.93 48.18 88.0 ;
    RECT 47.97 88.29 48.18 88.36 ;
    RECT 47.97 88.65 48.18 88.72 ;
    RECT 48.43 87.93 48.64 88.0 ;
    RECT 48.43 88.29 48.64 88.36 ;
    RECT 48.43 88.65 48.64 88.72 ;
    RECT 44.65 87.93 44.86 88.0 ;
    RECT 44.65 88.29 44.86 88.36 ;
    RECT 44.65 88.65 44.86 88.72 ;
    RECT 45.11 87.93 45.32 88.0 ;
    RECT 45.11 88.29 45.32 88.36 ;
    RECT 45.11 88.65 45.32 88.72 ;
    RECT 41.33 87.93 41.54 88.0 ;
    RECT 41.33 88.29 41.54 88.36 ;
    RECT 41.33 88.65 41.54 88.72 ;
    RECT 41.79 87.93 42.0 88.0 ;
    RECT 41.79 88.29 42.0 88.36 ;
    RECT 41.79 88.65 42.0 88.72 ;
    RECT 38.01 87.93 38.22 88.0 ;
    RECT 38.01 88.29 38.22 88.36 ;
    RECT 38.01 88.65 38.22 88.72 ;
    RECT 38.47 87.93 38.68 88.0 ;
    RECT 38.47 88.29 38.68 88.36 ;
    RECT 38.47 88.65 38.68 88.72 ;
    RECT 0.4 88.29 0.47 88.36 ;
    RECT 34.69 87.93 34.9 88.0 ;
    RECT 34.69 88.29 34.9 88.36 ;
    RECT 34.69 88.65 34.9 88.72 ;
    RECT 35.15 87.93 35.36 88.0 ;
    RECT 35.15 88.29 35.36 88.36 ;
    RECT 35.15 88.65 35.36 88.72 ;
    RECT 117.69 87.93 117.9 88.0 ;
    RECT 117.69 88.29 117.9 88.36 ;
    RECT 117.69 88.65 117.9 88.72 ;
    RECT 118.15 87.93 118.36 88.0 ;
    RECT 118.15 88.29 118.36 88.36 ;
    RECT 118.15 88.65 118.36 88.72 ;
    RECT 114.37 87.93 114.58 88.0 ;
    RECT 114.37 88.29 114.58 88.36 ;
    RECT 114.37 88.65 114.58 88.72 ;
    RECT 114.83 87.93 115.04 88.0 ;
    RECT 114.83 88.29 115.04 88.36 ;
    RECT 114.83 88.65 115.04 88.72 ;
    RECT 111.05 87.93 111.26 88.0 ;
    RECT 111.05 88.29 111.26 88.36 ;
    RECT 111.05 88.65 111.26 88.72 ;
    RECT 111.51 87.93 111.72 88.0 ;
    RECT 111.51 88.29 111.72 88.36 ;
    RECT 111.51 88.65 111.72 88.72 ;
    RECT 107.73 87.93 107.94 88.0 ;
    RECT 107.73 88.29 107.94 88.36 ;
    RECT 107.73 88.65 107.94 88.72 ;
    RECT 108.19 87.93 108.4 88.0 ;
    RECT 108.19 88.29 108.4 88.36 ;
    RECT 108.19 88.65 108.4 88.72 ;
    RECT 104.41 87.93 104.62 88.0 ;
    RECT 104.41 88.29 104.62 88.36 ;
    RECT 104.41 88.65 104.62 88.72 ;
    RECT 104.87 87.93 105.08 88.0 ;
    RECT 104.87 88.29 105.08 88.36 ;
    RECT 104.87 88.65 105.08 88.72 ;
    RECT 101.09 87.93 101.3 88.0 ;
    RECT 101.09 88.29 101.3 88.36 ;
    RECT 101.09 88.65 101.3 88.72 ;
    RECT 101.55 87.93 101.76 88.0 ;
    RECT 101.55 88.29 101.76 88.36 ;
    RECT 101.55 88.65 101.76 88.72 ;
    RECT 97.77 87.93 97.98 88.0 ;
    RECT 97.77 88.29 97.98 88.36 ;
    RECT 97.77 88.65 97.98 88.72 ;
    RECT 98.23 87.93 98.44 88.0 ;
    RECT 98.23 88.29 98.44 88.36 ;
    RECT 98.23 88.65 98.44 88.72 ;
    RECT 94.45 87.93 94.66 88.0 ;
    RECT 94.45 88.29 94.66 88.36 ;
    RECT 94.45 88.65 94.66 88.72 ;
    RECT 94.91 87.93 95.12 88.0 ;
    RECT 94.91 88.29 95.12 88.36 ;
    RECT 94.91 88.65 95.12 88.72 ;
    RECT 91.13 87.93 91.34 88.0 ;
    RECT 91.13 88.29 91.34 88.36 ;
    RECT 91.13 88.65 91.34 88.72 ;
    RECT 91.59 87.93 91.8 88.0 ;
    RECT 91.59 88.29 91.8 88.36 ;
    RECT 91.59 88.65 91.8 88.72 ;
    RECT 87.81 87.93 88.02 88.0 ;
    RECT 87.81 88.29 88.02 88.36 ;
    RECT 87.81 88.65 88.02 88.72 ;
    RECT 88.27 87.93 88.48 88.0 ;
    RECT 88.27 88.29 88.48 88.36 ;
    RECT 88.27 88.65 88.48 88.72 ;
    RECT 84.49 87.93 84.7 88.0 ;
    RECT 84.49 88.29 84.7 88.36 ;
    RECT 84.49 88.65 84.7 88.72 ;
    RECT 84.95 87.93 85.16 88.0 ;
    RECT 84.95 88.29 85.16 88.36 ;
    RECT 84.95 88.65 85.16 88.72 ;
    RECT 81.17 87.93 81.38 88.0 ;
    RECT 81.17 88.29 81.38 88.36 ;
    RECT 81.17 88.65 81.38 88.72 ;
    RECT 81.63 87.93 81.84 88.0 ;
    RECT 81.63 88.29 81.84 88.36 ;
    RECT 81.63 88.65 81.84 88.72 ;
    RECT 77.85 87.93 78.06 88.0 ;
    RECT 77.85 88.29 78.06 88.36 ;
    RECT 77.85 88.65 78.06 88.72 ;
    RECT 78.31 87.93 78.52 88.0 ;
    RECT 78.31 88.29 78.52 88.36 ;
    RECT 78.31 88.65 78.52 88.72 ;
    RECT 74.53 87.93 74.74 88.0 ;
    RECT 74.53 88.29 74.74 88.36 ;
    RECT 74.53 88.65 74.74 88.72 ;
    RECT 74.99 87.93 75.2 88.0 ;
    RECT 74.99 88.29 75.2 88.36 ;
    RECT 74.99 88.65 75.2 88.72 ;
    RECT 71.21 87.93 71.42 88.0 ;
    RECT 71.21 88.29 71.42 88.36 ;
    RECT 71.21 88.65 71.42 88.72 ;
    RECT 71.67 87.93 71.88 88.0 ;
    RECT 71.67 88.29 71.88 88.36 ;
    RECT 71.67 88.65 71.88 88.72 ;
    RECT 31.37 87.93 31.58 88.0 ;
    RECT 31.37 88.29 31.58 88.36 ;
    RECT 31.37 88.65 31.58 88.72 ;
    RECT 31.83 87.93 32.04 88.0 ;
    RECT 31.83 88.29 32.04 88.36 ;
    RECT 31.83 88.65 32.04 88.72 ;
    RECT 67.89 87.93 68.1 88.0 ;
    RECT 67.89 88.29 68.1 88.36 ;
    RECT 67.89 88.65 68.1 88.72 ;
    RECT 68.35 87.93 68.56 88.0 ;
    RECT 68.35 88.29 68.56 88.36 ;
    RECT 68.35 88.65 68.56 88.72 ;
    RECT 28.05 87.93 28.26 88.0 ;
    RECT 28.05 88.29 28.26 88.36 ;
    RECT 28.05 88.65 28.26 88.72 ;
    RECT 28.51 87.93 28.72 88.0 ;
    RECT 28.51 88.29 28.72 88.36 ;
    RECT 28.51 88.65 28.72 88.72 ;
    RECT 24.73 87.93 24.94 88.0 ;
    RECT 24.73 88.29 24.94 88.36 ;
    RECT 24.73 88.65 24.94 88.72 ;
    RECT 25.19 87.93 25.4 88.0 ;
    RECT 25.19 88.29 25.4 88.36 ;
    RECT 25.19 88.65 25.4 88.72 ;
    RECT 21.41 87.93 21.62 88.0 ;
    RECT 21.41 88.29 21.62 88.36 ;
    RECT 21.41 88.65 21.62 88.72 ;
    RECT 21.87 87.93 22.08 88.0 ;
    RECT 21.87 88.29 22.08 88.36 ;
    RECT 21.87 88.65 22.08 88.72 ;
    RECT 18.09 87.93 18.3 88.0 ;
    RECT 18.09 88.29 18.3 88.36 ;
    RECT 18.09 88.65 18.3 88.72 ;
    RECT 18.55 87.93 18.76 88.0 ;
    RECT 18.55 88.29 18.76 88.36 ;
    RECT 18.55 88.65 18.76 88.72 ;
    RECT 120.825 88.29 120.895 88.36 ;
    RECT 14.77 87.93 14.98 88.0 ;
    RECT 14.77 88.29 14.98 88.36 ;
    RECT 14.77 88.65 14.98 88.72 ;
    RECT 15.23 87.93 15.44 88.0 ;
    RECT 15.23 88.29 15.44 88.36 ;
    RECT 15.23 88.65 15.44 88.72 ;
    RECT 11.45 87.93 11.66 88.0 ;
    RECT 11.45 88.29 11.66 88.36 ;
    RECT 11.45 88.65 11.66 88.72 ;
    RECT 11.91 87.93 12.12 88.0 ;
    RECT 11.91 88.29 12.12 88.36 ;
    RECT 11.91 88.65 12.12 88.72 ;
    RECT 8.13 87.93 8.34 88.0 ;
    RECT 8.13 88.29 8.34 88.36 ;
    RECT 8.13 88.65 8.34 88.72 ;
    RECT 8.59 87.93 8.8 88.0 ;
    RECT 8.59 88.29 8.8 88.36 ;
    RECT 8.59 88.65 8.8 88.72 ;
    RECT 4.81 87.93 5.02 88.0 ;
    RECT 4.81 88.29 5.02 88.36 ;
    RECT 4.81 88.65 5.02 88.72 ;
    RECT 5.27 87.93 5.48 88.0 ;
    RECT 5.27 88.29 5.48 88.36 ;
    RECT 5.27 88.65 5.48 88.72 ;
    RECT 1.49 87.93 1.7 88.0 ;
    RECT 1.49 88.29 1.7 88.36 ;
    RECT 1.49 88.65 1.7 88.72 ;
    RECT 1.95 87.93 2.16 88.0 ;
    RECT 1.95 88.29 2.16 88.36 ;
    RECT 1.95 88.65 2.16 88.72 ;
    RECT 64.57 87.93 64.78 88.0 ;
    RECT 64.57 88.29 64.78 88.36 ;
    RECT 64.57 88.65 64.78 88.72 ;
    RECT 65.03 87.93 65.24 88.0 ;
    RECT 65.03 88.29 65.24 88.36 ;
    RECT 65.03 88.65 65.24 88.72 ;
    RECT 61.25 20.23 61.46 20.3 ;
    RECT 61.25 20.59 61.46 20.66 ;
    RECT 61.25 20.95 61.46 21.02 ;
    RECT 61.71 20.23 61.92 20.3 ;
    RECT 61.71 20.59 61.92 20.66 ;
    RECT 61.71 20.95 61.92 21.02 ;
    RECT 57.93 20.23 58.14 20.3 ;
    RECT 57.93 20.59 58.14 20.66 ;
    RECT 57.93 20.95 58.14 21.02 ;
    RECT 58.39 20.23 58.6 20.3 ;
    RECT 58.39 20.59 58.6 20.66 ;
    RECT 58.39 20.95 58.6 21.02 ;
    RECT 54.61 20.23 54.82 20.3 ;
    RECT 54.61 20.59 54.82 20.66 ;
    RECT 54.61 20.95 54.82 21.02 ;
    RECT 55.07 20.23 55.28 20.3 ;
    RECT 55.07 20.59 55.28 20.66 ;
    RECT 55.07 20.95 55.28 21.02 ;
    RECT 51.29 20.23 51.5 20.3 ;
    RECT 51.29 20.59 51.5 20.66 ;
    RECT 51.29 20.95 51.5 21.02 ;
    RECT 51.75 20.23 51.96 20.3 ;
    RECT 51.75 20.59 51.96 20.66 ;
    RECT 51.75 20.95 51.96 21.02 ;
    RECT 47.97 20.23 48.18 20.3 ;
    RECT 47.97 20.59 48.18 20.66 ;
    RECT 47.97 20.95 48.18 21.02 ;
    RECT 48.43 20.23 48.64 20.3 ;
    RECT 48.43 20.59 48.64 20.66 ;
    RECT 48.43 20.95 48.64 21.02 ;
    RECT 44.65 20.23 44.86 20.3 ;
    RECT 44.65 20.59 44.86 20.66 ;
    RECT 44.65 20.95 44.86 21.02 ;
    RECT 45.11 20.23 45.32 20.3 ;
    RECT 45.11 20.59 45.32 20.66 ;
    RECT 45.11 20.95 45.32 21.02 ;
    RECT 41.33 20.23 41.54 20.3 ;
    RECT 41.33 20.59 41.54 20.66 ;
    RECT 41.33 20.95 41.54 21.02 ;
    RECT 41.79 20.23 42.0 20.3 ;
    RECT 41.79 20.59 42.0 20.66 ;
    RECT 41.79 20.95 42.0 21.02 ;
    RECT 38.01 20.23 38.22 20.3 ;
    RECT 38.01 20.59 38.22 20.66 ;
    RECT 38.01 20.95 38.22 21.02 ;
    RECT 38.47 20.23 38.68 20.3 ;
    RECT 38.47 20.59 38.68 20.66 ;
    RECT 38.47 20.95 38.68 21.02 ;
    RECT 0.4 20.59 0.47 20.66 ;
    RECT 34.69 20.23 34.9 20.3 ;
    RECT 34.69 20.59 34.9 20.66 ;
    RECT 34.69 20.95 34.9 21.02 ;
    RECT 35.15 20.23 35.36 20.3 ;
    RECT 35.15 20.59 35.36 20.66 ;
    RECT 35.15 20.95 35.36 21.02 ;
    RECT 117.69 20.23 117.9 20.3 ;
    RECT 117.69 20.59 117.9 20.66 ;
    RECT 117.69 20.95 117.9 21.02 ;
    RECT 118.15 20.23 118.36 20.3 ;
    RECT 118.15 20.59 118.36 20.66 ;
    RECT 118.15 20.95 118.36 21.02 ;
    RECT 114.37 20.23 114.58 20.3 ;
    RECT 114.37 20.59 114.58 20.66 ;
    RECT 114.37 20.95 114.58 21.02 ;
    RECT 114.83 20.23 115.04 20.3 ;
    RECT 114.83 20.59 115.04 20.66 ;
    RECT 114.83 20.95 115.04 21.02 ;
    RECT 111.05 20.23 111.26 20.3 ;
    RECT 111.05 20.59 111.26 20.66 ;
    RECT 111.05 20.95 111.26 21.02 ;
    RECT 111.51 20.23 111.72 20.3 ;
    RECT 111.51 20.59 111.72 20.66 ;
    RECT 111.51 20.95 111.72 21.02 ;
    RECT 107.73 20.23 107.94 20.3 ;
    RECT 107.73 20.59 107.94 20.66 ;
    RECT 107.73 20.95 107.94 21.02 ;
    RECT 108.19 20.23 108.4 20.3 ;
    RECT 108.19 20.59 108.4 20.66 ;
    RECT 108.19 20.95 108.4 21.02 ;
    RECT 104.41 20.23 104.62 20.3 ;
    RECT 104.41 20.59 104.62 20.66 ;
    RECT 104.41 20.95 104.62 21.02 ;
    RECT 104.87 20.23 105.08 20.3 ;
    RECT 104.87 20.59 105.08 20.66 ;
    RECT 104.87 20.95 105.08 21.02 ;
    RECT 101.09 20.23 101.3 20.3 ;
    RECT 101.09 20.59 101.3 20.66 ;
    RECT 101.09 20.95 101.3 21.02 ;
    RECT 101.55 20.23 101.76 20.3 ;
    RECT 101.55 20.59 101.76 20.66 ;
    RECT 101.55 20.95 101.76 21.02 ;
    RECT 97.77 20.23 97.98 20.3 ;
    RECT 97.77 20.59 97.98 20.66 ;
    RECT 97.77 20.95 97.98 21.02 ;
    RECT 98.23 20.23 98.44 20.3 ;
    RECT 98.23 20.59 98.44 20.66 ;
    RECT 98.23 20.95 98.44 21.02 ;
    RECT 94.45 20.23 94.66 20.3 ;
    RECT 94.45 20.59 94.66 20.66 ;
    RECT 94.45 20.95 94.66 21.02 ;
    RECT 94.91 20.23 95.12 20.3 ;
    RECT 94.91 20.59 95.12 20.66 ;
    RECT 94.91 20.95 95.12 21.02 ;
    RECT 91.13 20.23 91.34 20.3 ;
    RECT 91.13 20.59 91.34 20.66 ;
    RECT 91.13 20.95 91.34 21.02 ;
    RECT 91.59 20.23 91.8 20.3 ;
    RECT 91.59 20.59 91.8 20.66 ;
    RECT 91.59 20.95 91.8 21.02 ;
    RECT 87.81 20.23 88.02 20.3 ;
    RECT 87.81 20.59 88.02 20.66 ;
    RECT 87.81 20.95 88.02 21.02 ;
    RECT 88.27 20.23 88.48 20.3 ;
    RECT 88.27 20.59 88.48 20.66 ;
    RECT 88.27 20.95 88.48 21.02 ;
    RECT 84.49 20.23 84.7 20.3 ;
    RECT 84.49 20.59 84.7 20.66 ;
    RECT 84.49 20.95 84.7 21.02 ;
    RECT 84.95 20.23 85.16 20.3 ;
    RECT 84.95 20.59 85.16 20.66 ;
    RECT 84.95 20.95 85.16 21.02 ;
    RECT 81.17 20.23 81.38 20.3 ;
    RECT 81.17 20.59 81.38 20.66 ;
    RECT 81.17 20.95 81.38 21.02 ;
    RECT 81.63 20.23 81.84 20.3 ;
    RECT 81.63 20.59 81.84 20.66 ;
    RECT 81.63 20.95 81.84 21.02 ;
    RECT 77.85 20.23 78.06 20.3 ;
    RECT 77.85 20.59 78.06 20.66 ;
    RECT 77.85 20.95 78.06 21.02 ;
    RECT 78.31 20.23 78.52 20.3 ;
    RECT 78.31 20.59 78.52 20.66 ;
    RECT 78.31 20.95 78.52 21.02 ;
    RECT 74.53 20.23 74.74 20.3 ;
    RECT 74.53 20.59 74.74 20.66 ;
    RECT 74.53 20.95 74.74 21.02 ;
    RECT 74.99 20.23 75.2 20.3 ;
    RECT 74.99 20.59 75.2 20.66 ;
    RECT 74.99 20.95 75.2 21.02 ;
    RECT 71.21 20.23 71.42 20.3 ;
    RECT 71.21 20.59 71.42 20.66 ;
    RECT 71.21 20.95 71.42 21.02 ;
    RECT 71.67 20.23 71.88 20.3 ;
    RECT 71.67 20.59 71.88 20.66 ;
    RECT 71.67 20.95 71.88 21.02 ;
    RECT 31.37 20.23 31.58 20.3 ;
    RECT 31.37 20.59 31.58 20.66 ;
    RECT 31.37 20.95 31.58 21.02 ;
    RECT 31.83 20.23 32.04 20.3 ;
    RECT 31.83 20.59 32.04 20.66 ;
    RECT 31.83 20.95 32.04 21.02 ;
    RECT 67.89 20.23 68.1 20.3 ;
    RECT 67.89 20.59 68.1 20.66 ;
    RECT 67.89 20.95 68.1 21.02 ;
    RECT 68.35 20.23 68.56 20.3 ;
    RECT 68.35 20.59 68.56 20.66 ;
    RECT 68.35 20.95 68.56 21.02 ;
    RECT 28.05 20.23 28.26 20.3 ;
    RECT 28.05 20.59 28.26 20.66 ;
    RECT 28.05 20.95 28.26 21.02 ;
    RECT 28.51 20.23 28.72 20.3 ;
    RECT 28.51 20.59 28.72 20.66 ;
    RECT 28.51 20.95 28.72 21.02 ;
    RECT 24.73 20.23 24.94 20.3 ;
    RECT 24.73 20.59 24.94 20.66 ;
    RECT 24.73 20.95 24.94 21.02 ;
    RECT 25.19 20.23 25.4 20.3 ;
    RECT 25.19 20.59 25.4 20.66 ;
    RECT 25.19 20.95 25.4 21.02 ;
    RECT 21.41 20.23 21.62 20.3 ;
    RECT 21.41 20.59 21.62 20.66 ;
    RECT 21.41 20.95 21.62 21.02 ;
    RECT 21.87 20.23 22.08 20.3 ;
    RECT 21.87 20.59 22.08 20.66 ;
    RECT 21.87 20.95 22.08 21.02 ;
    RECT 18.09 20.23 18.3 20.3 ;
    RECT 18.09 20.59 18.3 20.66 ;
    RECT 18.09 20.95 18.3 21.02 ;
    RECT 18.55 20.23 18.76 20.3 ;
    RECT 18.55 20.59 18.76 20.66 ;
    RECT 18.55 20.95 18.76 21.02 ;
    RECT 120.825 20.59 120.895 20.66 ;
    RECT 14.77 20.23 14.98 20.3 ;
    RECT 14.77 20.59 14.98 20.66 ;
    RECT 14.77 20.95 14.98 21.02 ;
    RECT 15.23 20.23 15.44 20.3 ;
    RECT 15.23 20.59 15.44 20.66 ;
    RECT 15.23 20.95 15.44 21.02 ;
    RECT 11.45 20.23 11.66 20.3 ;
    RECT 11.45 20.59 11.66 20.66 ;
    RECT 11.45 20.95 11.66 21.02 ;
    RECT 11.91 20.23 12.12 20.3 ;
    RECT 11.91 20.59 12.12 20.66 ;
    RECT 11.91 20.95 12.12 21.02 ;
    RECT 8.13 20.23 8.34 20.3 ;
    RECT 8.13 20.59 8.34 20.66 ;
    RECT 8.13 20.95 8.34 21.02 ;
    RECT 8.59 20.23 8.8 20.3 ;
    RECT 8.59 20.59 8.8 20.66 ;
    RECT 8.59 20.95 8.8 21.02 ;
    RECT 4.81 20.23 5.02 20.3 ;
    RECT 4.81 20.59 5.02 20.66 ;
    RECT 4.81 20.95 5.02 21.02 ;
    RECT 5.27 20.23 5.48 20.3 ;
    RECT 5.27 20.59 5.48 20.66 ;
    RECT 5.27 20.95 5.48 21.02 ;
    RECT 1.49 20.23 1.7 20.3 ;
    RECT 1.49 20.59 1.7 20.66 ;
    RECT 1.49 20.95 1.7 21.02 ;
    RECT 1.95 20.23 2.16 20.3 ;
    RECT 1.95 20.59 2.16 20.66 ;
    RECT 1.95 20.95 2.16 21.02 ;
    RECT 64.57 20.23 64.78 20.3 ;
    RECT 64.57 20.59 64.78 20.66 ;
    RECT 64.57 20.95 64.78 21.02 ;
    RECT 65.03 20.23 65.24 20.3 ;
    RECT 65.03 20.59 65.24 20.66 ;
    RECT 65.03 20.95 65.24 21.02 ;
    RECT 61.25 87.21 61.46 87.28 ;
    RECT 61.25 87.57 61.46 87.64 ;
    RECT 61.25 87.93 61.46 88.0 ;
    RECT 61.71 87.21 61.92 87.28 ;
    RECT 61.71 87.57 61.92 87.64 ;
    RECT 61.71 87.93 61.92 88.0 ;
    RECT 57.93 87.21 58.14 87.28 ;
    RECT 57.93 87.57 58.14 87.64 ;
    RECT 57.93 87.93 58.14 88.0 ;
    RECT 58.39 87.21 58.6 87.28 ;
    RECT 58.39 87.57 58.6 87.64 ;
    RECT 58.39 87.93 58.6 88.0 ;
    RECT 54.61 87.21 54.82 87.28 ;
    RECT 54.61 87.57 54.82 87.64 ;
    RECT 54.61 87.93 54.82 88.0 ;
    RECT 55.07 87.21 55.28 87.28 ;
    RECT 55.07 87.57 55.28 87.64 ;
    RECT 55.07 87.93 55.28 88.0 ;
    RECT 51.29 87.21 51.5 87.28 ;
    RECT 51.29 87.57 51.5 87.64 ;
    RECT 51.29 87.93 51.5 88.0 ;
    RECT 51.75 87.21 51.96 87.28 ;
    RECT 51.75 87.57 51.96 87.64 ;
    RECT 51.75 87.93 51.96 88.0 ;
    RECT 47.97 87.21 48.18 87.28 ;
    RECT 47.97 87.57 48.18 87.64 ;
    RECT 47.97 87.93 48.18 88.0 ;
    RECT 48.43 87.21 48.64 87.28 ;
    RECT 48.43 87.57 48.64 87.64 ;
    RECT 48.43 87.93 48.64 88.0 ;
    RECT 44.65 87.21 44.86 87.28 ;
    RECT 44.65 87.57 44.86 87.64 ;
    RECT 44.65 87.93 44.86 88.0 ;
    RECT 45.11 87.21 45.32 87.28 ;
    RECT 45.11 87.57 45.32 87.64 ;
    RECT 45.11 87.93 45.32 88.0 ;
    RECT 41.33 87.21 41.54 87.28 ;
    RECT 41.33 87.57 41.54 87.64 ;
    RECT 41.33 87.93 41.54 88.0 ;
    RECT 41.79 87.21 42.0 87.28 ;
    RECT 41.79 87.57 42.0 87.64 ;
    RECT 41.79 87.93 42.0 88.0 ;
    RECT 38.01 87.21 38.22 87.28 ;
    RECT 38.01 87.57 38.22 87.64 ;
    RECT 38.01 87.93 38.22 88.0 ;
    RECT 38.47 87.21 38.68 87.28 ;
    RECT 38.47 87.57 38.68 87.64 ;
    RECT 38.47 87.93 38.68 88.0 ;
    RECT 0.4 87.57 0.47 87.64 ;
    RECT 34.69 87.21 34.9 87.28 ;
    RECT 34.69 87.57 34.9 87.64 ;
    RECT 34.69 87.93 34.9 88.0 ;
    RECT 35.15 87.21 35.36 87.28 ;
    RECT 35.15 87.57 35.36 87.64 ;
    RECT 35.15 87.93 35.36 88.0 ;
    RECT 117.69 87.21 117.9 87.28 ;
    RECT 117.69 87.57 117.9 87.64 ;
    RECT 117.69 87.93 117.9 88.0 ;
    RECT 118.15 87.21 118.36 87.28 ;
    RECT 118.15 87.57 118.36 87.64 ;
    RECT 118.15 87.93 118.36 88.0 ;
    RECT 114.37 87.21 114.58 87.28 ;
    RECT 114.37 87.57 114.58 87.64 ;
    RECT 114.37 87.93 114.58 88.0 ;
    RECT 114.83 87.21 115.04 87.28 ;
    RECT 114.83 87.57 115.04 87.64 ;
    RECT 114.83 87.93 115.04 88.0 ;
    RECT 111.05 87.21 111.26 87.28 ;
    RECT 111.05 87.57 111.26 87.64 ;
    RECT 111.05 87.93 111.26 88.0 ;
    RECT 111.51 87.21 111.72 87.28 ;
    RECT 111.51 87.57 111.72 87.64 ;
    RECT 111.51 87.93 111.72 88.0 ;
    RECT 107.73 87.21 107.94 87.28 ;
    RECT 107.73 87.57 107.94 87.64 ;
    RECT 107.73 87.93 107.94 88.0 ;
    RECT 108.19 87.21 108.4 87.28 ;
    RECT 108.19 87.57 108.4 87.64 ;
    RECT 108.19 87.93 108.4 88.0 ;
    RECT 104.41 87.21 104.62 87.28 ;
    RECT 104.41 87.57 104.62 87.64 ;
    RECT 104.41 87.93 104.62 88.0 ;
    RECT 104.87 87.21 105.08 87.28 ;
    RECT 104.87 87.57 105.08 87.64 ;
    RECT 104.87 87.93 105.08 88.0 ;
    RECT 101.09 87.21 101.3 87.28 ;
    RECT 101.09 87.57 101.3 87.64 ;
    RECT 101.09 87.93 101.3 88.0 ;
    RECT 101.55 87.21 101.76 87.28 ;
    RECT 101.55 87.57 101.76 87.64 ;
    RECT 101.55 87.93 101.76 88.0 ;
    RECT 97.77 87.21 97.98 87.28 ;
    RECT 97.77 87.57 97.98 87.64 ;
    RECT 97.77 87.93 97.98 88.0 ;
    RECT 98.23 87.21 98.44 87.28 ;
    RECT 98.23 87.57 98.44 87.64 ;
    RECT 98.23 87.93 98.44 88.0 ;
    RECT 94.45 87.21 94.66 87.28 ;
    RECT 94.45 87.57 94.66 87.64 ;
    RECT 94.45 87.93 94.66 88.0 ;
    RECT 94.91 87.21 95.12 87.28 ;
    RECT 94.91 87.57 95.12 87.64 ;
    RECT 94.91 87.93 95.12 88.0 ;
    RECT 91.13 87.21 91.34 87.28 ;
    RECT 91.13 87.57 91.34 87.64 ;
    RECT 91.13 87.93 91.34 88.0 ;
    RECT 91.59 87.21 91.8 87.28 ;
    RECT 91.59 87.57 91.8 87.64 ;
    RECT 91.59 87.93 91.8 88.0 ;
    RECT 87.81 87.21 88.02 87.28 ;
    RECT 87.81 87.57 88.02 87.64 ;
    RECT 87.81 87.93 88.02 88.0 ;
    RECT 88.27 87.21 88.48 87.28 ;
    RECT 88.27 87.57 88.48 87.64 ;
    RECT 88.27 87.93 88.48 88.0 ;
    RECT 84.49 87.21 84.7 87.28 ;
    RECT 84.49 87.57 84.7 87.64 ;
    RECT 84.49 87.93 84.7 88.0 ;
    RECT 84.95 87.21 85.16 87.28 ;
    RECT 84.95 87.57 85.16 87.64 ;
    RECT 84.95 87.93 85.16 88.0 ;
    RECT 81.17 87.21 81.38 87.28 ;
    RECT 81.17 87.57 81.38 87.64 ;
    RECT 81.17 87.93 81.38 88.0 ;
    RECT 81.63 87.21 81.84 87.28 ;
    RECT 81.63 87.57 81.84 87.64 ;
    RECT 81.63 87.93 81.84 88.0 ;
    RECT 77.85 87.21 78.06 87.28 ;
    RECT 77.85 87.57 78.06 87.64 ;
    RECT 77.85 87.93 78.06 88.0 ;
    RECT 78.31 87.21 78.52 87.28 ;
    RECT 78.31 87.57 78.52 87.64 ;
    RECT 78.31 87.93 78.52 88.0 ;
    RECT 74.53 87.21 74.74 87.28 ;
    RECT 74.53 87.57 74.74 87.64 ;
    RECT 74.53 87.93 74.74 88.0 ;
    RECT 74.99 87.21 75.2 87.28 ;
    RECT 74.99 87.57 75.2 87.64 ;
    RECT 74.99 87.93 75.2 88.0 ;
    RECT 71.21 87.21 71.42 87.28 ;
    RECT 71.21 87.57 71.42 87.64 ;
    RECT 71.21 87.93 71.42 88.0 ;
    RECT 71.67 87.21 71.88 87.28 ;
    RECT 71.67 87.57 71.88 87.64 ;
    RECT 71.67 87.93 71.88 88.0 ;
    RECT 31.37 87.21 31.58 87.28 ;
    RECT 31.37 87.57 31.58 87.64 ;
    RECT 31.37 87.93 31.58 88.0 ;
    RECT 31.83 87.21 32.04 87.28 ;
    RECT 31.83 87.57 32.04 87.64 ;
    RECT 31.83 87.93 32.04 88.0 ;
    RECT 67.89 87.21 68.1 87.28 ;
    RECT 67.89 87.57 68.1 87.64 ;
    RECT 67.89 87.93 68.1 88.0 ;
    RECT 68.35 87.21 68.56 87.28 ;
    RECT 68.35 87.57 68.56 87.64 ;
    RECT 68.35 87.93 68.56 88.0 ;
    RECT 28.05 87.21 28.26 87.28 ;
    RECT 28.05 87.57 28.26 87.64 ;
    RECT 28.05 87.93 28.26 88.0 ;
    RECT 28.51 87.21 28.72 87.28 ;
    RECT 28.51 87.57 28.72 87.64 ;
    RECT 28.51 87.93 28.72 88.0 ;
    RECT 24.73 87.21 24.94 87.28 ;
    RECT 24.73 87.57 24.94 87.64 ;
    RECT 24.73 87.93 24.94 88.0 ;
    RECT 25.19 87.21 25.4 87.28 ;
    RECT 25.19 87.57 25.4 87.64 ;
    RECT 25.19 87.93 25.4 88.0 ;
    RECT 21.41 87.21 21.62 87.28 ;
    RECT 21.41 87.57 21.62 87.64 ;
    RECT 21.41 87.93 21.62 88.0 ;
    RECT 21.87 87.21 22.08 87.28 ;
    RECT 21.87 87.57 22.08 87.64 ;
    RECT 21.87 87.93 22.08 88.0 ;
    RECT 18.09 87.21 18.3 87.28 ;
    RECT 18.09 87.57 18.3 87.64 ;
    RECT 18.09 87.93 18.3 88.0 ;
    RECT 18.55 87.21 18.76 87.28 ;
    RECT 18.55 87.57 18.76 87.64 ;
    RECT 18.55 87.93 18.76 88.0 ;
    RECT 120.825 87.57 120.895 87.64 ;
    RECT 14.77 87.21 14.98 87.28 ;
    RECT 14.77 87.57 14.98 87.64 ;
    RECT 14.77 87.93 14.98 88.0 ;
    RECT 15.23 87.21 15.44 87.28 ;
    RECT 15.23 87.57 15.44 87.64 ;
    RECT 15.23 87.93 15.44 88.0 ;
    RECT 11.45 87.21 11.66 87.28 ;
    RECT 11.45 87.57 11.66 87.64 ;
    RECT 11.45 87.93 11.66 88.0 ;
    RECT 11.91 87.21 12.12 87.28 ;
    RECT 11.91 87.57 12.12 87.64 ;
    RECT 11.91 87.93 12.12 88.0 ;
    RECT 8.13 87.21 8.34 87.28 ;
    RECT 8.13 87.57 8.34 87.64 ;
    RECT 8.13 87.93 8.34 88.0 ;
    RECT 8.59 87.21 8.8 87.28 ;
    RECT 8.59 87.57 8.8 87.64 ;
    RECT 8.59 87.93 8.8 88.0 ;
    RECT 4.81 87.21 5.02 87.28 ;
    RECT 4.81 87.57 5.02 87.64 ;
    RECT 4.81 87.93 5.02 88.0 ;
    RECT 5.27 87.21 5.48 87.28 ;
    RECT 5.27 87.57 5.48 87.64 ;
    RECT 5.27 87.93 5.48 88.0 ;
    RECT 1.49 87.21 1.7 87.28 ;
    RECT 1.49 87.57 1.7 87.64 ;
    RECT 1.49 87.93 1.7 88.0 ;
    RECT 1.95 87.21 2.16 87.28 ;
    RECT 1.95 87.57 2.16 87.64 ;
    RECT 1.95 87.93 2.16 88.0 ;
    RECT 64.57 87.21 64.78 87.28 ;
    RECT 64.57 87.57 64.78 87.64 ;
    RECT 64.57 87.93 64.78 88.0 ;
    RECT 65.03 87.21 65.24 87.28 ;
    RECT 65.03 87.57 65.24 87.64 ;
    RECT 65.03 87.93 65.24 88.0 ;
    RECT 61.25 19.51 61.46 19.58 ;
    RECT 61.25 19.87 61.46 19.94 ;
    RECT 61.25 20.23 61.46 20.3 ;
    RECT 61.71 19.51 61.92 19.58 ;
    RECT 61.71 19.87 61.92 19.94 ;
    RECT 61.71 20.23 61.92 20.3 ;
    RECT 57.93 19.51 58.14 19.58 ;
    RECT 57.93 19.87 58.14 19.94 ;
    RECT 57.93 20.23 58.14 20.3 ;
    RECT 58.39 19.51 58.6 19.58 ;
    RECT 58.39 19.87 58.6 19.94 ;
    RECT 58.39 20.23 58.6 20.3 ;
    RECT 54.61 19.51 54.82 19.58 ;
    RECT 54.61 19.87 54.82 19.94 ;
    RECT 54.61 20.23 54.82 20.3 ;
    RECT 55.07 19.51 55.28 19.58 ;
    RECT 55.07 19.87 55.28 19.94 ;
    RECT 55.07 20.23 55.28 20.3 ;
    RECT 51.29 19.51 51.5 19.58 ;
    RECT 51.29 19.87 51.5 19.94 ;
    RECT 51.29 20.23 51.5 20.3 ;
    RECT 51.75 19.51 51.96 19.58 ;
    RECT 51.75 19.87 51.96 19.94 ;
    RECT 51.75 20.23 51.96 20.3 ;
    RECT 47.97 19.51 48.18 19.58 ;
    RECT 47.97 19.87 48.18 19.94 ;
    RECT 47.97 20.23 48.18 20.3 ;
    RECT 48.43 19.51 48.64 19.58 ;
    RECT 48.43 19.87 48.64 19.94 ;
    RECT 48.43 20.23 48.64 20.3 ;
    RECT 44.65 19.51 44.86 19.58 ;
    RECT 44.65 19.87 44.86 19.94 ;
    RECT 44.65 20.23 44.86 20.3 ;
    RECT 45.11 19.51 45.32 19.58 ;
    RECT 45.11 19.87 45.32 19.94 ;
    RECT 45.11 20.23 45.32 20.3 ;
    RECT 41.33 19.51 41.54 19.58 ;
    RECT 41.33 19.87 41.54 19.94 ;
    RECT 41.33 20.23 41.54 20.3 ;
    RECT 41.79 19.51 42.0 19.58 ;
    RECT 41.79 19.87 42.0 19.94 ;
    RECT 41.79 20.23 42.0 20.3 ;
    RECT 38.01 19.51 38.22 19.58 ;
    RECT 38.01 19.87 38.22 19.94 ;
    RECT 38.01 20.23 38.22 20.3 ;
    RECT 38.47 19.51 38.68 19.58 ;
    RECT 38.47 19.87 38.68 19.94 ;
    RECT 38.47 20.23 38.68 20.3 ;
    RECT 0.4 19.87 0.47 19.94 ;
    RECT 34.69 19.51 34.9 19.58 ;
    RECT 34.69 19.87 34.9 19.94 ;
    RECT 34.69 20.23 34.9 20.3 ;
    RECT 35.15 19.51 35.36 19.58 ;
    RECT 35.15 19.87 35.36 19.94 ;
    RECT 35.15 20.23 35.36 20.3 ;
    RECT 117.69 19.51 117.9 19.58 ;
    RECT 117.69 19.87 117.9 19.94 ;
    RECT 117.69 20.23 117.9 20.3 ;
    RECT 118.15 19.51 118.36 19.58 ;
    RECT 118.15 19.87 118.36 19.94 ;
    RECT 118.15 20.23 118.36 20.3 ;
    RECT 114.37 19.51 114.58 19.58 ;
    RECT 114.37 19.87 114.58 19.94 ;
    RECT 114.37 20.23 114.58 20.3 ;
    RECT 114.83 19.51 115.04 19.58 ;
    RECT 114.83 19.87 115.04 19.94 ;
    RECT 114.83 20.23 115.04 20.3 ;
    RECT 111.05 19.51 111.26 19.58 ;
    RECT 111.05 19.87 111.26 19.94 ;
    RECT 111.05 20.23 111.26 20.3 ;
    RECT 111.51 19.51 111.72 19.58 ;
    RECT 111.51 19.87 111.72 19.94 ;
    RECT 111.51 20.23 111.72 20.3 ;
    RECT 107.73 19.51 107.94 19.58 ;
    RECT 107.73 19.87 107.94 19.94 ;
    RECT 107.73 20.23 107.94 20.3 ;
    RECT 108.19 19.51 108.4 19.58 ;
    RECT 108.19 19.87 108.4 19.94 ;
    RECT 108.19 20.23 108.4 20.3 ;
    RECT 104.41 19.51 104.62 19.58 ;
    RECT 104.41 19.87 104.62 19.94 ;
    RECT 104.41 20.23 104.62 20.3 ;
    RECT 104.87 19.51 105.08 19.58 ;
    RECT 104.87 19.87 105.08 19.94 ;
    RECT 104.87 20.23 105.08 20.3 ;
    RECT 101.09 19.51 101.3 19.58 ;
    RECT 101.09 19.87 101.3 19.94 ;
    RECT 101.09 20.23 101.3 20.3 ;
    RECT 101.55 19.51 101.76 19.58 ;
    RECT 101.55 19.87 101.76 19.94 ;
    RECT 101.55 20.23 101.76 20.3 ;
    RECT 97.77 19.51 97.98 19.58 ;
    RECT 97.77 19.87 97.98 19.94 ;
    RECT 97.77 20.23 97.98 20.3 ;
    RECT 98.23 19.51 98.44 19.58 ;
    RECT 98.23 19.87 98.44 19.94 ;
    RECT 98.23 20.23 98.44 20.3 ;
    RECT 94.45 19.51 94.66 19.58 ;
    RECT 94.45 19.87 94.66 19.94 ;
    RECT 94.45 20.23 94.66 20.3 ;
    RECT 94.91 19.51 95.12 19.58 ;
    RECT 94.91 19.87 95.12 19.94 ;
    RECT 94.91 20.23 95.12 20.3 ;
    RECT 91.13 19.51 91.34 19.58 ;
    RECT 91.13 19.87 91.34 19.94 ;
    RECT 91.13 20.23 91.34 20.3 ;
    RECT 91.59 19.51 91.8 19.58 ;
    RECT 91.59 19.87 91.8 19.94 ;
    RECT 91.59 20.23 91.8 20.3 ;
    RECT 87.81 19.51 88.02 19.58 ;
    RECT 87.81 19.87 88.02 19.94 ;
    RECT 87.81 20.23 88.02 20.3 ;
    RECT 88.27 19.51 88.48 19.58 ;
    RECT 88.27 19.87 88.48 19.94 ;
    RECT 88.27 20.23 88.48 20.3 ;
    RECT 84.49 19.51 84.7 19.58 ;
    RECT 84.49 19.87 84.7 19.94 ;
    RECT 84.49 20.23 84.7 20.3 ;
    RECT 84.95 19.51 85.16 19.58 ;
    RECT 84.95 19.87 85.16 19.94 ;
    RECT 84.95 20.23 85.16 20.3 ;
    RECT 81.17 19.51 81.38 19.58 ;
    RECT 81.17 19.87 81.38 19.94 ;
    RECT 81.17 20.23 81.38 20.3 ;
    RECT 81.63 19.51 81.84 19.58 ;
    RECT 81.63 19.87 81.84 19.94 ;
    RECT 81.63 20.23 81.84 20.3 ;
    RECT 77.85 19.51 78.06 19.58 ;
    RECT 77.85 19.87 78.06 19.94 ;
    RECT 77.85 20.23 78.06 20.3 ;
    RECT 78.31 19.51 78.52 19.58 ;
    RECT 78.31 19.87 78.52 19.94 ;
    RECT 78.31 20.23 78.52 20.3 ;
    RECT 74.53 19.51 74.74 19.58 ;
    RECT 74.53 19.87 74.74 19.94 ;
    RECT 74.53 20.23 74.74 20.3 ;
    RECT 74.99 19.51 75.2 19.58 ;
    RECT 74.99 19.87 75.2 19.94 ;
    RECT 74.99 20.23 75.2 20.3 ;
    RECT 71.21 19.51 71.42 19.58 ;
    RECT 71.21 19.87 71.42 19.94 ;
    RECT 71.21 20.23 71.42 20.3 ;
    RECT 71.67 19.51 71.88 19.58 ;
    RECT 71.67 19.87 71.88 19.94 ;
    RECT 71.67 20.23 71.88 20.3 ;
    RECT 31.37 19.51 31.58 19.58 ;
    RECT 31.37 19.87 31.58 19.94 ;
    RECT 31.37 20.23 31.58 20.3 ;
    RECT 31.83 19.51 32.04 19.58 ;
    RECT 31.83 19.87 32.04 19.94 ;
    RECT 31.83 20.23 32.04 20.3 ;
    RECT 67.89 19.51 68.1 19.58 ;
    RECT 67.89 19.87 68.1 19.94 ;
    RECT 67.89 20.23 68.1 20.3 ;
    RECT 68.35 19.51 68.56 19.58 ;
    RECT 68.35 19.87 68.56 19.94 ;
    RECT 68.35 20.23 68.56 20.3 ;
    RECT 28.05 19.51 28.26 19.58 ;
    RECT 28.05 19.87 28.26 19.94 ;
    RECT 28.05 20.23 28.26 20.3 ;
    RECT 28.51 19.51 28.72 19.58 ;
    RECT 28.51 19.87 28.72 19.94 ;
    RECT 28.51 20.23 28.72 20.3 ;
    RECT 24.73 19.51 24.94 19.58 ;
    RECT 24.73 19.87 24.94 19.94 ;
    RECT 24.73 20.23 24.94 20.3 ;
    RECT 25.19 19.51 25.4 19.58 ;
    RECT 25.19 19.87 25.4 19.94 ;
    RECT 25.19 20.23 25.4 20.3 ;
    RECT 21.41 19.51 21.62 19.58 ;
    RECT 21.41 19.87 21.62 19.94 ;
    RECT 21.41 20.23 21.62 20.3 ;
    RECT 21.87 19.51 22.08 19.58 ;
    RECT 21.87 19.87 22.08 19.94 ;
    RECT 21.87 20.23 22.08 20.3 ;
    RECT 18.09 19.51 18.3 19.58 ;
    RECT 18.09 19.87 18.3 19.94 ;
    RECT 18.09 20.23 18.3 20.3 ;
    RECT 18.55 19.51 18.76 19.58 ;
    RECT 18.55 19.87 18.76 19.94 ;
    RECT 18.55 20.23 18.76 20.3 ;
    RECT 120.825 19.87 120.895 19.94 ;
    RECT 14.77 19.51 14.98 19.58 ;
    RECT 14.77 19.87 14.98 19.94 ;
    RECT 14.77 20.23 14.98 20.3 ;
    RECT 15.23 19.51 15.44 19.58 ;
    RECT 15.23 19.87 15.44 19.94 ;
    RECT 15.23 20.23 15.44 20.3 ;
    RECT 11.45 19.51 11.66 19.58 ;
    RECT 11.45 19.87 11.66 19.94 ;
    RECT 11.45 20.23 11.66 20.3 ;
    RECT 11.91 19.51 12.12 19.58 ;
    RECT 11.91 19.87 12.12 19.94 ;
    RECT 11.91 20.23 12.12 20.3 ;
    RECT 8.13 19.51 8.34 19.58 ;
    RECT 8.13 19.87 8.34 19.94 ;
    RECT 8.13 20.23 8.34 20.3 ;
    RECT 8.59 19.51 8.8 19.58 ;
    RECT 8.59 19.87 8.8 19.94 ;
    RECT 8.59 20.23 8.8 20.3 ;
    RECT 4.81 19.51 5.02 19.58 ;
    RECT 4.81 19.87 5.02 19.94 ;
    RECT 4.81 20.23 5.02 20.3 ;
    RECT 5.27 19.51 5.48 19.58 ;
    RECT 5.27 19.87 5.48 19.94 ;
    RECT 5.27 20.23 5.48 20.3 ;
    RECT 1.49 19.51 1.7 19.58 ;
    RECT 1.49 19.87 1.7 19.94 ;
    RECT 1.49 20.23 1.7 20.3 ;
    RECT 1.95 19.51 2.16 19.58 ;
    RECT 1.95 19.87 2.16 19.94 ;
    RECT 1.95 20.23 2.16 20.3 ;
    RECT 64.57 19.51 64.78 19.58 ;
    RECT 64.57 19.87 64.78 19.94 ;
    RECT 64.57 20.23 64.78 20.3 ;
    RECT 65.03 19.51 65.24 19.58 ;
    RECT 65.03 19.87 65.24 19.94 ;
    RECT 65.03 20.23 65.24 20.3 ;
    RECT 61.25 18.79 61.46 18.86 ;
    RECT 61.25 19.15 61.46 19.22 ;
    RECT 61.25 19.51 61.46 19.58 ;
    RECT 61.71 18.79 61.92 18.86 ;
    RECT 61.71 19.15 61.92 19.22 ;
    RECT 61.71 19.51 61.92 19.58 ;
    RECT 57.93 18.79 58.14 18.86 ;
    RECT 57.93 19.15 58.14 19.22 ;
    RECT 57.93 19.51 58.14 19.58 ;
    RECT 58.39 18.79 58.6 18.86 ;
    RECT 58.39 19.15 58.6 19.22 ;
    RECT 58.39 19.51 58.6 19.58 ;
    RECT 54.61 18.79 54.82 18.86 ;
    RECT 54.61 19.15 54.82 19.22 ;
    RECT 54.61 19.51 54.82 19.58 ;
    RECT 55.07 18.79 55.28 18.86 ;
    RECT 55.07 19.15 55.28 19.22 ;
    RECT 55.07 19.51 55.28 19.58 ;
    RECT 51.29 18.79 51.5 18.86 ;
    RECT 51.29 19.15 51.5 19.22 ;
    RECT 51.29 19.51 51.5 19.58 ;
    RECT 51.75 18.79 51.96 18.86 ;
    RECT 51.75 19.15 51.96 19.22 ;
    RECT 51.75 19.51 51.96 19.58 ;
    RECT 47.97 18.79 48.18 18.86 ;
    RECT 47.97 19.15 48.18 19.22 ;
    RECT 47.97 19.51 48.18 19.58 ;
    RECT 48.43 18.79 48.64 18.86 ;
    RECT 48.43 19.15 48.64 19.22 ;
    RECT 48.43 19.51 48.64 19.58 ;
    RECT 44.65 18.79 44.86 18.86 ;
    RECT 44.65 19.15 44.86 19.22 ;
    RECT 44.65 19.51 44.86 19.58 ;
    RECT 45.11 18.79 45.32 18.86 ;
    RECT 45.11 19.15 45.32 19.22 ;
    RECT 45.11 19.51 45.32 19.58 ;
    RECT 41.33 18.79 41.54 18.86 ;
    RECT 41.33 19.15 41.54 19.22 ;
    RECT 41.33 19.51 41.54 19.58 ;
    RECT 41.79 18.79 42.0 18.86 ;
    RECT 41.79 19.15 42.0 19.22 ;
    RECT 41.79 19.51 42.0 19.58 ;
    RECT 38.01 18.79 38.22 18.86 ;
    RECT 38.01 19.15 38.22 19.22 ;
    RECT 38.01 19.51 38.22 19.58 ;
    RECT 38.47 18.79 38.68 18.86 ;
    RECT 38.47 19.15 38.68 19.22 ;
    RECT 38.47 19.51 38.68 19.58 ;
    RECT 0.4 19.15 0.47 19.22 ;
    RECT 34.69 18.79 34.9 18.86 ;
    RECT 34.69 19.15 34.9 19.22 ;
    RECT 34.69 19.51 34.9 19.58 ;
    RECT 35.15 18.79 35.36 18.86 ;
    RECT 35.15 19.15 35.36 19.22 ;
    RECT 35.15 19.51 35.36 19.58 ;
    RECT 117.69 18.79 117.9 18.86 ;
    RECT 117.69 19.15 117.9 19.22 ;
    RECT 117.69 19.51 117.9 19.58 ;
    RECT 118.15 18.79 118.36 18.86 ;
    RECT 118.15 19.15 118.36 19.22 ;
    RECT 118.15 19.51 118.36 19.58 ;
    RECT 114.37 18.79 114.58 18.86 ;
    RECT 114.37 19.15 114.58 19.22 ;
    RECT 114.37 19.51 114.58 19.58 ;
    RECT 114.83 18.79 115.04 18.86 ;
    RECT 114.83 19.15 115.04 19.22 ;
    RECT 114.83 19.51 115.04 19.58 ;
    RECT 111.05 18.79 111.26 18.86 ;
    RECT 111.05 19.15 111.26 19.22 ;
    RECT 111.05 19.51 111.26 19.58 ;
    RECT 111.51 18.79 111.72 18.86 ;
    RECT 111.51 19.15 111.72 19.22 ;
    RECT 111.51 19.51 111.72 19.58 ;
    RECT 107.73 18.79 107.94 18.86 ;
    RECT 107.73 19.15 107.94 19.22 ;
    RECT 107.73 19.51 107.94 19.58 ;
    RECT 108.19 18.79 108.4 18.86 ;
    RECT 108.19 19.15 108.4 19.22 ;
    RECT 108.19 19.51 108.4 19.58 ;
    RECT 104.41 18.79 104.62 18.86 ;
    RECT 104.41 19.15 104.62 19.22 ;
    RECT 104.41 19.51 104.62 19.58 ;
    RECT 104.87 18.79 105.08 18.86 ;
    RECT 104.87 19.15 105.08 19.22 ;
    RECT 104.87 19.51 105.08 19.58 ;
    RECT 101.09 18.79 101.3 18.86 ;
    RECT 101.09 19.15 101.3 19.22 ;
    RECT 101.09 19.51 101.3 19.58 ;
    RECT 101.55 18.79 101.76 18.86 ;
    RECT 101.55 19.15 101.76 19.22 ;
    RECT 101.55 19.51 101.76 19.58 ;
    RECT 97.77 18.79 97.98 18.86 ;
    RECT 97.77 19.15 97.98 19.22 ;
    RECT 97.77 19.51 97.98 19.58 ;
    RECT 98.23 18.79 98.44 18.86 ;
    RECT 98.23 19.15 98.44 19.22 ;
    RECT 98.23 19.51 98.44 19.58 ;
    RECT 94.45 18.79 94.66 18.86 ;
    RECT 94.45 19.15 94.66 19.22 ;
    RECT 94.45 19.51 94.66 19.58 ;
    RECT 94.91 18.79 95.12 18.86 ;
    RECT 94.91 19.15 95.12 19.22 ;
    RECT 94.91 19.51 95.12 19.58 ;
    RECT 91.13 18.79 91.34 18.86 ;
    RECT 91.13 19.15 91.34 19.22 ;
    RECT 91.13 19.51 91.34 19.58 ;
    RECT 91.59 18.79 91.8 18.86 ;
    RECT 91.59 19.15 91.8 19.22 ;
    RECT 91.59 19.51 91.8 19.58 ;
    RECT 87.81 18.79 88.02 18.86 ;
    RECT 87.81 19.15 88.02 19.22 ;
    RECT 87.81 19.51 88.02 19.58 ;
    RECT 88.27 18.79 88.48 18.86 ;
    RECT 88.27 19.15 88.48 19.22 ;
    RECT 88.27 19.51 88.48 19.58 ;
    RECT 84.49 18.79 84.7 18.86 ;
    RECT 84.49 19.15 84.7 19.22 ;
    RECT 84.49 19.51 84.7 19.58 ;
    RECT 84.95 18.79 85.16 18.86 ;
    RECT 84.95 19.15 85.16 19.22 ;
    RECT 84.95 19.51 85.16 19.58 ;
    RECT 81.17 18.79 81.38 18.86 ;
    RECT 81.17 19.15 81.38 19.22 ;
    RECT 81.17 19.51 81.38 19.58 ;
    RECT 81.63 18.79 81.84 18.86 ;
    RECT 81.63 19.15 81.84 19.22 ;
    RECT 81.63 19.51 81.84 19.58 ;
    RECT 77.85 18.79 78.06 18.86 ;
    RECT 77.85 19.15 78.06 19.22 ;
    RECT 77.85 19.51 78.06 19.58 ;
    RECT 78.31 18.79 78.52 18.86 ;
    RECT 78.31 19.15 78.52 19.22 ;
    RECT 78.31 19.51 78.52 19.58 ;
    RECT 74.53 18.79 74.74 18.86 ;
    RECT 74.53 19.15 74.74 19.22 ;
    RECT 74.53 19.51 74.74 19.58 ;
    RECT 74.99 18.79 75.2 18.86 ;
    RECT 74.99 19.15 75.2 19.22 ;
    RECT 74.99 19.51 75.2 19.58 ;
    RECT 71.21 18.79 71.42 18.86 ;
    RECT 71.21 19.15 71.42 19.22 ;
    RECT 71.21 19.51 71.42 19.58 ;
    RECT 71.67 18.79 71.88 18.86 ;
    RECT 71.67 19.15 71.88 19.22 ;
    RECT 71.67 19.51 71.88 19.58 ;
    RECT 31.37 18.79 31.58 18.86 ;
    RECT 31.37 19.15 31.58 19.22 ;
    RECT 31.37 19.51 31.58 19.58 ;
    RECT 31.83 18.79 32.04 18.86 ;
    RECT 31.83 19.15 32.04 19.22 ;
    RECT 31.83 19.51 32.04 19.58 ;
    RECT 67.89 18.79 68.1 18.86 ;
    RECT 67.89 19.15 68.1 19.22 ;
    RECT 67.89 19.51 68.1 19.58 ;
    RECT 68.35 18.79 68.56 18.86 ;
    RECT 68.35 19.15 68.56 19.22 ;
    RECT 68.35 19.51 68.56 19.58 ;
    RECT 28.05 18.79 28.26 18.86 ;
    RECT 28.05 19.15 28.26 19.22 ;
    RECT 28.05 19.51 28.26 19.58 ;
    RECT 28.51 18.79 28.72 18.86 ;
    RECT 28.51 19.15 28.72 19.22 ;
    RECT 28.51 19.51 28.72 19.58 ;
    RECT 24.73 18.79 24.94 18.86 ;
    RECT 24.73 19.15 24.94 19.22 ;
    RECT 24.73 19.51 24.94 19.58 ;
    RECT 25.19 18.79 25.4 18.86 ;
    RECT 25.19 19.15 25.4 19.22 ;
    RECT 25.19 19.51 25.4 19.58 ;
    RECT 21.41 18.79 21.62 18.86 ;
    RECT 21.41 19.15 21.62 19.22 ;
    RECT 21.41 19.51 21.62 19.58 ;
    RECT 21.87 18.79 22.08 18.86 ;
    RECT 21.87 19.15 22.08 19.22 ;
    RECT 21.87 19.51 22.08 19.58 ;
    RECT 18.09 18.79 18.3 18.86 ;
    RECT 18.09 19.15 18.3 19.22 ;
    RECT 18.09 19.51 18.3 19.58 ;
    RECT 18.55 18.79 18.76 18.86 ;
    RECT 18.55 19.15 18.76 19.22 ;
    RECT 18.55 19.51 18.76 19.58 ;
    RECT 120.825 19.15 120.895 19.22 ;
    RECT 14.77 18.79 14.98 18.86 ;
    RECT 14.77 19.15 14.98 19.22 ;
    RECT 14.77 19.51 14.98 19.58 ;
    RECT 15.23 18.79 15.44 18.86 ;
    RECT 15.23 19.15 15.44 19.22 ;
    RECT 15.23 19.51 15.44 19.58 ;
    RECT 11.45 18.79 11.66 18.86 ;
    RECT 11.45 19.15 11.66 19.22 ;
    RECT 11.45 19.51 11.66 19.58 ;
    RECT 11.91 18.79 12.12 18.86 ;
    RECT 11.91 19.15 12.12 19.22 ;
    RECT 11.91 19.51 12.12 19.58 ;
    RECT 8.13 18.79 8.34 18.86 ;
    RECT 8.13 19.15 8.34 19.22 ;
    RECT 8.13 19.51 8.34 19.58 ;
    RECT 8.59 18.79 8.8 18.86 ;
    RECT 8.59 19.15 8.8 19.22 ;
    RECT 8.59 19.51 8.8 19.58 ;
    RECT 4.81 18.79 5.02 18.86 ;
    RECT 4.81 19.15 5.02 19.22 ;
    RECT 4.81 19.51 5.02 19.58 ;
    RECT 5.27 18.79 5.48 18.86 ;
    RECT 5.27 19.15 5.48 19.22 ;
    RECT 5.27 19.51 5.48 19.58 ;
    RECT 1.49 18.79 1.7 18.86 ;
    RECT 1.49 19.15 1.7 19.22 ;
    RECT 1.49 19.51 1.7 19.58 ;
    RECT 1.95 18.79 2.16 18.86 ;
    RECT 1.95 19.15 2.16 19.22 ;
    RECT 1.95 19.51 2.16 19.58 ;
    RECT 64.57 18.79 64.78 18.86 ;
    RECT 64.57 19.15 64.78 19.22 ;
    RECT 64.57 19.51 64.78 19.58 ;
    RECT 65.03 18.79 65.24 18.86 ;
    RECT 65.03 19.15 65.24 19.22 ;
    RECT 65.03 19.51 65.24 19.58 ;
    RECT 61.25 49.75 61.46 49.82 ;
    RECT 61.25 50.11 61.46 50.18 ;
    RECT 61.25 50.47 61.46 50.54 ;
    RECT 61.71 49.75 61.92 49.82 ;
    RECT 61.71 50.11 61.92 50.18 ;
    RECT 61.71 50.47 61.92 50.54 ;
    RECT 57.93 49.75 58.14 49.82 ;
    RECT 57.93 50.11 58.14 50.18 ;
    RECT 57.93 50.47 58.14 50.54 ;
    RECT 58.39 49.75 58.6 49.82 ;
    RECT 58.39 50.11 58.6 50.18 ;
    RECT 58.39 50.47 58.6 50.54 ;
    RECT 54.61 49.75 54.82 49.82 ;
    RECT 54.61 50.11 54.82 50.18 ;
    RECT 54.61 50.47 54.82 50.54 ;
    RECT 55.07 49.75 55.28 49.82 ;
    RECT 55.07 50.11 55.28 50.18 ;
    RECT 55.07 50.47 55.28 50.54 ;
    RECT 51.29 49.75 51.5 49.82 ;
    RECT 51.29 50.11 51.5 50.18 ;
    RECT 51.29 50.47 51.5 50.54 ;
    RECT 51.75 49.75 51.96 49.82 ;
    RECT 51.75 50.11 51.96 50.18 ;
    RECT 51.75 50.47 51.96 50.54 ;
    RECT 47.97 49.75 48.18 49.82 ;
    RECT 47.97 50.11 48.18 50.18 ;
    RECT 47.97 50.47 48.18 50.54 ;
    RECT 48.43 49.75 48.64 49.82 ;
    RECT 48.43 50.11 48.64 50.18 ;
    RECT 48.43 50.47 48.64 50.54 ;
    RECT 44.65 49.75 44.86 49.82 ;
    RECT 44.65 50.11 44.86 50.18 ;
    RECT 44.65 50.47 44.86 50.54 ;
    RECT 45.11 49.75 45.32 49.82 ;
    RECT 45.11 50.11 45.32 50.18 ;
    RECT 45.11 50.47 45.32 50.54 ;
    RECT 41.33 49.75 41.54 49.82 ;
    RECT 41.33 50.11 41.54 50.18 ;
    RECT 41.33 50.47 41.54 50.54 ;
    RECT 41.79 49.75 42.0 49.82 ;
    RECT 41.79 50.11 42.0 50.18 ;
    RECT 41.79 50.47 42.0 50.54 ;
    RECT 38.01 49.75 38.22 49.82 ;
    RECT 38.01 50.11 38.22 50.18 ;
    RECT 38.01 50.47 38.22 50.54 ;
    RECT 38.47 49.75 38.68 49.82 ;
    RECT 38.47 50.11 38.68 50.18 ;
    RECT 38.47 50.47 38.68 50.54 ;
    RECT 0.4 50.11 0.47 50.18 ;
    RECT 34.69 49.75 34.9 49.82 ;
    RECT 34.69 50.11 34.9 50.18 ;
    RECT 34.69 50.47 34.9 50.54 ;
    RECT 35.15 49.75 35.36 49.82 ;
    RECT 35.15 50.11 35.36 50.18 ;
    RECT 35.15 50.47 35.36 50.54 ;
    RECT 117.69 49.75 117.9 49.82 ;
    RECT 117.69 50.11 117.9 50.18 ;
    RECT 117.69 50.47 117.9 50.54 ;
    RECT 118.15 49.75 118.36 49.82 ;
    RECT 118.15 50.11 118.36 50.18 ;
    RECT 118.15 50.47 118.36 50.54 ;
    RECT 114.37 49.75 114.58 49.82 ;
    RECT 114.37 50.11 114.58 50.18 ;
    RECT 114.37 50.47 114.58 50.54 ;
    RECT 114.83 49.75 115.04 49.82 ;
    RECT 114.83 50.11 115.04 50.18 ;
    RECT 114.83 50.47 115.04 50.54 ;
    RECT 111.05 49.75 111.26 49.82 ;
    RECT 111.05 50.11 111.26 50.18 ;
    RECT 111.05 50.47 111.26 50.54 ;
    RECT 111.51 49.75 111.72 49.82 ;
    RECT 111.51 50.11 111.72 50.18 ;
    RECT 111.51 50.47 111.72 50.54 ;
    RECT 107.73 49.75 107.94 49.82 ;
    RECT 107.73 50.11 107.94 50.18 ;
    RECT 107.73 50.47 107.94 50.54 ;
    RECT 108.19 49.75 108.4 49.82 ;
    RECT 108.19 50.11 108.4 50.18 ;
    RECT 108.19 50.47 108.4 50.54 ;
    RECT 104.41 49.75 104.62 49.82 ;
    RECT 104.41 50.11 104.62 50.18 ;
    RECT 104.41 50.47 104.62 50.54 ;
    RECT 104.87 49.75 105.08 49.82 ;
    RECT 104.87 50.11 105.08 50.18 ;
    RECT 104.87 50.47 105.08 50.54 ;
    RECT 101.09 49.75 101.3 49.82 ;
    RECT 101.09 50.11 101.3 50.18 ;
    RECT 101.09 50.47 101.3 50.54 ;
    RECT 101.55 49.75 101.76 49.82 ;
    RECT 101.55 50.11 101.76 50.18 ;
    RECT 101.55 50.47 101.76 50.54 ;
    RECT 97.77 49.75 97.98 49.82 ;
    RECT 97.77 50.11 97.98 50.18 ;
    RECT 97.77 50.47 97.98 50.54 ;
    RECT 98.23 49.75 98.44 49.82 ;
    RECT 98.23 50.11 98.44 50.18 ;
    RECT 98.23 50.47 98.44 50.54 ;
    RECT 94.45 49.75 94.66 49.82 ;
    RECT 94.45 50.11 94.66 50.18 ;
    RECT 94.45 50.47 94.66 50.54 ;
    RECT 94.91 49.75 95.12 49.82 ;
    RECT 94.91 50.11 95.12 50.18 ;
    RECT 94.91 50.47 95.12 50.54 ;
    RECT 91.13 49.75 91.34 49.82 ;
    RECT 91.13 50.11 91.34 50.18 ;
    RECT 91.13 50.47 91.34 50.54 ;
    RECT 91.59 49.75 91.8 49.82 ;
    RECT 91.59 50.11 91.8 50.18 ;
    RECT 91.59 50.47 91.8 50.54 ;
    RECT 87.81 49.75 88.02 49.82 ;
    RECT 87.81 50.11 88.02 50.18 ;
    RECT 87.81 50.47 88.02 50.54 ;
    RECT 88.27 49.75 88.48 49.82 ;
    RECT 88.27 50.11 88.48 50.18 ;
    RECT 88.27 50.47 88.48 50.54 ;
    RECT 84.49 49.75 84.7 49.82 ;
    RECT 84.49 50.11 84.7 50.18 ;
    RECT 84.49 50.47 84.7 50.54 ;
    RECT 84.95 49.75 85.16 49.82 ;
    RECT 84.95 50.11 85.16 50.18 ;
    RECT 84.95 50.47 85.16 50.54 ;
    RECT 81.17 49.75 81.38 49.82 ;
    RECT 81.17 50.11 81.38 50.18 ;
    RECT 81.17 50.47 81.38 50.54 ;
    RECT 81.63 49.75 81.84 49.82 ;
    RECT 81.63 50.11 81.84 50.18 ;
    RECT 81.63 50.47 81.84 50.54 ;
    RECT 77.85 49.75 78.06 49.82 ;
    RECT 77.85 50.11 78.06 50.18 ;
    RECT 77.85 50.47 78.06 50.54 ;
    RECT 78.31 49.75 78.52 49.82 ;
    RECT 78.31 50.11 78.52 50.18 ;
    RECT 78.31 50.47 78.52 50.54 ;
    RECT 74.53 49.75 74.74 49.82 ;
    RECT 74.53 50.11 74.74 50.18 ;
    RECT 74.53 50.47 74.74 50.54 ;
    RECT 74.99 49.75 75.2 49.82 ;
    RECT 74.99 50.11 75.2 50.18 ;
    RECT 74.99 50.47 75.2 50.54 ;
    RECT 71.21 49.75 71.42 49.82 ;
    RECT 71.21 50.11 71.42 50.18 ;
    RECT 71.21 50.47 71.42 50.54 ;
    RECT 71.67 49.75 71.88 49.82 ;
    RECT 71.67 50.11 71.88 50.18 ;
    RECT 71.67 50.47 71.88 50.54 ;
    RECT 31.37 49.75 31.58 49.82 ;
    RECT 31.37 50.11 31.58 50.18 ;
    RECT 31.37 50.47 31.58 50.54 ;
    RECT 31.83 49.75 32.04 49.82 ;
    RECT 31.83 50.11 32.04 50.18 ;
    RECT 31.83 50.47 32.04 50.54 ;
    RECT 67.89 49.75 68.1 49.82 ;
    RECT 67.89 50.11 68.1 50.18 ;
    RECT 67.89 50.47 68.1 50.54 ;
    RECT 68.35 49.75 68.56 49.82 ;
    RECT 68.35 50.11 68.56 50.18 ;
    RECT 68.35 50.47 68.56 50.54 ;
    RECT 28.05 49.75 28.26 49.82 ;
    RECT 28.05 50.11 28.26 50.18 ;
    RECT 28.05 50.47 28.26 50.54 ;
    RECT 28.51 49.75 28.72 49.82 ;
    RECT 28.51 50.11 28.72 50.18 ;
    RECT 28.51 50.47 28.72 50.54 ;
    RECT 24.73 49.75 24.94 49.82 ;
    RECT 24.73 50.11 24.94 50.18 ;
    RECT 24.73 50.47 24.94 50.54 ;
    RECT 25.19 49.75 25.4 49.82 ;
    RECT 25.19 50.11 25.4 50.18 ;
    RECT 25.19 50.47 25.4 50.54 ;
    RECT 21.41 49.75 21.62 49.82 ;
    RECT 21.41 50.11 21.62 50.18 ;
    RECT 21.41 50.47 21.62 50.54 ;
    RECT 21.87 49.75 22.08 49.82 ;
    RECT 21.87 50.11 22.08 50.18 ;
    RECT 21.87 50.47 22.08 50.54 ;
    RECT 18.09 49.75 18.3 49.82 ;
    RECT 18.09 50.11 18.3 50.18 ;
    RECT 18.09 50.47 18.3 50.54 ;
    RECT 18.55 49.75 18.76 49.82 ;
    RECT 18.55 50.11 18.76 50.18 ;
    RECT 18.55 50.47 18.76 50.54 ;
    RECT 120.825 50.11 120.895 50.18 ;
    RECT 14.77 49.75 14.98 49.82 ;
    RECT 14.77 50.11 14.98 50.18 ;
    RECT 14.77 50.47 14.98 50.54 ;
    RECT 15.23 49.75 15.44 49.82 ;
    RECT 15.23 50.11 15.44 50.18 ;
    RECT 15.23 50.47 15.44 50.54 ;
    RECT 11.45 49.75 11.66 49.82 ;
    RECT 11.45 50.11 11.66 50.18 ;
    RECT 11.45 50.47 11.66 50.54 ;
    RECT 11.91 49.75 12.12 49.82 ;
    RECT 11.91 50.11 12.12 50.18 ;
    RECT 11.91 50.47 12.12 50.54 ;
    RECT 8.13 49.75 8.34 49.82 ;
    RECT 8.13 50.11 8.34 50.18 ;
    RECT 8.13 50.47 8.34 50.54 ;
    RECT 8.59 49.75 8.8 49.82 ;
    RECT 8.59 50.11 8.8 50.18 ;
    RECT 8.59 50.47 8.8 50.54 ;
    RECT 4.81 49.75 5.02 49.82 ;
    RECT 4.81 50.11 5.02 50.18 ;
    RECT 4.81 50.47 5.02 50.54 ;
    RECT 5.27 49.75 5.48 49.82 ;
    RECT 5.27 50.11 5.48 50.18 ;
    RECT 5.27 50.47 5.48 50.54 ;
    RECT 1.49 49.75 1.7 49.82 ;
    RECT 1.49 50.11 1.7 50.18 ;
    RECT 1.49 50.47 1.7 50.54 ;
    RECT 1.95 49.75 2.16 49.82 ;
    RECT 1.95 50.11 2.16 50.18 ;
    RECT 1.95 50.47 2.16 50.54 ;
    RECT 64.57 49.75 64.78 49.82 ;
    RECT 64.57 50.11 64.78 50.18 ;
    RECT 64.57 50.47 64.78 50.54 ;
    RECT 65.03 49.75 65.24 49.82 ;
    RECT 65.03 50.11 65.24 50.18 ;
    RECT 65.03 50.47 65.24 50.54 ;
    RECT 61.25 18.07 61.46 18.14 ;
    RECT 61.25 18.43 61.46 18.5 ;
    RECT 61.25 18.79 61.46 18.86 ;
    RECT 61.71 18.07 61.92 18.14 ;
    RECT 61.71 18.43 61.92 18.5 ;
    RECT 61.71 18.79 61.92 18.86 ;
    RECT 57.93 18.07 58.14 18.14 ;
    RECT 57.93 18.43 58.14 18.5 ;
    RECT 57.93 18.79 58.14 18.86 ;
    RECT 58.39 18.07 58.6 18.14 ;
    RECT 58.39 18.43 58.6 18.5 ;
    RECT 58.39 18.79 58.6 18.86 ;
    RECT 54.61 18.07 54.82 18.14 ;
    RECT 54.61 18.43 54.82 18.5 ;
    RECT 54.61 18.79 54.82 18.86 ;
    RECT 55.07 18.07 55.28 18.14 ;
    RECT 55.07 18.43 55.28 18.5 ;
    RECT 55.07 18.79 55.28 18.86 ;
    RECT 51.29 18.07 51.5 18.14 ;
    RECT 51.29 18.43 51.5 18.5 ;
    RECT 51.29 18.79 51.5 18.86 ;
    RECT 51.75 18.07 51.96 18.14 ;
    RECT 51.75 18.43 51.96 18.5 ;
    RECT 51.75 18.79 51.96 18.86 ;
    RECT 47.97 18.07 48.18 18.14 ;
    RECT 47.97 18.43 48.18 18.5 ;
    RECT 47.97 18.79 48.18 18.86 ;
    RECT 48.43 18.07 48.64 18.14 ;
    RECT 48.43 18.43 48.64 18.5 ;
    RECT 48.43 18.79 48.64 18.86 ;
    RECT 44.65 18.07 44.86 18.14 ;
    RECT 44.65 18.43 44.86 18.5 ;
    RECT 44.65 18.79 44.86 18.86 ;
    RECT 45.11 18.07 45.32 18.14 ;
    RECT 45.11 18.43 45.32 18.5 ;
    RECT 45.11 18.79 45.32 18.86 ;
    RECT 41.33 18.07 41.54 18.14 ;
    RECT 41.33 18.43 41.54 18.5 ;
    RECT 41.33 18.79 41.54 18.86 ;
    RECT 41.79 18.07 42.0 18.14 ;
    RECT 41.79 18.43 42.0 18.5 ;
    RECT 41.79 18.79 42.0 18.86 ;
    RECT 38.01 18.07 38.22 18.14 ;
    RECT 38.01 18.43 38.22 18.5 ;
    RECT 38.01 18.79 38.22 18.86 ;
    RECT 38.47 18.07 38.68 18.14 ;
    RECT 38.47 18.43 38.68 18.5 ;
    RECT 38.47 18.79 38.68 18.86 ;
    RECT 0.4 18.43 0.47 18.5 ;
    RECT 34.69 18.07 34.9 18.14 ;
    RECT 34.69 18.43 34.9 18.5 ;
    RECT 34.69 18.79 34.9 18.86 ;
    RECT 35.15 18.07 35.36 18.14 ;
    RECT 35.15 18.43 35.36 18.5 ;
    RECT 35.15 18.79 35.36 18.86 ;
    RECT 117.69 18.07 117.9 18.14 ;
    RECT 117.69 18.43 117.9 18.5 ;
    RECT 117.69 18.79 117.9 18.86 ;
    RECT 118.15 18.07 118.36 18.14 ;
    RECT 118.15 18.43 118.36 18.5 ;
    RECT 118.15 18.79 118.36 18.86 ;
    RECT 114.37 18.07 114.58 18.14 ;
    RECT 114.37 18.43 114.58 18.5 ;
    RECT 114.37 18.79 114.58 18.86 ;
    RECT 114.83 18.07 115.04 18.14 ;
    RECT 114.83 18.43 115.04 18.5 ;
    RECT 114.83 18.79 115.04 18.86 ;
    RECT 111.05 18.07 111.26 18.14 ;
    RECT 111.05 18.43 111.26 18.5 ;
    RECT 111.05 18.79 111.26 18.86 ;
    RECT 111.51 18.07 111.72 18.14 ;
    RECT 111.51 18.43 111.72 18.5 ;
    RECT 111.51 18.79 111.72 18.86 ;
    RECT 107.73 18.07 107.94 18.14 ;
    RECT 107.73 18.43 107.94 18.5 ;
    RECT 107.73 18.79 107.94 18.86 ;
    RECT 108.19 18.07 108.4 18.14 ;
    RECT 108.19 18.43 108.4 18.5 ;
    RECT 108.19 18.79 108.4 18.86 ;
    RECT 104.41 18.07 104.62 18.14 ;
    RECT 104.41 18.43 104.62 18.5 ;
    RECT 104.41 18.79 104.62 18.86 ;
    RECT 104.87 18.07 105.08 18.14 ;
    RECT 104.87 18.43 105.08 18.5 ;
    RECT 104.87 18.79 105.08 18.86 ;
    RECT 101.09 18.07 101.3 18.14 ;
    RECT 101.09 18.43 101.3 18.5 ;
    RECT 101.09 18.79 101.3 18.86 ;
    RECT 101.55 18.07 101.76 18.14 ;
    RECT 101.55 18.43 101.76 18.5 ;
    RECT 101.55 18.79 101.76 18.86 ;
    RECT 97.77 18.07 97.98 18.14 ;
    RECT 97.77 18.43 97.98 18.5 ;
    RECT 97.77 18.79 97.98 18.86 ;
    RECT 98.23 18.07 98.44 18.14 ;
    RECT 98.23 18.43 98.44 18.5 ;
    RECT 98.23 18.79 98.44 18.86 ;
    RECT 94.45 18.07 94.66 18.14 ;
    RECT 94.45 18.43 94.66 18.5 ;
    RECT 94.45 18.79 94.66 18.86 ;
    RECT 94.91 18.07 95.12 18.14 ;
    RECT 94.91 18.43 95.12 18.5 ;
    RECT 94.91 18.79 95.12 18.86 ;
    RECT 91.13 18.07 91.34 18.14 ;
    RECT 91.13 18.43 91.34 18.5 ;
    RECT 91.13 18.79 91.34 18.86 ;
    RECT 91.59 18.07 91.8 18.14 ;
    RECT 91.59 18.43 91.8 18.5 ;
    RECT 91.59 18.79 91.8 18.86 ;
    RECT 87.81 18.07 88.02 18.14 ;
    RECT 87.81 18.43 88.02 18.5 ;
    RECT 87.81 18.79 88.02 18.86 ;
    RECT 88.27 18.07 88.48 18.14 ;
    RECT 88.27 18.43 88.48 18.5 ;
    RECT 88.27 18.79 88.48 18.86 ;
    RECT 84.49 18.07 84.7 18.14 ;
    RECT 84.49 18.43 84.7 18.5 ;
    RECT 84.49 18.79 84.7 18.86 ;
    RECT 84.95 18.07 85.16 18.14 ;
    RECT 84.95 18.43 85.16 18.5 ;
    RECT 84.95 18.79 85.16 18.86 ;
    RECT 81.17 18.07 81.38 18.14 ;
    RECT 81.17 18.43 81.38 18.5 ;
    RECT 81.17 18.79 81.38 18.86 ;
    RECT 81.63 18.07 81.84 18.14 ;
    RECT 81.63 18.43 81.84 18.5 ;
    RECT 81.63 18.79 81.84 18.86 ;
    RECT 77.85 18.07 78.06 18.14 ;
    RECT 77.85 18.43 78.06 18.5 ;
    RECT 77.85 18.79 78.06 18.86 ;
    RECT 78.31 18.07 78.52 18.14 ;
    RECT 78.31 18.43 78.52 18.5 ;
    RECT 78.31 18.79 78.52 18.86 ;
    RECT 74.53 18.07 74.74 18.14 ;
    RECT 74.53 18.43 74.74 18.5 ;
    RECT 74.53 18.79 74.74 18.86 ;
    RECT 74.99 18.07 75.2 18.14 ;
    RECT 74.99 18.43 75.2 18.5 ;
    RECT 74.99 18.79 75.2 18.86 ;
    RECT 71.21 18.07 71.42 18.14 ;
    RECT 71.21 18.43 71.42 18.5 ;
    RECT 71.21 18.79 71.42 18.86 ;
    RECT 71.67 18.07 71.88 18.14 ;
    RECT 71.67 18.43 71.88 18.5 ;
    RECT 71.67 18.79 71.88 18.86 ;
    RECT 31.37 18.07 31.58 18.14 ;
    RECT 31.37 18.43 31.58 18.5 ;
    RECT 31.37 18.79 31.58 18.86 ;
    RECT 31.83 18.07 32.04 18.14 ;
    RECT 31.83 18.43 32.04 18.5 ;
    RECT 31.83 18.79 32.04 18.86 ;
    RECT 67.89 18.07 68.1 18.14 ;
    RECT 67.89 18.43 68.1 18.5 ;
    RECT 67.89 18.79 68.1 18.86 ;
    RECT 68.35 18.07 68.56 18.14 ;
    RECT 68.35 18.43 68.56 18.5 ;
    RECT 68.35 18.79 68.56 18.86 ;
    RECT 28.05 18.07 28.26 18.14 ;
    RECT 28.05 18.43 28.26 18.5 ;
    RECT 28.05 18.79 28.26 18.86 ;
    RECT 28.51 18.07 28.72 18.14 ;
    RECT 28.51 18.43 28.72 18.5 ;
    RECT 28.51 18.79 28.72 18.86 ;
    RECT 24.73 18.07 24.94 18.14 ;
    RECT 24.73 18.43 24.94 18.5 ;
    RECT 24.73 18.79 24.94 18.86 ;
    RECT 25.19 18.07 25.4 18.14 ;
    RECT 25.19 18.43 25.4 18.5 ;
    RECT 25.19 18.79 25.4 18.86 ;
    RECT 21.41 18.07 21.62 18.14 ;
    RECT 21.41 18.43 21.62 18.5 ;
    RECT 21.41 18.79 21.62 18.86 ;
    RECT 21.87 18.07 22.08 18.14 ;
    RECT 21.87 18.43 22.08 18.5 ;
    RECT 21.87 18.79 22.08 18.86 ;
    RECT 18.09 18.07 18.3 18.14 ;
    RECT 18.09 18.43 18.3 18.5 ;
    RECT 18.09 18.79 18.3 18.86 ;
    RECT 18.55 18.07 18.76 18.14 ;
    RECT 18.55 18.43 18.76 18.5 ;
    RECT 18.55 18.79 18.76 18.86 ;
    RECT 120.825 18.43 120.895 18.5 ;
    RECT 14.77 18.07 14.98 18.14 ;
    RECT 14.77 18.43 14.98 18.5 ;
    RECT 14.77 18.79 14.98 18.86 ;
    RECT 15.23 18.07 15.44 18.14 ;
    RECT 15.23 18.43 15.44 18.5 ;
    RECT 15.23 18.79 15.44 18.86 ;
    RECT 11.45 18.07 11.66 18.14 ;
    RECT 11.45 18.43 11.66 18.5 ;
    RECT 11.45 18.79 11.66 18.86 ;
    RECT 11.91 18.07 12.12 18.14 ;
    RECT 11.91 18.43 12.12 18.5 ;
    RECT 11.91 18.79 12.12 18.86 ;
    RECT 8.13 18.07 8.34 18.14 ;
    RECT 8.13 18.43 8.34 18.5 ;
    RECT 8.13 18.79 8.34 18.86 ;
    RECT 8.59 18.07 8.8 18.14 ;
    RECT 8.59 18.43 8.8 18.5 ;
    RECT 8.59 18.79 8.8 18.86 ;
    RECT 4.81 18.07 5.02 18.14 ;
    RECT 4.81 18.43 5.02 18.5 ;
    RECT 4.81 18.79 5.02 18.86 ;
    RECT 5.27 18.07 5.48 18.14 ;
    RECT 5.27 18.43 5.48 18.5 ;
    RECT 5.27 18.79 5.48 18.86 ;
    RECT 1.49 18.07 1.7 18.14 ;
    RECT 1.49 18.43 1.7 18.5 ;
    RECT 1.49 18.79 1.7 18.86 ;
    RECT 1.95 18.07 2.16 18.14 ;
    RECT 1.95 18.43 2.16 18.5 ;
    RECT 1.95 18.79 2.16 18.86 ;
    RECT 64.57 18.07 64.78 18.14 ;
    RECT 64.57 18.43 64.78 18.5 ;
    RECT 64.57 18.79 64.78 18.86 ;
    RECT 65.03 18.07 65.24 18.14 ;
    RECT 65.03 18.43 65.24 18.5 ;
    RECT 65.03 18.79 65.24 18.86 ;
    RECT 61.25 49.03 61.46 49.1 ;
    RECT 61.25 49.39 61.46 49.46 ;
    RECT 61.25 49.75 61.46 49.82 ;
    RECT 61.71 49.03 61.92 49.1 ;
    RECT 61.71 49.39 61.92 49.46 ;
    RECT 61.71 49.75 61.92 49.82 ;
    RECT 57.93 49.03 58.14 49.1 ;
    RECT 57.93 49.39 58.14 49.46 ;
    RECT 57.93 49.75 58.14 49.82 ;
    RECT 58.39 49.03 58.6 49.1 ;
    RECT 58.39 49.39 58.6 49.46 ;
    RECT 58.39 49.75 58.6 49.82 ;
    RECT 54.61 49.03 54.82 49.1 ;
    RECT 54.61 49.39 54.82 49.46 ;
    RECT 54.61 49.75 54.82 49.82 ;
    RECT 55.07 49.03 55.28 49.1 ;
    RECT 55.07 49.39 55.28 49.46 ;
    RECT 55.07 49.75 55.28 49.82 ;
    RECT 51.29 49.03 51.5 49.1 ;
    RECT 51.29 49.39 51.5 49.46 ;
    RECT 51.29 49.75 51.5 49.82 ;
    RECT 51.75 49.03 51.96 49.1 ;
    RECT 51.75 49.39 51.96 49.46 ;
    RECT 51.75 49.75 51.96 49.82 ;
    RECT 47.97 49.03 48.18 49.1 ;
    RECT 47.97 49.39 48.18 49.46 ;
    RECT 47.97 49.75 48.18 49.82 ;
    RECT 48.43 49.03 48.64 49.1 ;
    RECT 48.43 49.39 48.64 49.46 ;
    RECT 48.43 49.75 48.64 49.82 ;
    RECT 44.65 49.03 44.86 49.1 ;
    RECT 44.65 49.39 44.86 49.46 ;
    RECT 44.65 49.75 44.86 49.82 ;
    RECT 45.11 49.03 45.32 49.1 ;
    RECT 45.11 49.39 45.32 49.46 ;
    RECT 45.11 49.75 45.32 49.82 ;
    RECT 41.33 49.03 41.54 49.1 ;
    RECT 41.33 49.39 41.54 49.46 ;
    RECT 41.33 49.75 41.54 49.82 ;
    RECT 41.79 49.03 42.0 49.1 ;
    RECT 41.79 49.39 42.0 49.46 ;
    RECT 41.79 49.75 42.0 49.82 ;
    RECT 38.01 49.03 38.22 49.1 ;
    RECT 38.01 49.39 38.22 49.46 ;
    RECT 38.01 49.75 38.22 49.82 ;
    RECT 38.47 49.03 38.68 49.1 ;
    RECT 38.47 49.39 38.68 49.46 ;
    RECT 38.47 49.75 38.68 49.82 ;
    RECT 0.4 49.39 0.47 49.46 ;
    RECT 34.69 49.03 34.9 49.1 ;
    RECT 34.69 49.39 34.9 49.46 ;
    RECT 34.69 49.75 34.9 49.82 ;
    RECT 35.15 49.03 35.36 49.1 ;
    RECT 35.15 49.39 35.36 49.46 ;
    RECT 35.15 49.75 35.36 49.82 ;
    RECT 117.69 49.03 117.9 49.1 ;
    RECT 117.69 49.39 117.9 49.46 ;
    RECT 117.69 49.75 117.9 49.82 ;
    RECT 118.15 49.03 118.36 49.1 ;
    RECT 118.15 49.39 118.36 49.46 ;
    RECT 118.15 49.75 118.36 49.82 ;
    RECT 114.37 49.03 114.58 49.1 ;
    RECT 114.37 49.39 114.58 49.46 ;
    RECT 114.37 49.75 114.58 49.82 ;
    RECT 114.83 49.03 115.04 49.1 ;
    RECT 114.83 49.39 115.04 49.46 ;
    RECT 114.83 49.75 115.04 49.82 ;
    RECT 111.05 49.03 111.26 49.1 ;
    RECT 111.05 49.39 111.26 49.46 ;
    RECT 111.05 49.75 111.26 49.82 ;
    RECT 111.51 49.03 111.72 49.1 ;
    RECT 111.51 49.39 111.72 49.46 ;
    RECT 111.51 49.75 111.72 49.82 ;
    RECT 107.73 49.03 107.94 49.1 ;
    RECT 107.73 49.39 107.94 49.46 ;
    RECT 107.73 49.75 107.94 49.82 ;
    RECT 108.19 49.03 108.4 49.1 ;
    RECT 108.19 49.39 108.4 49.46 ;
    RECT 108.19 49.75 108.4 49.82 ;
    RECT 104.41 49.03 104.62 49.1 ;
    RECT 104.41 49.39 104.62 49.46 ;
    RECT 104.41 49.75 104.62 49.82 ;
    RECT 104.87 49.03 105.08 49.1 ;
    RECT 104.87 49.39 105.08 49.46 ;
    RECT 104.87 49.75 105.08 49.82 ;
    RECT 101.09 49.03 101.3 49.1 ;
    RECT 101.09 49.39 101.3 49.46 ;
    RECT 101.09 49.75 101.3 49.82 ;
    RECT 101.55 49.03 101.76 49.1 ;
    RECT 101.55 49.39 101.76 49.46 ;
    RECT 101.55 49.75 101.76 49.82 ;
    RECT 97.77 49.03 97.98 49.1 ;
    RECT 97.77 49.39 97.98 49.46 ;
    RECT 97.77 49.75 97.98 49.82 ;
    RECT 98.23 49.03 98.44 49.1 ;
    RECT 98.23 49.39 98.44 49.46 ;
    RECT 98.23 49.75 98.44 49.82 ;
    RECT 94.45 49.03 94.66 49.1 ;
    RECT 94.45 49.39 94.66 49.46 ;
    RECT 94.45 49.75 94.66 49.82 ;
    RECT 94.91 49.03 95.12 49.1 ;
    RECT 94.91 49.39 95.12 49.46 ;
    RECT 94.91 49.75 95.12 49.82 ;
    RECT 91.13 49.03 91.34 49.1 ;
    RECT 91.13 49.39 91.34 49.46 ;
    RECT 91.13 49.75 91.34 49.82 ;
    RECT 91.59 49.03 91.8 49.1 ;
    RECT 91.59 49.39 91.8 49.46 ;
    RECT 91.59 49.75 91.8 49.82 ;
    RECT 87.81 49.03 88.02 49.1 ;
    RECT 87.81 49.39 88.02 49.46 ;
    RECT 87.81 49.75 88.02 49.82 ;
    RECT 88.27 49.03 88.48 49.1 ;
    RECT 88.27 49.39 88.48 49.46 ;
    RECT 88.27 49.75 88.48 49.82 ;
    RECT 84.49 49.03 84.7 49.1 ;
    RECT 84.49 49.39 84.7 49.46 ;
    RECT 84.49 49.75 84.7 49.82 ;
    RECT 84.95 49.03 85.16 49.1 ;
    RECT 84.95 49.39 85.16 49.46 ;
    RECT 84.95 49.75 85.16 49.82 ;
    RECT 81.17 49.03 81.38 49.1 ;
    RECT 81.17 49.39 81.38 49.46 ;
    RECT 81.17 49.75 81.38 49.82 ;
    RECT 81.63 49.03 81.84 49.1 ;
    RECT 81.63 49.39 81.84 49.46 ;
    RECT 81.63 49.75 81.84 49.82 ;
    RECT 77.85 49.03 78.06 49.1 ;
    RECT 77.85 49.39 78.06 49.46 ;
    RECT 77.85 49.75 78.06 49.82 ;
    RECT 78.31 49.03 78.52 49.1 ;
    RECT 78.31 49.39 78.52 49.46 ;
    RECT 78.31 49.75 78.52 49.82 ;
    RECT 74.53 49.03 74.74 49.1 ;
    RECT 74.53 49.39 74.74 49.46 ;
    RECT 74.53 49.75 74.74 49.82 ;
    RECT 74.99 49.03 75.2 49.1 ;
    RECT 74.99 49.39 75.2 49.46 ;
    RECT 74.99 49.75 75.2 49.82 ;
    RECT 71.21 49.03 71.42 49.1 ;
    RECT 71.21 49.39 71.42 49.46 ;
    RECT 71.21 49.75 71.42 49.82 ;
    RECT 71.67 49.03 71.88 49.1 ;
    RECT 71.67 49.39 71.88 49.46 ;
    RECT 71.67 49.75 71.88 49.82 ;
    RECT 31.37 49.03 31.58 49.1 ;
    RECT 31.37 49.39 31.58 49.46 ;
    RECT 31.37 49.75 31.58 49.82 ;
    RECT 31.83 49.03 32.04 49.1 ;
    RECT 31.83 49.39 32.04 49.46 ;
    RECT 31.83 49.75 32.04 49.82 ;
    RECT 67.89 49.03 68.1 49.1 ;
    RECT 67.89 49.39 68.1 49.46 ;
    RECT 67.89 49.75 68.1 49.82 ;
    RECT 68.35 49.03 68.56 49.1 ;
    RECT 68.35 49.39 68.56 49.46 ;
    RECT 68.35 49.75 68.56 49.82 ;
    RECT 28.05 49.03 28.26 49.1 ;
    RECT 28.05 49.39 28.26 49.46 ;
    RECT 28.05 49.75 28.26 49.82 ;
    RECT 28.51 49.03 28.72 49.1 ;
    RECT 28.51 49.39 28.72 49.46 ;
    RECT 28.51 49.75 28.72 49.82 ;
    RECT 24.73 49.03 24.94 49.1 ;
    RECT 24.73 49.39 24.94 49.46 ;
    RECT 24.73 49.75 24.94 49.82 ;
    RECT 25.19 49.03 25.4 49.1 ;
    RECT 25.19 49.39 25.4 49.46 ;
    RECT 25.19 49.75 25.4 49.82 ;
    RECT 21.41 49.03 21.62 49.1 ;
    RECT 21.41 49.39 21.62 49.46 ;
    RECT 21.41 49.75 21.62 49.82 ;
    RECT 21.87 49.03 22.08 49.1 ;
    RECT 21.87 49.39 22.08 49.46 ;
    RECT 21.87 49.75 22.08 49.82 ;
    RECT 18.09 49.03 18.3 49.1 ;
    RECT 18.09 49.39 18.3 49.46 ;
    RECT 18.09 49.75 18.3 49.82 ;
    RECT 18.55 49.03 18.76 49.1 ;
    RECT 18.55 49.39 18.76 49.46 ;
    RECT 18.55 49.75 18.76 49.82 ;
    RECT 120.825 49.39 120.895 49.46 ;
    RECT 14.77 49.03 14.98 49.1 ;
    RECT 14.77 49.39 14.98 49.46 ;
    RECT 14.77 49.75 14.98 49.82 ;
    RECT 15.23 49.03 15.44 49.1 ;
    RECT 15.23 49.39 15.44 49.46 ;
    RECT 15.23 49.75 15.44 49.82 ;
    RECT 11.45 49.03 11.66 49.1 ;
    RECT 11.45 49.39 11.66 49.46 ;
    RECT 11.45 49.75 11.66 49.82 ;
    RECT 11.91 49.03 12.12 49.1 ;
    RECT 11.91 49.39 12.12 49.46 ;
    RECT 11.91 49.75 12.12 49.82 ;
    RECT 8.13 49.03 8.34 49.1 ;
    RECT 8.13 49.39 8.34 49.46 ;
    RECT 8.13 49.75 8.34 49.82 ;
    RECT 8.59 49.03 8.8 49.1 ;
    RECT 8.59 49.39 8.8 49.46 ;
    RECT 8.59 49.75 8.8 49.82 ;
    RECT 4.81 49.03 5.02 49.1 ;
    RECT 4.81 49.39 5.02 49.46 ;
    RECT 4.81 49.75 5.02 49.82 ;
    RECT 5.27 49.03 5.48 49.1 ;
    RECT 5.27 49.39 5.48 49.46 ;
    RECT 5.27 49.75 5.48 49.82 ;
    RECT 1.49 49.03 1.7 49.1 ;
    RECT 1.49 49.39 1.7 49.46 ;
    RECT 1.49 49.75 1.7 49.82 ;
    RECT 1.95 49.03 2.16 49.1 ;
    RECT 1.95 49.39 2.16 49.46 ;
    RECT 1.95 49.75 2.16 49.82 ;
    RECT 64.57 49.03 64.78 49.1 ;
    RECT 64.57 49.39 64.78 49.46 ;
    RECT 64.57 49.75 64.78 49.82 ;
    RECT 65.03 49.03 65.24 49.1 ;
    RECT 65.03 49.39 65.24 49.46 ;
    RECT 65.03 49.75 65.24 49.82 ;
    RECT 61.25 17.35 61.46 17.42 ;
    RECT 61.25 17.71 61.46 17.78 ;
    RECT 61.25 18.07 61.46 18.14 ;
    RECT 61.71 17.35 61.92 17.42 ;
    RECT 61.71 17.71 61.92 17.78 ;
    RECT 61.71 18.07 61.92 18.14 ;
    RECT 57.93 17.35 58.14 17.42 ;
    RECT 57.93 17.71 58.14 17.78 ;
    RECT 57.93 18.07 58.14 18.14 ;
    RECT 58.39 17.35 58.6 17.42 ;
    RECT 58.39 17.71 58.6 17.78 ;
    RECT 58.39 18.07 58.6 18.14 ;
    RECT 54.61 17.35 54.82 17.42 ;
    RECT 54.61 17.71 54.82 17.78 ;
    RECT 54.61 18.07 54.82 18.14 ;
    RECT 55.07 17.35 55.28 17.42 ;
    RECT 55.07 17.71 55.28 17.78 ;
    RECT 55.07 18.07 55.28 18.14 ;
    RECT 51.29 17.35 51.5 17.42 ;
    RECT 51.29 17.71 51.5 17.78 ;
    RECT 51.29 18.07 51.5 18.14 ;
    RECT 51.75 17.35 51.96 17.42 ;
    RECT 51.75 17.71 51.96 17.78 ;
    RECT 51.75 18.07 51.96 18.14 ;
    RECT 47.97 17.35 48.18 17.42 ;
    RECT 47.97 17.71 48.18 17.78 ;
    RECT 47.97 18.07 48.18 18.14 ;
    RECT 48.43 17.35 48.64 17.42 ;
    RECT 48.43 17.71 48.64 17.78 ;
    RECT 48.43 18.07 48.64 18.14 ;
    RECT 44.65 17.35 44.86 17.42 ;
    RECT 44.65 17.71 44.86 17.78 ;
    RECT 44.65 18.07 44.86 18.14 ;
    RECT 45.11 17.35 45.32 17.42 ;
    RECT 45.11 17.71 45.32 17.78 ;
    RECT 45.11 18.07 45.32 18.14 ;
    RECT 41.33 17.35 41.54 17.42 ;
    RECT 41.33 17.71 41.54 17.78 ;
    RECT 41.33 18.07 41.54 18.14 ;
    RECT 41.79 17.35 42.0 17.42 ;
    RECT 41.79 17.71 42.0 17.78 ;
    RECT 41.79 18.07 42.0 18.14 ;
    RECT 38.01 17.35 38.22 17.42 ;
    RECT 38.01 17.71 38.22 17.78 ;
    RECT 38.01 18.07 38.22 18.14 ;
    RECT 38.47 17.35 38.68 17.42 ;
    RECT 38.47 17.71 38.68 17.78 ;
    RECT 38.47 18.07 38.68 18.14 ;
    RECT 0.4 17.71 0.47 17.78 ;
    RECT 34.69 17.35 34.9 17.42 ;
    RECT 34.69 17.71 34.9 17.78 ;
    RECT 34.69 18.07 34.9 18.14 ;
    RECT 35.15 17.35 35.36 17.42 ;
    RECT 35.15 17.71 35.36 17.78 ;
    RECT 35.15 18.07 35.36 18.14 ;
    RECT 117.69 17.35 117.9 17.42 ;
    RECT 117.69 17.71 117.9 17.78 ;
    RECT 117.69 18.07 117.9 18.14 ;
    RECT 118.15 17.35 118.36 17.42 ;
    RECT 118.15 17.71 118.36 17.78 ;
    RECT 118.15 18.07 118.36 18.14 ;
    RECT 114.37 17.35 114.58 17.42 ;
    RECT 114.37 17.71 114.58 17.78 ;
    RECT 114.37 18.07 114.58 18.14 ;
    RECT 114.83 17.35 115.04 17.42 ;
    RECT 114.83 17.71 115.04 17.78 ;
    RECT 114.83 18.07 115.04 18.14 ;
    RECT 111.05 17.35 111.26 17.42 ;
    RECT 111.05 17.71 111.26 17.78 ;
    RECT 111.05 18.07 111.26 18.14 ;
    RECT 111.51 17.35 111.72 17.42 ;
    RECT 111.51 17.71 111.72 17.78 ;
    RECT 111.51 18.07 111.72 18.14 ;
    RECT 107.73 17.35 107.94 17.42 ;
    RECT 107.73 17.71 107.94 17.78 ;
    RECT 107.73 18.07 107.94 18.14 ;
    RECT 108.19 17.35 108.4 17.42 ;
    RECT 108.19 17.71 108.4 17.78 ;
    RECT 108.19 18.07 108.4 18.14 ;
    RECT 104.41 17.35 104.62 17.42 ;
    RECT 104.41 17.71 104.62 17.78 ;
    RECT 104.41 18.07 104.62 18.14 ;
    RECT 104.87 17.35 105.08 17.42 ;
    RECT 104.87 17.71 105.08 17.78 ;
    RECT 104.87 18.07 105.08 18.14 ;
    RECT 101.09 17.35 101.3 17.42 ;
    RECT 101.09 17.71 101.3 17.78 ;
    RECT 101.09 18.07 101.3 18.14 ;
    RECT 101.55 17.35 101.76 17.42 ;
    RECT 101.55 17.71 101.76 17.78 ;
    RECT 101.55 18.07 101.76 18.14 ;
    RECT 97.77 17.35 97.98 17.42 ;
    RECT 97.77 17.71 97.98 17.78 ;
    RECT 97.77 18.07 97.98 18.14 ;
    RECT 98.23 17.35 98.44 17.42 ;
    RECT 98.23 17.71 98.44 17.78 ;
    RECT 98.23 18.07 98.44 18.14 ;
    RECT 94.45 17.35 94.66 17.42 ;
    RECT 94.45 17.71 94.66 17.78 ;
    RECT 94.45 18.07 94.66 18.14 ;
    RECT 94.91 17.35 95.12 17.42 ;
    RECT 94.91 17.71 95.12 17.78 ;
    RECT 94.91 18.07 95.12 18.14 ;
    RECT 91.13 17.35 91.34 17.42 ;
    RECT 91.13 17.71 91.34 17.78 ;
    RECT 91.13 18.07 91.34 18.14 ;
    RECT 91.59 17.35 91.8 17.42 ;
    RECT 91.59 17.71 91.8 17.78 ;
    RECT 91.59 18.07 91.8 18.14 ;
    RECT 87.81 17.35 88.02 17.42 ;
    RECT 87.81 17.71 88.02 17.78 ;
    RECT 87.81 18.07 88.02 18.14 ;
    RECT 88.27 17.35 88.48 17.42 ;
    RECT 88.27 17.71 88.48 17.78 ;
    RECT 88.27 18.07 88.48 18.14 ;
    RECT 84.49 17.35 84.7 17.42 ;
    RECT 84.49 17.71 84.7 17.78 ;
    RECT 84.49 18.07 84.7 18.14 ;
    RECT 84.95 17.35 85.16 17.42 ;
    RECT 84.95 17.71 85.16 17.78 ;
    RECT 84.95 18.07 85.16 18.14 ;
    RECT 81.17 17.35 81.38 17.42 ;
    RECT 81.17 17.71 81.38 17.78 ;
    RECT 81.17 18.07 81.38 18.14 ;
    RECT 81.63 17.35 81.84 17.42 ;
    RECT 81.63 17.71 81.84 17.78 ;
    RECT 81.63 18.07 81.84 18.14 ;
    RECT 77.85 17.35 78.06 17.42 ;
    RECT 77.85 17.71 78.06 17.78 ;
    RECT 77.85 18.07 78.06 18.14 ;
    RECT 78.31 17.35 78.52 17.42 ;
    RECT 78.31 17.71 78.52 17.78 ;
    RECT 78.31 18.07 78.52 18.14 ;
    RECT 74.53 17.35 74.74 17.42 ;
    RECT 74.53 17.71 74.74 17.78 ;
    RECT 74.53 18.07 74.74 18.14 ;
    RECT 74.99 17.35 75.2 17.42 ;
    RECT 74.99 17.71 75.2 17.78 ;
    RECT 74.99 18.07 75.2 18.14 ;
    RECT 71.21 17.35 71.42 17.42 ;
    RECT 71.21 17.71 71.42 17.78 ;
    RECT 71.21 18.07 71.42 18.14 ;
    RECT 71.67 17.35 71.88 17.42 ;
    RECT 71.67 17.71 71.88 17.78 ;
    RECT 71.67 18.07 71.88 18.14 ;
    RECT 31.37 17.35 31.58 17.42 ;
    RECT 31.37 17.71 31.58 17.78 ;
    RECT 31.37 18.07 31.58 18.14 ;
    RECT 31.83 17.35 32.04 17.42 ;
    RECT 31.83 17.71 32.04 17.78 ;
    RECT 31.83 18.07 32.04 18.14 ;
    RECT 67.89 17.35 68.1 17.42 ;
    RECT 67.89 17.71 68.1 17.78 ;
    RECT 67.89 18.07 68.1 18.14 ;
    RECT 68.35 17.35 68.56 17.42 ;
    RECT 68.35 17.71 68.56 17.78 ;
    RECT 68.35 18.07 68.56 18.14 ;
    RECT 28.05 17.35 28.26 17.42 ;
    RECT 28.05 17.71 28.26 17.78 ;
    RECT 28.05 18.07 28.26 18.14 ;
    RECT 28.51 17.35 28.72 17.42 ;
    RECT 28.51 17.71 28.72 17.78 ;
    RECT 28.51 18.07 28.72 18.14 ;
    RECT 24.73 17.35 24.94 17.42 ;
    RECT 24.73 17.71 24.94 17.78 ;
    RECT 24.73 18.07 24.94 18.14 ;
    RECT 25.19 17.35 25.4 17.42 ;
    RECT 25.19 17.71 25.4 17.78 ;
    RECT 25.19 18.07 25.4 18.14 ;
    RECT 21.41 17.35 21.62 17.42 ;
    RECT 21.41 17.71 21.62 17.78 ;
    RECT 21.41 18.07 21.62 18.14 ;
    RECT 21.87 17.35 22.08 17.42 ;
    RECT 21.87 17.71 22.08 17.78 ;
    RECT 21.87 18.07 22.08 18.14 ;
    RECT 18.09 17.35 18.3 17.42 ;
    RECT 18.09 17.71 18.3 17.78 ;
    RECT 18.09 18.07 18.3 18.14 ;
    RECT 18.55 17.35 18.76 17.42 ;
    RECT 18.55 17.71 18.76 17.78 ;
    RECT 18.55 18.07 18.76 18.14 ;
    RECT 120.825 17.71 120.895 17.78 ;
    RECT 14.77 17.35 14.98 17.42 ;
    RECT 14.77 17.71 14.98 17.78 ;
    RECT 14.77 18.07 14.98 18.14 ;
    RECT 15.23 17.35 15.44 17.42 ;
    RECT 15.23 17.71 15.44 17.78 ;
    RECT 15.23 18.07 15.44 18.14 ;
    RECT 11.45 17.35 11.66 17.42 ;
    RECT 11.45 17.71 11.66 17.78 ;
    RECT 11.45 18.07 11.66 18.14 ;
    RECT 11.91 17.35 12.12 17.42 ;
    RECT 11.91 17.71 12.12 17.78 ;
    RECT 11.91 18.07 12.12 18.14 ;
    RECT 8.13 17.35 8.34 17.42 ;
    RECT 8.13 17.71 8.34 17.78 ;
    RECT 8.13 18.07 8.34 18.14 ;
    RECT 8.59 17.35 8.8 17.42 ;
    RECT 8.59 17.71 8.8 17.78 ;
    RECT 8.59 18.07 8.8 18.14 ;
    RECT 4.81 17.35 5.02 17.42 ;
    RECT 4.81 17.71 5.02 17.78 ;
    RECT 4.81 18.07 5.02 18.14 ;
    RECT 5.27 17.35 5.48 17.42 ;
    RECT 5.27 17.71 5.48 17.78 ;
    RECT 5.27 18.07 5.48 18.14 ;
    RECT 1.49 17.35 1.7 17.42 ;
    RECT 1.49 17.71 1.7 17.78 ;
    RECT 1.49 18.07 1.7 18.14 ;
    RECT 1.95 17.35 2.16 17.42 ;
    RECT 1.95 17.71 2.16 17.78 ;
    RECT 1.95 18.07 2.16 18.14 ;
    RECT 64.57 17.35 64.78 17.42 ;
    RECT 64.57 17.71 64.78 17.78 ;
    RECT 64.57 18.07 64.78 18.14 ;
    RECT 65.03 17.35 65.24 17.42 ;
    RECT 65.03 17.71 65.24 17.78 ;
    RECT 65.03 18.07 65.24 18.14 ;
    RECT 61.25 48.31 61.46 48.38 ;
    RECT 61.25 48.67 61.46 48.74 ;
    RECT 61.25 49.03 61.46 49.1 ;
    RECT 61.71 48.31 61.92 48.38 ;
    RECT 61.71 48.67 61.92 48.74 ;
    RECT 61.71 49.03 61.92 49.1 ;
    RECT 57.93 48.31 58.14 48.38 ;
    RECT 57.93 48.67 58.14 48.74 ;
    RECT 57.93 49.03 58.14 49.1 ;
    RECT 58.39 48.31 58.6 48.38 ;
    RECT 58.39 48.67 58.6 48.74 ;
    RECT 58.39 49.03 58.6 49.1 ;
    RECT 54.61 48.31 54.82 48.38 ;
    RECT 54.61 48.67 54.82 48.74 ;
    RECT 54.61 49.03 54.82 49.1 ;
    RECT 55.07 48.31 55.28 48.38 ;
    RECT 55.07 48.67 55.28 48.74 ;
    RECT 55.07 49.03 55.28 49.1 ;
    RECT 51.29 48.31 51.5 48.38 ;
    RECT 51.29 48.67 51.5 48.74 ;
    RECT 51.29 49.03 51.5 49.1 ;
    RECT 51.75 48.31 51.96 48.38 ;
    RECT 51.75 48.67 51.96 48.74 ;
    RECT 51.75 49.03 51.96 49.1 ;
    RECT 47.97 48.31 48.18 48.38 ;
    RECT 47.97 48.67 48.18 48.74 ;
    RECT 47.97 49.03 48.18 49.1 ;
    RECT 48.43 48.31 48.64 48.38 ;
    RECT 48.43 48.67 48.64 48.74 ;
    RECT 48.43 49.03 48.64 49.1 ;
    RECT 44.65 48.31 44.86 48.38 ;
    RECT 44.65 48.67 44.86 48.74 ;
    RECT 44.65 49.03 44.86 49.1 ;
    RECT 45.11 48.31 45.32 48.38 ;
    RECT 45.11 48.67 45.32 48.74 ;
    RECT 45.11 49.03 45.32 49.1 ;
    RECT 41.33 48.31 41.54 48.38 ;
    RECT 41.33 48.67 41.54 48.74 ;
    RECT 41.33 49.03 41.54 49.1 ;
    RECT 41.79 48.31 42.0 48.38 ;
    RECT 41.79 48.67 42.0 48.74 ;
    RECT 41.79 49.03 42.0 49.1 ;
    RECT 38.01 48.31 38.22 48.38 ;
    RECT 38.01 48.67 38.22 48.74 ;
    RECT 38.01 49.03 38.22 49.1 ;
    RECT 38.47 48.31 38.68 48.38 ;
    RECT 38.47 48.67 38.68 48.74 ;
    RECT 38.47 49.03 38.68 49.1 ;
    RECT 0.4 48.67 0.47 48.74 ;
    RECT 34.69 48.31 34.9 48.38 ;
    RECT 34.69 48.67 34.9 48.74 ;
    RECT 34.69 49.03 34.9 49.1 ;
    RECT 35.15 48.31 35.36 48.38 ;
    RECT 35.15 48.67 35.36 48.74 ;
    RECT 35.15 49.03 35.36 49.1 ;
    RECT 117.69 48.31 117.9 48.38 ;
    RECT 117.69 48.67 117.9 48.74 ;
    RECT 117.69 49.03 117.9 49.1 ;
    RECT 118.15 48.31 118.36 48.38 ;
    RECT 118.15 48.67 118.36 48.74 ;
    RECT 118.15 49.03 118.36 49.1 ;
    RECT 114.37 48.31 114.58 48.38 ;
    RECT 114.37 48.67 114.58 48.74 ;
    RECT 114.37 49.03 114.58 49.1 ;
    RECT 114.83 48.31 115.04 48.38 ;
    RECT 114.83 48.67 115.04 48.74 ;
    RECT 114.83 49.03 115.04 49.1 ;
    RECT 111.05 48.31 111.26 48.38 ;
    RECT 111.05 48.67 111.26 48.74 ;
    RECT 111.05 49.03 111.26 49.1 ;
    RECT 111.51 48.31 111.72 48.38 ;
    RECT 111.51 48.67 111.72 48.74 ;
    RECT 111.51 49.03 111.72 49.1 ;
    RECT 107.73 48.31 107.94 48.38 ;
    RECT 107.73 48.67 107.94 48.74 ;
    RECT 107.73 49.03 107.94 49.1 ;
    RECT 108.19 48.31 108.4 48.38 ;
    RECT 108.19 48.67 108.4 48.74 ;
    RECT 108.19 49.03 108.4 49.1 ;
    RECT 104.41 48.31 104.62 48.38 ;
    RECT 104.41 48.67 104.62 48.74 ;
    RECT 104.41 49.03 104.62 49.1 ;
    RECT 104.87 48.31 105.08 48.38 ;
    RECT 104.87 48.67 105.08 48.74 ;
    RECT 104.87 49.03 105.08 49.1 ;
    RECT 101.09 48.31 101.3 48.38 ;
    RECT 101.09 48.67 101.3 48.74 ;
    RECT 101.09 49.03 101.3 49.1 ;
    RECT 101.55 48.31 101.76 48.38 ;
    RECT 101.55 48.67 101.76 48.74 ;
    RECT 101.55 49.03 101.76 49.1 ;
    RECT 97.77 48.31 97.98 48.38 ;
    RECT 97.77 48.67 97.98 48.74 ;
    RECT 97.77 49.03 97.98 49.1 ;
    RECT 98.23 48.31 98.44 48.38 ;
    RECT 98.23 48.67 98.44 48.74 ;
    RECT 98.23 49.03 98.44 49.1 ;
    RECT 94.45 48.31 94.66 48.38 ;
    RECT 94.45 48.67 94.66 48.74 ;
    RECT 94.45 49.03 94.66 49.1 ;
    RECT 94.91 48.31 95.12 48.38 ;
    RECT 94.91 48.67 95.12 48.74 ;
    RECT 94.91 49.03 95.12 49.1 ;
    RECT 91.13 48.31 91.34 48.38 ;
    RECT 91.13 48.67 91.34 48.74 ;
    RECT 91.13 49.03 91.34 49.1 ;
    RECT 91.59 48.31 91.8 48.38 ;
    RECT 91.59 48.67 91.8 48.74 ;
    RECT 91.59 49.03 91.8 49.1 ;
    RECT 87.81 48.31 88.02 48.38 ;
    RECT 87.81 48.67 88.02 48.74 ;
    RECT 87.81 49.03 88.02 49.1 ;
    RECT 88.27 48.31 88.48 48.38 ;
    RECT 88.27 48.67 88.48 48.74 ;
    RECT 88.27 49.03 88.48 49.1 ;
    RECT 84.49 48.31 84.7 48.38 ;
    RECT 84.49 48.67 84.7 48.74 ;
    RECT 84.49 49.03 84.7 49.1 ;
    RECT 84.95 48.31 85.16 48.38 ;
    RECT 84.95 48.67 85.16 48.74 ;
    RECT 84.95 49.03 85.16 49.1 ;
    RECT 81.17 48.31 81.38 48.38 ;
    RECT 81.17 48.67 81.38 48.74 ;
    RECT 81.17 49.03 81.38 49.1 ;
    RECT 81.63 48.31 81.84 48.38 ;
    RECT 81.63 48.67 81.84 48.74 ;
    RECT 81.63 49.03 81.84 49.1 ;
    RECT 77.85 48.31 78.06 48.38 ;
    RECT 77.85 48.67 78.06 48.74 ;
    RECT 77.85 49.03 78.06 49.1 ;
    RECT 78.31 48.31 78.52 48.38 ;
    RECT 78.31 48.67 78.52 48.74 ;
    RECT 78.31 49.03 78.52 49.1 ;
    RECT 74.53 48.31 74.74 48.38 ;
    RECT 74.53 48.67 74.74 48.74 ;
    RECT 74.53 49.03 74.74 49.1 ;
    RECT 74.99 48.31 75.2 48.38 ;
    RECT 74.99 48.67 75.2 48.74 ;
    RECT 74.99 49.03 75.2 49.1 ;
    RECT 71.21 48.31 71.42 48.38 ;
    RECT 71.21 48.67 71.42 48.74 ;
    RECT 71.21 49.03 71.42 49.1 ;
    RECT 71.67 48.31 71.88 48.38 ;
    RECT 71.67 48.67 71.88 48.74 ;
    RECT 71.67 49.03 71.88 49.1 ;
    RECT 31.37 48.31 31.58 48.38 ;
    RECT 31.37 48.67 31.58 48.74 ;
    RECT 31.37 49.03 31.58 49.1 ;
    RECT 31.83 48.31 32.04 48.38 ;
    RECT 31.83 48.67 32.04 48.74 ;
    RECT 31.83 49.03 32.04 49.1 ;
    RECT 67.89 48.31 68.1 48.38 ;
    RECT 67.89 48.67 68.1 48.74 ;
    RECT 67.89 49.03 68.1 49.1 ;
    RECT 68.35 48.31 68.56 48.38 ;
    RECT 68.35 48.67 68.56 48.74 ;
    RECT 68.35 49.03 68.56 49.1 ;
    RECT 28.05 48.31 28.26 48.38 ;
    RECT 28.05 48.67 28.26 48.74 ;
    RECT 28.05 49.03 28.26 49.1 ;
    RECT 28.51 48.31 28.72 48.38 ;
    RECT 28.51 48.67 28.72 48.74 ;
    RECT 28.51 49.03 28.72 49.1 ;
    RECT 24.73 48.31 24.94 48.38 ;
    RECT 24.73 48.67 24.94 48.74 ;
    RECT 24.73 49.03 24.94 49.1 ;
    RECT 25.19 48.31 25.4 48.38 ;
    RECT 25.19 48.67 25.4 48.74 ;
    RECT 25.19 49.03 25.4 49.1 ;
    RECT 21.41 48.31 21.62 48.38 ;
    RECT 21.41 48.67 21.62 48.74 ;
    RECT 21.41 49.03 21.62 49.1 ;
    RECT 21.87 48.31 22.08 48.38 ;
    RECT 21.87 48.67 22.08 48.74 ;
    RECT 21.87 49.03 22.08 49.1 ;
    RECT 18.09 48.31 18.3 48.38 ;
    RECT 18.09 48.67 18.3 48.74 ;
    RECT 18.09 49.03 18.3 49.1 ;
    RECT 18.55 48.31 18.76 48.38 ;
    RECT 18.55 48.67 18.76 48.74 ;
    RECT 18.55 49.03 18.76 49.1 ;
    RECT 120.825 48.67 120.895 48.74 ;
    RECT 14.77 48.31 14.98 48.38 ;
    RECT 14.77 48.67 14.98 48.74 ;
    RECT 14.77 49.03 14.98 49.1 ;
    RECT 15.23 48.31 15.44 48.38 ;
    RECT 15.23 48.67 15.44 48.74 ;
    RECT 15.23 49.03 15.44 49.1 ;
    RECT 11.45 48.31 11.66 48.38 ;
    RECT 11.45 48.67 11.66 48.74 ;
    RECT 11.45 49.03 11.66 49.1 ;
    RECT 11.91 48.31 12.12 48.38 ;
    RECT 11.91 48.67 12.12 48.74 ;
    RECT 11.91 49.03 12.12 49.1 ;
    RECT 8.13 48.31 8.34 48.38 ;
    RECT 8.13 48.67 8.34 48.74 ;
    RECT 8.13 49.03 8.34 49.1 ;
    RECT 8.59 48.31 8.8 48.38 ;
    RECT 8.59 48.67 8.8 48.74 ;
    RECT 8.59 49.03 8.8 49.1 ;
    RECT 4.81 48.31 5.02 48.38 ;
    RECT 4.81 48.67 5.02 48.74 ;
    RECT 4.81 49.03 5.02 49.1 ;
    RECT 5.27 48.31 5.48 48.38 ;
    RECT 5.27 48.67 5.48 48.74 ;
    RECT 5.27 49.03 5.48 49.1 ;
    RECT 1.49 48.31 1.7 48.38 ;
    RECT 1.49 48.67 1.7 48.74 ;
    RECT 1.49 49.03 1.7 49.1 ;
    RECT 1.95 48.31 2.16 48.38 ;
    RECT 1.95 48.67 2.16 48.74 ;
    RECT 1.95 49.03 2.16 49.1 ;
    RECT 64.57 48.31 64.78 48.38 ;
    RECT 64.57 48.67 64.78 48.74 ;
    RECT 64.57 49.03 64.78 49.1 ;
    RECT 65.03 48.31 65.24 48.38 ;
    RECT 65.03 48.67 65.24 48.74 ;
    RECT 65.03 49.03 65.24 49.1 ;
    RECT 61.25 16.63 61.46 16.7 ;
    RECT 61.25 16.99 61.46 17.06 ;
    RECT 61.25 17.35 61.46 17.42 ;
    RECT 61.71 16.63 61.92 16.7 ;
    RECT 61.71 16.99 61.92 17.06 ;
    RECT 61.71 17.35 61.92 17.42 ;
    RECT 57.93 16.63 58.14 16.7 ;
    RECT 57.93 16.99 58.14 17.06 ;
    RECT 57.93 17.35 58.14 17.42 ;
    RECT 58.39 16.63 58.6 16.7 ;
    RECT 58.39 16.99 58.6 17.06 ;
    RECT 58.39 17.35 58.6 17.42 ;
    RECT 54.61 16.63 54.82 16.7 ;
    RECT 54.61 16.99 54.82 17.06 ;
    RECT 54.61 17.35 54.82 17.42 ;
    RECT 55.07 16.63 55.28 16.7 ;
    RECT 55.07 16.99 55.28 17.06 ;
    RECT 55.07 17.35 55.28 17.42 ;
    RECT 51.29 16.63 51.5 16.7 ;
    RECT 51.29 16.99 51.5 17.06 ;
    RECT 51.29 17.35 51.5 17.42 ;
    RECT 51.75 16.63 51.96 16.7 ;
    RECT 51.75 16.99 51.96 17.06 ;
    RECT 51.75 17.35 51.96 17.42 ;
    RECT 47.97 16.63 48.18 16.7 ;
    RECT 47.97 16.99 48.18 17.06 ;
    RECT 47.97 17.35 48.18 17.42 ;
    RECT 48.43 16.63 48.64 16.7 ;
    RECT 48.43 16.99 48.64 17.06 ;
    RECT 48.43 17.35 48.64 17.42 ;
    RECT 44.65 16.63 44.86 16.7 ;
    RECT 44.65 16.99 44.86 17.06 ;
    RECT 44.65 17.35 44.86 17.42 ;
    RECT 45.11 16.63 45.32 16.7 ;
    RECT 45.11 16.99 45.32 17.06 ;
    RECT 45.11 17.35 45.32 17.42 ;
    RECT 41.33 16.63 41.54 16.7 ;
    RECT 41.33 16.99 41.54 17.06 ;
    RECT 41.33 17.35 41.54 17.42 ;
    RECT 41.79 16.63 42.0 16.7 ;
    RECT 41.79 16.99 42.0 17.06 ;
    RECT 41.79 17.35 42.0 17.42 ;
    RECT 38.01 16.63 38.22 16.7 ;
    RECT 38.01 16.99 38.22 17.06 ;
    RECT 38.01 17.35 38.22 17.42 ;
    RECT 38.47 16.63 38.68 16.7 ;
    RECT 38.47 16.99 38.68 17.06 ;
    RECT 38.47 17.35 38.68 17.42 ;
    RECT 0.4 16.99 0.47 17.06 ;
    RECT 34.69 16.63 34.9 16.7 ;
    RECT 34.69 16.99 34.9 17.06 ;
    RECT 34.69 17.35 34.9 17.42 ;
    RECT 35.15 16.63 35.36 16.7 ;
    RECT 35.15 16.99 35.36 17.06 ;
    RECT 35.15 17.35 35.36 17.42 ;
    RECT 117.69 16.63 117.9 16.7 ;
    RECT 117.69 16.99 117.9 17.06 ;
    RECT 117.69 17.35 117.9 17.42 ;
    RECT 118.15 16.63 118.36 16.7 ;
    RECT 118.15 16.99 118.36 17.06 ;
    RECT 118.15 17.35 118.36 17.42 ;
    RECT 114.37 16.63 114.58 16.7 ;
    RECT 114.37 16.99 114.58 17.06 ;
    RECT 114.37 17.35 114.58 17.42 ;
    RECT 114.83 16.63 115.04 16.7 ;
    RECT 114.83 16.99 115.04 17.06 ;
    RECT 114.83 17.35 115.04 17.42 ;
    RECT 111.05 16.63 111.26 16.7 ;
    RECT 111.05 16.99 111.26 17.06 ;
    RECT 111.05 17.35 111.26 17.42 ;
    RECT 111.51 16.63 111.72 16.7 ;
    RECT 111.51 16.99 111.72 17.06 ;
    RECT 111.51 17.35 111.72 17.42 ;
    RECT 107.73 16.63 107.94 16.7 ;
    RECT 107.73 16.99 107.94 17.06 ;
    RECT 107.73 17.35 107.94 17.42 ;
    RECT 108.19 16.63 108.4 16.7 ;
    RECT 108.19 16.99 108.4 17.06 ;
    RECT 108.19 17.35 108.4 17.42 ;
    RECT 104.41 16.63 104.62 16.7 ;
    RECT 104.41 16.99 104.62 17.06 ;
    RECT 104.41 17.35 104.62 17.42 ;
    RECT 104.87 16.63 105.08 16.7 ;
    RECT 104.87 16.99 105.08 17.06 ;
    RECT 104.87 17.35 105.08 17.42 ;
    RECT 101.09 16.63 101.3 16.7 ;
    RECT 101.09 16.99 101.3 17.06 ;
    RECT 101.09 17.35 101.3 17.42 ;
    RECT 101.55 16.63 101.76 16.7 ;
    RECT 101.55 16.99 101.76 17.06 ;
    RECT 101.55 17.35 101.76 17.42 ;
    RECT 97.77 16.63 97.98 16.7 ;
    RECT 97.77 16.99 97.98 17.06 ;
    RECT 97.77 17.35 97.98 17.42 ;
    RECT 98.23 16.63 98.44 16.7 ;
    RECT 98.23 16.99 98.44 17.06 ;
    RECT 98.23 17.35 98.44 17.42 ;
    RECT 94.45 16.63 94.66 16.7 ;
    RECT 94.45 16.99 94.66 17.06 ;
    RECT 94.45 17.35 94.66 17.42 ;
    RECT 94.91 16.63 95.12 16.7 ;
    RECT 94.91 16.99 95.12 17.06 ;
    RECT 94.91 17.35 95.12 17.42 ;
    RECT 91.13 16.63 91.34 16.7 ;
    RECT 91.13 16.99 91.34 17.06 ;
    RECT 91.13 17.35 91.34 17.42 ;
    RECT 91.59 16.63 91.8 16.7 ;
    RECT 91.59 16.99 91.8 17.06 ;
    RECT 91.59 17.35 91.8 17.42 ;
    RECT 87.81 16.63 88.02 16.7 ;
    RECT 87.81 16.99 88.02 17.06 ;
    RECT 87.81 17.35 88.02 17.42 ;
    RECT 88.27 16.63 88.48 16.7 ;
    RECT 88.27 16.99 88.48 17.06 ;
    RECT 88.27 17.35 88.48 17.42 ;
    RECT 84.49 16.63 84.7 16.7 ;
    RECT 84.49 16.99 84.7 17.06 ;
    RECT 84.49 17.35 84.7 17.42 ;
    RECT 84.95 16.63 85.16 16.7 ;
    RECT 84.95 16.99 85.16 17.06 ;
    RECT 84.95 17.35 85.16 17.42 ;
    RECT 81.17 16.63 81.38 16.7 ;
    RECT 81.17 16.99 81.38 17.06 ;
    RECT 81.17 17.35 81.38 17.42 ;
    RECT 81.63 16.63 81.84 16.7 ;
    RECT 81.63 16.99 81.84 17.06 ;
    RECT 81.63 17.35 81.84 17.42 ;
    RECT 77.85 16.63 78.06 16.7 ;
    RECT 77.85 16.99 78.06 17.06 ;
    RECT 77.85 17.35 78.06 17.42 ;
    RECT 78.31 16.63 78.52 16.7 ;
    RECT 78.31 16.99 78.52 17.06 ;
    RECT 78.31 17.35 78.52 17.42 ;
    RECT 74.53 16.63 74.74 16.7 ;
    RECT 74.53 16.99 74.74 17.06 ;
    RECT 74.53 17.35 74.74 17.42 ;
    RECT 74.99 16.63 75.2 16.7 ;
    RECT 74.99 16.99 75.2 17.06 ;
    RECT 74.99 17.35 75.2 17.42 ;
    RECT 71.21 16.63 71.42 16.7 ;
    RECT 71.21 16.99 71.42 17.06 ;
    RECT 71.21 17.35 71.42 17.42 ;
    RECT 71.67 16.63 71.88 16.7 ;
    RECT 71.67 16.99 71.88 17.06 ;
    RECT 71.67 17.35 71.88 17.42 ;
    RECT 31.37 16.63 31.58 16.7 ;
    RECT 31.37 16.99 31.58 17.06 ;
    RECT 31.37 17.35 31.58 17.42 ;
    RECT 31.83 16.63 32.04 16.7 ;
    RECT 31.83 16.99 32.04 17.06 ;
    RECT 31.83 17.35 32.04 17.42 ;
    RECT 67.89 16.63 68.1 16.7 ;
    RECT 67.89 16.99 68.1 17.06 ;
    RECT 67.89 17.35 68.1 17.42 ;
    RECT 68.35 16.63 68.56 16.7 ;
    RECT 68.35 16.99 68.56 17.06 ;
    RECT 68.35 17.35 68.56 17.42 ;
    RECT 28.05 16.63 28.26 16.7 ;
    RECT 28.05 16.99 28.26 17.06 ;
    RECT 28.05 17.35 28.26 17.42 ;
    RECT 28.51 16.63 28.72 16.7 ;
    RECT 28.51 16.99 28.72 17.06 ;
    RECT 28.51 17.35 28.72 17.42 ;
    RECT 24.73 16.63 24.94 16.7 ;
    RECT 24.73 16.99 24.94 17.06 ;
    RECT 24.73 17.35 24.94 17.42 ;
    RECT 25.19 16.63 25.4 16.7 ;
    RECT 25.19 16.99 25.4 17.06 ;
    RECT 25.19 17.35 25.4 17.42 ;
    RECT 21.41 16.63 21.62 16.7 ;
    RECT 21.41 16.99 21.62 17.06 ;
    RECT 21.41 17.35 21.62 17.42 ;
    RECT 21.87 16.63 22.08 16.7 ;
    RECT 21.87 16.99 22.08 17.06 ;
    RECT 21.87 17.35 22.08 17.42 ;
    RECT 18.09 16.63 18.3 16.7 ;
    RECT 18.09 16.99 18.3 17.06 ;
    RECT 18.09 17.35 18.3 17.42 ;
    RECT 18.55 16.63 18.76 16.7 ;
    RECT 18.55 16.99 18.76 17.06 ;
    RECT 18.55 17.35 18.76 17.42 ;
    RECT 120.825 16.99 120.895 17.06 ;
    RECT 14.77 16.63 14.98 16.7 ;
    RECT 14.77 16.99 14.98 17.06 ;
    RECT 14.77 17.35 14.98 17.42 ;
    RECT 15.23 16.63 15.44 16.7 ;
    RECT 15.23 16.99 15.44 17.06 ;
    RECT 15.23 17.35 15.44 17.42 ;
    RECT 11.45 16.63 11.66 16.7 ;
    RECT 11.45 16.99 11.66 17.06 ;
    RECT 11.45 17.35 11.66 17.42 ;
    RECT 11.91 16.63 12.12 16.7 ;
    RECT 11.91 16.99 12.12 17.06 ;
    RECT 11.91 17.35 12.12 17.42 ;
    RECT 8.13 16.63 8.34 16.7 ;
    RECT 8.13 16.99 8.34 17.06 ;
    RECT 8.13 17.35 8.34 17.42 ;
    RECT 8.59 16.63 8.8 16.7 ;
    RECT 8.59 16.99 8.8 17.06 ;
    RECT 8.59 17.35 8.8 17.42 ;
    RECT 4.81 16.63 5.02 16.7 ;
    RECT 4.81 16.99 5.02 17.06 ;
    RECT 4.81 17.35 5.02 17.42 ;
    RECT 5.27 16.63 5.48 16.7 ;
    RECT 5.27 16.99 5.48 17.06 ;
    RECT 5.27 17.35 5.48 17.42 ;
    RECT 1.49 16.63 1.7 16.7 ;
    RECT 1.49 16.99 1.7 17.06 ;
    RECT 1.49 17.35 1.7 17.42 ;
    RECT 1.95 16.63 2.16 16.7 ;
    RECT 1.95 16.99 2.16 17.06 ;
    RECT 1.95 17.35 2.16 17.42 ;
    RECT 64.57 16.63 64.78 16.7 ;
    RECT 64.57 16.99 64.78 17.06 ;
    RECT 64.57 17.35 64.78 17.42 ;
    RECT 65.03 16.63 65.24 16.7 ;
    RECT 65.03 16.99 65.24 17.06 ;
    RECT 65.03 17.35 65.24 17.42 ;
    RECT 61.25 47.59 61.46 47.66 ;
    RECT 61.25 47.95 61.46 48.02 ;
    RECT 61.25 48.31 61.46 48.38 ;
    RECT 61.71 47.59 61.92 47.66 ;
    RECT 61.71 47.95 61.92 48.02 ;
    RECT 61.71 48.31 61.92 48.38 ;
    RECT 57.93 47.59 58.14 47.66 ;
    RECT 57.93 47.95 58.14 48.02 ;
    RECT 57.93 48.31 58.14 48.38 ;
    RECT 58.39 47.59 58.6 47.66 ;
    RECT 58.39 47.95 58.6 48.02 ;
    RECT 58.39 48.31 58.6 48.38 ;
    RECT 54.61 47.59 54.82 47.66 ;
    RECT 54.61 47.95 54.82 48.02 ;
    RECT 54.61 48.31 54.82 48.38 ;
    RECT 55.07 47.59 55.28 47.66 ;
    RECT 55.07 47.95 55.28 48.02 ;
    RECT 55.07 48.31 55.28 48.38 ;
    RECT 51.29 47.59 51.5 47.66 ;
    RECT 51.29 47.95 51.5 48.02 ;
    RECT 51.29 48.31 51.5 48.38 ;
    RECT 51.75 47.59 51.96 47.66 ;
    RECT 51.75 47.95 51.96 48.02 ;
    RECT 51.75 48.31 51.96 48.38 ;
    RECT 47.97 47.59 48.18 47.66 ;
    RECT 47.97 47.95 48.18 48.02 ;
    RECT 47.97 48.31 48.18 48.38 ;
    RECT 48.43 47.59 48.64 47.66 ;
    RECT 48.43 47.95 48.64 48.02 ;
    RECT 48.43 48.31 48.64 48.38 ;
    RECT 44.65 47.59 44.86 47.66 ;
    RECT 44.65 47.95 44.86 48.02 ;
    RECT 44.65 48.31 44.86 48.38 ;
    RECT 45.11 47.59 45.32 47.66 ;
    RECT 45.11 47.95 45.32 48.02 ;
    RECT 45.11 48.31 45.32 48.38 ;
    RECT 41.33 47.59 41.54 47.66 ;
    RECT 41.33 47.95 41.54 48.02 ;
    RECT 41.33 48.31 41.54 48.38 ;
    RECT 41.79 47.59 42.0 47.66 ;
    RECT 41.79 47.95 42.0 48.02 ;
    RECT 41.79 48.31 42.0 48.38 ;
    RECT 38.01 47.59 38.22 47.66 ;
    RECT 38.01 47.95 38.22 48.02 ;
    RECT 38.01 48.31 38.22 48.38 ;
    RECT 38.47 47.59 38.68 47.66 ;
    RECT 38.47 47.95 38.68 48.02 ;
    RECT 38.47 48.31 38.68 48.38 ;
    RECT 0.4 47.95 0.47 48.02 ;
    RECT 34.69 47.59 34.9 47.66 ;
    RECT 34.69 47.95 34.9 48.02 ;
    RECT 34.69 48.31 34.9 48.38 ;
    RECT 35.15 47.59 35.36 47.66 ;
    RECT 35.15 47.95 35.36 48.02 ;
    RECT 35.15 48.31 35.36 48.38 ;
    RECT 117.69 47.59 117.9 47.66 ;
    RECT 117.69 47.95 117.9 48.02 ;
    RECT 117.69 48.31 117.9 48.38 ;
    RECT 118.15 47.59 118.36 47.66 ;
    RECT 118.15 47.95 118.36 48.02 ;
    RECT 118.15 48.31 118.36 48.38 ;
    RECT 114.37 47.59 114.58 47.66 ;
    RECT 114.37 47.95 114.58 48.02 ;
    RECT 114.37 48.31 114.58 48.38 ;
    RECT 114.83 47.59 115.04 47.66 ;
    RECT 114.83 47.95 115.04 48.02 ;
    RECT 114.83 48.31 115.04 48.38 ;
    RECT 111.05 47.59 111.26 47.66 ;
    RECT 111.05 47.95 111.26 48.02 ;
    RECT 111.05 48.31 111.26 48.38 ;
    RECT 111.51 47.59 111.72 47.66 ;
    RECT 111.51 47.95 111.72 48.02 ;
    RECT 111.51 48.31 111.72 48.38 ;
    RECT 107.73 47.59 107.94 47.66 ;
    RECT 107.73 47.95 107.94 48.02 ;
    RECT 107.73 48.31 107.94 48.38 ;
    RECT 108.19 47.59 108.4 47.66 ;
    RECT 108.19 47.95 108.4 48.02 ;
    RECT 108.19 48.31 108.4 48.38 ;
    RECT 104.41 47.59 104.62 47.66 ;
    RECT 104.41 47.95 104.62 48.02 ;
    RECT 104.41 48.31 104.62 48.38 ;
    RECT 104.87 47.59 105.08 47.66 ;
    RECT 104.87 47.95 105.08 48.02 ;
    RECT 104.87 48.31 105.08 48.38 ;
    RECT 101.09 47.59 101.3 47.66 ;
    RECT 101.09 47.95 101.3 48.02 ;
    RECT 101.09 48.31 101.3 48.38 ;
    RECT 101.55 47.59 101.76 47.66 ;
    RECT 101.55 47.95 101.76 48.02 ;
    RECT 101.55 48.31 101.76 48.38 ;
    RECT 97.77 47.59 97.98 47.66 ;
    RECT 97.77 47.95 97.98 48.02 ;
    RECT 97.77 48.31 97.98 48.38 ;
    RECT 98.23 47.59 98.44 47.66 ;
    RECT 98.23 47.95 98.44 48.02 ;
    RECT 98.23 48.31 98.44 48.38 ;
    RECT 94.45 47.59 94.66 47.66 ;
    RECT 94.45 47.95 94.66 48.02 ;
    RECT 94.45 48.31 94.66 48.38 ;
    RECT 94.91 47.59 95.12 47.66 ;
    RECT 94.91 47.95 95.12 48.02 ;
    RECT 94.91 48.31 95.12 48.38 ;
    RECT 91.13 47.59 91.34 47.66 ;
    RECT 91.13 47.95 91.34 48.02 ;
    RECT 91.13 48.31 91.34 48.38 ;
    RECT 91.59 47.59 91.8 47.66 ;
    RECT 91.59 47.95 91.8 48.02 ;
    RECT 91.59 48.31 91.8 48.38 ;
    RECT 87.81 47.59 88.02 47.66 ;
    RECT 87.81 47.95 88.02 48.02 ;
    RECT 87.81 48.31 88.02 48.38 ;
    RECT 88.27 47.59 88.48 47.66 ;
    RECT 88.27 47.95 88.48 48.02 ;
    RECT 88.27 48.31 88.48 48.38 ;
    RECT 84.49 47.59 84.7 47.66 ;
    RECT 84.49 47.95 84.7 48.02 ;
    RECT 84.49 48.31 84.7 48.38 ;
    RECT 84.95 47.59 85.16 47.66 ;
    RECT 84.95 47.95 85.16 48.02 ;
    RECT 84.95 48.31 85.16 48.38 ;
    RECT 81.17 47.59 81.38 47.66 ;
    RECT 81.17 47.95 81.38 48.02 ;
    RECT 81.17 48.31 81.38 48.38 ;
    RECT 81.63 47.59 81.84 47.66 ;
    RECT 81.63 47.95 81.84 48.02 ;
    RECT 81.63 48.31 81.84 48.38 ;
    RECT 77.85 47.59 78.06 47.66 ;
    RECT 77.85 47.95 78.06 48.02 ;
    RECT 77.85 48.31 78.06 48.38 ;
    RECT 78.31 47.59 78.52 47.66 ;
    RECT 78.31 47.95 78.52 48.02 ;
    RECT 78.31 48.31 78.52 48.38 ;
    RECT 74.53 47.59 74.74 47.66 ;
    RECT 74.53 47.95 74.74 48.02 ;
    RECT 74.53 48.31 74.74 48.38 ;
    RECT 74.99 47.59 75.2 47.66 ;
    RECT 74.99 47.95 75.2 48.02 ;
    RECT 74.99 48.31 75.2 48.38 ;
    RECT 71.21 47.59 71.42 47.66 ;
    RECT 71.21 47.95 71.42 48.02 ;
    RECT 71.21 48.31 71.42 48.38 ;
    RECT 71.67 47.59 71.88 47.66 ;
    RECT 71.67 47.95 71.88 48.02 ;
    RECT 71.67 48.31 71.88 48.38 ;
    RECT 31.37 47.59 31.58 47.66 ;
    RECT 31.37 47.95 31.58 48.02 ;
    RECT 31.37 48.31 31.58 48.38 ;
    RECT 31.83 47.59 32.04 47.66 ;
    RECT 31.83 47.95 32.04 48.02 ;
    RECT 31.83 48.31 32.04 48.38 ;
    RECT 67.89 47.59 68.1 47.66 ;
    RECT 67.89 47.95 68.1 48.02 ;
    RECT 67.89 48.31 68.1 48.38 ;
    RECT 68.35 47.59 68.56 47.66 ;
    RECT 68.35 47.95 68.56 48.02 ;
    RECT 68.35 48.31 68.56 48.38 ;
    RECT 28.05 47.59 28.26 47.66 ;
    RECT 28.05 47.95 28.26 48.02 ;
    RECT 28.05 48.31 28.26 48.38 ;
    RECT 28.51 47.59 28.72 47.66 ;
    RECT 28.51 47.95 28.72 48.02 ;
    RECT 28.51 48.31 28.72 48.38 ;
    RECT 24.73 47.59 24.94 47.66 ;
    RECT 24.73 47.95 24.94 48.02 ;
    RECT 24.73 48.31 24.94 48.38 ;
    RECT 25.19 47.59 25.4 47.66 ;
    RECT 25.19 47.95 25.4 48.02 ;
    RECT 25.19 48.31 25.4 48.38 ;
    RECT 21.41 47.59 21.62 47.66 ;
    RECT 21.41 47.95 21.62 48.02 ;
    RECT 21.41 48.31 21.62 48.38 ;
    RECT 21.87 47.59 22.08 47.66 ;
    RECT 21.87 47.95 22.08 48.02 ;
    RECT 21.87 48.31 22.08 48.38 ;
    RECT 18.09 47.59 18.3 47.66 ;
    RECT 18.09 47.95 18.3 48.02 ;
    RECT 18.09 48.31 18.3 48.38 ;
    RECT 18.55 47.59 18.76 47.66 ;
    RECT 18.55 47.95 18.76 48.02 ;
    RECT 18.55 48.31 18.76 48.38 ;
    RECT 120.825 47.95 120.895 48.02 ;
    RECT 14.77 47.59 14.98 47.66 ;
    RECT 14.77 47.95 14.98 48.02 ;
    RECT 14.77 48.31 14.98 48.38 ;
    RECT 15.23 47.59 15.44 47.66 ;
    RECT 15.23 47.95 15.44 48.02 ;
    RECT 15.23 48.31 15.44 48.38 ;
    RECT 11.45 47.59 11.66 47.66 ;
    RECT 11.45 47.95 11.66 48.02 ;
    RECT 11.45 48.31 11.66 48.38 ;
    RECT 11.91 47.59 12.12 47.66 ;
    RECT 11.91 47.95 12.12 48.02 ;
    RECT 11.91 48.31 12.12 48.38 ;
    RECT 8.13 47.59 8.34 47.66 ;
    RECT 8.13 47.95 8.34 48.02 ;
    RECT 8.13 48.31 8.34 48.38 ;
    RECT 8.59 47.59 8.8 47.66 ;
    RECT 8.59 47.95 8.8 48.02 ;
    RECT 8.59 48.31 8.8 48.38 ;
    RECT 4.81 47.59 5.02 47.66 ;
    RECT 4.81 47.95 5.02 48.02 ;
    RECT 4.81 48.31 5.02 48.38 ;
    RECT 5.27 47.59 5.48 47.66 ;
    RECT 5.27 47.95 5.48 48.02 ;
    RECT 5.27 48.31 5.48 48.38 ;
    RECT 1.49 47.59 1.7 47.66 ;
    RECT 1.49 47.95 1.7 48.02 ;
    RECT 1.49 48.31 1.7 48.38 ;
    RECT 1.95 47.59 2.16 47.66 ;
    RECT 1.95 47.95 2.16 48.02 ;
    RECT 1.95 48.31 2.16 48.38 ;
    RECT 64.57 47.59 64.78 47.66 ;
    RECT 64.57 47.95 64.78 48.02 ;
    RECT 64.57 48.31 64.78 48.38 ;
    RECT 65.03 47.59 65.24 47.66 ;
    RECT 65.03 47.95 65.24 48.02 ;
    RECT 65.03 48.31 65.24 48.38 ;
    RECT 61.25 15.91 61.46 15.98 ;
    RECT 61.25 16.27 61.46 16.34 ;
    RECT 61.25 16.63 61.46 16.7 ;
    RECT 61.71 15.91 61.92 15.98 ;
    RECT 61.71 16.27 61.92 16.34 ;
    RECT 61.71 16.63 61.92 16.7 ;
    RECT 57.93 15.91 58.14 15.98 ;
    RECT 57.93 16.27 58.14 16.34 ;
    RECT 57.93 16.63 58.14 16.7 ;
    RECT 58.39 15.91 58.6 15.98 ;
    RECT 58.39 16.27 58.6 16.34 ;
    RECT 58.39 16.63 58.6 16.7 ;
    RECT 54.61 15.91 54.82 15.98 ;
    RECT 54.61 16.27 54.82 16.34 ;
    RECT 54.61 16.63 54.82 16.7 ;
    RECT 55.07 15.91 55.28 15.98 ;
    RECT 55.07 16.27 55.28 16.34 ;
    RECT 55.07 16.63 55.28 16.7 ;
    RECT 51.29 15.91 51.5 15.98 ;
    RECT 51.29 16.27 51.5 16.34 ;
    RECT 51.29 16.63 51.5 16.7 ;
    RECT 51.75 15.91 51.96 15.98 ;
    RECT 51.75 16.27 51.96 16.34 ;
    RECT 51.75 16.63 51.96 16.7 ;
    RECT 47.97 15.91 48.18 15.98 ;
    RECT 47.97 16.27 48.18 16.34 ;
    RECT 47.97 16.63 48.18 16.7 ;
    RECT 48.43 15.91 48.64 15.98 ;
    RECT 48.43 16.27 48.64 16.34 ;
    RECT 48.43 16.63 48.64 16.7 ;
    RECT 44.65 15.91 44.86 15.98 ;
    RECT 44.65 16.27 44.86 16.34 ;
    RECT 44.65 16.63 44.86 16.7 ;
    RECT 45.11 15.91 45.32 15.98 ;
    RECT 45.11 16.27 45.32 16.34 ;
    RECT 45.11 16.63 45.32 16.7 ;
    RECT 41.33 15.91 41.54 15.98 ;
    RECT 41.33 16.27 41.54 16.34 ;
    RECT 41.33 16.63 41.54 16.7 ;
    RECT 41.79 15.91 42.0 15.98 ;
    RECT 41.79 16.27 42.0 16.34 ;
    RECT 41.79 16.63 42.0 16.7 ;
    RECT 38.01 15.91 38.22 15.98 ;
    RECT 38.01 16.27 38.22 16.34 ;
    RECT 38.01 16.63 38.22 16.7 ;
    RECT 38.47 15.91 38.68 15.98 ;
    RECT 38.47 16.27 38.68 16.34 ;
    RECT 38.47 16.63 38.68 16.7 ;
    RECT 0.4 16.27 0.47 16.34 ;
    RECT 34.69 15.91 34.9 15.98 ;
    RECT 34.69 16.27 34.9 16.34 ;
    RECT 34.69 16.63 34.9 16.7 ;
    RECT 35.15 15.91 35.36 15.98 ;
    RECT 35.15 16.27 35.36 16.34 ;
    RECT 35.15 16.63 35.36 16.7 ;
    RECT 117.69 15.91 117.9 15.98 ;
    RECT 117.69 16.27 117.9 16.34 ;
    RECT 117.69 16.63 117.9 16.7 ;
    RECT 118.15 15.91 118.36 15.98 ;
    RECT 118.15 16.27 118.36 16.34 ;
    RECT 118.15 16.63 118.36 16.7 ;
    RECT 114.37 15.91 114.58 15.98 ;
    RECT 114.37 16.27 114.58 16.34 ;
    RECT 114.37 16.63 114.58 16.7 ;
    RECT 114.83 15.91 115.04 15.98 ;
    RECT 114.83 16.27 115.04 16.34 ;
    RECT 114.83 16.63 115.04 16.7 ;
    RECT 111.05 15.91 111.26 15.98 ;
    RECT 111.05 16.27 111.26 16.34 ;
    RECT 111.05 16.63 111.26 16.7 ;
    RECT 111.51 15.91 111.72 15.98 ;
    RECT 111.51 16.27 111.72 16.34 ;
    RECT 111.51 16.63 111.72 16.7 ;
    RECT 107.73 15.91 107.94 15.98 ;
    RECT 107.73 16.27 107.94 16.34 ;
    RECT 107.73 16.63 107.94 16.7 ;
    RECT 108.19 15.91 108.4 15.98 ;
    RECT 108.19 16.27 108.4 16.34 ;
    RECT 108.19 16.63 108.4 16.7 ;
    RECT 104.41 15.91 104.62 15.98 ;
    RECT 104.41 16.27 104.62 16.34 ;
    RECT 104.41 16.63 104.62 16.7 ;
    RECT 104.87 15.91 105.08 15.98 ;
    RECT 104.87 16.27 105.08 16.34 ;
    RECT 104.87 16.63 105.08 16.7 ;
    RECT 101.09 15.91 101.3 15.98 ;
    RECT 101.09 16.27 101.3 16.34 ;
    RECT 101.09 16.63 101.3 16.7 ;
    RECT 101.55 15.91 101.76 15.98 ;
    RECT 101.55 16.27 101.76 16.34 ;
    RECT 101.55 16.63 101.76 16.7 ;
    RECT 97.77 15.91 97.98 15.98 ;
    RECT 97.77 16.27 97.98 16.34 ;
    RECT 97.77 16.63 97.98 16.7 ;
    RECT 98.23 15.91 98.44 15.98 ;
    RECT 98.23 16.27 98.44 16.34 ;
    RECT 98.23 16.63 98.44 16.7 ;
    RECT 94.45 15.91 94.66 15.98 ;
    RECT 94.45 16.27 94.66 16.34 ;
    RECT 94.45 16.63 94.66 16.7 ;
    RECT 94.91 15.91 95.12 15.98 ;
    RECT 94.91 16.27 95.12 16.34 ;
    RECT 94.91 16.63 95.12 16.7 ;
    RECT 91.13 15.91 91.34 15.98 ;
    RECT 91.13 16.27 91.34 16.34 ;
    RECT 91.13 16.63 91.34 16.7 ;
    RECT 91.59 15.91 91.8 15.98 ;
    RECT 91.59 16.27 91.8 16.34 ;
    RECT 91.59 16.63 91.8 16.7 ;
    RECT 87.81 15.91 88.02 15.98 ;
    RECT 87.81 16.27 88.02 16.34 ;
    RECT 87.81 16.63 88.02 16.7 ;
    RECT 88.27 15.91 88.48 15.98 ;
    RECT 88.27 16.27 88.48 16.34 ;
    RECT 88.27 16.63 88.48 16.7 ;
    RECT 84.49 15.91 84.7 15.98 ;
    RECT 84.49 16.27 84.7 16.34 ;
    RECT 84.49 16.63 84.7 16.7 ;
    RECT 84.95 15.91 85.16 15.98 ;
    RECT 84.95 16.27 85.16 16.34 ;
    RECT 84.95 16.63 85.16 16.7 ;
    RECT 81.17 15.91 81.38 15.98 ;
    RECT 81.17 16.27 81.38 16.34 ;
    RECT 81.17 16.63 81.38 16.7 ;
    RECT 81.63 15.91 81.84 15.98 ;
    RECT 81.63 16.27 81.84 16.34 ;
    RECT 81.63 16.63 81.84 16.7 ;
    RECT 77.85 15.91 78.06 15.98 ;
    RECT 77.85 16.27 78.06 16.34 ;
    RECT 77.85 16.63 78.06 16.7 ;
    RECT 78.31 15.91 78.52 15.98 ;
    RECT 78.31 16.27 78.52 16.34 ;
    RECT 78.31 16.63 78.52 16.7 ;
    RECT 74.53 15.91 74.74 15.98 ;
    RECT 74.53 16.27 74.74 16.34 ;
    RECT 74.53 16.63 74.74 16.7 ;
    RECT 74.99 15.91 75.2 15.98 ;
    RECT 74.99 16.27 75.2 16.34 ;
    RECT 74.99 16.63 75.2 16.7 ;
    RECT 71.21 15.91 71.42 15.98 ;
    RECT 71.21 16.27 71.42 16.34 ;
    RECT 71.21 16.63 71.42 16.7 ;
    RECT 71.67 15.91 71.88 15.98 ;
    RECT 71.67 16.27 71.88 16.34 ;
    RECT 71.67 16.63 71.88 16.7 ;
    RECT 31.37 15.91 31.58 15.98 ;
    RECT 31.37 16.27 31.58 16.34 ;
    RECT 31.37 16.63 31.58 16.7 ;
    RECT 31.83 15.91 32.04 15.98 ;
    RECT 31.83 16.27 32.04 16.34 ;
    RECT 31.83 16.63 32.04 16.7 ;
    RECT 67.89 15.91 68.1 15.98 ;
    RECT 67.89 16.27 68.1 16.34 ;
    RECT 67.89 16.63 68.1 16.7 ;
    RECT 68.35 15.91 68.56 15.98 ;
    RECT 68.35 16.27 68.56 16.34 ;
    RECT 68.35 16.63 68.56 16.7 ;
    RECT 28.05 15.91 28.26 15.98 ;
    RECT 28.05 16.27 28.26 16.34 ;
    RECT 28.05 16.63 28.26 16.7 ;
    RECT 28.51 15.91 28.72 15.98 ;
    RECT 28.51 16.27 28.72 16.34 ;
    RECT 28.51 16.63 28.72 16.7 ;
    RECT 24.73 15.91 24.94 15.98 ;
    RECT 24.73 16.27 24.94 16.34 ;
    RECT 24.73 16.63 24.94 16.7 ;
    RECT 25.19 15.91 25.4 15.98 ;
    RECT 25.19 16.27 25.4 16.34 ;
    RECT 25.19 16.63 25.4 16.7 ;
    RECT 21.41 15.91 21.62 15.98 ;
    RECT 21.41 16.27 21.62 16.34 ;
    RECT 21.41 16.63 21.62 16.7 ;
    RECT 21.87 15.91 22.08 15.98 ;
    RECT 21.87 16.27 22.08 16.34 ;
    RECT 21.87 16.63 22.08 16.7 ;
    RECT 18.09 15.91 18.3 15.98 ;
    RECT 18.09 16.27 18.3 16.34 ;
    RECT 18.09 16.63 18.3 16.7 ;
    RECT 18.55 15.91 18.76 15.98 ;
    RECT 18.55 16.27 18.76 16.34 ;
    RECT 18.55 16.63 18.76 16.7 ;
    RECT 120.825 16.27 120.895 16.34 ;
    RECT 14.77 15.91 14.98 15.98 ;
    RECT 14.77 16.27 14.98 16.34 ;
    RECT 14.77 16.63 14.98 16.7 ;
    RECT 15.23 15.91 15.44 15.98 ;
    RECT 15.23 16.27 15.44 16.34 ;
    RECT 15.23 16.63 15.44 16.7 ;
    RECT 11.45 15.91 11.66 15.98 ;
    RECT 11.45 16.27 11.66 16.34 ;
    RECT 11.45 16.63 11.66 16.7 ;
    RECT 11.91 15.91 12.12 15.98 ;
    RECT 11.91 16.27 12.12 16.34 ;
    RECT 11.91 16.63 12.12 16.7 ;
    RECT 8.13 15.91 8.34 15.98 ;
    RECT 8.13 16.27 8.34 16.34 ;
    RECT 8.13 16.63 8.34 16.7 ;
    RECT 8.59 15.91 8.8 15.98 ;
    RECT 8.59 16.27 8.8 16.34 ;
    RECT 8.59 16.63 8.8 16.7 ;
    RECT 4.81 15.91 5.02 15.98 ;
    RECT 4.81 16.27 5.02 16.34 ;
    RECT 4.81 16.63 5.02 16.7 ;
    RECT 5.27 15.91 5.48 15.98 ;
    RECT 5.27 16.27 5.48 16.34 ;
    RECT 5.27 16.63 5.48 16.7 ;
    RECT 1.49 15.91 1.7 15.98 ;
    RECT 1.49 16.27 1.7 16.34 ;
    RECT 1.49 16.63 1.7 16.7 ;
    RECT 1.95 15.91 2.16 15.98 ;
    RECT 1.95 16.27 2.16 16.34 ;
    RECT 1.95 16.63 2.16 16.7 ;
    RECT 64.57 15.91 64.78 15.98 ;
    RECT 64.57 16.27 64.78 16.34 ;
    RECT 64.57 16.63 64.78 16.7 ;
    RECT 65.03 15.91 65.24 15.98 ;
    RECT 65.03 16.27 65.24 16.34 ;
    RECT 65.03 16.63 65.24 16.7 ;
    RECT 61.25 46.87 61.46 46.94 ;
    RECT 61.25 47.23 61.46 47.3 ;
    RECT 61.25 47.59 61.46 47.66 ;
    RECT 61.71 46.87 61.92 46.94 ;
    RECT 61.71 47.23 61.92 47.3 ;
    RECT 61.71 47.59 61.92 47.66 ;
    RECT 57.93 46.87 58.14 46.94 ;
    RECT 57.93 47.23 58.14 47.3 ;
    RECT 57.93 47.59 58.14 47.66 ;
    RECT 58.39 46.87 58.6 46.94 ;
    RECT 58.39 47.23 58.6 47.3 ;
    RECT 58.39 47.59 58.6 47.66 ;
    RECT 54.61 46.87 54.82 46.94 ;
    RECT 54.61 47.23 54.82 47.3 ;
    RECT 54.61 47.59 54.82 47.66 ;
    RECT 55.07 46.87 55.28 46.94 ;
    RECT 55.07 47.23 55.28 47.3 ;
    RECT 55.07 47.59 55.28 47.66 ;
    RECT 51.29 46.87 51.5 46.94 ;
    RECT 51.29 47.23 51.5 47.3 ;
    RECT 51.29 47.59 51.5 47.66 ;
    RECT 51.75 46.87 51.96 46.94 ;
    RECT 51.75 47.23 51.96 47.3 ;
    RECT 51.75 47.59 51.96 47.66 ;
    RECT 47.97 46.87 48.18 46.94 ;
    RECT 47.97 47.23 48.18 47.3 ;
    RECT 47.97 47.59 48.18 47.66 ;
    RECT 48.43 46.87 48.64 46.94 ;
    RECT 48.43 47.23 48.64 47.3 ;
    RECT 48.43 47.59 48.64 47.66 ;
    RECT 44.65 46.87 44.86 46.94 ;
    RECT 44.65 47.23 44.86 47.3 ;
    RECT 44.65 47.59 44.86 47.66 ;
    RECT 45.11 46.87 45.32 46.94 ;
    RECT 45.11 47.23 45.32 47.3 ;
    RECT 45.11 47.59 45.32 47.66 ;
    RECT 41.33 46.87 41.54 46.94 ;
    RECT 41.33 47.23 41.54 47.3 ;
    RECT 41.33 47.59 41.54 47.66 ;
    RECT 41.79 46.87 42.0 46.94 ;
    RECT 41.79 47.23 42.0 47.3 ;
    RECT 41.79 47.59 42.0 47.66 ;
    RECT 38.01 46.87 38.22 46.94 ;
    RECT 38.01 47.23 38.22 47.3 ;
    RECT 38.01 47.59 38.22 47.66 ;
    RECT 38.47 46.87 38.68 46.94 ;
    RECT 38.47 47.23 38.68 47.3 ;
    RECT 38.47 47.59 38.68 47.66 ;
    RECT 0.4 47.23 0.47 47.3 ;
    RECT 34.69 46.87 34.9 46.94 ;
    RECT 34.69 47.23 34.9 47.3 ;
    RECT 34.69 47.59 34.9 47.66 ;
    RECT 35.15 46.87 35.36 46.94 ;
    RECT 35.15 47.23 35.36 47.3 ;
    RECT 35.15 47.59 35.36 47.66 ;
    RECT 117.69 46.87 117.9 46.94 ;
    RECT 117.69 47.23 117.9 47.3 ;
    RECT 117.69 47.59 117.9 47.66 ;
    RECT 118.15 46.87 118.36 46.94 ;
    RECT 118.15 47.23 118.36 47.3 ;
    RECT 118.15 47.59 118.36 47.66 ;
    RECT 114.37 46.87 114.58 46.94 ;
    RECT 114.37 47.23 114.58 47.3 ;
    RECT 114.37 47.59 114.58 47.66 ;
    RECT 114.83 46.87 115.04 46.94 ;
    RECT 114.83 47.23 115.04 47.3 ;
    RECT 114.83 47.59 115.04 47.66 ;
    RECT 111.05 46.87 111.26 46.94 ;
    RECT 111.05 47.23 111.26 47.3 ;
    RECT 111.05 47.59 111.26 47.66 ;
    RECT 111.51 46.87 111.72 46.94 ;
    RECT 111.51 47.23 111.72 47.3 ;
    RECT 111.51 47.59 111.72 47.66 ;
    RECT 107.73 46.87 107.94 46.94 ;
    RECT 107.73 47.23 107.94 47.3 ;
    RECT 107.73 47.59 107.94 47.66 ;
    RECT 108.19 46.87 108.4 46.94 ;
    RECT 108.19 47.23 108.4 47.3 ;
    RECT 108.19 47.59 108.4 47.66 ;
    RECT 104.41 46.87 104.62 46.94 ;
    RECT 104.41 47.23 104.62 47.3 ;
    RECT 104.41 47.59 104.62 47.66 ;
    RECT 104.87 46.87 105.08 46.94 ;
    RECT 104.87 47.23 105.08 47.3 ;
    RECT 104.87 47.59 105.08 47.66 ;
    RECT 101.09 46.87 101.3 46.94 ;
    RECT 101.09 47.23 101.3 47.3 ;
    RECT 101.09 47.59 101.3 47.66 ;
    RECT 101.55 46.87 101.76 46.94 ;
    RECT 101.55 47.23 101.76 47.3 ;
    RECT 101.55 47.59 101.76 47.66 ;
    RECT 97.77 46.87 97.98 46.94 ;
    RECT 97.77 47.23 97.98 47.3 ;
    RECT 97.77 47.59 97.98 47.66 ;
    RECT 98.23 46.87 98.44 46.94 ;
    RECT 98.23 47.23 98.44 47.3 ;
    RECT 98.23 47.59 98.44 47.66 ;
    RECT 94.45 46.87 94.66 46.94 ;
    RECT 94.45 47.23 94.66 47.3 ;
    RECT 94.45 47.59 94.66 47.66 ;
    RECT 94.91 46.87 95.12 46.94 ;
    RECT 94.91 47.23 95.12 47.3 ;
    RECT 94.91 47.59 95.12 47.66 ;
    RECT 91.13 46.87 91.34 46.94 ;
    RECT 91.13 47.23 91.34 47.3 ;
    RECT 91.13 47.59 91.34 47.66 ;
    RECT 91.59 46.87 91.8 46.94 ;
    RECT 91.59 47.23 91.8 47.3 ;
    RECT 91.59 47.59 91.8 47.66 ;
    RECT 87.81 46.87 88.02 46.94 ;
    RECT 87.81 47.23 88.02 47.3 ;
    RECT 87.81 47.59 88.02 47.66 ;
    RECT 88.27 46.87 88.48 46.94 ;
    RECT 88.27 47.23 88.48 47.3 ;
    RECT 88.27 47.59 88.48 47.66 ;
    RECT 84.49 46.87 84.7 46.94 ;
    RECT 84.49 47.23 84.7 47.3 ;
    RECT 84.49 47.59 84.7 47.66 ;
    RECT 84.95 46.87 85.16 46.94 ;
    RECT 84.95 47.23 85.16 47.3 ;
    RECT 84.95 47.59 85.16 47.66 ;
    RECT 81.17 46.87 81.38 46.94 ;
    RECT 81.17 47.23 81.38 47.3 ;
    RECT 81.17 47.59 81.38 47.66 ;
    RECT 81.63 46.87 81.84 46.94 ;
    RECT 81.63 47.23 81.84 47.3 ;
    RECT 81.63 47.59 81.84 47.66 ;
    RECT 77.85 46.87 78.06 46.94 ;
    RECT 77.85 47.23 78.06 47.3 ;
    RECT 77.85 47.59 78.06 47.66 ;
    RECT 78.31 46.87 78.52 46.94 ;
    RECT 78.31 47.23 78.52 47.3 ;
    RECT 78.31 47.59 78.52 47.66 ;
    RECT 74.53 46.87 74.74 46.94 ;
    RECT 74.53 47.23 74.74 47.3 ;
    RECT 74.53 47.59 74.74 47.66 ;
    RECT 74.99 46.87 75.2 46.94 ;
    RECT 74.99 47.23 75.2 47.3 ;
    RECT 74.99 47.59 75.2 47.66 ;
    RECT 71.21 46.87 71.42 46.94 ;
    RECT 71.21 47.23 71.42 47.3 ;
    RECT 71.21 47.59 71.42 47.66 ;
    RECT 71.67 46.87 71.88 46.94 ;
    RECT 71.67 47.23 71.88 47.3 ;
    RECT 71.67 47.59 71.88 47.66 ;
    RECT 31.37 46.87 31.58 46.94 ;
    RECT 31.37 47.23 31.58 47.3 ;
    RECT 31.37 47.59 31.58 47.66 ;
    RECT 31.83 46.87 32.04 46.94 ;
    RECT 31.83 47.23 32.04 47.3 ;
    RECT 31.83 47.59 32.04 47.66 ;
    RECT 67.89 46.87 68.1 46.94 ;
    RECT 67.89 47.23 68.1 47.3 ;
    RECT 67.89 47.59 68.1 47.66 ;
    RECT 68.35 46.87 68.56 46.94 ;
    RECT 68.35 47.23 68.56 47.3 ;
    RECT 68.35 47.59 68.56 47.66 ;
    RECT 28.05 46.87 28.26 46.94 ;
    RECT 28.05 47.23 28.26 47.3 ;
    RECT 28.05 47.59 28.26 47.66 ;
    RECT 28.51 46.87 28.72 46.94 ;
    RECT 28.51 47.23 28.72 47.3 ;
    RECT 28.51 47.59 28.72 47.66 ;
    RECT 24.73 46.87 24.94 46.94 ;
    RECT 24.73 47.23 24.94 47.3 ;
    RECT 24.73 47.59 24.94 47.66 ;
    RECT 25.19 46.87 25.4 46.94 ;
    RECT 25.19 47.23 25.4 47.3 ;
    RECT 25.19 47.59 25.4 47.66 ;
    RECT 21.41 46.87 21.62 46.94 ;
    RECT 21.41 47.23 21.62 47.3 ;
    RECT 21.41 47.59 21.62 47.66 ;
    RECT 21.87 46.87 22.08 46.94 ;
    RECT 21.87 47.23 22.08 47.3 ;
    RECT 21.87 47.59 22.08 47.66 ;
    RECT 18.09 46.87 18.3 46.94 ;
    RECT 18.09 47.23 18.3 47.3 ;
    RECT 18.09 47.59 18.3 47.66 ;
    RECT 18.55 46.87 18.76 46.94 ;
    RECT 18.55 47.23 18.76 47.3 ;
    RECT 18.55 47.59 18.76 47.66 ;
    RECT 120.825 47.23 120.895 47.3 ;
    RECT 14.77 46.87 14.98 46.94 ;
    RECT 14.77 47.23 14.98 47.3 ;
    RECT 14.77 47.59 14.98 47.66 ;
    RECT 15.23 46.87 15.44 46.94 ;
    RECT 15.23 47.23 15.44 47.3 ;
    RECT 15.23 47.59 15.44 47.66 ;
    RECT 11.45 46.87 11.66 46.94 ;
    RECT 11.45 47.23 11.66 47.3 ;
    RECT 11.45 47.59 11.66 47.66 ;
    RECT 11.91 46.87 12.12 46.94 ;
    RECT 11.91 47.23 12.12 47.3 ;
    RECT 11.91 47.59 12.12 47.66 ;
    RECT 8.13 46.87 8.34 46.94 ;
    RECT 8.13 47.23 8.34 47.3 ;
    RECT 8.13 47.59 8.34 47.66 ;
    RECT 8.59 46.87 8.8 46.94 ;
    RECT 8.59 47.23 8.8 47.3 ;
    RECT 8.59 47.59 8.8 47.66 ;
    RECT 4.81 46.87 5.02 46.94 ;
    RECT 4.81 47.23 5.02 47.3 ;
    RECT 4.81 47.59 5.02 47.66 ;
    RECT 5.27 46.87 5.48 46.94 ;
    RECT 5.27 47.23 5.48 47.3 ;
    RECT 5.27 47.59 5.48 47.66 ;
    RECT 1.49 46.87 1.7 46.94 ;
    RECT 1.49 47.23 1.7 47.3 ;
    RECT 1.49 47.59 1.7 47.66 ;
    RECT 1.95 46.87 2.16 46.94 ;
    RECT 1.95 47.23 2.16 47.3 ;
    RECT 1.95 47.59 2.16 47.66 ;
    RECT 64.57 46.87 64.78 46.94 ;
    RECT 64.57 47.23 64.78 47.3 ;
    RECT 64.57 47.59 64.78 47.66 ;
    RECT 65.03 46.87 65.24 46.94 ;
    RECT 65.03 47.23 65.24 47.3 ;
    RECT 65.03 47.59 65.24 47.66 ;
    RECT 61.25 86.49 61.46 86.56 ;
    RECT 61.25 86.85 61.46 86.92 ;
    RECT 61.25 87.21 61.46 87.28 ;
    RECT 61.71 86.49 61.92 86.56 ;
    RECT 61.71 86.85 61.92 86.92 ;
    RECT 61.71 87.21 61.92 87.28 ;
    RECT 57.93 86.49 58.14 86.56 ;
    RECT 57.93 86.85 58.14 86.92 ;
    RECT 57.93 87.21 58.14 87.28 ;
    RECT 58.39 86.49 58.6 86.56 ;
    RECT 58.39 86.85 58.6 86.92 ;
    RECT 58.39 87.21 58.6 87.28 ;
    RECT 54.61 86.49 54.82 86.56 ;
    RECT 54.61 86.85 54.82 86.92 ;
    RECT 54.61 87.21 54.82 87.28 ;
    RECT 55.07 86.49 55.28 86.56 ;
    RECT 55.07 86.85 55.28 86.92 ;
    RECT 55.07 87.21 55.28 87.28 ;
    RECT 51.29 86.49 51.5 86.56 ;
    RECT 51.29 86.85 51.5 86.92 ;
    RECT 51.29 87.21 51.5 87.28 ;
    RECT 51.75 86.49 51.96 86.56 ;
    RECT 51.75 86.85 51.96 86.92 ;
    RECT 51.75 87.21 51.96 87.28 ;
    RECT 47.97 86.49 48.18 86.56 ;
    RECT 47.97 86.85 48.18 86.92 ;
    RECT 47.97 87.21 48.18 87.28 ;
    RECT 48.43 86.49 48.64 86.56 ;
    RECT 48.43 86.85 48.64 86.92 ;
    RECT 48.43 87.21 48.64 87.28 ;
    RECT 44.65 86.49 44.86 86.56 ;
    RECT 44.65 86.85 44.86 86.92 ;
    RECT 44.65 87.21 44.86 87.28 ;
    RECT 45.11 86.49 45.32 86.56 ;
    RECT 45.11 86.85 45.32 86.92 ;
    RECT 45.11 87.21 45.32 87.28 ;
    RECT 41.33 86.49 41.54 86.56 ;
    RECT 41.33 86.85 41.54 86.92 ;
    RECT 41.33 87.21 41.54 87.28 ;
    RECT 41.79 86.49 42.0 86.56 ;
    RECT 41.79 86.85 42.0 86.92 ;
    RECT 41.79 87.21 42.0 87.28 ;
    RECT 38.01 86.49 38.22 86.56 ;
    RECT 38.01 86.85 38.22 86.92 ;
    RECT 38.01 87.21 38.22 87.28 ;
    RECT 38.47 86.49 38.68 86.56 ;
    RECT 38.47 86.85 38.68 86.92 ;
    RECT 38.47 87.21 38.68 87.28 ;
    RECT 0.4 86.85 0.47 86.92 ;
    RECT 34.69 86.49 34.9 86.56 ;
    RECT 34.69 86.85 34.9 86.92 ;
    RECT 34.69 87.21 34.9 87.28 ;
    RECT 35.15 86.49 35.36 86.56 ;
    RECT 35.15 86.85 35.36 86.92 ;
    RECT 35.15 87.21 35.36 87.28 ;
    RECT 117.69 86.49 117.9 86.56 ;
    RECT 117.69 86.85 117.9 86.92 ;
    RECT 117.69 87.21 117.9 87.28 ;
    RECT 118.15 86.49 118.36 86.56 ;
    RECT 118.15 86.85 118.36 86.92 ;
    RECT 118.15 87.21 118.36 87.28 ;
    RECT 114.37 86.49 114.58 86.56 ;
    RECT 114.37 86.85 114.58 86.92 ;
    RECT 114.37 87.21 114.58 87.28 ;
    RECT 114.83 86.49 115.04 86.56 ;
    RECT 114.83 86.85 115.04 86.92 ;
    RECT 114.83 87.21 115.04 87.28 ;
    RECT 111.05 86.49 111.26 86.56 ;
    RECT 111.05 86.85 111.26 86.92 ;
    RECT 111.05 87.21 111.26 87.28 ;
    RECT 111.51 86.49 111.72 86.56 ;
    RECT 111.51 86.85 111.72 86.92 ;
    RECT 111.51 87.21 111.72 87.28 ;
    RECT 107.73 86.49 107.94 86.56 ;
    RECT 107.73 86.85 107.94 86.92 ;
    RECT 107.73 87.21 107.94 87.28 ;
    RECT 108.19 86.49 108.4 86.56 ;
    RECT 108.19 86.85 108.4 86.92 ;
    RECT 108.19 87.21 108.4 87.28 ;
    RECT 104.41 86.49 104.62 86.56 ;
    RECT 104.41 86.85 104.62 86.92 ;
    RECT 104.41 87.21 104.62 87.28 ;
    RECT 104.87 86.49 105.08 86.56 ;
    RECT 104.87 86.85 105.08 86.92 ;
    RECT 104.87 87.21 105.08 87.28 ;
    RECT 101.09 86.49 101.3 86.56 ;
    RECT 101.09 86.85 101.3 86.92 ;
    RECT 101.09 87.21 101.3 87.28 ;
    RECT 101.55 86.49 101.76 86.56 ;
    RECT 101.55 86.85 101.76 86.92 ;
    RECT 101.55 87.21 101.76 87.28 ;
    RECT 97.77 86.49 97.98 86.56 ;
    RECT 97.77 86.85 97.98 86.92 ;
    RECT 97.77 87.21 97.98 87.28 ;
    RECT 98.23 86.49 98.44 86.56 ;
    RECT 98.23 86.85 98.44 86.92 ;
    RECT 98.23 87.21 98.44 87.28 ;
    RECT 94.45 86.49 94.66 86.56 ;
    RECT 94.45 86.85 94.66 86.92 ;
    RECT 94.45 87.21 94.66 87.28 ;
    RECT 94.91 86.49 95.12 86.56 ;
    RECT 94.91 86.85 95.12 86.92 ;
    RECT 94.91 87.21 95.12 87.28 ;
    RECT 91.13 86.49 91.34 86.56 ;
    RECT 91.13 86.85 91.34 86.92 ;
    RECT 91.13 87.21 91.34 87.28 ;
    RECT 91.59 86.49 91.8 86.56 ;
    RECT 91.59 86.85 91.8 86.92 ;
    RECT 91.59 87.21 91.8 87.28 ;
    RECT 87.81 86.49 88.02 86.56 ;
    RECT 87.81 86.85 88.02 86.92 ;
    RECT 87.81 87.21 88.02 87.28 ;
    RECT 88.27 86.49 88.48 86.56 ;
    RECT 88.27 86.85 88.48 86.92 ;
    RECT 88.27 87.21 88.48 87.28 ;
    RECT 84.49 86.49 84.7 86.56 ;
    RECT 84.49 86.85 84.7 86.92 ;
    RECT 84.49 87.21 84.7 87.28 ;
    RECT 84.95 86.49 85.16 86.56 ;
    RECT 84.95 86.85 85.16 86.92 ;
    RECT 84.95 87.21 85.16 87.28 ;
    RECT 81.17 86.49 81.38 86.56 ;
    RECT 81.17 86.85 81.38 86.92 ;
    RECT 81.17 87.21 81.38 87.28 ;
    RECT 81.63 86.49 81.84 86.56 ;
    RECT 81.63 86.85 81.84 86.92 ;
    RECT 81.63 87.21 81.84 87.28 ;
    RECT 77.85 86.49 78.06 86.56 ;
    RECT 77.85 86.85 78.06 86.92 ;
    RECT 77.85 87.21 78.06 87.28 ;
    RECT 78.31 86.49 78.52 86.56 ;
    RECT 78.31 86.85 78.52 86.92 ;
    RECT 78.31 87.21 78.52 87.28 ;
    RECT 74.53 86.49 74.74 86.56 ;
    RECT 74.53 86.85 74.74 86.92 ;
    RECT 74.53 87.21 74.74 87.28 ;
    RECT 74.99 86.49 75.2 86.56 ;
    RECT 74.99 86.85 75.2 86.92 ;
    RECT 74.99 87.21 75.2 87.28 ;
    RECT 71.21 86.49 71.42 86.56 ;
    RECT 71.21 86.85 71.42 86.92 ;
    RECT 71.21 87.21 71.42 87.28 ;
    RECT 71.67 86.49 71.88 86.56 ;
    RECT 71.67 86.85 71.88 86.92 ;
    RECT 71.67 87.21 71.88 87.28 ;
    RECT 31.37 86.49 31.58 86.56 ;
    RECT 31.37 86.85 31.58 86.92 ;
    RECT 31.37 87.21 31.58 87.28 ;
    RECT 31.83 86.49 32.04 86.56 ;
    RECT 31.83 86.85 32.04 86.92 ;
    RECT 31.83 87.21 32.04 87.28 ;
    RECT 67.89 86.49 68.1 86.56 ;
    RECT 67.89 86.85 68.1 86.92 ;
    RECT 67.89 87.21 68.1 87.28 ;
    RECT 68.35 86.49 68.56 86.56 ;
    RECT 68.35 86.85 68.56 86.92 ;
    RECT 68.35 87.21 68.56 87.28 ;
    RECT 28.05 86.49 28.26 86.56 ;
    RECT 28.05 86.85 28.26 86.92 ;
    RECT 28.05 87.21 28.26 87.28 ;
    RECT 28.51 86.49 28.72 86.56 ;
    RECT 28.51 86.85 28.72 86.92 ;
    RECT 28.51 87.21 28.72 87.28 ;
    RECT 24.73 86.49 24.94 86.56 ;
    RECT 24.73 86.85 24.94 86.92 ;
    RECT 24.73 87.21 24.94 87.28 ;
    RECT 25.19 86.49 25.4 86.56 ;
    RECT 25.19 86.85 25.4 86.92 ;
    RECT 25.19 87.21 25.4 87.28 ;
    RECT 21.41 86.49 21.62 86.56 ;
    RECT 21.41 86.85 21.62 86.92 ;
    RECT 21.41 87.21 21.62 87.28 ;
    RECT 21.87 86.49 22.08 86.56 ;
    RECT 21.87 86.85 22.08 86.92 ;
    RECT 21.87 87.21 22.08 87.28 ;
    RECT 18.09 86.49 18.3 86.56 ;
    RECT 18.09 86.85 18.3 86.92 ;
    RECT 18.09 87.21 18.3 87.28 ;
    RECT 18.55 86.49 18.76 86.56 ;
    RECT 18.55 86.85 18.76 86.92 ;
    RECT 18.55 87.21 18.76 87.28 ;
    RECT 120.825 86.85 120.895 86.92 ;
    RECT 14.77 86.49 14.98 86.56 ;
    RECT 14.77 86.85 14.98 86.92 ;
    RECT 14.77 87.21 14.98 87.28 ;
    RECT 15.23 86.49 15.44 86.56 ;
    RECT 15.23 86.85 15.44 86.92 ;
    RECT 15.23 87.21 15.44 87.28 ;
    RECT 11.45 86.49 11.66 86.56 ;
    RECT 11.45 86.85 11.66 86.92 ;
    RECT 11.45 87.21 11.66 87.28 ;
    RECT 11.91 86.49 12.12 86.56 ;
    RECT 11.91 86.85 12.12 86.92 ;
    RECT 11.91 87.21 12.12 87.28 ;
    RECT 8.13 86.49 8.34 86.56 ;
    RECT 8.13 86.85 8.34 86.92 ;
    RECT 8.13 87.21 8.34 87.28 ;
    RECT 8.59 86.49 8.8 86.56 ;
    RECT 8.59 86.85 8.8 86.92 ;
    RECT 8.59 87.21 8.8 87.28 ;
    RECT 4.81 86.49 5.02 86.56 ;
    RECT 4.81 86.85 5.02 86.92 ;
    RECT 4.81 87.21 5.02 87.28 ;
    RECT 5.27 86.49 5.48 86.56 ;
    RECT 5.27 86.85 5.48 86.92 ;
    RECT 5.27 87.21 5.48 87.28 ;
    RECT 1.49 86.49 1.7 86.56 ;
    RECT 1.49 86.85 1.7 86.92 ;
    RECT 1.49 87.21 1.7 87.28 ;
    RECT 1.95 86.49 2.16 86.56 ;
    RECT 1.95 86.85 2.16 86.92 ;
    RECT 1.95 87.21 2.16 87.28 ;
    RECT 64.57 86.49 64.78 86.56 ;
    RECT 64.57 86.85 64.78 86.92 ;
    RECT 64.57 87.21 64.78 87.28 ;
    RECT 65.03 86.49 65.24 86.56 ;
    RECT 65.03 86.85 65.24 86.92 ;
    RECT 65.03 87.21 65.24 87.28 ;
    RECT 61.25 15.19 61.46 15.26 ;
    RECT 61.25 15.55 61.46 15.62 ;
    RECT 61.25 15.91 61.46 15.98 ;
    RECT 61.71 15.19 61.92 15.26 ;
    RECT 61.71 15.55 61.92 15.62 ;
    RECT 61.71 15.91 61.92 15.98 ;
    RECT 57.93 15.19 58.14 15.26 ;
    RECT 57.93 15.55 58.14 15.62 ;
    RECT 57.93 15.91 58.14 15.98 ;
    RECT 58.39 15.19 58.6 15.26 ;
    RECT 58.39 15.55 58.6 15.62 ;
    RECT 58.39 15.91 58.6 15.98 ;
    RECT 54.61 15.19 54.82 15.26 ;
    RECT 54.61 15.55 54.82 15.62 ;
    RECT 54.61 15.91 54.82 15.98 ;
    RECT 55.07 15.19 55.28 15.26 ;
    RECT 55.07 15.55 55.28 15.62 ;
    RECT 55.07 15.91 55.28 15.98 ;
    RECT 51.29 15.19 51.5 15.26 ;
    RECT 51.29 15.55 51.5 15.62 ;
    RECT 51.29 15.91 51.5 15.98 ;
    RECT 51.75 15.19 51.96 15.26 ;
    RECT 51.75 15.55 51.96 15.62 ;
    RECT 51.75 15.91 51.96 15.98 ;
    RECT 47.97 15.19 48.18 15.26 ;
    RECT 47.97 15.55 48.18 15.62 ;
    RECT 47.97 15.91 48.18 15.98 ;
    RECT 48.43 15.19 48.64 15.26 ;
    RECT 48.43 15.55 48.64 15.62 ;
    RECT 48.43 15.91 48.64 15.98 ;
    RECT 44.65 15.19 44.86 15.26 ;
    RECT 44.65 15.55 44.86 15.62 ;
    RECT 44.65 15.91 44.86 15.98 ;
    RECT 45.11 15.19 45.32 15.26 ;
    RECT 45.11 15.55 45.32 15.62 ;
    RECT 45.11 15.91 45.32 15.98 ;
    RECT 41.33 15.19 41.54 15.26 ;
    RECT 41.33 15.55 41.54 15.62 ;
    RECT 41.33 15.91 41.54 15.98 ;
    RECT 41.79 15.19 42.0 15.26 ;
    RECT 41.79 15.55 42.0 15.62 ;
    RECT 41.79 15.91 42.0 15.98 ;
    RECT 38.01 15.19 38.22 15.26 ;
    RECT 38.01 15.55 38.22 15.62 ;
    RECT 38.01 15.91 38.22 15.98 ;
    RECT 38.47 15.19 38.68 15.26 ;
    RECT 38.47 15.55 38.68 15.62 ;
    RECT 38.47 15.91 38.68 15.98 ;
    RECT 0.4 15.55 0.47 15.62 ;
    RECT 34.69 15.19 34.9 15.26 ;
    RECT 34.69 15.55 34.9 15.62 ;
    RECT 34.69 15.91 34.9 15.98 ;
    RECT 35.15 15.19 35.36 15.26 ;
    RECT 35.15 15.55 35.36 15.62 ;
    RECT 35.15 15.91 35.36 15.98 ;
    RECT 117.69 15.19 117.9 15.26 ;
    RECT 117.69 15.55 117.9 15.62 ;
    RECT 117.69 15.91 117.9 15.98 ;
    RECT 118.15 15.19 118.36 15.26 ;
    RECT 118.15 15.55 118.36 15.62 ;
    RECT 118.15 15.91 118.36 15.98 ;
    RECT 114.37 15.19 114.58 15.26 ;
    RECT 114.37 15.55 114.58 15.62 ;
    RECT 114.37 15.91 114.58 15.98 ;
    RECT 114.83 15.19 115.04 15.26 ;
    RECT 114.83 15.55 115.04 15.62 ;
    RECT 114.83 15.91 115.04 15.98 ;
    RECT 111.05 15.19 111.26 15.26 ;
    RECT 111.05 15.55 111.26 15.62 ;
    RECT 111.05 15.91 111.26 15.98 ;
    RECT 111.51 15.19 111.72 15.26 ;
    RECT 111.51 15.55 111.72 15.62 ;
    RECT 111.51 15.91 111.72 15.98 ;
    RECT 107.73 15.19 107.94 15.26 ;
    RECT 107.73 15.55 107.94 15.62 ;
    RECT 107.73 15.91 107.94 15.98 ;
    RECT 108.19 15.19 108.4 15.26 ;
    RECT 108.19 15.55 108.4 15.62 ;
    RECT 108.19 15.91 108.4 15.98 ;
    RECT 104.41 15.19 104.62 15.26 ;
    RECT 104.41 15.55 104.62 15.62 ;
    RECT 104.41 15.91 104.62 15.98 ;
    RECT 104.87 15.19 105.08 15.26 ;
    RECT 104.87 15.55 105.08 15.62 ;
    RECT 104.87 15.91 105.08 15.98 ;
    RECT 101.09 15.19 101.3 15.26 ;
    RECT 101.09 15.55 101.3 15.62 ;
    RECT 101.09 15.91 101.3 15.98 ;
    RECT 101.55 15.19 101.76 15.26 ;
    RECT 101.55 15.55 101.76 15.62 ;
    RECT 101.55 15.91 101.76 15.98 ;
    RECT 97.77 15.19 97.98 15.26 ;
    RECT 97.77 15.55 97.98 15.62 ;
    RECT 97.77 15.91 97.98 15.98 ;
    RECT 98.23 15.19 98.44 15.26 ;
    RECT 98.23 15.55 98.44 15.62 ;
    RECT 98.23 15.91 98.44 15.98 ;
    RECT 94.45 15.19 94.66 15.26 ;
    RECT 94.45 15.55 94.66 15.62 ;
    RECT 94.45 15.91 94.66 15.98 ;
    RECT 94.91 15.19 95.12 15.26 ;
    RECT 94.91 15.55 95.12 15.62 ;
    RECT 94.91 15.91 95.12 15.98 ;
    RECT 91.13 15.19 91.34 15.26 ;
    RECT 91.13 15.55 91.34 15.62 ;
    RECT 91.13 15.91 91.34 15.98 ;
    RECT 91.59 15.19 91.8 15.26 ;
    RECT 91.59 15.55 91.8 15.62 ;
    RECT 91.59 15.91 91.8 15.98 ;
    RECT 87.81 15.19 88.02 15.26 ;
    RECT 87.81 15.55 88.02 15.62 ;
    RECT 87.81 15.91 88.02 15.98 ;
    RECT 88.27 15.19 88.48 15.26 ;
    RECT 88.27 15.55 88.48 15.62 ;
    RECT 88.27 15.91 88.48 15.98 ;
    RECT 84.49 15.19 84.7 15.26 ;
    RECT 84.49 15.55 84.7 15.62 ;
    RECT 84.49 15.91 84.7 15.98 ;
    RECT 84.95 15.19 85.16 15.26 ;
    RECT 84.95 15.55 85.16 15.62 ;
    RECT 84.95 15.91 85.16 15.98 ;
    RECT 81.17 15.19 81.38 15.26 ;
    RECT 81.17 15.55 81.38 15.62 ;
    RECT 81.17 15.91 81.38 15.98 ;
    RECT 81.63 15.19 81.84 15.26 ;
    RECT 81.63 15.55 81.84 15.62 ;
    RECT 81.63 15.91 81.84 15.98 ;
    RECT 77.85 15.19 78.06 15.26 ;
    RECT 77.85 15.55 78.06 15.62 ;
    RECT 77.85 15.91 78.06 15.98 ;
    RECT 78.31 15.19 78.52 15.26 ;
    RECT 78.31 15.55 78.52 15.62 ;
    RECT 78.31 15.91 78.52 15.98 ;
    RECT 74.53 15.19 74.74 15.26 ;
    RECT 74.53 15.55 74.74 15.62 ;
    RECT 74.53 15.91 74.74 15.98 ;
    RECT 74.99 15.19 75.2 15.26 ;
    RECT 74.99 15.55 75.2 15.62 ;
    RECT 74.99 15.91 75.2 15.98 ;
    RECT 71.21 15.19 71.42 15.26 ;
    RECT 71.21 15.55 71.42 15.62 ;
    RECT 71.21 15.91 71.42 15.98 ;
    RECT 71.67 15.19 71.88 15.26 ;
    RECT 71.67 15.55 71.88 15.62 ;
    RECT 71.67 15.91 71.88 15.98 ;
    RECT 31.37 15.19 31.58 15.26 ;
    RECT 31.37 15.55 31.58 15.62 ;
    RECT 31.37 15.91 31.58 15.98 ;
    RECT 31.83 15.19 32.04 15.26 ;
    RECT 31.83 15.55 32.04 15.62 ;
    RECT 31.83 15.91 32.04 15.98 ;
    RECT 67.89 15.19 68.1 15.26 ;
    RECT 67.89 15.55 68.1 15.62 ;
    RECT 67.89 15.91 68.1 15.98 ;
    RECT 68.35 15.19 68.56 15.26 ;
    RECT 68.35 15.55 68.56 15.62 ;
    RECT 68.35 15.91 68.56 15.98 ;
    RECT 28.05 15.19 28.26 15.26 ;
    RECT 28.05 15.55 28.26 15.62 ;
    RECT 28.05 15.91 28.26 15.98 ;
    RECT 28.51 15.19 28.72 15.26 ;
    RECT 28.51 15.55 28.72 15.62 ;
    RECT 28.51 15.91 28.72 15.98 ;
    RECT 24.73 15.19 24.94 15.26 ;
    RECT 24.73 15.55 24.94 15.62 ;
    RECT 24.73 15.91 24.94 15.98 ;
    RECT 25.19 15.19 25.4 15.26 ;
    RECT 25.19 15.55 25.4 15.62 ;
    RECT 25.19 15.91 25.4 15.98 ;
    RECT 21.41 15.19 21.62 15.26 ;
    RECT 21.41 15.55 21.62 15.62 ;
    RECT 21.41 15.91 21.62 15.98 ;
    RECT 21.87 15.19 22.08 15.26 ;
    RECT 21.87 15.55 22.08 15.62 ;
    RECT 21.87 15.91 22.08 15.98 ;
    RECT 18.09 15.19 18.3 15.26 ;
    RECT 18.09 15.55 18.3 15.62 ;
    RECT 18.09 15.91 18.3 15.98 ;
    RECT 18.55 15.19 18.76 15.26 ;
    RECT 18.55 15.55 18.76 15.62 ;
    RECT 18.55 15.91 18.76 15.98 ;
    RECT 120.825 15.55 120.895 15.62 ;
    RECT 14.77 15.19 14.98 15.26 ;
    RECT 14.77 15.55 14.98 15.62 ;
    RECT 14.77 15.91 14.98 15.98 ;
    RECT 15.23 15.19 15.44 15.26 ;
    RECT 15.23 15.55 15.44 15.62 ;
    RECT 15.23 15.91 15.44 15.98 ;
    RECT 11.45 15.19 11.66 15.26 ;
    RECT 11.45 15.55 11.66 15.62 ;
    RECT 11.45 15.91 11.66 15.98 ;
    RECT 11.91 15.19 12.12 15.26 ;
    RECT 11.91 15.55 12.12 15.62 ;
    RECT 11.91 15.91 12.12 15.98 ;
    RECT 8.13 15.19 8.34 15.26 ;
    RECT 8.13 15.55 8.34 15.62 ;
    RECT 8.13 15.91 8.34 15.98 ;
    RECT 8.59 15.19 8.8 15.26 ;
    RECT 8.59 15.55 8.8 15.62 ;
    RECT 8.59 15.91 8.8 15.98 ;
    RECT 4.81 15.19 5.02 15.26 ;
    RECT 4.81 15.55 5.02 15.62 ;
    RECT 4.81 15.91 5.02 15.98 ;
    RECT 5.27 15.19 5.48 15.26 ;
    RECT 5.27 15.55 5.48 15.62 ;
    RECT 5.27 15.91 5.48 15.98 ;
    RECT 1.49 15.19 1.7 15.26 ;
    RECT 1.49 15.55 1.7 15.62 ;
    RECT 1.49 15.91 1.7 15.98 ;
    RECT 1.95 15.19 2.16 15.26 ;
    RECT 1.95 15.55 2.16 15.62 ;
    RECT 1.95 15.91 2.16 15.98 ;
    RECT 64.57 15.19 64.78 15.26 ;
    RECT 64.57 15.55 64.78 15.62 ;
    RECT 64.57 15.91 64.78 15.98 ;
    RECT 65.03 15.19 65.24 15.26 ;
    RECT 65.03 15.55 65.24 15.62 ;
    RECT 65.03 15.91 65.24 15.98 ;
    RECT 61.25 46.15 61.46 46.22 ;
    RECT 61.25 46.51 61.46 46.58 ;
    RECT 61.25 46.87 61.46 46.94 ;
    RECT 61.71 46.15 61.92 46.22 ;
    RECT 61.71 46.51 61.92 46.58 ;
    RECT 61.71 46.87 61.92 46.94 ;
    RECT 57.93 46.15 58.14 46.22 ;
    RECT 57.93 46.51 58.14 46.58 ;
    RECT 57.93 46.87 58.14 46.94 ;
    RECT 58.39 46.15 58.6 46.22 ;
    RECT 58.39 46.51 58.6 46.58 ;
    RECT 58.39 46.87 58.6 46.94 ;
    RECT 54.61 46.15 54.82 46.22 ;
    RECT 54.61 46.51 54.82 46.58 ;
    RECT 54.61 46.87 54.82 46.94 ;
    RECT 55.07 46.15 55.28 46.22 ;
    RECT 55.07 46.51 55.28 46.58 ;
    RECT 55.07 46.87 55.28 46.94 ;
    RECT 51.29 46.15 51.5 46.22 ;
    RECT 51.29 46.51 51.5 46.58 ;
    RECT 51.29 46.87 51.5 46.94 ;
    RECT 51.75 46.15 51.96 46.22 ;
    RECT 51.75 46.51 51.96 46.58 ;
    RECT 51.75 46.87 51.96 46.94 ;
    RECT 47.97 46.15 48.18 46.22 ;
    RECT 47.97 46.51 48.18 46.58 ;
    RECT 47.97 46.87 48.18 46.94 ;
    RECT 48.43 46.15 48.64 46.22 ;
    RECT 48.43 46.51 48.64 46.58 ;
    RECT 48.43 46.87 48.64 46.94 ;
    RECT 44.65 46.15 44.86 46.22 ;
    RECT 44.65 46.51 44.86 46.58 ;
    RECT 44.65 46.87 44.86 46.94 ;
    RECT 45.11 46.15 45.32 46.22 ;
    RECT 45.11 46.51 45.32 46.58 ;
    RECT 45.11 46.87 45.32 46.94 ;
    RECT 41.33 46.15 41.54 46.22 ;
    RECT 41.33 46.51 41.54 46.58 ;
    RECT 41.33 46.87 41.54 46.94 ;
    RECT 41.79 46.15 42.0 46.22 ;
    RECT 41.79 46.51 42.0 46.58 ;
    RECT 41.79 46.87 42.0 46.94 ;
    RECT 38.01 46.15 38.22 46.22 ;
    RECT 38.01 46.51 38.22 46.58 ;
    RECT 38.01 46.87 38.22 46.94 ;
    RECT 38.47 46.15 38.68 46.22 ;
    RECT 38.47 46.51 38.68 46.58 ;
    RECT 38.47 46.87 38.68 46.94 ;
    RECT 0.4 46.51 0.47 46.58 ;
    RECT 34.69 46.15 34.9 46.22 ;
    RECT 34.69 46.51 34.9 46.58 ;
    RECT 34.69 46.87 34.9 46.94 ;
    RECT 35.15 46.15 35.36 46.22 ;
    RECT 35.15 46.51 35.36 46.58 ;
    RECT 35.15 46.87 35.36 46.94 ;
    RECT 117.69 46.15 117.9 46.22 ;
    RECT 117.69 46.51 117.9 46.58 ;
    RECT 117.69 46.87 117.9 46.94 ;
    RECT 118.15 46.15 118.36 46.22 ;
    RECT 118.15 46.51 118.36 46.58 ;
    RECT 118.15 46.87 118.36 46.94 ;
    RECT 114.37 46.15 114.58 46.22 ;
    RECT 114.37 46.51 114.58 46.58 ;
    RECT 114.37 46.87 114.58 46.94 ;
    RECT 114.83 46.15 115.04 46.22 ;
    RECT 114.83 46.51 115.04 46.58 ;
    RECT 114.83 46.87 115.04 46.94 ;
    RECT 111.05 46.15 111.26 46.22 ;
    RECT 111.05 46.51 111.26 46.58 ;
    RECT 111.05 46.87 111.26 46.94 ;
    RECT 111.51 46.15 111.72 46.22 ;
    RECT 111.51 46.51 111.72 46.58 ;
    RECT 111.51 46.87 111.72 46.94 ;
    RECT 107.73 46.15 107.94 46.22 ;
    RECT 107.73 46.51 107.94 46.58 ;
    RECT 107.73 46.87 107.94 46.94 ;
    RECT 108.19 46.15 108.4 46.22 ;
    RECT 108.19 46.51 108.4 46.58 ;
    RECT 108.19 46.87 108.4 46.94 ;
    RECT 104.41 46.15 104.62 46.22 ;
    RECT 104.41 46.51 104.62 46.58 ;
    RECT 104.41 46.87 104.62 46.94 ;
    RECT 104.87 46.15 105.08 46.22 ;
    RECT 104.87 46.51 105.08 46.58 ;
    RECT 104.87 46.87 105.08 46.94 ;
    RECT 101.09 46.15 101.3 46.22 ;
    RECT 101.09 46.51 101.3 46.58 ;
    RECT 101.09 46.87 101.3 46.94 ;
    RECT 101.55 46.15 101.76 46.22 ;
    RECT 101.55 46.51 101.76 46.58 ;
    RECT 101.55 46.87 101.76 46.94 ;
    RECT 97.77 46.15 97.98 46.22 ;
    RECT 97.77 46.51 97.98 46.58 ;
    RECT 97.77 46.87 97.98 46.94 ;
    RECT 98.23 46.15 98.44 46.22 ;
    RECT 98.23 46.51 98.44 46.58 ;
    RECT 98.23 46.87 98.44 46.94 ;
    RECT 94.45 46.15 94.66 46.22 ;
    RECT 94.45 46.51 94.66 46.58 ;
    RECT 94.45 46.87 94.66 46.94 ;
    RECT 94.91 46.15 95.12 46.22 ;
    RECT 94.91 46.51 95.12 46.58 ;
    RECT 94.91 46.87 95.12 46.94 ;
    RECT 91.13 46.15 91.34 46.22 ;
    RECT 91.13 46.51 91.34 46.58 ;
    RECT 91.13 46.87 91.34 46.94 ;
    RECT 91.59 46.15 91.8 46.22 ;
    RECT 91.59 46.51 91.8 46.58 ;
    RECT 91.59 46.87 91.8 46.94 ;
    RECT 87.81 46.15 88.02 46.22 ;
    RECT 87.81 46.51 88.02 46.58 ;
    RECT 87.81 46.87 88.02 46.94 ;
    RECT 88.27 46.15 88.48 46.22 ;
    RECT 88.27 46.51 88.48 46.58 ;
    RECT 88.27 46.87 88.48 46.94 ;
    RECT 84.49 46.15 84.7 46.22 ;
    RECT 84.49 46.51 84.7 46.58 ;
    RECT 84.49 46.87 84.7 46.94 ;
    RECT 84.95 46.15 85.16 46.22 ;
    RECT 84.95 46.51 85.16 46.58 ;
    RECT 84.95 46.87 85.16 46.94 ;
    RECT 81.17 46.15 81.38 46.22 ;
    RECT 81.17 46.51 81.38 46.58 ;
    RECT 81.17 46.87 81.38 46.94 ;
    RECT 81.63 46.15 81.84 46.22 ;
    RECT 81.63 46.51 81.84 46.58 ;
    RECT 81.63 46.87 81.84 46.94 ;
    RECT 77.85 46.15 78.06 46.22 ;
    RECT 77.85 46.51 78.06 46.58 ;
    RECT 77.85 46.87 78.06 46.94 ;
    RECT 78.31 46.15 78.52 46.22 ;
    RECT 78.31 46.51 78.52 46.58 ;
    RECT 78.31 46.87 78.52 46.94 ;
    RECT 74.53 46.15 74.74 46.22 ;
    RECT 74.53 46.51 74.74 46.58 ;
    RECT 74.53 46.87 74.74 46.94 ;
    RECT 74.99 46.15 75.2 46.22 ;
    RECT 74.99 46.51 75.2 46.58 ;
    RECT 74.99 46.87 75.2 46.94 ;
    RECT 71.21 46.15 71.42 46.22 ;
    RECT 71.21 46.51 71.42 46.58 ;
    RECT 71.21 46.87 71.42 46.94 ;
    RECT 71.67 46.15 71.88 46.22 ;
    RECT 71.67 46.51 71.88 46.58 ;
    RECT 71.67 46.87 71.88 46.94 ;
    RECT 31.37 46.15 31.58 46.22 ;
    RECT 31.37 46.51 31.58 46.58 ;
    RECT 31.37 46.87 31.58 46.94 ;
    RECT 31.83 46.15 32.04 46.22 ;
    RECT 31.83 46.51 32.04 46.58 ;
    RECT 31.83 46.87 32.04 46.94 ;
    RECT 67.89 46.15 68.1 46.22 ;
    RECT 67.89 46.51 68.1 46.58 ;
    RECT 67.89 46.87 68.1 46.94 ;
    RECT 68.35 46.15 68.56 46.22 ;
    RECT 68.35 46.51 68.56 46.58 ;
    RECT 68.35 46.87 68.56 46.94 ;
    RECT 28.05 46.15 28.26 46.22 ;
    RECT 28.05 46.51 28.26 46.58 ;
    RECT 28.05 46.87 28.26 46.94 ;
    RECT 28.51 46.15 28.72 46.22 ;
    RECT 28.51 46.51 28.72 46.58 ;
    RECT 28.51 46.87 28.72 46.94 ;
    RECT 24.73 46.15 24.94 46.22 ;
    RECT 24.73 46.51 24.94 46.58 ;
    RECT 24.73 46.87 24.94 46.94 ;
    RECT 25.19 46.15 25.4 46.22 ;
    RECT 25.19 46.51 25.4 46.58 ;
    RECT 25.19 46.87 25.4 46.94 ;
    RECT 21.41 46.15 21.62 46.22 ;
    RECT 21.41 46.51 21.62 46.58 ;
    RECT 21.41 46.87 21.62 46.94 ;
    RECT 21.87 46.15 22.08 46.22 ;
    RECT 21.87 46.51 22.08 46.58 ;
    RECT 21.87 46.87 22.08 46.94 ;
    RECT 18.09 46.15 18.3 46.22 ;
    RECT 18.09 46.51 18.3 46.58 ;
    RECT 18.09 46.87 18.3 46.94 ;
    RECT 18.55 46.15 18.76 46.22 ;
    RECT 18.55 46.51 18.76 46.58 ;
    RECT 18.55 46.87 18.76 46.94 ;
    RECT 120.825 46.51 120.895 46.58 ;
    RECT 14.77 46.15 14.98 46.22 ;
    RECT 14.77 46.51 14.98 46.58 ;
    RECT 14.77 46.87 14.98 46.94 ;
    RECT 15.23 46.15 15.44 46.22 ;
    RECT 15.23 46.51 15.44 46.58 ;
    RECT 15.23 46.87 15.44 46.94 ;
    RECT 11.45 46.15 11.66 46.22 ;
    RECT 11.45 46.51 11.66 46.58 ;
    RECT 11.45 46.87 11.66 46.94 ;
    RECT 11.91 46.15 12.12 46.22 ;
    RECT 11.91 46.51 12.12 46.58 ;
    RECT 11.91 46.87 12.12 46.94 ;
    RECT 8.13 46.15 8.34 46.22 ;
    RECT 8.13 46.51 8.34 46.58 ;
    RECT 8.13 46.87 8.34 46.94 ;
    RECT 8.59 46.15 8.8 46.22 ;
    RECT 8.59 46.51 8.8 46.58 ;
    RECT 8.59 46.87 8.8 46.94 ;
    RECT 4.81 46.15 5.02 46.22 ;
    RECT 4.81 46.51 5.02 46.58 ;
    RECT 4.81 46.87 5.02 46.94 ;
    RECT 5.27 46.15 5.48 46.22 ;
    RECT 5.27 46.51 5.48 46.58 ;
    RECT 5.27 46.87 5.48 46.94 ;
    RECT 1.49 46.15 1.7 46.22 ;
    RECT 1.49 46.51 1.7 46.58 ;
    RECT 1.49 46.87 1.7 46.94 ;
    RECT 1.95 46.15 2.16 46.22 ;
    RECT 1.95 46.51 2.16 46.58 ;
    RECT 1.95 46.87 2.16 46.94 ;
    RECT 64.57 46.15 64.78 46.22 ;
    RECT 64.57 46.51 64.78 46.58 ;
    RECT 64.57 46.87 64.78 46.94 ;
    RECT 65.03 46.15 65.24 46.22 ;
    RECT 65.03 46.51 65.24 46.58 ;
    RECT 65.03 46.87 65.24 46.94 ;
    RECT 61.25 85.77 61.46 85.84 ;
    RECT 61.25 86.13 61.46 86.2 ;
    RECT 61.25 86.49 61.46 86.56 ;
    RECT 61.71 85.77 61.92 85.84 ;
    RECT 61.71 86.13 61.92 86.2 ;
    RECT 61.71 86.49 61.92 86.56 ;
    RECT 57.93 85.77 58.14 85.84 ;
    RECT 57.93 86.13 58.14 86.2 ;
    RECT 57.93 86.49 58.14 86.56 ;
    RECT 58.39 85.77 58.6 85.84 ;
    RECT 58.39 86.13 58.6 86.2 ;
    RECT 58.39 86.49 58.6 86.56 ;
    RECT 54.61 85.77 54.82 85.84 ;
    RECT 54.61 86.13 54.82 86.2 ;
    RECT 54.61 86.49 54.82 86.56 ;
    RECT 55.07 85.77 55.28 85.84 ;
    RECT 55.07 86.13 55.28 86.2 ;
    RECT 55.07 86.49 55.28 86.56 ;
    RECT 51.29 85.77 51.5 85.84 ;
    RECT 51.29 86.13 51.5 86.2 ;
    RECT 51.29 86.49 51.5 86.56 ;
    RECT 51.75 85.77 51.96 85.84 ;
    RECT 51.75 86.13 51.96 86.2 ;
    RECT 51.75 86.49 51.96 86.56 ;
    RECT 47.97 85.77 48.18 85.84 ;
    RECT 47.97 86.13 48.18 86.2 ;
    RECT 47.97 86.49 48.18 86.56 ;
    RECT 48.43 85.77 48.64 85.84 ;
    RECT 48.43 86.13 48.64 86.2 ;
    RECT 48.43 86.49 48.64 86.56 ;
    RECT 44.65 85.77 44.86 85.84 ;
    RECT 44.65 86.13 44.86 86.2 ;
    RECT 44.65 86.49 44.86 86.56 ;
    RECT 45.11 85.77 45.32 85.84 ;
    RECT 45.11 86.13 45.32 86.2 ;
    RECT 45.11 86.49 45.32 86.56 ;
    RECT 41.33 85.77 41.54 85.84 ;
    RECT 41.33 86.13 41.54 86.2 ;
    RECT 41.33 86.49 41.54 86.56 ;
    RECT 41.79 85.77 42.0 85.84 ;
    RECT 41.79 86.13 42.0 86.2 ;
    RECT 41.79 86.49 42.0 86.56 ;
    RECT 38.01 85.77 38.22 85.84 ;
    RECT 38.01 86.13 38.22 86.2 ;
    RECT 38.01 86.49 38.22 86.56 ;
    RECT 38.47 85.77 38.68 85.84 ;
    RECT 38.47 86.13 38.68 86.2 ;
    RECT 38.47 86.49 38.68 86.56 ;
    RECT 0.4 86.13 0.47 86.2 ;
    RECT 34.69 85.77 34.9 85.84 ;
    RECT 34.69 86.13 34.9 86.2 ;
    RECT 34.69 86.49 34.9 86.56 ;
    RECT 35.15 85.77 35.36 85.84 ;
    RECT 35.15 86.13 35.36 86.2 ;
    RECT 35.15 86.49 35.36 86.56 ;
    RECT 117.69 85.77 117.9 85.84 ;
    RECT 117.69 86.13 117.9 86.2 ;
    RECT 117.69 86.49 117.9 86.56 ;
    RECT 118.15 85.77 118.36 85.84 ;
    RECT 118.15 86.13 118.36 86.2 ;
    RECT 118.15 86.49 118.36 86.56 ;
    RECT 114.37 85.77 114.58 85.84 ;
    RECT 114.37 86.13 114.58 86.2 ;
    RECT 114.37 86.49 114.58 86.56 ;
    RECT 114.83 85.77 115.04 85.84 ;
    RECT 114.83 86.13 115.04 86.2 ;
    RECT 114.83 86.49 115.04 86.56 ;
    RECT 111.05 85.77 111.26 85.84 ;
    RECT 111.05 86.13 111.26 86.2 ;
    RECT 111.05 86.49 111.26 86.56 ;
    RECT 111.51 85.77 111.72 85.84 ;
    RECT 111.51 86.13 111.72 86.2 ;
    RECT 111.51 86.49 111.72 86.56 ;
    RECT 107.73 85.77 107.94 85.84 ;
    RECT 107.73 86.13 107.94 86.2 ;
    RECT 107.73 86.49 107.94 86.56 ;
    RECT 108.19 85.77 108.4 85.84 ;
    RECT 108.19 86.13 108.4 86.2 ;
    RECT 108.19 86.49 108.4 86.56 ;
    RECT 104.41 85.77 104.62 85.84 ;
    RECT 104.41 86.13 104.62 86.2 ;
    RECT 104.41 86.49 104.62 86.56 ;
    RECT 104.87 85.77 105.08 85.84 ;
    RECT 104.87 86.13 105.08 86.2 ;
    RECT 104.87 86.49 105.08 86.56 ;
    RECT 101.09 85.77 101.3 85.84 ;
    RECT 101.09 86.13 101.3 86.2 ;
    RECT 101.09 86.49 101.3 86.56 ;
    RECT 101.55 85.77 101.76 85.84 ;
    RECT 101.55 86.13 101.76 86.2 ;
    RECT 101.55 86.49 101.76 86.56 ;
    RECT 97.77 85.77 97.98 85.84 ;
    RECT 97.77 86.13 97.98 86.2 ;
    RECT 97.77 86.49 97.98 86.56 ;
    RECT 98.23 85.77 98.44 85.84 ;
    RECT 98.23 86.13 98.44 86.2 ;
    RECT 98.23 86.49 98.44 86.56 ;
    RECT 94.45 85.77 94.66 85.84 ;
    RECT 94.45 86.13 94.66 86.2 ;
    RECT 94.45 86.49 94.66 86.56 ;
    RECT 94.91 85.77 95.12 85.84 ;
    RECT 94.91 86.13 95.12 86.2 ;
    RECT 94.91 86.49 95.12 86.56 ;
    RECT 91.13 85.77 91.34 85.84 ;
    RECT 91.13 86.13 91.34 86.2 ;
    RECT 91.13 86.49 91.34 86.56 ;
    RECT 91.59 85.77 91.8 85.84 ;
    RECT 91.59 86.13 91.8 86.2 ;
    RECT 91.59 86.49 91.8 86.56 ;
    RECT 87.81 85.77 88.02 85.84 ;
    RECT 87.81 86.13 88.02 86.2 ;
    RECT 87.81 86.49 88.02 86.56 ;
    RECT 88.27 85.77 88.48 85.84 ;
    RECT 88.27 86.13 88.48 86.2 ;
    RECT 88.27 86.49 88.48 86.56 ;
    RECT 84.49 85.77 84.7 85.84 ;
    RECT 84.49 86.13 84.7 86.2 ;
    RECT 84.49 86.49 84.7 86.56 ;
    RECT 84.95 85.77 85.16 85.84 ;
    RECT 84.95 86.13 85.16 86.2 ;
    RECT 84.95 86.49 85.16 86.56 ;
    RECT 81.17 85.77 81.38 85.84 ;
    RECT 81.17 86.13 81.38 86.2 ;
    RECT 81.17 86.49 81.38 86.56 ;
    RECT 81.63 85.77 81.84 85.84 ;
    RECT 81.63 86.13 81.84 86.2 ;
    RECT 81.63 86.49 81.84 86.56 ;
    RECT 77.85 85.77 78.06 85.84 ;
    RECT 77.85 86.13 78.06 86.2 ;
    RECT 77.85 86.49 78.06 86.56 ;
    RECT 78.31 85.77 78.52 85.84 ;
    RECT 78.31 86.13 78.52 86.2 ;
    RECT 78.31 86.49 78.52 86.56 ;
    RECT 74.53 85.77 74.74 85.84 ;
    RECT 74.53 86.13 74.74 86.2 ;
    RECT 74.53 86.49 74.74 86.56 ;
    RECT 74.99 85.77 75.2 85.84 ;
    RECT 74.99 86.13 75.2 86.2 ;
    RECT 74.99 86.49 75.2 86.56 ;
    RECT 71.21 85.77 71.42 85.84 ;
    RECT 71.21 86.13 71.42 86.2 ;
    RECT 71.21 86.49 71.42 86.56 ;
    RECT 71.67 85.77 71.88 85.84 ;
    RECT 71.67 86.13 71.88 86.2 ;
    RECT 71.67 86.49 71.88 86.56 ;
    RECT 31.37 85.77 31.58 85.84 ;
    RECT 31.37 86.13 31.58 86.2 ;
    RECT 31.37 86.49 31.58 86.56 ;
    RECT 31.83 85.77 32.04 85.84 ;
    RECT 31.83 86.13 32.04 86.2 ;
    RECT 31.83 86.49 32.04 86.56 ;
    RECT 67.89 85.77 68.1 85.84 ;
    RECT 67.89 86.13 68.1 86.2 ;
    RECT 67.89 86.49 68.1 86.56 ;
    RECT 68.35 85.77 68.56 85.84 ;
    RECT 68.35 86.13 68.56 86.2 ;
    RECT 68.35 86.49 68.56 86.56 ;
    RECT 28.05 85.77 28.26 85.84 ;
    RECT 28.05 86.13 28.26 86.2 ;
    RECT 28.05 86.49 28.26 86.56 ;
    RECT 28.51 85.77 28.72 85.84 ;
    RECT 28.51 86.13 28.72 86.2 ;
    RECT 28.51 86.49 28.72 86.56 ;
    RECT 24.73 85.77 24.94 85.84 ;
    RECT 24.73 86.13 24.94 86.2 ;
    RECT 24.73 86.49 24.94 86.56 ;
    RECT 25.19 85.77 25.4 85.84 ;
    RECT 25.19 86.13 25.4 86.2 ;
    RECT 25.19 86.49 25.4 86.56 ;
    RECT 21.41 85.77 21.62 85.84 ;
    RECT 21.41 86.13 21.62 86.2 ;
    RECT 21.41 86.49 21.62 86.56 ;
    RECT 21.87 85.77 22.08 85.84 ;
    RECT 21.87 86.13 22.08 86.2 ;
    RECT 21.87 86.49 22.08 86.56 ;
    RECT 18.09 85.77 18.3 85.84 ;
    RECT 18.09 86.13 18.3 86.2 ;
    RECT 18.09 86.49 18.3 86.56 ;
    RECT 18.55 85.77 18.76 85.84 ;
    RECT 18.55 86.13 18.76 86.2 ;
    RECT 18.55 86.49 18.76 86.56 ;
    RECT 120.825 86.13 120.895 86.2 ;
    RECT 14.77 85.77 14.98 85.84 ;
    RECT 14.77 86.13 14.98 86.2 ;
    RECT 14.77 86.49 14.98 86.56 ;
    RECT 15.23 85.77 15.44 85.84 ;
    RECT 15.23 86.13 15.44 86.2 ;
    RECT 15.23 86.49 15.44 86.56 ;
    RECT 11.45 85.77 11.66 85.84 ;
    RECT 11.45 86.13 11.66 86.2 ;
    RECT 11.45 86.49 11.66 86.56 ;
    RECT 11.91 85.77 12.12 85.84 ;
    RECT 11.91 86.13 12.12 86.2 ;
    RECT 11.91 86.49 12.12 86.56 ;
    RECT 8.13 85.77 8.34 85.84 ;
    RECT 8.13 86.13 8.34 86.2 ;
    RECT 8.13 86.49 8.34 86.56 ;
    RECT 8.59 85.77 8.8 85.84 ;
    RECT 8.59 86.13 8.8 86.2 ;
    RECT 8.59 86.49 8.8 86.56 ;
    RECT 4.81 85.77 5.02 85.84 ;
    RECT 4.81 86.13 5.02 86.2 ;
    RECT 4.81 86.49 5.02 86.56 ;
    RECT 5.27 85.77 5.48 85.84 ;
    RECT 5.27 86.13 5.48 86.2 ;
    RECT 5.27 86.49 5.48 86.56 ;
    RECT 1.49 85.77 1.7 85.84 ;
    RECT 1.49 86.13 1.7 86.2 ;
    RECT 1.49 86.49 1.7 86.56 ;
    RECT 1.95 85.77 2.16 85.84 ;
    RECT 1.95 86.13 2.16 86.2 ;
    RECT 1.95 86.49 2.16 86.56 ;
    RECT 64.57 85.77 64.78 85.84 ;
    RECT 64.57 86.13 64.78 86.2 ;
    RECT 64.57 86.49 64.78 86.56 ;
    RECT 65.03 85.77 65.24 85.84 ;
    RECT 65.03 86.13 65.24 86.2 ;
    RECT 65.03 86.49 65.24 86.56 ;
    RECT 61.25 45.43 61.46 45.5 ;
    RECT 61.25 45.79 61.46 45.86 ;
    RECT 61.25 46.15 61.46 46.22 ;
    RECT 61.71 45.43 61.92 45.5 ;
    RECT 61.71 45.79 61.92 45.86 ;
    RECT 61.71 46.15 61.92 46.22 ;
    RECT 57.93 45.43 58.14 45.5 ;
    RECT 57.93 45.79 58.14 45.86 ;
    RECT 57.93 46.15 58.14 46.22 ;
    RECT 58.39 45.43 58.6 45.5 ;
    RECT 58.39 45.79 58.6 45.86 ;
    RECT 58.39 46.15 58.6 46.22 ;
    RECT 54.61 45.43 54.82 45.5 ;
    RECT 54.61 45.79 54.82 45.86 ;
    RECT 54.61 46.15 54.82 46.22 ;
    RECT 55.07 45.43 55.28 45.5 ;
    RECT 55.07 45.79 55.28 45.86 ;
    RECT 55.07 46.15 55.28 46.22 ;
    RECT 51.29 45.43 51.5 45.5 ;
    RECT 51.29 45.79 51.5 45.86 ;
    RECT 51.29 46.15 51.5 46.22 ;
    RECT 51.75 45.43 51.96 45.5 ;
    RECT 51.75 45.79 51.96 45.86 ;
    RECT 51.75 46.15 51.96 46.22 ;
    RECT 47.97 45.43 48.18 45.5 ;
    RECT 47.97 45.79 48.18 45.86 ;
    RECT 47.97 46.15 48.18 46.22 ;
    RECT 48.43 45.43 48.64 45.5 ;
    RECT 48.43 45.79 48.64 45.86 ;
    RECT 48.43 46.15 48.64 46.22 ;
    RECT 44.65 45.43 44.86 45.5 ;
    RECT 44.65 45.79 44.86 45.86 ;
    RECT 44.65 46.15 44.86 46.22 ;
    RECT 45.11 45.43 45.32 45.5 ;
    RECT 45.11 45.79 45.32 45.86 ;
    RECT 45.11 46.15 45.32 46.22 ;
    RECT 41.33 45.43 41.54 45.5 ;
    RECT 41.33 45.79 41.54 45.86 ;
    RECT 41.33 46.15 41.54 46.22 ;
    RECT 41.79 45.43 42.0 45.5 ;
    RECT 41.79 45.79 42.0 45.86 ;
    RECT 41.79 46.15 42.0 46.22 ;
    RECT 38.01 45.43 38.22 45.5 ;
    RECT 38.01 45.79 38.22 45.86 ;
    RECT 38.01 46.15 38.22 46.22 ;
    RECT 38.47 45.43 38.68 45.5 ;
    RECT 38.47 45.79 38.68 45.86 ;
    RECT 38.47 46.15 38.68 46.22 ;
    RECT 0.4 45.79 0.47 45.86 ;
    RECT 34.69 45.43 34.9 45.5 ;
    RECT 34.69 45.79 34.9 45.86 ;
    RECT 34.69 46.15 34.9 46.22 ;
    RECT 35.15 45.43 35.36 45.5 ;
    RECT 35.15 45.79 35.36 45.86 ;
    RECT 35.15 46.15 35.36 46.22 ;
    RECT 117.69 45.43 117.9 45.5 ;
    RECT 117.69 45.79 117.9 45.86 ;
    RECT 117.69 46.15 117.9 46.22 ;
    RECT 118.15 45.43 118.36 45.5 ;
    RECT 118.15 45.79 118.36 45.86 ;
    RECT 118.15 46.15 118.36 46.22 ;
    RECT 114.37 45.43 114.58 45.5 ;
    RECT 114.37 45.79 114.58 45.86 ;
    RECT 114.37 46.15 114.58 46.22 ;
    RECT 114.83 45.43 115.04 45.5 ;
    RECT 114.83 45.79 115.04 45.86 ;
    RECT 114.83 46.15 115.04 46.22 ;
    RECT 111.05 45.43 111.26 45.5 ;
    RECT 111.05 45.79 111.26 45.86 ;
    RECT 111.05 46.15 111.26 46.22 ;
    RECT 111.51 45.43 111.72 45.5 ;
    RECT 111.51 45.79 111.72 45.86 ;
    RECT 111.51 46.15 111.72 46.22 ;
    RECT 107.73 45.43 107.94 45.5 ;
    RECT 107.73 45.79 107.94 45.86 ;
    RECT 107.73 46.15 107.94 46.22 ;
    RECT 108.19 45.43 108.4 45.5 ;
    RECT 108.19 45.79 108.4 45.86 ;
    RECT 108.19 46.15 108.4 46.22 ;
    RECT 104.41 45.43 104.62 45.5 ;
    RECT 104.41 45.79 104.62 45.86 ;
    RECT 104.41 46.15 104.62 46.22 ;
    RECT 104.87 45.43 105.08 45.5 ;
    RECT 104.87 45.79 105.08 45.86 ;
    RECT 104.87 46.15 105.08 46.22 ;
    RECT 101.09 45.43 101.3 45.5 ;
    RECT 101.09 45.79 101.3 45.86 ;
    RECT 101.09 46.15 101.3 46.22 ;
    RECT 101.55 45.43 101.76 45.5 ;
    RECT 101.55 45.79 101.76 45.86 ;
    RECT 101.55 46.15 101.76 46.22 ;
    RECT 97.77 45.43 97.98 45.5 ;
    RECT 97.77 45.79 97.98 45.86 ;
    RECT 97.77 46.15 97.98 46.22 ;
    RECT 98.23 45.43 98.44 45.5 ;
    RECT 98.23 45.79 98.44 45.86 ;
    RECT 98.23 46.15 98.44 46.22 ;
    RECT 94.45 45.43 94.66 45.5 ;
    RECT 94.45 45.79 94.66 45.86 ;
    RECT 94.45 46.15 94.66 46.22 ;
    RECT 94.91 45.43 95.12 45.5 ;
    RECT 94.91 45.79 95.12 45.86 ;
    RECT 94.91 46.15 95.12 46.22 ;
    RECT 91.13 45.43 91.34 45.5 ;
    RECT 91.13 45.79 91.34 45.86 ;
    RECT 91.13 46.15 91.34 46.22 ;
    RECT 91.59 45.43 91.8 45.5 ;
    RECT 91.59 45.79 91.8 45.86 ;
    RECT 91.59 46.15 91.8 46.22 ;
    RECT 87.81 45.43 88.02 45.5 ;
    RECT 87.81 45.79 88.02 45.86 ;
    RECT 87.81 46.15 88.02 46.22 ;
    RECT 88.27 45.43 88.48 45.5 ;
    RECT 88.27 45.79 88.48 45.86 ;
    RECT 88.27 46.15 88.48 46.22 ;
    RECT 84.49 45.43 84.7 45.5 ;
    RECT 84.49 45.79 84.7 45.86 ;
    RECT 84.49 46.15 84.7 46.22 ;
    RECT 84.95 45.43 85.16 45.5 ;
    RECT 84.95 45.79 85.16 45.86 ;
    RECT 84.95 46.15 85.16 46.22 ;
    RECT 81.17 45.43 81.38 45.5 ;
    RECT 81.17 45.79 81.38 45.86 ;
    RECT 81.17 46.15 81.38 46.22 ;
    RECT 81.63 45.43 81.84 45.5 ;
    RECT 81.63 45.79 81.84 45.86 ;
    RECT 81.63 46.15 81.84 46.22 ;
    RECT 77.85 45.43 78.06 45.5 ;
    RECT 77.85 45.79 78.06 45.86 ;
    RECT 77.85 46.15 78.06 46.22 ;
    RECT 78.31 45.43 78.52 45.5 ;
    RECT 78.31 45.79 78.52 45.86 ;
    RECT 78.31 46.15 78.52 46.22 ;
    RECT 74.53 45.43 74.74 45.5 ;
    RECT 74.53 45.79 74.74 45.86 ;
    RECT 74.53 46.15 74.74 46.22 ;
    RECT 74.99 45.43 75.2 45.5 ;
    RECT 74.99 45.79 75.2 45.86 ;
    RECT 74.99 46.15 75.2 46.22 ;
    RECT 71.21 45.43 71.42 45.5 ;
    RECT 71.21 45.79 71.42 45.86 ;
    RECT 71.21 46.15 71.42 46.22 ;
    RECT 71.67 45.43 71.88 45.5 ;
    RECT 71.67 45.79 71.88 45.86 ;
    RECT 71.67 46.15 71.88 46.22 ;
    RECT 31.37 45.43 31.58 45.5 ;
    RECT 31.37 45.79 31.58 45.86 ;
    RECT 31.37 46.15 31.58 46.22 ;
    RECT 31.83 45.43 32.04 45.5 ;
    RECT 31.83 45.79 32.04 45.86 ;
    RECT 31.83 46.15 32.04 46.22 ;
    RECT 67.89 45.43 68.1 45.5 ;
    RECT 67.89 45.79 68.1 45.86 ;
    RECT 67.89 46.15 68.1 46.22 ;
    RECT 68.35 45.43 68.56 45.5 ;
    RECT 68.35 45.79 68.56 45.86 ;
    RECT 68.35 46.15 68.56 46.22 ;
    RECT 28.05 45.43 28.26 45.5 ;
    RECT 28.05 45.79 28.26 45.86 ;
    RECT 28.05 46.15 28.26 46.22 ;
    RECT 28.51 45.43 28.72 45.5 ;
    RECT 28.51 45.79 28.72 45.86 ;
    RECT 28.51 46.15 28.72 46.22 ;
    RECT 24.73 45.43 24.94 45.5 ;
    RECT 24.73 45.79 24.94 45.86 ;
    RECT 24.73 46.15 24.94 46.22 ;
    RECT 25.19 45.43 25.4 45.5 ;
    RECT 25.19 45.79 25.4 45.86 ;
    RECT 25.19 46.15 25.4 46.22 ;
    RECT 21.41 45.43 21.62 45.5 ;
    RECT 21.41 45.79 21.62 45.86 ;
    RECT 21.41 46.15 21.62 46.22 ;
    RECT 21.87 45.43 22.08 45.5 ;
    RECT 21.87 45.79 22.08 45.86 ;
    RECT 21.87 46.15 22.08 46.22 ;
    RECT 18.09 45.43 18.3 45.5 ;
    RECT 18.09 45.79 18.3 45.86 ;
    RECT 18.09 46.15 18.3 46.22 ;
    RECT 18.55 45.43 18.76 45.5 ;
    RECT 18.55 45.79 18.76 45.86 ;
    RECT 18.55 46.15 18.76 46.22 ;
    RECT 120.825 45.79 120.895 45.86 ;
    RECT 14.77 45.43 14.98 45.5 ;
    RECT 14.77 45.79 14.98 45.86 ;
    RECT 14.77 46.15 14.98 46.22 ;
    RECT 15.23 45.43 15.44 45.5 ;
    RECT 15.23 45.79 15.44 45.86 ;
    RECT 15.23 46.15 15.44 46.22 ;
    RECT 11.45 45.43 11.66 45.5 ;
    RECT 11.45 45.79 11.66 45.86 ;
    RECT 11.45 46.15 11.66 46.22 ;
    RECT 11.91 45.43 12.12 45.5 ;
    RECT 11.91 45.79 12.12 45.86 ;
    RECT 11.91 46.15 12.12 46.22 ;
    RECT 8.13 45.43 8.34 45.5 ;
    RECT 8.13 45.79 8.34 45.86 ;
    RECT 8.13 46.15 8.34 46.22 ;
    RECT 8.59 45.43 8.8 45.5 ;
    RECT 8.59 45.79 8.8 45.86 ;
    RECT 8.59 46.15 8.8 46.22 ;
    RECT 4.81 45.43 5.02 45.5 ;
    RECT 4.81 45.79 5.02 45.86 ;
    RECT 4.81 46.15 5.02 46.22 ;
    RECT 5.27 45.43 5.48 45.5 ;
    RECT 5.27 45.79 5.48 45.86 ;
    RECT 5.27 46.15 5.48 46.22 ;
    RECT 1.49 45.43 1.7 45.5 ;
    RECT 1.49 45.79 1.7 45.86 ;
    RECT 1.49 46.15 1.7 46.22 ;
    RECT 1.95 45.43 2.16 45.5 ;
    RECT 1.95 45.79 2.16 45.86 ;
    RECT 1.95 46.15 2.16 46.22 ;
    RECT 64.57 45.43 64.78 45.5 ;
    RECT 64.57 45.79 64.78 45.86 ;
    RECT 64.57 46.15 64.78 46.22 ;
    RECT 65.03 45.43 65.24 45.5 ;
    RECT 65.03 45.79 65.24 45.86 ;
    RECT 65.03 46.15 65.24 46.22 ;
    RECT 61.25 85.05 61.46 85.12 ;
    RECT 61.25 85.41 61.46 85.48 ;
    RECT 61.25 85.77 61.46 85.84 ;
    RECT 61.71 85.05 61.92 85.12 ;
    RECT 61.71 85.41 61.92 85.48 ;
    RECT 61.71 85.77 61.92 85.84 ;
    RECT 57.93 85.05 58.14 85.12 ;
    RECT 57.93 85.41 58.14 85.48 ;
    RECT 57.93 85.77 58.14 85.84 ;
    RECT 58.39 85.05 58.6 85.12 ;
    RECT 58.39 85.41 58.6 85.48 ;
    RECT 58.39 85.77 58.6 85.84 ;
    RECT 54.61 85.05 54.82 85.12 ;
    RECT 54.61 85.41 54.82 85.48 ;
    RECT 54.61 85.77 54.82 85.84 ;
    RECT 55.07 85.05 55.28 85.12 ;
    RECT 55.07 85.41 55.28 85.48 ;
    RECT 55.07 85.77 55.28 85.84 ;
    RECT 51.29 85.05 51.5 85.12 ;
    RECT 51.29 85.41 51.5 85.48 ;
    RECT 51.29 85.77 51.5 85.84 ;
    RECT 51.75 85.05 51.96 85.12 ;
    RECT 51.75 85.41 51.96 85.48 ;
    RECT 51.75 85.77 51.96 85.84 ;
    RECT 47.97 85.05 48.18 85.12 ;
    RECT 47.97 85.41 48.18 85.48 ;
    RECT 47.97 85.77 48.18 85.84 ;
    RECT 48.43 85.05 48.64 85.12 ;
    RECT 48.43 85.41 48.64 85.48 ;
    RECT 48.43 85.77 48.64 85.84 ;
    RECT 44.65 85.05 44.86 85.12 ;
    RECT 44.65 85.41 44.86 85.48 ;
    RECT 44.65 85.77 44.86 85.84 ;
    RECT 45.11 85.05 45.32 85.12 ;
    RECT 45.11 85.41 45.32 85.48 ;
    RECT 45.11 85.77 45.32 85.84 ;
    RECT 41.33 85.05 41.54 85.12 ;
    RECT 41.33 85.41 41.54 85.48 ;
    RECT 41.33 85.77 41.54 85.84 ;
    RECT 41.79 85.05 42.0 85.12 ;
    RECT 41.79 85.41 42.0 85.48 ;
    RECT 41.79 85.77 42.0 85.84 ;
    RECT 38.01 85.05 38.22 85.12 ;
    RECT 38.01 85.41 38.22 85.48 ;
    RECT 38.01 85.77 38.22 85.84 ;
    RECT 38.47 85.05 38.68 85.12 ;
    RECT 38.47 85.41 38.68 85.48 ;
    RECT 38.47 85.77 38.68 85.84 ;
    RECT 0.4 85.41 0.47 85.48 ;
    RECT 34.69 85.05 34.9 85.12 ;
    RECT 34.69 85.41 34.9 85.48 ;
    RECT 34.69 85.77 34.9 85.84 ;
    RECT 35.15 85.05 35.36 85.12 ;
    RECT 35.15 85.41 35.36 85.48 ;
    RECT 35.15 85.77 35.36 85.84 ;
    RECT 117.69 85.05 117.9 85.12 ;
    RECT 117.69 85.41 117.9 85.48 ;
    RECT 117.69 85.77 117.9 85.84 ;
    RECT 118.15 85.05 118.36 85.12 ;
    RECT 118.15 85.41 118.36 85.48 ;
    RECT 118.15 85.77 118.36 85.84 ;
    RECT 114.37 85.05 114.58 85.12 ;
    RECT 114.37 85.41 114.58 85.48 ;
    RECT 114.37 85.77 114.58 85.84 ;
    RECT 114.83 85.05 115.04 85.12 ;
    RECT 114.83 85.41 115.04 85.48 ;
    RECT 114.83 85.77 115.04 85.84 ;
    RECT 111.05 85.05 111.26 85.12 ;
    RECT 111.05 85.41 111.26 85.48 ;
    RECT 111.05 85.77 111.26 85.84 ;
    RECT 111.51 85.05 111.72 85.12 ;
    RECT 111.51 85.41 111.72 85.48 ;
    RECT 111.51 85.77 111.72 85.84 ;
    RECT 107.73 85.05 107.94 85.12 ;
    RECT 107.73 85.41 107.94 85.48 ;
    RECT 107.73 85.77 107.94 85.84 ;
    RECT 108.19 85.05 108.4 85.12 ;
    RECT 108.19 85.41 108.4 85.48 ;
    RECT 108.19 85.77 108.4 85.84 ;
    RECT 104.41 85.05 104.62 85.12 ;
    RECT 104.41 85.41 104.62 85.48 ;
    RECT 104.41 85.77 104.62 85.84 ;
    RECT 104.87 85.05 105.08 85.12 ;
    RECT 104.87 85.41 105.08 85.48 ;
    RECT 104.87 85.77 105.08 85.84 ;
    RECT 101.09 85.05 101.3 85.12 ;
    RECT 101.09 85.41 101.3 85.48 ;
    RECT 101.09 85.77 101.3 85.84 ;
    RECT 101.55 85.05 101.76 85.12 ;
    RECT 101.55 85.41 101.76 85.48 ;
    RECT 101.55 85.77 101.76 85.84 ;
    RECT 97.77 85.05 97.98 85.12 ;
    RECT 97.77 85.41 97.98 85.48 ;
    RECT 97.77 85.77 97.98 85.84 ;
    RECT 98.23 85.05 98.44 85.12 ;
    RECT 98.23 85.41 98.44 85.48 ;
    RECT 98.23 85.77 98.44 85.84 ;
    RECT 94.45 85.05 94.66 85.12 ;
    RECT 94.45 85.41 94.66 85.48 ;
    RECT 94.45 85.77 94.66 85.84 ;
    RECT 94.91 85.05 95.12 85.12 ;
    RECT 94.91 85.41 95.12 85.48 ;
    RECT 94.91 85.77 95.12 85.84 ;
    RECT 91.13 85.05 91.34 85.12 ;
    RECT 91.13 85.41 91.34 85.48 ;
    RECT 91.13 85.77 91.34 85.84 ;
    RECT 91.59 85.05 91.8 85.12 ;
    RECT 91.59 85.41 91.8 85.48 ;
    RECT 91.59 85.77 91.8 85.84 ;
    RECT 87.81 85.05 88.02 85.12 ;
    RECT 87.81 85.41 88.02 85.48 ;
    RECT 87.81 85.77 88.02 85.84 ;
    RECT 88.27 85.05 88.48 85.12 ;
    RECT 88.27 85.41 88.48 85.48 ;
    RECT 88.27 85.77 88.48 85.84 ;
    RECT 84.49 85.05 84.7 85.12 ;
    RECT 84.49 85.41 84.7 85.48 ;
    RECT 84.49 85.77 84.7 85.84 ;
    RECT 84.95 85.05 85.16 85.12 ;
    RECT 84.95 85.41 85.16 85.48 ;
    RECT 84.95 85.77 85.16 85.84 ;
    RECT 81.17 85.05 81.38 85.12 ;
    RECT 81.17 85.41 81.38 85.48 ;
    RECT 81.17 85.77 81.38 85.84 ;
    RECT 81.63 85.05 81.84 85.12 ;
    RECT 81.63 85.41 81.84 85.48 ;
    RECT 81.63 85.77 81.84 85.84 ;
    RECT 77.85 85.05 78.06 85.12 ;
    RECT 77.85 85.41 78.06 85.48 ;
    RECT 77.85 85.77 78.06 85.84 ;
    RECT 78.31 85.05 78.52 85.12 ;
    RECT 78.31 85.41 78.52 85.48 ;
    RECT 78.31 85.77 78.52 85.84 ;
    RECT 74.53 85.05 74.74 85.12 ;
    RECT 74.53 85.41 74.74 85.48 ;
    RECT 74.53 85.77 74.74 85.84 ;
    RECT 74.99 85.05 75.2 85.12 ;
    RECT 74.99 85.41 75.2 85.48 ;
    RECT 74.99 85.77 75.2 85.84 ;
    RECT 71.21 85.05 71.42 85.12 ;
    RECT 71.21 85.41 71.42 85.48 ;
    RECT 71.21 85.77 71.42 85.84 ;
    RECT 71.67 85.05 71.88 85.12 ;
    RECT 71.67 85.41 71.88 85.48 ;
    RECT 71.67 85.77 71.88 85.84 ;
    RECT 31.37 85.05 31.58 85.12 ;
    RECT 31.37 85.41 31.58 85.48 ;
    RECT 31.37 85.77 31.58 85.84 ;
    RECT 31.83 85.05 32.04 85.12 ;
    RECT 31.83 85.41 32.04 85.48 ;
    RECT 31.83 85.77 32.04 85.84 ;
    RECT 67.89 85.05 68.1 85.12 ;
    RECT 67.89 85.41 68.1 85.48 ;
    RECT 67.89 85.77 68.1 85.84 ;
    RECT 68.35 85.05 68.56 85.12 ;
    RECT 68.35 85.41 68.56 85.48 ;
    RECT 68.35 85.77 68.56 85.84 ;
    RECT 28.05 85.05 28.26 85.12 ;
    RECT 28.05 85.41 28.26 85.48 ;
    RECT 28.05 85.77 28.26 85.84 ;
    RECT 28.51 85.05 28.72 85.12 ;
    RECT 28.51 85.41 28.72 85.48 ;
    RECT 28.51 85.77 28.72 85.84 ;
    RECT 24.73 85.05 24.94 85.12 ;
    RECT 24.73 85.41 24.94 85.48 ;
    RECT 24.73 85.77 24.94 85.84 ;
    RECT 25.19 85.05 25.4 85.12 ;
    RECT 25.19 85.41 25.4 85.48 ;
    RECT 25.19 85.77 25.4 85.84 ;
    RECT 21.41 85.05 21.62 85.12 ;
    RECT 21.41 85.41 21.62 85.48 ;
    RECT 21.41 85.77 21.62 85.84 ;
    RECT 21.87 85.05 22.08 85.12 ;
    RECT 21.87 85.41 22.08 85.48 ;
    RECT 21.87 85.77 22.08 85.84 ;
    RECT 18.09 85.05 18.3 85.12 ;
    RECT 18.09 85.41 18.3 85.48 ;
    RECT 18.09 85.77 18.3 85.84 ;
    RECT 18.55 85.05 18.76 85.12 ;
    RECT 18.55 85.41 18.76 85.48 ;
    RECT 18.55 85.77 18.76 85.84 ;
    RECT 120.825 85.41 120.895 85.48 ;
    RECT 14.77 85.05 14.98 85.12 ;
    RECT 14.77 85.41 14.98 85.48 ;
    RECT 14.77 85.77 14.98 85.84 ;
    RECT 15.23 85.05 15.44 85.12 ;
    RECT 15.23 85.41 15.44 85.48 ;
    RECT 15.23 85.77 15.44 85.84 ;
    RECT 11.45 85.05 11.66 85.12 ;
    RECT 11.45 85.41 11.66 85.48 ;
    RECT 11.45 85.77 11.66 85.84 ;
    RECT 11.91 85.05 12.12 85.12 ;
    RECT 11.91 85.41 12.12 85.48 ;
    RECT 11.91 85.77 12.12 85.84 ;
    RECT 8.13 85.05 8.34 85.12 ;
    RECT 8.13 85.41 8.34 85.48 ;
    RECT 8.13 85.77 8.34 85.84 ;
    RECT 8.59 85.05 8.8 85.12 ;
    RECT 8.59 85.41 8.8 85.48 ;
    RECT 8.59 85.77 8.8 85.84 ;
    RECT 4.81 85.05 5.02 85.12 ;
    RECT 4.81 85.41 5.02 85.48 ;
    RECT 4.81 85.77 5.02 85.84 ;
    RECT 5.27 85.05 5.48 85.12 ;
    RECT 5.27 85.41 5.48 85.48 ;
    RECT 5.27 85.77 5.48 85.84 ;
    RECT 1.49 85.05 1.7 85.12 ;
    RECT 1.49 85.41 1.7 85.48 ;
    RECT 1.49 85.77 1.7 85.84 ;
    RECT 1.95 85.05 2.16 85.12 ;
    RECT 1.95 85.41 2.16 85.48 ;
    RECT 1.95 85.77 2.16 85.84 ;
    RECT 64.57 85.05 64.78 85.12 ;
    RECT 64.57 85.41 64.78 85.48 ;
    RECT 64.57 85.77 64.78 85.84 ;
    RECT 65.03 85.05 65.24 85.12 ;
    RECT 65.03 85.41 65.24 85.48 ;
    RECT 65.03 85.77 65.24 85.84 ;
    RECT 61.25 44.71 61.46 44.78 ;
    RECT 61.25 45.07 61.46 45.14 ;
    RECT 61.25 45.43 61.46 45.5 ;
    RECT 61.71 44.71 61.92 44.78 ;
    RECT 61.71 45.07 61.92 45.14 ;
    RECT 61.71 45.43 61.92 45.5 ;
    RECT 57.93 44.71 58.14 44.78 ;
    RECT 57.93 45.07 58.14 45.14 ;
    RECT 57.93 45.43 58.14 45.5 ;
    RECT 58.39 44.71 58.6 44.78 ;
    RECT 58.39 45.07 58.6 45.14 ;
    RECT 58.39 45.43 58.6 45.5 ;
    RECT 54.61 44.71 54.82 44.78 ;
    RECT 54.61 45.07 54.82 45.14 ;
    RECT 54.61 45.43 54.82 45.5 ;
    RECT 55.07 44.71 55.28 44.78 ;
    RECT 55.07 45.07 55.28 45.14 ;
    RECT 55.07 45.43 55.28 45.5 ;
    RECT 51.29 44.71 51.5 44.78 ;
    RECT 51.29 45.07 51.5 45.14 ;
    RECT 51.29 45.43 51.5 45.5 ;
    RECT 51.75 44.71 51.96 44.78 ;
    RECT 51.75 45.07 51.96 45.14 ;
    RECT 51.75 45.43 51.96 45.5 ;
    RECT 47.97 44.71 48.18 44.78 ;
    RECT 47.97 45.07 48.18 45.14 ;
    RECT 47.97 45.43 48.18 45.5 ;
    RECT 48.43 44.71 48.64 44.78 ;
    RECT 48.43 45.07 48.64 45.14 ;
    RECT 48.43 45.43 48.64 45.5 ;
    RECT 44.65 44.71 44.86 44.78 ;
    RECT 44.65 45.07 44.86 45.14 ;
    RECT 44.65 45.43 44.86 45.5 ;
    RECT 45.11 44.71 45.32 44.78 ;
    RECT 45.11 45.07 45.32 45.14 ;
    RECT 45.11 45.43 45.32 45.5 ;
    RECT 41.33 44.71 41.54 44.78 ;
    RECT 41.33 45.07 41.54 45.14 ;
    RECT 41.33 45.43 41.54 45.5 ;
    RECT 41.79 44.71 42.0 44.78 ;
    RECT 41.79 45.07 42.0 45.14 ;
    RECT 41.79 45.43 42.0 45.5 ;
    RECT 38.01 44.71 38.22 44.78 ;
    RECT 38.01 45.07 38.22 45.14 ;
    RECT 38.01 45.43 38.22 45.5 ;
    RECT 38.47 44.71 38.68 44.78 ;
    RECT 38.47 45.07 38.68 45.14 ;
    RECT 38.47 45.43 38.68 45.5 ;
    RECT 0.4 45.07 0.47 45.14 ;
    RECT 34.69 44.71 34.9 44.78 ;
    RECT 34.69 45.07 34.9 45.14 ;
    RECT 34.69 45.43 34.9 45.5 ;
    RECT 35.15 44.71 35.36 44.78 ;
    RECT 35.15 45.07 35.36 45.14 ;
    RECT 35.15 45.43 35.36 45.5 ;
    RECT 117.69 44.71 117.9 44.78 ;
    RECT 117.69 45.07 117.9 45.14 ;
    RECT 117.69 45.43 117.9 45.5 ;
    RECT 118.15 44.71 118.36 44.78 ;
    RECT 118.15 45.07 118.36 45.14 ;
    RECT 118.15 45.43 118.36 45.5 ;
    RECT 114.37 44.71 114.58 44.78 ;
    RECT 114.37 45.07 114.58 45.14 ;
    RECT 114.37 45.43 114.58 45.5 ;
    RECT 114.83 44.71 115.04 44.78 ;
    RECT 114.83 45.07 115.04 45.14 ;
    RECT 114.83 45.43 115.04 45.5 ;
    RECT 111.05 44.71 111.26 44.78 ;
    RECT 111.05 45.07 111.26 45.14 ;
    RECT 111.05 45.43 111.26 45.5 ;
    RECT 111.51 44.71 111.72 44.78 ;
    RECT 111.51 45.07 111.72 45.14 ;
    RECT 111.51 45.43 111.72 45.5 ;
    RECT 107.73 44.71 107.94 44.78 ;
    RECT 107.73 45.07 107.94 45.14 ;
    RECT 107.73 45.43 107.94 45.5 ;
    RECT 108.19 44.71 108.4 44.78 ;
    RECT 108.19 45.07 108.4 45.14 ;
    RECT 108.19 45.43 108.4 45.5 ;
    RECT 104.41 44.71 104.62 44.78 ;
    RECT 104.41 45.07 104.62 45.14 ;
    RECT 104.41 45.43 104.62 45.5 ;
    RECT 104.87 44.71 105.08 44.78 ;
    RECT 104.87 45.07 105.08 45.14 ;
    RECT 104.87 45.43 105.08 45.5 ;
    RECT 101.09 44.71 101.3 44.78 ;
    RECT 101.09 45.07 101.3 45.14 ;
    RECT 101.09 45.43 101.3 45.5 ;
    RECT 101.55 44.71 101.76 44.78 ;
    RECT 101.55 45.07 101.76 45.14 ;
    RECT 101.55 45.43 101.76 45.5 ;
    RECT 97.77 44.71 97.98 44.78 ;
    RECT 97.77 45.07 97.98 45.14 ;
    RECT 97.77 45.43 97.98 45.5 ;
    RECT 98.23 44.71 98.44 44.78 ;
    RECT 98.23 45.07 98.44 45.14 ;
    RECT 98.23 45.43 98.44 45.5 ;
    RECT 94.45 44.71 94.66 44.78 ;
    RECT 94.45 45.07 94.66 45.14 ;
    RECT 94.45 45.43 94.66 45.5 ;
    RECT 94.91 44.71 95.12 44.78 ;
    RECT 94.91 45.07 95.12 45.14 ;
    RECT 94.91 45.43 95.12 45.5 ;
    RECT 91.13 44.71 91.34 44.78 ;
    RECT 91.13 45.07 91.34 45.14 ;
    RECT 91.13 45.43 91.34 45.5 ;
    RECT 91.59 44.71 91.8 44.78 ;
    RECT 91.59 45.07 91.8 45.14 ;
    RECT 91.59 45.43 91.8 45.5 ;
    RECT 87.81 44.71 88.02 44.78 ;
    RECT 87.81 45.07 88.02 45.14 ;
    RECT 87.81 45.43 88.02 45.5 ;
    RECT 88.27 44.71 88.48 44.78 ;
    RECT 88.27 45.07 88.48 45.14 ;
    RECT 88.27 45.43 88.48 45.5 ;
    RECT 84.49 44.71 84.7 44.78 ;
    RECT 84.49 45.07 84.7 45.14 ;
    RECT 84.49 45.43 84.7 45.5 ;
    RECT 84.95 44.71 85.16 44.78 ;
    RECT 84.95 45.07 85.16 45.14 ;
    RECT 84.95 45.43 85.16 45.5 ;
    RECT 81.17 44.71 81.38 44.78 ;
    RECT 81.17 45.07 81.38 45.14 ;
    RECT 81.17 45.43 81.38 45.5 ;
    RECT 81.63 44.71 81.84 44.78 ;
    RECT 81.63 45.07 81.84 45.14 ;
    RECT 81.63 45.43 81.84 45.5 ;
    RECT 77.85 44.71 78.06 44.78 ;
    RECT 77.85 45.07 78.06 45.14 ;
    RECT 77.85 45.43 78.06 45.5 ;
    RECT 78.31 44.71 78.52 44.78 ;
    RECT 78.31 45.07 78.52 45.14 ;
    RECT 78.31 45.43 78.52 45.5 ;
    RECT 74.53 44.71 74.74 44.78 ;
    RECT 74.53 45.07 74.74 45.14 ;
    RECT 74.53 45.43 74.74 45.5 ;
    RECT 74.99 44.71 75.2 44.78 ;
    RECT 74.99 45.07 75.2 45.14 ;
    RECT 74.99 45.43 75.2 45.5 ;
    RECT 71.21 44.71 71.42 44.78 ;
    RECT 71.21 45.07 71.42 45.14 ;
    RECT 71.21 45.43 71.42 45.5 ;
    RECT 71.67 44.71 71.88 44.78 ;
    RECT 71.67 45.07 71.88 45.14 ;
    RECT 71.67 45.43 71.88 45.5 ;
    RECT 31.37 44.71 31.58 44.78 ;
    RECT 31.37 45.07 31.58 45.14 ;
    RECT 31.37 45.43 31.58 45.5 ;
    RECT 31.83 44.71 32.04 44.78 ;
    RECT 31.83 45.07 32.04 45.14 ;
    RECT 31.83 45.43 32.04 45.5 ;
    RECT 67.89 44.71 68.1 44.78 ;
    RECT 67.89 45.07 68.1 45.14 ;
    RECT 67.89 45.43 68.1 45.5 ;
    RECT 68.35 44.71 68.56 44.78 ;
    RECT 68.35 45.07 68.56 45.14 ;
    RECT 68.35 45.43 68.56 45.5 ;
    RECT 28.05 44.71 28.26 44.78 ;
    RECT 28.05 45.07 28.26 45.14 ;
    RECT 28.05 45.43 28.26 45.5 ;
    RECT 28.51 44.71 28.72 44.78 ;
    RECT 28.51 45.07 28.72 45.14 ;
    RECT 28.51 45.43 28.72 45.5 ;
    RECT 24.73 44.71 24.94 44.78 ;
    RECT 24.73 45.07 24.94 45.14 ;
    RECT 24.73 45.43 24.94 45.5 ;
    RECT 25.19 44.71 25.4 44.78 ;
    RECT 25.19 45.07 25.4 45.14 ;
    RECT 25.19 45.43 25.4 45.5 ;
    RECT 21.41 44.71 21.62 44.78 ;
    RECT 21.41 45.07 21.62 45.14 ;
    RECT 21.41 45.43 21.62 45.5 ;
    RECT 21.87 44.71 22.08 44.78 ;
    RECT 21.87 45.07 22.08 45.14 ;
    RECT 21.87 45.43 22.08 45.5 ;
    RECT 18.09 44.71 18.3 44.78 ;
    RECT 18.09 45.07 18.3 45.14 ;
    RECT 18.09 45.43 18.3 45.5 ;
    RECT 18.55 44.71 18.76 44.78 ;
    RECT 18.55 45.07 18.76 45.14 ;
    RECT 18.55 45.43 18.76 45.5 ;
    RECT 120.825 45.07 120.895 45.14 ;
    RECT 14.77 44.71 14.98 44.78 ;
    RECT 14.77 45.07 14.98 45.14 ;
    RECT 14.77 45.43 14.98 45.5 ;
    RECT 15.23 44.71 15.44 44.78 ;
    RECT 15.23 45.07 15.44 45.14 ;
    RECT 15.23 45.43 15.44 45.5 ;
    RECT 11.45 44.71 11.66 44.78 ;
    RECT 11.45 45.07 11.66 45.14 ;
    RECT 11.45 45.43 11.66 45.5 ;
    RECT 11.91 44.71 12.12 44.78 ;
    RECT 11.91 45.07 12.12 45.14 ;
    RECT 11.91 45.43 12.12 45.5 ;
    RECT 8.13 44.71 8.34 44.78 ;
    RECT 8.13 45.07 8.34 45.14 ;
    RECT 8.13 45.43 8.34 45.5 ;
    RECT 8.59 44.71 8.8 44.78 ;
    RECT 8.59 45.07 8.8 45.14 ;
    RECT 8.59 45.43 8.8 45.5 ;
    RECT 4.81 44.71 5.02 44.78 ;
    RECT 4.81 45.07 5.02 45.14 ;
    RECT 4.81 45.43 5.02 45.5 ;
    RECT 5.27 44.71 5.48 44.78 ;
    RECT 5.27 45.07 5.48 45.14 ;
    RECT 5.27 45.43 5.48 45.5 ;
    RECT 1.49 44.71 1.7 44.78 ;
    RECT 1.49 45.07 1.7 45.14 ;
    RECT 1.49 45.43 1.7 45.5 ;
    RECT 1.95 44.71 2.16 44.78 ;
    RECT 1.95 45.07 2.16 45.14 ;
    RECT 1.95 45.43 2.16 45.5 ;
    RECT 64.57 44.71 64.78 44.78 ;
    RECT 64.57 45.07 64.78 45.14 ;
    RECT 64.57 45.43 64.78 45.5 ;
    RECT 65.03 44.71 65.24 44.78 ;
    RECT 65.03 45.07 65.24 45.14 ;
    RECT 65.03 45.43 65.24 45.5 ;
    RECT 61.25 84.33 61.46 84.4 ;
    RECT 61.25 84.69 61.46 84.76 ;
    RECT 61.25 85.05 61.46 85.12 ;
    RECT 61.71 84.33 61.92 84.4 ;
    RECT 61.71 84.69 61.92 84.76 ;
    RECT 61.71 85.05 61.92 85.12 ;
    RECT 57.93 84.33 58.14 84.4 ;
    RECT 57.93 84.69 58.14 84.76 ;
    RECT 57.93 85.05 58.14 85.12 ;
    RECT 58.39 84.33 58.6 84.4 ;
    RECT 58.39 84.69 58.6 84.76 ;
    RECT 58.39 85.05 58.6 85.12 ;
    RECT 54.61 84.33 54.82 84.4 ;
    RECT 54.61 84.69 54.82 84.76 ;
    RECT 54.61 85.05 54.82 85.12 ;
    RECT 55.07 84.33 55.28 84.4 ;
    RECT 55.07 84.69 55.28 84.76 ;
    RECT 55.07 85.05 55.28 85.12 ;
    RECT 51.29 84.33 51.5 84.4 ;
    RECT 51.29 84.69 51.5 84.76 ;
    RECT 51.29 85.05 51.5 85.12 ;
    RECT 51.75 84.33 51.96 84.4 ;
    RECT 51.75 84.69 51.96 84.76 ;
    RECT 51.75 85.05 51.96 85.12 ;
    RECT 47.97 84.33 48.18 84.4 ;
    RECT 47.97 84.69 48.18 84.76 ;
    RECT 47.97 85.05 48.18 85.12 ;
    RECT 48.43 84.33 48.64 84.4 ;
    RECT 48.43 84.69 48.64 84.76 ;
    RECT 48.43 85.05 48.64 85.12 ;
    RECT 44.65 84.33 44.86 84.4 ;
    RECT 44.65 84.69 44.86 84.76 ;
    RECT 44.65 85.05 44.86 85.12 ;
    RECT 45.11 84.33 45.32 84.4 ;
    RECT 45.11 84.69 45.32 84.76 ;
    RECT 45.11 85.05 45.32 85.12 ;
    RECT 41.33 84.33 41.54 84.4 ;
    RECT 41.33 84.69 41.54 84.76 ;
    RECT 41.33 85.05 41.54 85.12 ;
    RECT 41.79 84.33 42.0 84.4 ;
    RECT 41.79 84.69 42.0 84.76 ;
    RECT 41.79 85.05 42.0 85.12 ;
    RECT 38.01 84.33 38.22 84.4 ;
    RECT 38.01 84.69 38.22 84.76 ;
    RECT 38.01 85.05 38.22 85.12 ;
    RECT 38.47 84.33 38.68 84.4 ;
    RECT 38.47 84.69 38.68 84.76 ;
    RECT 38.47 85.05 38.68 85.12 ;
    RECT 0.4 84.69 0.47 84.76 ;
    RECT 34.69 84.33 34.9 84.4 ;
    RECT 34.69 84.69 34.9 84.76 ;
    RECT 34.69 85.05 34.9 85.12 ;
    RECT 35.15 84.33 35.36 84.4 ;
    RECT 35.15 84.69 35.36 84.76 ;
    RECT 35.15 85.05 35.36 85.12 ;
    RECT 117.69 84.33 117.9 84.4 ;
    RECT 117.69 84.69 117.9 84.76 ;
    RECT 117.69 85.05 117.9 85.12 ;
    RECT 118.15 84.33 118.36 84.4 ;
    RECT 118.15 84.69 118.36 84.76 ;
    RECT 118.15 85.05 118.36 85.12 ;
    RECT 114.37 84.33 114.58 84.4 ;
    RECT 114.37 84.69 114.58 84.76 ;
    RECT 114.37 85.05 114.58 85.12 ;
    RECT 114.83 84.33 115.04 84.4 ;
    RECT 114.83 84.69 115.04 84.76 ;
    RECT 114.83 85.05 115.04 85.12 ;
    RECT 111.05 84.33 111.26 84.4 ;
    RECT 111.05 84.69 111.26 84.76 ;
    RECT 111.05 85.05 111.26 85.12 ;
    RECT 111.51 84.33 111.72 84.4 ;
    RECT 111.51 84.69 111.72 84.76 ;
    RECT 111.51 85.05 111.72 85.12 ;
    RECT 107.73 84.33 107.94 84.4 ;
    RECT 107.73 84.69 107.94 84.76 ;
    RECT 107.73 85.05 107.94 85.12 ;
    RECT 108.19 84.33 108.4 84.4 ;
    RECT 108.19 84.69 108.4 84.76 ;
    RECT 108.19 85.05 108.4 85.12 ;
    RECT 104.41 84.33 104.62 84.4 ;
    RECT 104.41 84.69 104.62 84.76 ;
    RECT 104.41 85.05 104.62 85.12 ;
    RECT 104.87 84.33 105.08 84.4 ;
    RECT 104.87 84.69 105.08 84.76 ;
    RECT 104.87 85.05 105.08 85.12 ;
    RECT 101.09 84.33 101.3 84.4 ;
    RECT 101.09 84.69 101.3 84.76 ;
    RECT 101.09 85.05 101.3 85.12 ;
    RECT 101.55 84.33 101.76 84.4 ;
    RECT 101.55 84.69 101.76 84.76 ;
    RECT 101.55 85.05 101.76 85.12 ;
    RECT 97.77 84.33 97.98 84.4 ;
    RECT 97.77 84.69 97.98 84.76 ;
    RECT 97.77 85.05 97.98 85.12 ;
    RECT 98.23 84.33 98.44 84.4 ;
    RECT 98.23 84.69 98.44 84.76 ;
    RECT 98.23 85.05 98.44 85.12 ;
    RECT 94.45 84.33 94.66 84.4 ;
    RECT 94.45 84.69 94.66 84.76 ;
    RECT 94.45 85.05 94.66 85.12 ;
    RECT 94.91 84.33 95.12 84.4 ;
    RECT 94.91 84.69 95.12 84.76 ;
    RECT 94.91 85.05 95.12 85.12 ;
    RECT 91.13 84.33 91.34 84.4 ;
    RECT 91.13 84.69 91.34 84.76 ;
    RECT 91.13 85.05 91.34 85.12 ;
    RECT 91.59 84.33 91.8 84.4 ;
    RECT 91.59 84.69 91.8 84.76 ;
    RECT 91.59 85.05 91.8 85.12 ;
    RECT 87.81 84.33 88.02 84.4 ;
    RECT 87.81 84.69 88.02 84.76 ;
    RECT 87.81 85.05 88.02 85.12 ;
    RECT 88.27 84.33 88.48 84.4 ;
    RECT 88.27 84.69 88.48 84.76 ;
    RECT 88.27 85.05 88.48 85.12 ;
    RECT 84.49 84.33 84.7 84.4 ;
    RECT 84.49 84.69 84.7 84.76 ;
    RECT 84.49 85.05 84.7 85.12 ;
    RECT 84.95 84.33 85.16 84.4 ;
    RECT 84.95 84.69 85.16 84.76 ;
    RECT 84.95 85.05 85.16 85.12 ;
    RECT 81.17 84.33 81.38 84.4 ;
    RECT 81.17 84.69 81.38 84.76 ;
    RECT 81.17 85.05 81.38 85.12 ;
    RECT 81.63 84.33 81.84 84.4 ;
    RECT 81.63 84.69 81.84 84.76 ;
    RECT 81.63 85.05 81.84 85.12 ;
    RECT 77.85 84.33 78.06 84.4 ;
    RECT 77.85 84.69 78.06 84.76 ;
    RECT 77.85 85.05 78.06 85.12 ;
    RECT 78.31 84.33 78.52 84.4 ;
    RECT 78.31 84.69 78.52 84.76 ;
    RECT 78.31 85.05 78.52 85.12 ;
    RECT 74.53 84.33 74.74 84.4 ;
    RECT 74.53 84.69 74.74 84.76 ;
    RECT 74.53 85.05 74.74 85.12 ;
    RECT 74.99 84.33 75.2 84.4 ;
    RECT 74.99 84.69 75.2 84.76 ;
    RECT 74.99 85.05 75.2 85.12 ;
    RECT 71.21 84.33 71.42 84.4 ;
    RECT 71.21 84.69 71.42 84.76 ;
    RECT 71.21 85.05 71.42 85.12 ;
    RECT 71.67 84.33 71.88 84.4 ;
    RECT 71.67 84.69 71.88 84.76 ;
    RECT 71.67 85.05 71.88 85.12 ;
    RECT 31.37 84.33 31.58 84.4 ;
    RECT 31.37 84.69 31.58 84.76 ;
    RECT 31.37 85.05 31.58 85.12 ;
    RECT 31.83 84.33 32.04 84.4 ;
    RECT 31.83 84.69 32.04 84.76 ;
    RECT 31.83 85.05 32.04 85.12 ;
    RECT 67.89 84.33 68.1 84.4 ;
    RECT 67.89 84.69 68.1 84.76 ;
    RECT 67.89 85.05 68.1 85.12 ;
    RECT 68.35 84.33 68.56 84.4 ;
    RECT 68.35 84.69 68.56 84.76 ;
    RECT 68.35 85.05 68.56 85.12 ;
    RECT 28.05 84.33 28.26 84.4 ;
    RECT 28.05 84.69 28.26 84.76 ;
    RECT 28.05 85.05 28.26 85.12 ;
    RECT 28.51 84.33 28.72 84.4 ;
    RECT 28.51 84.69 28.72 84.76 ;
    RECT 28.51 85.05 28.72 85.12 ;
    RECT 24.73 84.33 24.94 84.4 ;
    RECT 24.73 84.69 24.94 84.76 ;
    RECT 24.73 85.05 24.94 85.12 ;
    RECT 25.19 84.33 25.4 84.4 ;
    RECT 25.19 84.69 25.4 84.76 ;
    RECT 25.19 85.05 25.4 85.12 ;
    RECT 21.41 84.33 21.62 84.4 ;
    RECT 21.41 84.69 21.62 84.76 ;
    RECT 21.41 85.05 21.62 85.12 ;
    RECT 21.87 84.33 22.08 84.4 ;
    RECT 21.87 84.69 22.08 84.76 ;
    RECT 21.87 85.05 22.08 85.12 ;
    RECT 18.09 84.33 18.3 84.4 ;
    RECT 18.09 84.69 18.3 84.76 ;
    RECT 18.09 85.05 18.3 85.12 ;
    RECT 18.55 84.33 18.76 84.4 ;
    RECT 18.55 84.69 18.76 84.76 ;
    RECT 18.55 85.05 18.76 85.12 ;
    RECT 120.825 84.69 120.895 84.76 ;
    RECT 14.77 84.33 14.98 84.4 ;
    RECT 14.77 84.69 14.98 84.76 ;
    RECT 14.77 85.05 14.98 85.12 ;
    RECT 15.23 84.33 15.44 84.4 ;
    RECT 15.23 84.69 15.44 84.76 ;
    RECT 15.23 85.05 15.44 85.12 ;
    RECT 11.45 84.33 11.66 84.4 ;
    RECT 11.45 84.69 11.66 84.76 ;
    RECT 11.45 85.05 11.66 85.12 ;
    RECT 11.91 84.33 12.12 84.4 ;
    RECT 11.91 84.69 12.12 84.76 ;
    RECT 11.91 85.05 12.12 85.12 ;
    RECT 8.13 84.33 8.34 84.4 ;
    RECT 8.13 84.69 8.34 84.76 ;
    RECT 8.13 85.05 8.34 85.12 ;
    RECT 8.59 84.33 8.8 84.4 ;
    RECT 8.59 84.69 8.8 84.76 ;
    RECT 8.59 85.05 8.8 85.12 ;
    RECT 4.81 84.33 5.02 84.4 ;
    RECT 4.81 84.69 5.02 84.76 ;
    RECT 4.81 85.05 5.02 85.12 ;
    RECT 5.27 84.33 5.48 84.4 ;
    RECT 5.27 84.69 5.48 84.76 ;
    RECT 5.27 85.05 5.48 85.12 ;
    RECT 1.49 84.33 1.7 84.4 ;
    RECT 1.49 84.69 1.7 84.76 ;
    RECT 1.49 85.05 1.7 85.12 ;
    RECT 1.95 84.33 2.16 84.4 ;
    RECT 1.95 84.69 2.16 84.76 ;
    RECT 1.95 85.05 2.16 85.12 ;
    RECT 64.57 84.33 64.78 84.4 ;
    RECT 64.57 84.69 64.78 84.76 ;
    RECT 64.57 85.05 64.78 85.12 ;
    RECT 65.03 84.33 65.24 84.4 ;
    RECT 65.03 84.69 65.24 84.76 ;
    RECT 65.03 85.05 65.24 85.12 ;
    RECT 61.25 43.99 61.46 44.06 ;
    RECT 61.25 44.35 61.46 44.42 ;
    RECT 61.25 44.71 61.46 44.78 ;
    RECT 61.71 43.99 61.92 44.06 ;
    RECT 61.71 44.35 61.92 44.42 ;
    RECT 61.71 44.71 61.92 44.78 ;
    RECT 57.93 43.99 58.14 44.06 ;
    RECT 57.93 44.35 58.14 44.42 ;
    RECT 57.93 44.71 58.14 44.78 ;
    RECT 58.39 43.99 58.6 44.06 ;
    RECT 58.39 44.35 58.6 44.42 ;
    RECT 58.39 44.71 58.6 44.78 ;
    RECT 54.61 43.99 54.82 44.06 ;
    RECT 54.61 44.35 54.82 44.42 ;
    RECT 54.61 44.71 54.82 44.78 ;
    RECT 55.07 43.99 55.28 44.06 ;
    RECT 55.07 44.35 55.28 44.42 ;
    RECT 55.07 44.71 55.28 44.78 ;
    RECT 51.29 43.99 51.5 44.06 ;
    RECT 51.29 44.35 51.5 44.42 ;
    RECT 51.29 44.71 51.5 44.78 ;
    RECT 51.75 43.99 51.96 44.06 ;
    RECT 51.75 44.35 51.96 44.42 ;
    RECT 51.75 44.71 51.96 44.78 ;
    RECT 47.97 43.99 48.18 44.06 ;
    RECT 47.97 44.35 48.18 44.42 ;
    RECT 47.97 44.71 48.18 44.78 ;
    RECT 48.43 43.99 48.64 44.06 ;
    RECT 48.43 44.35 48.64 44.42 ;
    RECT 48.43 44.71 48.64 44.78 ;
    RECT 44.65 43.99 44.86 44.06 ;
    RECT 44.65 44.35 44.86 44.42 ;
    RECT 44.65 44.71 44.86 44.78 ;
    RECT 45.11 43.99 45.32 44.06 ;
    RECT 45.11 44.35 45.32 44.42 ;
    RECT 45.11 44.71 45.32 44.78 ;
    RECT 41.33 43.99 41.54 44.06 ;
    RECT 41.33 44.35 41.54 44.42 ;
    RECT 41.33 44.71 41.54 44.78 ;
    RECT 41.79 43.99 42.0 44.06 ;
    RECT 41.79 44.35 42.0 44.42 ;
    RECT 41.79 44.71 42.0 44.78 ;
    RECT 38.01 43.99 38.22 44.06 ;
    RECT 38.01 44.35 38.22 44.42 ;
    RECT 38.01 44.71 38.22 44.78 ;
    RECT 38.47 43.99 38.68 44.06 ;
    RECT 38.47 44.35 38.68 44.42 ;
    RECT 38.47 44.71 38.68 44.78 ;
    RECT 0.4 44.35 0.47 44.42 ;
    RECT 34.69 43.99 34.9 44.06 ;
    RECT 34.69 44.35 34.9 44.42 ;
    RECT 34.69 44.71 34.9 44.78 ;
    RECT 35.15 43.99 35.36 44.06 ;
    RECT 35.15 44.35 35.36 44.42 ;
    RECT 35.15 44.71 35.36 44.78 ;
    RECT 117.69 43.99 117.9 44.06 ;
    RECT 117.69 44.35 117.9 44.42 ;
    RECT 117.69 44.71 117.9 44.78 ;
    RECT 118.15 43.99 118.36 44.06 ;
    RECT 118.15 44.35 118.36 44.42 ;
    RECT 118.15 44.71 118.36 44.78 ;
    RECT 114.37 43.99 114.58 44.06 ;
    RECT 114.37 44.35 114.58 44.42 ;
    RECT 114.37 44.71 114.58 44.78 ;
    RECT 114.83 43.99 115.04 44.06 ;
    RECT 114.83 44.35 115.04 44.42 ;
    RECT 114.83 44.71 115.04 44.78 ;
    RECT 111.05 43.99 111.26 44.06 ;
    RECT 111.05 44.35 111.26 44.42 ;
    RECT 111.05 44.71 111.26 44.78 ;
    RECT 111.51 43.99 111.72 44.06 ;
    RECT 111.51 44.35 111.72 44.42 ;
    RECT 111.51 44.71 111.72 44.78 ;
    RECT 107.73 43.99 107.94 44.06 ;
    RECT 107.73 44.35 107.94 44.42 ;
    RECT 107.73 44.71 107.94 44.78 ;
    RECT 108.19 43.99 108.4 44.06 ;
    RECT 108.19 44.35 108.4 44.42 ;
    RECT 108.19 44.71 108.4 44.78 ;
    RECT 104.41 43.99 104.62 44.06 ;
    RECT 104.41 44.35 104.62 44.42 ;
    RECT 104.41 44.71 104.62 44.78 ;
    RECT 104.87 43.99 105.08 44.06 ;
    RECT 104.87 44.35 105.08 44.42 ;
    RECT 104.87 44.71 105.08 44.78 ;
    RECT 101.09 43.99 101.3 44.06 ;
    RECT 101.09 44.35 101.3 44.42 ;
    RECT 101.09 44.71 101.3 44.78 ;
    RECT 101.55 43.99 101.76 44.06 ;
    RECT 101.55 44.35 101.76 44.42 ;
    RECT 101.55 44.71 101.76 44.78 ;
    RECT 97.77 43.99 97.98 44.06 ;
    RECT 97.77 44.35 97.98 44.42 ;
    RECT 97.77 44.71 97.98 44.78 ;
    RECT 98.23 43.99 98.44 44.06 ;
    RECT 98.23 44.35 98.44 44.42 ;
    RECT 98.23 44.71 98.44 44.78 ;
    RECT 94.45 43.99 94.66 44.06 ;
    RECT 94.45 44.35 94.66 44.42 ;
    RECT 94.45 44.71 94.66 44.78 ;
    RECT 94.91 43.99 95.12 44.06 ;
    RECT 94.91 44.35 95.12 44.42 ;
    RECT 94.91 44.71 95.12 44.78 ;
    RECT 91.13 43.99 91.34 44.06 ;
    RECT 91.13 44.35 91.34 44.42 ;
    RECT 91.13 44.71 91.34 44.78 ;
    RECT 91.59 43.99 91.8 44.06 ;
    RECT 91.59 44.35 91.8 44.42 ;
    RECT 91.59 44.71 91.8 44.78 ;
    RECT 87.81 43.99 88.02 44.06 ;
    RECT 87.81 44.35 88.02 44.42 ;
    RECT 87.81 44.71 88.02 44.78 ;
    RECT 88.27 43.99 88.48 44.06 ;
    RECT 88.27 44.35 88.48 44.42 ;
    RECT 88.27 44.71 88.48 44.78 ;
    RECT 84.49 43.99 84.7 44.06 ;
    RECT 84.49 44.35 84.7 44.42 ;
    RECT 84.49 44.71 84.7 44.78 ;
    RECT 84.95 43.99 85.16 44.06 ;
    RECT 84.95 44.35 85.16 44.42 ;
    RECT 84.95 44.71 85.16 44.78 ;
    RECT 81.17 43.99 81.38 44.06 ;
    RECT 81.17 44.35 81.38 44.42 ;
    RECT 81.17 44.71 81.38 44.78 ;
    RECT 81.63 43.99 81.84 44.06 ;
    RECT 81.63 44.35 81.84 44.42 ;
    RECT 81.63 44.71 81.84 44.78 ;
    RECT 77.85 43.99 78.06 44.06 ;
    RECT 77.85 44.35 78.06 44.42 ;
    RECT 77.85 44.71 78.06 44.78 ;
    RECT 78.31 43.99 78.52 44.06 ;
    RECT 78.31 44.35 78.52 44.42 ;
    RECT 78.31 44.71 78.52 44.78 ;
    RECT 74.53 43.99 74.74 44.06 ;
    RECT 74.53 44.35 74.74 44.42 ;
    RECT 74.53 44.71 74.74 44.78 ;
    RECT 74.99 43.99 75.2 44.06 ;
    RECT 74.99 44.35 75.2 44.42 ;
    RECT 74.99 44.71 75.2 44.78 ;
    RECT 71.21 43.99 71.42 44.06 ;
    RECT 71.21 44.35 71.42 44.42 ;
    RECT 71.21 44.71 71.42 44.78 ;
    RECT 71.67 43.99 71.88 44.06 ;
    RECT 71.67 44.35 71.88 44.42 ;
    RECT 71.67 44.71 71.88 44.78 ;
    RECT 31.37 43.99 31.58 44.06 ;
    RECT 31.37 44.35 31.58 44.42 ;
    RECT 31.37 44.71 31.58 44.78 ;
    RECT 31.83 43.99 32.04 44.06 ;
    RECT 31.83 44.35 32.04 44.42 ;
    RECT 31.83 44.71 32.04 44.78 ;
    RECT 67.89 43.99 68.1 44.06 ;
    RECT 67.89 44.35 68.1 44.42 ;
    RECT 67.89 44.71 68.1 44.78 ;
    RECT 68.35 43.99 68.56 44.06 ;
    RECT 68.35 44.35 68.56 44.42 ;
    RECT 68.35 44.71 68.56 44.78 ;
    RECT 28.05 43.99 28.26 44.06 ;
    RECT 28.05 44.35 28.26 44.42 ;
    RECT 28.05 44.71 28.26 44.78 ;
    RECT 28.51 43.99 28.72 44.06 ;
    RECT 28.51 44.35 28.72 44.42 ;
    RECT 28.51 44.71 28.72 44.78 ;
    RECT 24.73 43.99 24.94 44.06 ;
    RECT 24.73 44.35 24.94 44.42 ;
    RECT 24.73 44.71 24.94 44.78 ;
    RECT 25.19 43.99 25.4 44.06 ;
    RECT 25.19 44.35 25.4 44.42 ;
    RECT 25.19 44.71 25.4 44.78 ;
    RECT 21.41 43.99 21.62 44.06 ;
    RECT 21.41 44.35 21.62 44.42 ;
    RECT 21.41 44.71 21.62 44.78 ;
    RECT 21.87 43.99 22.08 44.06 ;
    RECT 21.87 44.35 22.08 44.42 ;
    RECT 21.87 44.71 22.08 44.78 ;
    RECT 18.09 43.99 18.3 44.06 ;
    RECT 18.09 44.35 18.3 44.42 ;
    RECT 18.09 44.71 18.3 44.78 ;
    RECT 18.55 43.99 18.76 44.06 ;
    RECT 18.55 44.35 18.76 44.42 ;
    RECT 18.55 44.71 18.76 44.78 ;
    RECT 120.825 44.35 120.895 44.42 ;
    RECT 14.77 43.99 14.98 44.06 ;
    RECT 14.77 44.35 14.98 44.42 ;
    RECT 14.77 44.71 14.98 44.78 ;
    RECT 15.23 43.99 15.44 44.06 ;
    RECT 15.23 44.35 15.44 44.42 ;
    RECT 15.23 44.71 15.44 44.78 ;
    RECT 11.45 43.99 11.66 44.06 ;
    RECT 11.45 44.35 11.66 44.42 ;
    RECT 11.45 44.71 11.66 44.78 ;
    RECT 11.91 43.99 12.12 44.06 ;
    RECT 11.91 44.35 12.12 44.42 ;
    RECT 11.91 44.71 12.12 44.78 ;
    RECT 8.13 43.99 8.34 44.06 ;
    RECT 8.13 44.35 8.34 44.42 ;
    RECT 8.13 44.71 8.34 44.78 ;
    RECT 8.59 43.99 8.8 44.06 ;
    RECT 8.59 44.35 8.8 44.42 ;
    RECT 8.59 44.71 8.8 44.78 ;
    RECT 4.81 43.99 5.02 44.06 ;
    RECT 4.81 44.35 5.02 44.42 ;
    RECT 4.81 44.71 5.02 44.78 ;
    RECT 5.27 43.99 5.48 44.06 ;
    RECT 5.27 44.35 5.48 44.42 ;
    RECT 5.27 44.71 5.48 44.78 ;
    RECT 1.49 43.99 1.7 44.06 ;
    RECT 1.49 44.35 1.7 44.42 ;
    RECT 1.49 44.71 1.7 44.78 ;
    RECT 1.95 43.99 2.16 44.06 ;
    RECT 1.95 44.35 2.16 44.42 ;
    RECT 1.95 44.71 2.16 44.78 ;
    RECT 64.57 43.99 64.78 44.06 ;
    RECT 64.57 44.35 64.78 44.42 ;
    RECT 64.57 44.71 64.78 44.78 ;
    RECT 65.03 43.99 65.24 44.06 ;
    RECT 65.03 44.35 65.24 44.42 ;
    RECT 65.03 44.71 65.24 44.78 ;
    RECT 61.25 83.61 61.46 83.68 ;
    RECT 61.25 83.97 61.46 84.04 ;
    RECT 61.25 84.33 61.46 84.4 ;
    RECT 61.71 83.61 61.92 83.68 ;
    RECT 61.71 83.97 61.92 84.04 ;
    RECT 61.71 84.33 61.92 84.4 ;
    RECT 57.93 83.61 58.14 83.68 ;
    RECT 57.93 83.97 58.14 84.04 ;
    RECT 57.93 84.33 58.14 84.4 ;
    RECT 58.39 83.61 58.6 83.68 ;
    RECT 58.39 83.97 58.6 84.04 ;
    RECT 58.39 84.33 58.6 84.4 ;
    RECT 54.61 83.61 54.82 83.68 ;
    RECT 54.61 83.97 54.82 84.04 ;
    RECT 54.61 84.33 54.82 84.4 ;
    RECT 55.07 83.61 55.28 83.68 ;
    RECT 55.07 83.97 55.28 84.04 ;
    RECT 55.07 84.33 55.28 84.4 ;
    RECT 51.29 83.61 51.5 83.68 ;
    RECT 51.29 83.97 51.5 84.04 ;
    RECT 51.29 84.33 51.5 84.4 ;
    RECT 51.75 83.61 51.96 83.68 ;
    RECT 51.75 83.97 51.96 84.04 ;
    RECT 51.75 84.33 51.96 84.4 ;
    RECT 47.97 83.61 48.18 83.68 ;
    RECT 47.97 83.97 48.18 84.04 ;
    RECT 47.97 84.33 48.18 84.4 ;
    RECT 48.43 83.61 48.64 83.68 ;
    RECT 48.43 83.97 48.64 84.04 ;
    RECT 48.43 84.33 48.64 84.4 ;
    RECT 44.65 83.61 44.86 83.68 ;
    RECT 44.65 83.97 44.86 84.04 ;
    RECT 44.65 84.33 44.86 84.4 ;
    RECT 45.11 83.61 45.32 83.68 ;
    RECT 45.11 83.97 45.32 84.04 ;
    RECT 45.11 84.33 45.32 84.4 ;
    RECT 41.33 83.61 41.54 83.68 ;
    RECT 41.33 83.97 41.54 84.04 ;
    RECT 41.33 84.33 41.54 84.4 ;
    RECT 41.79 83.61 42.0 83.68 ;
    RECT 41.79 83.97 42.0 84.04 ;
    RECT 41.79 84.33 42.0 84.4 ;
    RECT 38.01 83.61 38.22 83.68 ;
    RECT 38.01 83.97 38.22 84.04 ;
    RECT 38.01 84.33 38.22 84.4 ;
    RECT 38.47 83.61 38.68 83.68 ;
    RECT 38.47 83.97 38.68 84.04 ;
    RECT 38.47 84.33 38.68 84.4 ;
    RECT 0.4 83.97 0.47 84.04 ;
    RECT 34.69 83.61 34.9 83.68 ;
    RECT 34.69 83.97 34.9 84.04 ;
    RECT 34.69 84.33 34.9 84.4 ;
    RECT 35.15 83.61 35.36 83.68 ;
    RECT 35.15 83.97 35.36 84.04 ;
    RECT 35.15 84.33 35.36 84.4 ;
    RECT 117.69 83.61 117.9 83.68 ;
    RECT 117.69 83.97 117.9 84.04 ;
    RECT 117.69 84.33 117.9 84.4 ;
    RECT 118.15 83.61 118.36 83.68 ;
    RECT 118.15 83.97 118.36 84.04 ;
    RECT 118.15 84.33 118.36 84.4 ;
    RECT 114.37 83.61 114.58 83.68 ;
    RECT 114.37 83.97 114.58 84.04 ;
    RECT 114.37 84.33 114.58 84.4 ;
    RECT 114.83 83.61 115.04 83.68 ;
    RECT 114.83 83.97 115.04 84.04 ;
    RECT 114.83 84.33 115.04 84.4 ;
    RECT 111.05 83.61 111.26 83.68 ;
    RECT 111.05 83.97 111.26 84.04 ;
    RECT 111.05 84.33 111.26 84.4 ;
    RECT 111.51 83.61 111.72 83.68 ;
    RECT 111.51 83.97 111.72 84.04 ;
    RECT 111.51 84.33 111.72 84.4 ;
    RECT 107.73 83.61 107.94 83.68 ;
    RECT 107.73 83.97 107.94 84.04 ;
    RECT 107.73 84.33 107.94 84.4 ;
    RECT 108.19 83.61 108.4 83.68 ;
    RECT 108.19 83.97 108.4 84.04 ;
    RECT 108.19 84.33 108.4 84.4 ;
    RECT 104.41 83.61 104.62 83.68 ;
    RECT 104.41 83.97 104.62 84.04 ;
    RECT 104.41 84.33 104.62 84.4 ;
    RECT 104.87 83.61 105.08 83.68 ;
    RECT 104.87 83.97 105.08 84.04 ;
    RECT 104.87 84.33 105.08 84.4 ;
    RECT 101.09 83.61 101.3 83.68 ;
    RECT 101.09 83.97 101.3 84.04 ;
    RECT 101.09 84.33 101.3 84.4 ;
    RECT 101.55 83.61 101.76 83.68 ;
    RECT 101.55 83.97 101.76 84.04 ;
    RECT 101.55 84.33 101.76 84.4 ;
    RECT 97.77 83.61 97.98 83.68 ;
    RECT 97.77 83.97 97.98 84.04 ;
    RECT 97.77 84.33 97.98 84.4 ;
    RECT 98.23 83.61 98.44 83.68 ;
    RECT 98.23 83.97 98.44 84.04 ;
    RECT 98.23 84.33 98.44 84.4 ;
    RECT 94.45 83.61 94.66 83.68 ;
    RECT 94.45 83.97 94.66 84.04 ;
    RECT 94.45 84.33 94.66 84.4 ;
    RECT 94.91 83.61 95.12 83.68 ;
    RECT 94.91 83.97 95.12 84.04 ;
    RECT 94.91 84.33 95.12 84.4 ;
    RECT 91.13 83.61 91.34 83.68 ;
    RECT 91.13 83.97 91.34 84.04 ;
    RECT 91.13 84.33 91.34 84.4 ;
    RECT 91.59 83.61 91.8 83.68 ;
    RECT 91.59 83.97 91.8 84.04 ;
    RECT 91.59 84.33 91.8 84.4 ;
    RECT 87.81 83.61 88.02 83.68 ;
    RECT 87.81 83.97 88.02 84.04 ;
    RECT 87.81 84.33 88.02 84.4 ;
    RECT 88.27 83.61 88.48 83.68 ;
    RECT 88.27 83.97 88.48 84.04 ;
    RECT 88.27 84.33 88.48 84.4 ;
    RECT 84.49 83.61 84.7 83.68 ;
    RECT 84.49 83.97 84.7 84.04 ;
    RECT 84.49 84.33 84.7 84.4 ;
    RECT 84.95 83.61 85.16 83.68 ;
    RECT 84.95 83.97 85.16 84.04 ;
    RECT 84.95 84.33 85.16 84.4 ;
    RECT 81.17 83.61 81.38 83.68 ;
    RECT 81.17 83.97 81.38 84.04 ;
    RECT 81.17 84.33 81.38 84.4 ;
    RECT 81.63 83.61 81.84 83.68 ;
    RECT 81.63 83.97 81.84 84.04 ;
    RECT 81.63 84.33 81.84 84.4 ;
    RECT 77.85 83.61 78.06 83.68 ;
    RECT 77.85 83.97 78.06 84.04 ;
    RECT 77.85 84.33 78.06 84.4 ;
    RECT 78.31 83.61 78.52 83.68 ;
    RECT 78.31 83.97 78.52 84.04 ;
    RECT 78.31 84.33 78.52 84.4 ;
    RECT 74.53 83.61 74.74 83.68 ;
    RECT 74.53 83.97 74.74 84.04 ;
    RECT 74.53 84.33 74.74 84.4 ;
    RECT 74.99 83.61 75.2 83.68 ;
    RECT 74.99 83.97 75.2 84.04 ;
    RECT 74.99 84.33 75.2 84.4 ;
    RECT 71.21 83.61 71.42 83.68 ;
    RECT 71.21 83.97 71.42 84.04 ;
    RECT 71.21 84.33 71.42 84.4 ;
    RECT 71.67 83.61 71.88 83.68 ;
    RECT 71.67 83.97 71.88 84.04 ;
    RECT 71.67 84.33 71.88 84.4 ;
    RECT 31.37 83.61 31.58 83.68 ;
    RECT 31.37 83.97 31.58 84.04 ;
    RECT 31.37 84.33 31.58 84.4 ;
    RECT 31.83 83.61 32.04 83.68 ;
    RECT 31.83 83.97 32.04 84.04 ;
    RECT 31.83 84.33 32.04 84.4 ;
    RECT 67.89 83.61 68.1 83.68 ;
    RECT 67.89 83.97 68.1 84.04 ;
    RECT 67.89 84.33 68.1 84.4 ;
    RECT 68.35 83.61 68.56 83.68 ;
    RECT 68.35 83.97 68.56 84.04 ;
    RECT 68.35 84.33 68.56 84.4 ;
    RECT 28.05 83.61 28.26 83.68 ;
    RECT 28.05 83.97 28.26 84.04 ;
    RECT 28.05 84.33 28.26 84.4 ;
    RECT 28.51 83.61 28.72 83.68 ;
    RECT 28.51 83.97 28.72 84.04 ;
    RECT 28.51 84.33 28.72 84.4 ;
    RECT 24.73 83.61 24.94 83.68 ;
    RECT 24.73 83.97 24.94 84.04 ;
    RECT 24.73 84.33 24.94 84.4 ;
    RECT 25.19 83.61 25.4 83.68 ;
    RECT 25.19 83.97 25.4 84.04 ;
    RECT 25.19 84.33 25.4 84.4 ;
    RECT 21.41 83.61 21.62 83.68 ;
    RECT 21.41 83.97 21.62 84.04 ;
    RECT 21.41 84.33 21.62 84.4 ;
    RECT 21.87 83.61 22.08 83.68 ;
    RECT 21.87 83.97 22.08 84.04 ;
    RECT 21.87 84.33 22.08 84.4 ;
    RECT 18.09 83.61 18.3 83.68 ;
    RECT 18.09 83.97 18.3 84.04 ;
    RECT 18.09 84.33 18.3 84.4 ;
    RECT 18.55 83.61 18.76 83.68 ;
    RECT 18.55 83.97 18.76 84.04 ;
    RECT 18.55 84.33 18.76 84.4 ;
    RECT 120.825 83.97 120.895 84.04 ;
    RECT 14.77 83.61 14.98 83.68 ;
    RECT 14.77 83.97 14.98 84.04 ;
    RECT 14.77 84.33 14.98 84.4 ;
    RECT 15.23 83.61 15.44 83.68 ;
    RECT 15.23 83.97 15.44 84.04 ;
    RECT 15.23 84.33 15.44 84.4 ;
    RECT 11.45 83.61 11.66 83.68 ;
    RECT 11.45 83.97 11.66 84.04 ;
    RECT 11.45 84.33 11.66 84.4 ;
    RECT 11.91 83.61 12.12 83.68 ;
    RECT 11.91 83.97 12.12 84.04 ;
    RECT 11.91 84.33 12.12 84.4 ;
    RECT 8.13 83.61 8.34 83.68 ;
    RECT 8.13 83.97 8.34 84.04 ;
    RECT 8.13 84.33 8.34 84.4 ;
    RECT 8.59 83.61 8.8 83.68 ;
    RECT 8.59 83.97 8.8 84.04 ;
    RECT 8.59 84.33 8.8 84.4 ;
    RECT 4.81 83.61 5.02 83.68 ;
    RECT 4.81 83.97 5.02 84.04 ;
    RECT 4.81 84.33 5.02 84.4 ;
    RECT 5.27 83.61 5.48 83.68 ;
    RECT 5.27 83.97 5.48 84.04 ;
    RECT 5.27 84.33 5.48 84.4 ;
    RECT 1.49 83.61 1.7 83.68 ;
    RECT 1.49 83.97 1.7 84.04 ;
    RECT 1.49 84.33 1.7 84.4 ;
    RECT 1.95 83.61 2.16 83.68 ;
    RECT 1.95 83.97 2.16 84.04 ;
    RECT 1.95 84.33 2.16 84.4 ;
    RECT 64.57 83.61 64.78 83.68 ;
    RECT 64.57 83.97 64.78 84.04 ;
    RECT 64.57 84.33 64.78 84.4 ;
    RECT 65.03 83.61 65.24 83.68 ;
    RECT 65.03 83.97 65.24 84.04 ;
    RECT 65.03 84.33 65.24 84.4 ;
    RECT 61.25 43.27 61.46 43.34 ;
    RECT 61.25 43.63 61.46 43.7 ;
    RECT 61.25 43.99 61.46 44.06 ;
    RECT 61.71 43.27 61.92 43.34 ;
    RECT 61.71 43.63 61.92 43.7 ;
    RECT 61.71 43.99 61.92 44.06 ;
    RECT 57.93 43.27 58.14 43.34 ;
    RECT 57.93 43.63 58.14 43.7 ;
    RECT 57.93 43.99 58.14 44.06 ;
    RECT 58.39 43.27 58.6 43.34 ;
    RECT 58.39 43.63 58.6 43.7 ;
    RECT 58.39 43.99 58.6 44.06 ;
    RECT 54.61 43.27 54.82 43.34 ;
    RECT 54.61 43.63 54.82 43.7 ;
    RECT 54.61 43.99 54.82 44.06 ;
    RECT 55.07 43.27 55.28 43.34 ;
    RECT 55.07 43.63 55.28 43.7 ;
    RECT 55.07 43.99 55.28 44.06 ;
    RECT 51.29 43.27 51.5 43.34 ;
    RECT 51.29 43.63 51.5 43.7 ;
    RECT 51.29 43.99 51.5 44.06 ;
    RECT 51.75 43.27 51.96 43.34 ;
    RECT 51.75 43.63 51.96 43.7 ;
    RECT 51.75 43.99 51.96 44.06 ;
    RECT 47.97 43.27 48.18 43.34 ;
    RECT 47.97 43.63 48.18 43.7 ;
    RECT 47.97 43.99 48.18 44.06 ;
    RECT 48.43 43.27 48.64 43.34 ;
    RECT 48.43 43.63 48.64 43.7 ;
    RECT 48.43 43.99 48.64 44.06 ;
    RECT 44.65 43.27 44.86 43.34 ;
    RECT 44.65 43.63 44.86 43.7 ;
    RECT 44.65 43.99 44.86 44.06 ;
    RECT 45.11 43.27 45.32 43.34 ;
    RECT 45.11 43.63 45.32 43.7 ;
    RECT 45.11 43.99 45.32 44.06 ;
    RECT 41.33 43.27 41.54 43.34 ;
    RECT 41.33 43.63 41.54 43.7 ;
    RECT 41.33 43.99 41.54 44.06 ;
    RECT 41.79 43.27 42.0 43.34 ;
    RECT 41.79 43.63 42.0 43.7 ;
    RECT 41.79 43.99 42.0 44.06 ;
    RECT 38.01 43.27 38.22 43.34 ;
    RECT 38.01 43.63 38.22 43.7 ;
    RECT 38.01 43.99 38.22 44.06 ;
    RECT 38.47 43.27 38.68 43.34 ;
    RECT 38.47 43.63 38.68 43.7 ;
    RECT 38.47 43.99 38.68 44.06 ;
    RECT 0.4 43.63 0.47 43.7 ;
    RECT 34.69 43.27 34.9 43.34 ;
    RECT 34.69 43.63 34.9 43.7 ;
    RECT 34.69 43.99 34.9 44.06 ;
    RECT 35.15 43.27 35.36 43.34 ;
    RECT 35.15 43.63 35.36 43.7 ;
    RECT 35.15 43.99 35.36 44.06 ;
    RECT 117.69 43.27 117.9 43.34 ;
    RECT 117.69 43.63 117.9 43.7 ;
    RECT 117.69 43.99 117.9 44.06 ;
    RECT 118.15 43.27 118.36 43.34 ;
    RECT 118.15 43.63 118.36 43.7 ;
    RECT 118.15 43.99 118.36 44.06 ;
    RECT 114.37 43.27 114.58 43.34 ;
    RECT 114.37 43.63 114.58 43.7 ;
    RECT 114.37 43.99 114.58 44.06 ;
    RECT 114.83 43.27 115.04 43.34 ;
    RECT 114.83 43.63 115.04 43.7 ;
    RECT 114.83 43.99 115.04 44.06 ;
    RECT 111.05 43.27 111.26 43.34 ;
    RECT 111.05 43.63 111.26 43.7 ;
    RECT 111.05 43.99 111.26 44.06 ;
    RECT 111.51 43.27 111.72 43.34 ;
    RECT 111.51 43.63 111.72 43.7 ;
    RECT 111.51 43.99 111.72 44.06 ;
    RECT 107.73 43.27 107.94 43.34 ;
    RECT 107.73 43.63 107.94 43.7 ;
    RECT 107.73 43.99 107.94 44.06 ;
    RECT 108.19 43.27 108.4 43.34 ;
    RECT 108.19 43.63 108.4 43.7 ;
    RECT 108.19 43.99 108.4 44.06 ;
    RECT 104.41 43.27 104.62 43.34 ;
    RECT 104.41 43.63 104.62 43.7 ;
    RECT 104.41 43.99 104.62 44.06 ;
    RECT 104.87 43.27 105.08 43.34 ;
    RECT 104.87 43.63 105.08 43.7 ;
    RECT 104.87 43.99 105.08 44.06 ;
    RECT 101.09 43.27 101.3 43.34 ;
    RECT 101.09 43.63 101.3 43.7 ;
    RECT 101.09 43.99 101.3 44.06 ;
    RECT 101.55 43.27 101.76 43.34 ;
    RECT 101.55 43.63 101.76 43.7 ;
    RECT 101.55 43.99 101.76 44.06 ;
    RECT 97.77 43.27 97.98 43.34 ;
    RECT 97.77 43.63 97.98 43.7 ;
    RECT 97.77 43.99 97.98 44.06 ;
    RECT 98.23 43.27 98.44 43.34 ;
    RECT 98.23 43.63 98.44 43.7 ;
    RECT 98.23 43.99 98.44 44.06 ;
    RECT 94.45 43.27 94.66 43.34 ;
    RECT 94.45 43.63 94.66 43.7 ;
    RECT 94.45 43.99 94.66 44.06 ;
    RECT 94.91 43.27 95.12 43.34 ;
    RECT 94.91 43.63 95.12 43.7 ;
    RECT 94.91 43.99 95.12 44.06 ;
    RECT 91.13 43.27 91.34 43.34 ;
    RECT 91.13 43.63 91.34 43.7 ;
    RECT 91.13 43.99 91.34 44.06 ;
    RECT 91.59 43.27 91.8 43.34 ;
    RECT 91.59 43.63 91.8 43.7 ;
    RECT 91.59 43.99 91.8 44.06 ;
    RECT 87.81 43.27 88.02 43.34 ;
    RECT 87.81 43.63 88.02 43.7 ;
    RECT 87.81 43.99 88.02 44.06 ;
    RECT 88.27 43.27 88.48 43.34 ;
    RECT 88.27 43.63 88.48 43.7 ;
    RECT 88.27 43.99 88.48 44.06 ;
    RECT 84.49 43.27 84.7 43.34 ;
    RECT 84.49 43.63 84.7 43.7 ;
    RECT 84.49 43.99 84.7 44.06 ;
    RECT 84.95 43.27 85.16 43.34 ;
    RECT 84.95 43.63 85.16 43.7 ;
    RECT 84.95 43.99 85.16 44.06 ;
    RECT 81.17 43.27 81.38 43.34 ;
    RECT 81.17 43.63 81.38 43.7 ;
    RECT 81.17 43.99 81.38 44.06 ;
    RECT 81.63 43.27 81.84 43.34 ;
    RECT 81.63 43.63 81.84 43.7 ;
    RECT 81.63 43.99 81.84 44.06 ;
    RECT 77.85 43.27 78.06 43.34 ;
    RECT 77.85 43.63 78.06 43.7 ;
    RECT 77.85 43.99 78.06 44.06 ;
    RECT 78.31 43.27 78.52 43.34 ;
    RECT 78.31 43.63 78.52 43.7 ;
    RECT 78.31 43.99 78.52 44.06 ;
    RECT 74.53 43.27 74.74 43.34 ;
    RECT 74.53 43.63 74.74 43.7 ;
    RECT 74.53 43.99 74.74 44.06 ;
    RECT 74.99 43.27 75.2 43.34 ;
    RECT 74.99 43.63 75.2 43.7 ;
    RECT 74.99 43.99 75.2 44.06 ;
    RECT 71.21 43.27 71.42 43.34 ;
    RECT 71.21 43.63 71.42 43.7 ;
    RECT 71.21 43.99 71.42 44.06 ;
    RECT 71.67 43.27 71.88 43.34 ;
    RECT 71.67 43.63 71.88 43.7 ;
    RECT 71.67 43.99 71.88 44.06 ;
    RECT 31.37 43.27 31.58 43.34 ;
    RECT 31.37 43.63 31.58 43.7 ;
    RECT 31.37 43.99 31.58 44.06 ;
    RECT 31.83 43.27 32.04 43.34 ;
    RECT 31.83 43.63 32.04 43.7 ;
    RECT 31.83 43.99 32.04 44.06 ;
    RECT 67.89 43.27 68.1 43.34 ;
    RECT 67.89 43.63 68.1 43.7 ;
    RECT 67.89 43.99 68.1 44.06 ;
    RECT 68.35 43.27 68.56 43.34 ;
    RECT 68.35 43.63 68.56 43.7 ;
    RECT 68.35 43.99 68.56 44.06 ;
    RECT 28.05 43.27 28.26 43.34 ;
    RECT 28.05 43.63 28.26 43.7 ;
    RECT 28.05 43.99 28.26 44.06 ;
    RECT 28.51 43.27 28.72 43.34 ;
    RECT 28.51 43.63 28.72 43.7 ;
    RECT 28.51 43.99 28.72 44.06 ;
    RECT 24.73 43.27 24.94 43.34 ;
    RECT 24.73 43.63 24.94 43.7 ;
    RECT 24.73 43.99 24.94 44.06 ;
    RECT 25.19 43.27 25.4 43.34 ;
    RECT 25.19 43.63 25.4 43.7 ;
    RECT 25.19 43.99 25.4 44.06 ;
    RECT 21.41 43.27 21.62 43.34 ;
    RECT 21.41 43.63 21.62 43.7 ;
    RECT 21.41 43.99 21.62 44.06 ;
    RECT 21.87 43.27 22.08 43.34 ;
    RECT 21.87 43.63 22.08 43.7 ;
    RECT 21.87 43.99 22.08 44.06 ;
    RECT 18.09 43.27 18.3 43.34 ;
    RECT 18.09 43.63 18.3 43.7 ;
    RECT 18.09 43.99 18.3 44.06 ;
    RECT 18.55 43.27 18.76 43.34 ;
    RECT 18.55 43.63 18.76 43.7 ;
    RECT 18.55 43.99 18.76 44.06 ;
    RECT 120.825 43.63 120.895 43.7 ;
    RECT 14.77 43.27 14.98 43.34 ;
    RECT 14.77 43.63 14.98 43.7 ;
    RECT 14.77 43.99 14.98 44.06 ;
    RECT 15.23 43.27 15.44 43.34 ;
    RECT 15.23 43.63 15.44 43.7 ;
    RECT 15.23 43.99 15.44 44.06 ;
    RECT 11.45 43.27 11.66 43.34 ;
    RECT 11.45 43.63 11.66 43.7 ;
    RECT 11.45 43.99 11.66 44.06 ;
    RECT 11.91 43.27 12.12 43.34 ;
    RECT 11.91 43.63 12.12 43.7 ;
    RECT 11.91 43.99 12.12 44.06 ;
    RECT 8.13 43.27 8.34 43.34 ;
    RECT 8.13 43.63 8.34 43.7 ;
    RECT 8.13 43.99 8.34 44.06 ;
    RECT 8.59 43.27 8.8 43.34 ;
    RECT 8.59 43.63 8.8 43.7 ;
    RECT 8.59 43.99 8.8 44.06 ;
    RECT 4.81 43.27 5.02 43.34 ;
    RECT 4.81 43.63 5.02 43.7 ;
    RECT 4.81 43.99 5.02 44.06 ;
    RECT 5.27 43.27 5.48 43.34 ;
    RECT 5.27 43.63 5.48 43.7 ;
    RECT 5.27 43.99 5.48 44.06 ;
    RECT 1.49 43.27 1.7 43.34 ;
    RECT 1.49 43.63 1.7 43.7 ;
    RECT 1.49 43.99 1.7 44.06 ;
    RECT 1.95 43.27 2.16 43.34 ;
    RECT 1.95 43.63 2.16 43.7 ;
    RECT 1.95 43.99 2.16 44.06 ;
    RECT 64.57 43.27 64.78 43.34 ;
    RECT 64.57 43.63 64.78 43.7 ;
    RECT 64.57 43.99 64.78 44.06 ;
    RECT 65.03 43.27 65.24 43.34 ;
    RECT 65.03 43.63 65.24 43.7 ;
    RECT 65.03 43.99 65.24 44.06 ;
    RECT 61.25 82.89 61.46 82.96 ;
    RECT 61.25 83.25 61.46 83.32 ;
    RECT 61.25 83.61 61.46 83.68 ;
    RECT 61.71 82.89 61.92 82.96 ;
    RECT 61.71 83.25 61.92 83.32 ;
    RECT 61.71 83.61 61.92 83.68 ;
    RECT 57.93 82.89 58.14 82.96 ;
    RECT 57.93 83.25 58.14 83.32 ;
    RECT 57.93 83.61 58.14 83.68 ;
    RECT 58.39 82.89 58.6 82.96 ;
    RECT 58.39 83.25 58.6 83.32 ;
    RECT 58.39 83.61 58.6 83.68 ;
    RECT 54.61 82.89 54.82 82.96 ;
    RECT 54.61 83.25 54.82 83.32 ;
    RECT 54.61 83.61 54.82 83.68 ;
    RECT 55.07 82.89 55.28 82.96 ;
    RECT 55.07 83.25 55.28 83.32 ;
    RECT 55.07 83.61 55.28 83.68 ;
    RECT 51.29 82.89 51.5 82.96 ;
    RECT 51.29 83.25 51.5 83.32 ;
    RECT 51.29 83.61 51.5 83.68 ;
    RECT 51.75 82.89 51.96 82.96 ;
    RECT 51.75 83.25 51.96 83.32 ;
    RECT 51.75 83.61 51.96 83.68 ;
    RECT 47.97 82.89 48.18 82.96 ;
    RECT 47.97 83.25 48.18 83.32 ;
    RECT 47.97 83.61 48.18 83.68 ;
    RECT 48.43 82.89 48.64 82.96 ;
    RECT 48.43 83.25 48.64 83.32 ;
    RECT 48.43 83.61 48.64 83.68 ;
    RECT 44.65 82.89 44.86 82.96 ;
    RECT 44.65 83.25 44.86 83.32 ;
    RECT 44.65 83.61 44.86 83.68 ;
    RECT 45.11 82.89 45.32 82.96 ;
    RECT 45.11 83.25 45.32 83.32 ;
    RECT 45.11 83.61 45.32 83.68 ;
    RECT 41.33 82.89 41.54 82.96 ;
    RECT 41.33 83.25 41.54 83.32 ;
    RECT 41.33 83.61 41.54 83.68 ;
    RECT 41.79 82.89 42.0 82.96 ;
    RECT 41.79 83.25 42.0 83.32 ;
    RECT 41.79 83.61 42.0 83.68 ;
    RECT 38.01 82.89 38.22 82.96 ;
    RECT 38.01 83.25 38.22 83.32 ;
    RECT 38.01 83.61 38.22 83.68 ;
    RECT 38.47 82.89 38.68 82.96 ;
    RECT 38.47 83.25 38.68 83.32 ;
    RECT 38.47 83.61 38.68 83.68 ;
    RECT 0.4 83.25 0.47 83.32 ;
    RECT 34.69 82.89 34.9 82.96 ;
    RECT 34.69 83.25 34.9 83.32 ;
    RECT 34.69 83.61 34.9 83.68 ;
    RECT 35.15 82.89 35.36 82.96 ;
    RECT 35.15 83.25 35.36 83.32 ;
    RECT 35.15 83.61 35.36 83.68 ;
    RECT 117.69 82.89 117.9 82.96 ;
    RECT 117.69 83.25 117.9 83.32 ;
    RECT 117.69 83.61 117.9 83.68 ;
    RECT 118.15 82.89 118.36 82.96 ;
    RECT 118.15 83.25 118.36 83.32 ;
    RECT 118.15 83.61 118.36 83.68 ;
    RECT 114.37 82.89 114.58 82.96 ;
    RECT 114.37 83.25 114.58 83.32 ;
    RECT 114.37 83.61 114.58 83.68 ;
    RECT 114.83 82.89 115.04 82.96 ;
    RECT 114.83 83.25 115.04 83.32 ;
    RECT 114.83 83.61 115.04 83.68 ;
    RECT 111.05 82.89 111.26 82.96 ;
    RECT 111.05 83.25 111.26 83.32 ;
    RECT 111.05 83.61 111.26 83.68 ;
    RECT 111.51 82.89 111.72 82.96 ;
    RECT 111.51 83.25 111.72 83.32 ;
    RECT 111.51 83.61 111.72 83.68 ;
    RECT 107.73 82.89 107.94 82.96 ;
    RECT 107.73 83.25 107.94 83.32 ;
    RECT 107.73 83.61 107.94 83.68 ;
    RECT 108.19 82.89 108.4 82.96 ;
    RECT 108.19 83.25 108.4 83.32 ;
    RECT 108.19 83.61 108.4 83.68 ;
    RECT 104.41 82.89 104.62 82.96 ;
    RECT 104.41 83.25 104.62 83.32 ;
    RECT 104.41 83.61 104.62 83.68 ;
    RECT 104.87 82.89 105.08 82.96 ;
    RECT 104.87 83.25 105.08 83.32 ;
    RECT 104.87 83.61 105.08 83.68 ;
    RECT 101.09 82.89 101.3 82.96 ;
    RECT 101.09 83.25 101.3 83.32 ;
    RECT 101.09 83.61 101.3 83.68 ;
    RECT 101.55 82.89 101.76 82.96 ;
    RECT 101.55 83.25 101.76 83.32 ;
    RECT 101.55 83.61 101.76 83.68 ;
    RECT 97.77 82.89 97.98 82.96 ;
    RECT 97.77 83.25 97.98 83.32 ;
    RECT 97.77 83.61 97.98 83.68 ;
    RECT 98.23 82.89 98.44 82.96 ;
    RECT 98.23 83.25 98.44 83.32 ;
    RECT 98.23 83.61 98.44 83.68 ;
    RECT 94.45 82.89 94.66 82.96 ;
    RECT 94.45 83.25 94.66 83.32 ;
    RECT 94.45 83.61 94.66 83.68 ;
    RECT 94.91 82.89 95.12 82.96 ;
    RECT 94.91 83.25 95.12 83.32 ;
    RECT 94.91 83.61 95.12 83.68 ;
    RECT 91.13 82.89 91.34 82.96 ;
    RECT 91.13 83.25 91.34 83.32 ;
    RECT 91.13 83.61 91.34 83.68 ;
    RECT 91.59 82.89 91.8 82.96 ;
    RECT 91.59 83.25 91.8 83.32 ;
    RECT 91.59 83.61 91.8 83.68 ;
    RECT 87.81 82.89 88.02 82.96 ;
    RECT 87.81 83.25 88.02 83.32 ;
    RECT 87.81 83.61 88.02 83.68 ;
    RECT 88.27 82.89 88.48 82.96 ;
    RECT 88.27 83.25 88.48 83.32 ;
    RECT 88.27 83.61 88.48 83.68 ;
    RECT 84.49 82.89 84.7 82.96 ;
    RECT 84.49 83.25 84.7 83.32 ;
    RECT 84.49 83.61 84.7 83.68 ;
    RECT 84.95 82.89 85.16 82.96 ;
    RECT 84.95 83.25 85.16 83.32 ;
    RECT 84.95 83.61 85.16 83.68 ;
    RECT 81.17 82.89 81.38 82.96 ;
    RECT 81.17 83.25 81.38 83.32 ;
    RECT 81.17 83.61 81.38 83.68 ;
    RECT 81.63 82.89 81.84 82.96 ;
    RECT 81.63 83.25 81.84 83.32 ;
    RECT 81.63 83.61 81.84 83.68 ;
    RECT 77.85 82.89 78.06 82.96 ;
    RECT 77.85 83.25 78.06 83.32 ;
    RECT 77.85 83.61 78.06 83.68 ;
    RECT 78.31 82.89 78.52 82.96 ;
    RECT 78.31 83.25 78.52 83.32 ;
    RECT 78.31 83.61 78.52 83.68 ;
    RECT 74.53 82.89 74.74 82.96 ;
    RECT 74.53 83.25 74.74 83.32 ;
    RECT 74.53 83.61 74.74 83.68 ;
    RECT 74.99 82.89 75.2 82.96 ;
    RECT 74.99 83.25 75.2 83.32 ;
    RECT 74.99 83.61 75.2 83.68 ;
    RECT 71.21 82.89 71.42 82.96 ;
    RECT 71.21 83.25 71.42 83.32 ;
    RECT 71.21 83.61 71.42 83.68 ;
    RECT 71.67 82.89 71.88 82.96 ;
    RECT 71.67 83.25 71.88 83.32 ;
    RECT 71.67 83.61 71.88 83.68 ;
    RECT 31.37 82.89 31.58 82.96 ;
    RECT 31.37 83.25 31.58 83.32 ;
    RECT 31.37 83.61 31.58 83.68 ;
    RECT 31.83 82.89 32.04 82.96 ;
    RECT 31.83 83.25 32.04 83.32 ;
    RECT 31.83 83.61 32.04 83.68 ;
    RECT 67.89 82.89 68.1 82.96 ;
    RECT 67.89 83.25 68.1 83.32 ;
    RECT 67.89 83.61 68.1 83.68 ;
    RECT 68.35 82.89 68.56 82.96 ;
    RECT 68.35 83.25 68.56 83.32 ;
    RECT 68.35 83.61 68.56 83.68 ;
    RECT 28.05 82.89 28.26 82.96 ;
    RECT 28.05 83.25 28.26 83.32 ;
    RECT 28.05 83.61 28.26 83.68 ;
    RECT 28.51 82.89 28.72 82.96 ;
    RECT 28.51 83.25 28.72 83.32 ;
    RECT 28.51 83.61 28.72 83.68 ;
    RECT 24.73 82.89 24.94 82.96 ;
    RECT 24.73 83.25 24.94 83.32 ;
    RECT 24.73 83.61 24.94 83.68 ;
    RECT 25.19 82.89 25.4 82.96 ;
    RECT 25.19 83.25 25.4 83.32 ;
    RECT 25.19 83.61 25.4 83.68 ;
    RECT 21.41 82.89 21.62 82.96 ;
    RECT 21.41 83.25 21.62 83.32 ;
    RECT 21.41 83.61 21.62 83.68 ;
    RECT 21.87 82.89 22.08 82.96 ;
    RECT 21.87 83.25 22.08 83.32 ;
    RECT 21.87 83.61 22.08 83.68 ;
    RECT 18.09 82.89 18.3 82.96 ;
    RECT 18.09 83.25 18.3 83.32 ;
    RECT 18.09 83.61 18.3 83.68 ;
    RECT 18.55 82.89 18.76 82.96 ;
    RECT 18.55 83.25 18.76 83.32 ;
    RECT 18.55 83.61 18.76 83.68 ;
    RECT 120.825 83.25 120.895 83.32 ;
    RECT 14.77 82.89 14.98 82.96 ;
    RECT 14.77 83.25 14.98 83.32 ;
    RECT 14.77 83.61 14.98 83.68 ;
    RECT 15.23 82.89 15.44 82.96 ;
    RECT 15.23 83.25 15.44 83.32 ;
    RECT 15.23 83.61 15.44 83.68 ;
    RECT 11.45 82.89 11.66 82.96 ;
    RECT 11.45 83.25 11.66 83.32 ;
    RECT 11.45 83.61 11.66 83.68 ;
    RECT 11.91 82.89 12.12 82.96 ;
    RECT 11.91 83.25 12.12 83.32 ;
    RECT 11.91 83.61 12.12 83.68 ;
    RECT 8.13 82.89 8.34 82.96 ;
    RECT 8.13 83.25 8.34 83.32 ;
    RECT 8.13 83.61 8.34 83.68 ;
    RECT 8.59 82.89 8.8 82.96 ;
    RECT 8.59 83.25 8.8 83.32 ;
    RECT 8.59 83.61 8.8 83.68 ;
    RECT 4.81 82.89 5.02 82.96 ;
    RECT 4.81 83.25 5.02 83.32 ;
    RECT 4.81 83.61 5.02 83.68 ;
    RECT 5.27 82.89 5.48 82.96 ;
    RECT 5.27 83.25 5.48 83.32 ;
    RECT 5.27 83.61 5.48 83.68 ;
    RECT 1.49 82.89 1.7 82.96 ;
    RECT 1.49 83.25 1.7 83.32 ;
    RECT 1.49 83.61 1.7 83.68 ;
    RECT 1.95 82.89 2.16 82.96 ;
    RECT 1.95 83.25 2.16 83.32 ;
    RECT 1.95 83.61 2.16 83.68 ;
    RECT 64.57 82.89 64.78 82.96 ;
    RECT 64.57 83.25 64.78 83.32 ;
    RECT 64.57 83.61 64.78 83.68 ;
    RECT 65.03 82.89 65.24 82.96 ;
    RECT 65.03 83.25 65.24 83.32 ;
    RECT 65.03 83.61 65.24 83.68 ;
    RECT 61.25 82.17 61.46 82.24 ;
    RECT 61.25 82.53 61.46 82.6 ;
    RECT 61.25 82.89 61.46 82.96 ;
    RECT 61.71 82.17 61.92 82.24 ;
    RECT 61.71 82.53 61.92 82.6 ;
    RECT 61.71 82.89 61.92 82.96 ;
    RECT 57.93 82.17 58.14 82.24 ;
    RECT 57.93 82.53 58.14 82.6 ;
    RECT 57.93 82.89 58.14 82.96 ;
    RECT 58.39 82.17 58.6 82.24 ;
    RECT 58.39 82.53 58.6 82.6 ;
    RECT 58.39 82.89 58.6 82.96 ;
    RECT 54.61 82.17 54.82 82.24 ;
    RECT 54.61 82.53 54.82 82.6 ;
    RECT 54.61 82.89 54.82 82.96 ;
    RECT 55.07 82.17 55.28 82.24 ;
    RECT 55.07 82.53 55.28 82.6 ;
    RECT 55.07 82.89 55.28 82.96 ;
    RECT 51.29 82.17 51.5 82.24 ;
    RECT 51.29 82.53 51.5 82.6 ;
    RECT 51.29 82.89 51.5 82.96 ;
    RECT 51.75 82.17 51.96 82.24 ;
    RECT 51.75 82.53 51.96 82.6 ;
    RECT 51.75 82.89 51.96 82.96 ;
    RECT 47.97 82.17 48.18 82.24 ;
    RECT 47.97 82.53 48.18 82.6 ;
    RECT 47.97 82.89 48.18 82.96 ;
    RECT 48.43 82.17 48.64 82.24 ;
    RECT 48.43 82.53 48.64 82.6 ;
    RECT 48.43 82.89 48.64 82.96 ;
    RECT 44.65 82.17 44.86 82.24 ;
    RECT 44.65 82.53 44.86 82.6 ;
    RECT 44.65 82.89 44.86 82.96 ;
    RECT 45.11 82.17 45.32 82.24 ;
    RECT 45.11 82.53 45.32 82.6 ;
    RECT 45.11 82.89 45.32 82.96 ;
    RECT 41.33 82.17 41.54 82.24 ;
    RECT 41.33 82.53 41.54 82.6 ;
    RECT 41.33 82.89 41.54 82.96 ;
    RECT 41.79 82.17 42.0 82.24 ;
    RECT 41.79 82.53 42.0 82.6 ;
    RECT 41.79 82.89 42.0 82.96 ;
    RECT 38.01 82.17 38.22 82.24 ;
    RECT 38.01 82.53 38.22 82.6 ;
    RECT 38.01 82.89 38.22 82.96 ;
    RECT 38.47 82.17 38.68 82.24 ;
    RECT 38.47 82.53 38.68 82.6 ;
    RECT 38.47 82.89 38.68 82.96 ;
    RECT 0.4 82.53 0.47 82.6 ;
    RECT 34.69 82.17 34.9 82.24 ;
    RECT 34.69 82.53 34.9 82.6 ;
    RECT 34.69 82.89 34.9 82.96 ;
    RECT 35.15 82.17 35.36 82.24 ;
    RECT 35.15 82.53 35.36 82.6 ;
    RECT 35.15 82.89 35.36 82.96 ;
    RECT 117.69 82.17 117.9 82.24 ;
    RECT 117.69 82.53 117.9 82.6 ;
    RECT 117.69 82.89 117.9 82.96 ;
    RECT 118.15 82.17 118.36 82.24 ;
    RECT 118.15 82.53 118.36 82.6 ;
    RECT 118.15 82.89 118.36 82.96 ;
    RECT 114.37 82.17 114.58 82.24 ;
    RECT 114.37 82.53 114.58 82.6 ;
    RECT 114.37 82.89 114.58 82.96 ;
    RECT 114.83 82.17 115.04 82.24 ;
    RECT 114.83 82.53 115.04 82.6 ;
    RECT 114.83 82.89 115.04 82.96 ;
    RECT 111.05 82.17 111.26 82.24 ;
    RECT 111.05 82.53 111.26 82.6 ;
    RECT 111.05 82.89 111.26 82.96 ;
    RECT 111.51 82.17 111.72 82.24 ;
    RECT 111.51 82.53 111.72 82.6 ;
    RECT 111.51 82.89 111.72 82.96 ;
    RECT 107.73 82.17 107.94 82.24 ;
    RECT 107.73 82.53 107.94 82.6 ;
    RECT 107.73 82.89 107.94 82.96 ;
    RECT 108.19 82.17 108.4 82.24 ;
    RECT 108.19 82.53 108.4 82.6 ;
    RECT 108.19 82.89 108.4 82.96 ;
    RECT 104.41 82.17 104.62 82.24 ;
    RECT 104.41 82.53 104.62 82.6 ;
    RECT 104.41 82.89 104.62 82.96 ;
    RECT 104.87 82.17 105.08 82.24 ;
    RECT 104.87 82.53 105.08 82.6 ;
    RECT 104.87 82.89 105.08 82.96 ;
    RECT 101.09 82.17 101.3 82.24 ;
    RECT 101.09 82.53 101.3 82.6 ;
    RECT 101.09 82.89 101.3 82.96 ;
    RECT 101.55 82.17 101.76 82.24 ;
    RECT 101.55 82.53 101.76 82.6 ;
    RECT 101.55 82.89 101.76 82.96 ;
    RECT 97.77 82.17 97.98 82.24 ;
    RECT 97.77 82.53 97.98 82.6 ;
    RECT 97.77 82.89 97.98 82.96 ;
    RECT 98.23 82.17 98.44 82.24 ;
    RECT 98.23 82.53 98.44 82.6 ;
    RECT 98.23 82.89 98.44 82.96 ;
    RECT 94.45 82.17 94.66 82.24 ;
    RECT 94.45 82.53 94.66 82.6 ;
    RECT 94.45 82.89 94.66 82.96 ;
    RECT 94.91 82.17 95.12 82.24 ;
    RECT 94.91 82.53 95.12 82.6 ;
    RECT 94.91 82.89 95.12 82.96 ;
    RECT 91.13 82.17 91.34 82.24 ;
    RECT 91.13 82.53 91.34 82.6 ;
    RECT 91.13 82.89 91.34 82.96 ;
    RECT 91.59 82.17 91.8 82.24 ;
    RECT 91.59 82.53 91.8 82.6 ;
    RECT 91.59 82.89 91.8 82.96 ;
    RECT 87.81 82.17 88.02 82.24 ;
    RECT 87.81 82.53 88.02 82.6 ;
    RECT 87.81 82.89 88.02 82.96 ;
    RECT 88.27 82.17 88.48 82.24 ;
    RECT 88.27 82.53 88.48 82.6 ;
    RECT 88.27 82.89 88.48 82.96 ;
    RECT 84.49 82.17 84.7 82.24 ;
    RECT 84.49 82.53 84.7 82.6 ;
    RECT 84.49 82.89 84.7 82.96 ;
    RECT 84.95 82.17 85.16 82.24 ;
    RECT 84.95 82.53 85.16 82.6 ;
    RECT 84.95 82.89 85.16 82.96 ;
    RECT 81.17 82.17 81.38 82.24 ;
    RECT 81.17 82.53 81.38 82.6 ;
    RECT 81.17 82.89 81.38 82.96 ;
    RECT 81.63 82.17 81.84 82.24 ;
    RECT 81.63 82.53 81.84 82.6 ;
    RECT 81.63 82.89 81.84 82.96 ;
    RECT 77.85 82.17 78.06 82.24 ;
    RECT 77.85 82.53 78.06 82.6 ;
    RECT 77.85 82.89 78.06 82.96 ;
    RECT 78.31 82.17 78.52 82.24 ;
    RECT 78.31 82.53 78.52 82.6 ;
    RECT 78.31 82.89 78.52 82.96 ;
    RECT 74.53 82.17 74.74 82.24 ;
    RECT 74.53 82.53 74.74 82.6 ;
    RECT 74.53 82.89 74.74 82.96 ;
    RECT 74.99 82.17 75.2 82.24 ;
    RECT 74.99 82.53 75.2 82.6 ;
    RECT 74.99 82.89 75.2 82.96 ;
    RECT 71.21 82.17 71.42 82.24 ;
    RECT 71.21 82.53 71.42 82.6 ;
    RECT 71.21 82.89 71.42 82.96 ;
    RECT 71.67 82.17 71.88 82.24 ;
    RECT 71.67 82.53 71.88 82.6 ;
    RECT 71.67 82.89 71.88 82.96 ;
    RECT 31.37 82.17 31.58 82.24 ;
    RECT 31.37 82.53 31.58 82.6 ;
    RECT 31.37 82.89 31.58 82.96 ;
    RECT 31.83 82.17 32.04 82.24 ;
    RECT 31.83 82.53 32.04 82.6 ;
    RECT 31.83 82.89 32.04 82.96 ;
    RECT 67.89 82.17 68.1 82.24 ;
    RECT 67.89 82.53 68.1 82.6 ;
    RECT 67.89 82.89 68.1 82.96 ;
    RECT 68.35 82.17 68.56 82.24 ;
    RECT 68.35 82.53 68.56 82.6 ;
    RECT 68.35 82.89 68.56 82.96 ;
    RECT 28.05 82.17 28.26 82.24 ;
    RECT 28.05 82.53 28.26 82.6 ;
    RECT 28.05 82.89 28.26 82.96 ;
    RECT 28.51 82.17 28.72 82.24 ;
    RECT 28.51 82.53 28.72 82.6 ;
    RECT 28.51 82.89 28.72 82.96 ;
    RECT 24.73 82.17 24.94 82.24 ;
    RECT 24.73 82.53 24.94 82.6 ;
    RECT 24.73 82.89 24.94 82.96 ;
    RECT 25.19 82.17 25.4 82.24 ;
    RECT 25.19 82.53 25.4 82.6 ;
    RECT 25.19 82.89 25.4 82.96 ;
    RECT 21.41 82.17 21.62 82.24 ;
    RECT 21.41 82.53 21.62 82.6 ;
    RECT 21.41 82.89 21.62 82.96 ;
    RECT 21.87 82.17 22.08 82.24 ;
    RECT 21.87 82.53 22.08 82.6 ;
    RECT 21.87 82.89 22.08 82.96 ;
    RECT 18.09 82.17 18.3 82.24 ;
    RECT 18.09 82.53 18.3 82.6 ;
    RECT 18.09 82.89 18.3 82.96 ;
    RECT 18.55 82.17 18.76 82.24 ;
    RECT 18.55 82.53 18.76 82.6 ;
    RECT 18.55 82.89 18.76 82.96 ;
    RECT 120.825 82.53 120.895 82.6 ;
    RECT 14.77 82.17 14.98 82.24 ;
    RECT 14.77 82.53 14.98 82.6 ;
    RECT 14.77 82.89 14.98 82.96 ;
    RECT 15.23 82.17 15.44 82.24 ;
    RECT 15.23 82.53 15.44 82.6 ;
    RECT 15.23 82.89 15.44 82.96 ;
    RECT 11.45 82.17 11.66 82.24 ;
    RECT 11.45 82.53 11.66 82.6 ;
    RECT 11.45 82.89 11.66 82.96 ;
    RECT 11.91 82.17 12.12 82.24 ;
    RECT 11.91 82.53 12.12 82.6 ;
    RECT 11.91 82.89 12.12 82.96 ;
    RECT 8.13 82.17 8.34 82.24 ;
    RECT 8.13 82.53 8.34 82.6 ;
    RECT 8.13 82.89 8.34 82.96 ;
    RECT 8.59 82.17 8.8 82.24 ;
    RECT 8.59 82.53 8.8 82.6 ;
    RECT 8.59 82.89 8.8 82.96 ;
    RECT 4.81 82.17 5.02 82.24 ;
    RECT 4.81 82.53 5.02 82.6 ;
    RECT 4.81 82.89 5.02 82.96 ;
    RECT 5.27 82.17 5.48 82.24 ;
    RECT 5.27 82.53 5.48 82.6 ;
    RECT 5.27 82.89 5.48 82.96 ;
    RECT 1.49 82.17 1.7 82.24 ;
    RECT 1.49 82.53 1.7 82.6 ;
    RECT 1.49 82.89 1.7 82.96 ;
    RECT 1.95 82.17 2.16 82.24 ;
    RECT 1.95 82.53 2.16 82.6 ;
    RECT 1.95 82.89 2.16 82.96 ;
    RECT 64.57 82.17 64.78 82.24 ;
    RECT 64.57 82.53 64.78 82.6 ;
    RECT 64.57 82.89 64.78 82.96 ;
    RECT 65.03 82.17 65.24 82.24 ;
    RECT 65.03 82.53 65.24 82.6 ;
    RECT 65.03 82.89 65.24 82.96 ;
    RECT 61.25 81.45 61.46 81.52 ;
    RECT 61.25 81.81 61.46 81.88 ;
    RECT 61.25 82.17 61.46 82.24 ;
    RECT 61.71 81.45 61.92 81.52 ;
    RECT 61.71 81.81 61.92 81.88 ;
    RECT 61.71 82.17 61.92 82.24 ;
    RECT 57.93 81.45 58.14 81.52 ;
    RECT 57.93 81.81 58.14 81.88 ;
    RECT 57.93 82.17 58.14 82.24 ;
    RECT 58.39 81.45 58.6 81.52 ;
    RECT 58.39 81.81 58.6 81.88 ;
    RECT 58.39 82.17 58.6 82.24 ;
    RECT 54.61 81.45 54.82 81.52 ;
    RECT 54.61 81.81 54.82 81.88 ;
    RECT 54.61 82.17 54.82 82.24 ;
    RECT 55.07 81.45 55.28 81.52 ;
    RECT 55.07 81.81 55.28 81.88 ;
    RECT 55.07 82.17 55.28 82.24 ;
    RECT 51.29 81.45 51.5 81.52 ;
    RECT 51.29 81.81 51.5 81.88 ;
    RECT 51.29 82.17 51.5 82.24 ;
    RECT 51.75 81.45 51.96 81.52 ;
    RECT 51.75 81.81 51.96 81.88 ;
    RECT 51.75 82.17 51.96 82.24 ;
    RECT 47.97 81.45 48.18 81.52 ;
    RECT 47.97 81.81 48.18 81.88 ;
    RECT 47.97 82.17 48.18 82.24 ;
    RECT 48.43 81.45 48.64 81.52 ;
    RECT 48.43 81.81 48.64 81.88 ;
    RECT 48.43 82.17 48.64 82.24 ;
    RECT 44.65 81.45 44.86 81.52 ;
    RECT 44.65 81.81 44.86 81.88 ;
    RECT 44.65 82.17 44.86 82.24 ;
    RECT 45.11 81.45 45.32 81.52 ;
    RECT 45.11 81.81 45.32 81.88 ;
    RECT 45.11 82.17 45.32 82.24 ;
    RECT 41.33 81.45 41.54 81.52 ;
    RECT 41.33 81.81 41.54 81.88 ;
    RECT 41.33 82.17 41.54 82.24 ;
    RECT 41.79 81.45 42.0 81.52 ;
    RECT 41.79 81.81 42.0 81.88 ;
    RECT 41.79 82.17 42.0 82.24 ;
    RECT 38.01 81.45 38.22 81.52 ;
    RECT 38.01 81.81 38.22 81.88 ;
    RECT 38.01 82.17 38.22 82.24 ;
    RECT 38.47 81.45 38.68 81.52 ;
    RECT 38.47 81.81 38.68 81.88 ;
    RECT 38.47 82.17 38.68 82.24 ;
    RECT 0.4 81.81 0.47 81.88 ;
    RECT 34.69 81.45 34.9 81.52 ;
    RECT 34.69 81.81 34.9 81.88 ;
    RECT 34.69 82.17 34.9 82.24 ;
    RECT 35.15 81.45 35.36 81.52 ;
    RECT 35.15 81.81 35.36 81.88 ;
    RECT 35.15 82.17 35.36 82.24 ;
    RECT 117.69 81.45 117.9 81.52 ;
    RECT 117.69 81.81 117.9 81.88 ;
    RECT 117.69 82.17 117.9 82.24 ;
    RECT 118.15 81.45 118.36 81.52 ;
    RECT 118.15 81.81 118.36 81.88 ;
    RECT 118.15 82.17 118.36 82.24 ;
    RECT 114.37 81.45 114.58 81.52 ;
    RECT 114.37 81.81 114.58 81.88 ;
    RECT 114.37 82.17 114.58 82.24 ;
    RECT 114.83 81.45 115.04 81.52 ;
    RECT 114.83 81.81 115.04 81.88 ;
    RECT 114.83 82.17 115.04 82.24 ;
    RECT 111.05 81.45 111.26 81.52 ;
    RECT 111.05 81.81 111.26 81.88 ;
    RECT 111.05 82.17 111.26 82.24 ;
    RECT 111.51 81.45 111.72 81.52 ;
    RECT 111.51 81.81 111.72 81.88 ;
    RECT 111.51 82.17 111.72 82.24 ;
    RECT 107.73 81.45 107.94 81.52 ;
    RECT 107.73 81.81 107.94 81.88 ;
    RECT 107.73 82.17 107.94 82.24 ;
    RECT 108.19 81.45 108.4 81.52 ;
    RECT 108.19 81.81 108.4 81.88 ;
    RECT 108.19 82.17 108.4 82.24 ;
    RECT 104.41 81.45 104.62 81.52 ;
    RECT 104.41 81.81 104.62 81.88 ;
    RECT 104.41 82.17 104.62 82.24 ;
    RECT 104.87 81.45 105.08 81.52 ;
    RECT 104.87 81.81 105.08 81.88 ;
    RECT 104.87 82.17 105.08 82.24 ;
    RECT 101.09 81.45 101.3 81.52 ;
    RECT 101.09 81.81 101.3 81.88 ;
    RECT 101.09 82.17 101.3 82.24 ;
    RECT 101.55 81.45 101.76 81.52 ;
    RECT 101.55 81.81 101.76 81.88 ;
    RECT 101.55 82.17 101.76 82.24 ;
    RECT 97.77 81.45 97.98 81.52 ;
    RECT 97.77 81.81 97.98 81.88 ;
    RECT 97.77 82.17 97.98 82.24 ;
    RECT 98.23 81.45 98.44 81.52 ;
    RECT 98.23 81.81 98.44 81.88 ;
    RECT 98.23 82.17 98.44 82.24 ;
    RECT 94.45 81.45 94.66 81.52 ;
    RECT 94.45 81.81 94.66 81.88 ;
    RECT 94.45 82.17 94.66 82.24 ;
    RECT 94.91 81.45 95.12 81.52 ;
    RECT 94.91 81.81 95.12 81.88 ;
    RECT 94.91 82.17 95.12 82.24 ;
    RECT 91.13 81.45 91.34 81.52 ;
    RECT 91.13 81.81 91.34 81.88 ;
    RECT 91.13 82.17 91.34 82.24 ;
    RECT 91.59 81.45 91.8 81.52 ;
    RECT 91.59 81.81 91.8 81.88 ;
    RECT 91.59 82.17 91.8 82.24 ;
    RECT 87.81 81.45 88.02 81.52 ;
    RECT 87.81 81.81 88.02 81.88 ;
    RECT 87.81 82.17 88.02 82.24 ;
    RECT 88.27 81.45 88.48 81.52 ;
    RECT 88.27 81.81 88.48 81.88 ;
    RECT 88.27 82.17 88.48 82.24 ;
    RECT 84.49 81.45 84.7 81.52 ;
    RECT 84.49 81.81 84.7 81.88 ;
    RECT 84.49 82.17 84.7 82.24 ;
    RECT 84.95 81.45 85.16 81.52 ;
    RECT 84.95 81.81 85.16 81.88 ;
    RECT 84.95 82.17 85.16 82.24 ;
    RECT 81.17 81.45 81.38 81.52 ;
    RECT 81.17 81.81 81.38 81.88 ;
    RECT 81.17 82.17 81.38 82.24 ;
    RECT 81.63 81.45 81.84 81.52 ;
    RECT 81.63 81.81 81.84 81.88 ;
    RECT 81.63 82.17 81.84 82.24 ;
    RECT 77.85 81.45 78.06 81.52 ;
    RECT 77.85 81.81 78.06 81.88 ;
    RECT 77.85 82.17 78.06 82.24 ;
    RECT 78.31 81.45 78.52 81.52 ;
    RECT 78.31 81.81 78.52 81.88 ;
    RECT 78.31 82.17 78.52 82.24 ;
    RECT 74.53 81.45 74.74 81.52 ;
    RECT 74.53 81.81 74.74 81.88 ;
    RECT 74.53 82.17 74.74 82.24 ;
    RECT 74.99 81.45 75.2 81.52 ;
    RECT 74.99 81.81 75.2 81.88 ;
    RECT 74.99 82.17 75.2 82.24 ;
    RECT 71.21 81.45 71.42 81.52 ;
    RECT 71.21 81.81 71.42 81.88 ;
    RECT 71.21 82.17 71.42 82.24 ;
    RECT 71.67 81.45 71.88 81.52 ;
    RECT 71.67 81.81 71.88 81.88 ;
    RECT 71.67 82.17 71.88 82.24 ;
    RECT 31.37 81.45 31.58 81.52 ;
    RECT 31.37 81.81 31.58 81.88 ;
    RECT 31.37 82.17 31.58 82.24 ;
    RECT 31.83 81.45 32.04 81.52 ;
    RECT 31.83 81.81 32.04 81.88 ;
    RECT 31.83 82.17 32.04 82.24 ;
    RECT 67.89 81.45 68.1 81.52 ;
    RECT 67.89 81.81 68.1 81.88 ;
    RECT 67.89 82.17 68.1 82.24 ;
    RECT 68.35 81.45 68.56 81.52 ;
    RECT 68.35 81.81 68.56 81.88 ;
    RECT 68.35 82.17 68.56 82.24 ;
    RECT 28.05 81.45 28.26 81.52 ;
    RECT 28.05 81.81 28.26 81.88 ;
    RECT 28.05 82.17 28.26 82.24 ;
    RECT 28.51 81.45 28.72 81.52 ;
    RECT 28.51 81.81 28.72 81.88 ;
    RECT 28.51 82.17 28.72 82.24 ;
    RECT 24.73 81.45 24.94 81.52 ;
    RECT 24.73 81.81 24.94 81.88 ;
    RECT 24.73 82.17 24.94 82.24 ;
    RECT 25.19 81.45 25.4 81.52 ;
    RECT 25.19 81.81 25.4 81.88 ;
    RECT 25.19 82.17 25.4 82.24 ;
    RECT 21.41 81.45 21.62 81.52 ;
    RECT 21.41 81.81 21.62 81.88 ;
    RECT 21.41 82.17 21.62 82.24 ;
    RECT 21.87 81.45 22.08 81.52 ;
    RECT 21.87 81.81 22.08 81.88 ;
    RECT 21.87 82.17 22.08 82.24 ;
    RECT 18.09 81.45 18.3 81.52 ;
    RECT 18.09 81.81 18.3 81.88 ;
    RECT 18.09 82.17 18.3 82.24 ;
    RECT 18.55 81.45 18.76 81.52 ;
    RECT 18.55 81.81 18.76 81.88 ;
    RECT 18.55 82.17 18.76 82.24 ;
    RECT 120.825 81.81 120.895 81.88 ;
    RECT 14.77 81.45 14.98 81.52 ;
    RECT 14.77 81.81 14.98 81.88 ;
    RECT 14.77 82.17 14.98 82.24 ;
    RECT 15.23 81.45 15.44 81.52 ;
    RECT 15.23 81.81 15.44 81.88 ;
    RECT 15.23 82.17 15.44 82.24 ;
    RECT 11.45 81.45 11.66 81.52 ;
    RECT 11.45 81.81 11.66 81.88 ;
    RECT 11.45 82.17 11.66 82.24 ;
    RECT 11.91 81.45 12.12 81.52 ;
    RECT 11.91 81.81 12.12 81.88 ;
    RECT 11.91 82.17 12.12 82.24 ;
    RECT 8.13 81.45 8.34 81.52 ;
    RECT 8.13 81.81 8.34 81.88 ;
    RECT 8.13 82.17 8.34 82.24 ;
    RECT 8.59 81.45 8.8 81.52 ;
    RECT 8.59 81.81 8.8 81.88 ;
    RECT 8.59 82.17 8.8 82.24 ;
    RECT 4.81 81.45 5.02 81.52 ;
    RECT 4.81 81.81 5.02 81.88 ;
    RECT 4.81 82.17 5.02 82.24 ;
    RECT 5.27 81.45 5.48 81.52 ;
    RECT 5.27 81.81 5.48 81.88 ;
    RECT 5.27 82.17 5.48 82.24 ;
    RECT 1.49 81.45 1.7 81.52 ;
    RECT 1.49 81.81 1.7 81.88 ;
    RECT 1.49 82.17 1.7 82.24 ;
    RECT 1.95 81.45 2.16 81.52 ;
    RECT 1.95 81.81 2.16 81.88 ;
    RECT 1.95 82.17 2.16 82.24 ;
    RECT 64.57 81.45 64.78 81.52 ;
    RECT 64.57 81.81 64.78 81.88 ;
    RECT 64.57 82.17 64.78 82.24 ;
    RECT 65.03 81.45 65.24 81.52 ;
    RECT 65.03 81.81 65.24 81.88 ;
    RECT 65.03 82.17 65.24 82.24 ;
    RECT 61.25 80.73 61.46 80.8 ;
    RECT 61.25 81.09 61.46 81.16 ;
    RECT 61.25 81.45 61.46 81.52 ;
    RECT 61.71 80.73 61.92 80.8 ;
    RECT 61.71 81.09 61.92 81.16 ;
    RECT 61.71 81.45 61.92 81.52 ;
    RECT 57.93 80.73 58.14 80.8 ;
    RECT 57.93 81.09 58.14 81.16 ;
    RECT 57.93 81.45 58.14 81.52 ;
    RECT 58.39 80.73 58.6 80.8 ;
    RECT 58.39 81.09 58.6 81.16 ;
    RECT 58.39 81.45 58.6 81.52 ;
    RECT 54.61 80.73 54.82 80.8 ;
    RECT 54.61 81.09 54.82 81.16 ;
    RECT 54.61 81.45 54.82 81.52 ;
    RECT 55.07 80.73 55.28 80.8 ;
    RECT 55.07 81.09 55.28 81.16 ;
    RECT 55.07 81.45 55.28 81.52 ;
    RECT 51.29 80.73 51.5 80.8 ;
    RECT 51.29 81.09 51.5 81.16 ;
    RECT 51.29 81.45 51.5 81.52 ;
    RECT 51.75 80.73 51.96 80.8 ;
    RECT 51.75 81.09 51.96 81.16 ;
    RECT 51.75 81.45 51.96 81.52 ;
    RECT 47.97 80.73 48.18 80.8 ;
    RECT 47.97 81.09 48.18 81.16 ;
    RECT 47.97 81.45 48.18 81.52 ;
    RECT 48.43 80.73 48.64 80.8 ;
    RECT 48.43 81.09 48.64 81.16 ;
    RECT 48.43 81.45 48.64 81.52 ;
    RECT 44.65 80.73 44.86 80.8 ;
    RECT 44.65 81.09 44.86 81.16 ;
    RECT 44.65 81.45 44.86 81.52 ;
    RECT 45.11 80.73 45.32 80.8 ;
    RECT 45.11 81.09 45.32 81.16 ;
    RECT 45.11 81.45 45.32 81.52 ;
    RECT 41.33 80.73 41.54 80.8 ;
    RECT 41.33 81.09 41.54 81.16 ;
    RECT 41.33 81.45 41.54 81.52 ;
    RECT 41.79 80.73 42.0 80.8 ;
    RECT 41.79 81.09 42.0 81.16 ;
    RECT 41.79 81.45 42.0 81.52 ;
    RECT 38.01 80.73 38.22 80.8 ;
    RECT 38.01 81.09 38.22 81.16 ;
    RECT 38.01 81.45 38.22 81.52 ;
    RECT 38.47 80.73 38.68 80.8 ;
    RECT 38.47 81.09 38.68 81.16 ;
    RECT 38.47 81.45 38.68 81.52 ;
    RECT 0.4 81.09 0.47 81.16 ;
    RECT 34.69 80.73 34.9 80.8 ;
    RECT 34.69 81.09 34.9 81.16 ;
    RECT 34.69 81.45 34.9 81.52 ;
    RECT 35.15 80.73 35.36 80.8 ;
    RECT 35.15 81.09 35.36 81.16 ;
    RECT 35.15 81.45 35.36 81.52 ;
    RECT 117.69 80.73 117.9 80.8 ;
    RECT 117.69 81.09 117.9 81.16 ;
    RECT 117.69 81.45 117.9 81.52 ;
    RECT 118.15 80.73 118.36 80.8 ;
    RECT 118.15 81.09 118.36 81.16 ;
    RECT 118.15 81.45 118.36 81.52 ;
    RECT 114.37 80.73 114.58 80.8 ;
    RECT 114.37 81.09 114.58 81.16 ;
    RECT 114.37 81.45 114.58 81.52 ;
    RECT 114.83 80.73 115.04 80.8 ;
    RECT 114.83 81.09 115.04 81.16 ;
    RECT 114.83 81.45 115.04 81.52 ;
    RECT 111.05 80.73 111.26 80.8 ;
    RECT 111.05 81.09 111.26 81.16 ;
    RECT 111.05 81.45 111.26 81.52 ;
    RECT 111.51 80.73 111.72 80.8 ;
    RECT 111.51 81.09 111.72 81.16 ;
    RECT 111.51 81.45 111.72 81.52 ;
    RECT 107.73 80.73 107.94 80.8 ;
    RECT 107.73 81.09 107.94 81.16 ;
    RECT 107.73 81.45 107.94 81.52 ;
    RECT 108.19 80.73 108.4 80.8 ;
    RECT 108.19 81.09 108.4 81.16 ;
    RECT 108.19 81.45 108.4 81.52 ;
    RECT 104.41 80.73 104.62 80.8 ;
    RECT 104.41 81.09 104.62 81.16 ;
    RECT 104.41 81.45 104.62 81.52 ;
    RECT 104.87 80.73 105.08 80.8 ;
    RECT 104.87 81.09 105.08 81.16 ;
    RECT 104.87 81.45 105.08 81.52 ;
    RECT 101.09 80.73 101.3 80.8 ;
    RECT 101.09 81.09 101.3 81.16 ;
    RECT 101.09 81.45 101.3 81.52 ;
    RECT 101.55 80.73 101.76 80.8 ;
    RECT 101.55 81.09 101.76 81.16 ;
    RECT 101.55 81.45 101.76 81.52 ;
    RECT 97.77 80.73 97.98 80.8 ;
    RECT 97.77 81.09 97.98 81.16 ;
    RECT 97.77 81.45 97.98 81.52 ;
    RECT 98.23 80.73 98.44 80.8 ;
    RECT 98.23 81.09 98.44 81.16 ;
    RECT 98.23 81.45 98.44 81.52 ;
    RECT 94.45 80.73 94.66 80.8 ;
    RECT 94.45 81.09 94.66 81.16 ;
    RECT 94.45 81.45 94.66 81.52 ;
    RECT 94.91 80.73 95.12 80.8 ;
    RECT 94.91 81.09 95.12 81.16 ;
    RECT 94.91 81.45 95.12 81.52 ;
    RECT 91.13 80.73 91.34 80.8 ;
    RECT 91.13 81.09 91.34 81.16 ;
    RECT 91.13 81.45 91.34 81.52 ;
    RECT 91.59 80.73 91.8 80.8 ;
    RECT 91.59 81.09 91.8 81.16 ;
    RECT 91.59 81.45 91.8 81.52 ;
    RECT 87.81 80.73 88.02 80.8 ;
    RECT 87.81 81.09 88.02 81.16 ;
    RECT 87.81 81.45 88.02 81.52 ;
    RECT 88.27 80.73 88.48 80.8 ;
    RECT 88.27 81.09 88.48 81.16 ;
    RECT 88.27 81.45 88.48 81.52 ;
    RECT 84.49 80.73 84.7 80.8 ;
    RECT 84.49 81.09 84.7 81.16 ;
    RECT 84.49 81.45 84.7 81.52 ;
    RECT 84.95 80.73 85.16 80.8 ;
    RECT 84.95 81.09 85.16 81.16 ;
    RECT 84.95 81.45 85.16 81.52 ;
    RECT 81.17 80.73 81.38 80.8 ;
    RECT 81.17 81.09 81.38 81.16 ;
    RECT 81.17 81.45 81.38 81.52 ;
    RECT 81.63 80.73 81.84 80.8 ;
    RECT 81.63 81.09 81.84 81.16 ;
    RECT 81.63 81.45 81.84 81.52 ;
    RECT 77.85 80.73 78.06 80.8 ;
    RECT 77.85 81.09 78.06 81.16 ;
    RECT 77.85 81.45 78.06 81.52 ;
    RECT 78.31 80.73 78.52 80.8 ;
    RECT 78.31 81.09 78.52 81.16 ;
    RECT 78.31 81.45 78.52 81.52 ;
    RECT 74.53 80.73 74.74 80.8 ;
    RECT 74.53 81.09 74.74 81.16 ;
    RECT 74.53 81.45 74.74 81.52 ;
    RECT 74.99 80.73 75.2 80.8 ;
    RECT 74.99 81.09 75.2 81.16 ;
    RECT 74.99 81.45 75.2 81.52 ;
    RECT 71.21 80.73 71.42 80.8 ;
    RECT 71.21 81.09 71.42 81.16 ;
    RECT 71.21 81.45 71.42 81.52 ;
    RECT 71.67 80.73 71.88 80.8 ;
    RECT 71.67 81.09 71.88 81.16 ;
    RECT 71.67 81.45 71.88 81.52 ;
    RECT 31.37 80.73 31.58 80.8 ;
    RECT 31.37 81.09 31.58 81.16 ;
    RECT 31.37 81.45 31.58 81.52 ;
    RECT 31.83 80.73 32.04 80.8 ;
    RECT 31.83 81.09 32.04 81.16 ;
    RECT 31.83 81.45 32.04 81.52 ;
    RECT 67.89 80.73 68.1 80.8 ;
    RECT 67.89 81.09 68.1 81.16 ;
    RECT 67.89 81.45 68.1 81.52 ;
    RECT 68.35 80.73 68.56 80.8 ;
    RECT 68.35 81.09 68.56 81.16 ;
    RECT 68.35 81.45 68.56 81.52 ;
    RECT 28.05 80.73 28.26 80.8 ;
    RECT 28.05 81.09 28.26 81.16 ;
    RECT 28.05 81.45 28.26 81.52 ;
    RECT 28.51 80.73 28.72 80.8 ;
    RECT 28.51 81.09 28.72 81.16 ;
    RECT 28.51 81.45 28.72 81.52 ;
    RECT 24.73 80.73 24.94 80.8 ;
    RECT 24.73 81.09 24.94 81.16 ;
    RECT 24.73 81.45 24.94 81.52 ;
    RECT 25.19 80.73 25.4 80.8 ;
    RECT 25.19 81.09 25.4 81.16 ;
    RECT 25.19 81.45 25.4 81.52 ;
    RECT 21.41 80.73 21.62 80.8 ;
    RECT 21.41 81.09 21.62 81.16 ;
    RECT 21.41 81.45 21.62 81.52 ;
    RECT 21.87 80.73 22.08 80.8 ;
    RECT 21.87 81.09 22.08 81.16 ;
    RECT 21.87 81.45 22.08 81.52 ;
    RECT 18.09 80.73 18.3 80.8 ;
    RECT 18.09 81.09 18.3 81.16 ;
    RECT 18.09 81.45 18.3 81.52 ;
    RECT 18.55 80.73 18.76 80.8 ;
    RECT 18.55 81.09 18.76 81.16 ;
    RECT 18.55 81.45 18.76 81.52 ;
    RECT 120.825 81.09 120.895 81.16 ;
    RECT 14.77 80.73 14.98 80.8 ;
    RECT 14.77 81.09 14.98 81.16 ;
    RECT 14.77 81.45 14.98 81.52 ;
    RECT 15.23 80.73 15.44 80.8 ;
    RECT 15.23 81.09 15.44 81.16 ;
    RECT 15.23 81.45 15.44 81.52 ;
    RECT 11.45 80.73 11.66 80.8 ;
    RECT 11.45 81.09 11.66 81.16 ;
    RECT 11.45 81.45 11.66 81.52 ;
    RECT 11.91 80.73 12.12 80.8 ;
    RECT 11.91 81.09 12.12 81.16 ;
    RECT 11.91 81.45 12.12 81.52 ;
    RECT 8.13 80.73 8.34 80.8 ;
    RECT 8.13 81.09 8.34 81.16 ;
    RECT 8.13 81.45 8.34 81.52 ;
    RECT 8.59 80.73 8.8 80.8 ;
    RECT 8.59 81.09 8.8 81.16 ;
    RECT 8.59 81.45 8.8 81.52 ;
    RECT 4.81 80.73 5.02 80.8 ;
    RECT 4.81 81.09 5.02 81.16 ;
    RECT 4.81 81.45 5.02 81.52 ;
    RECT 5.27 80.73 5.48 80.8 ;
    RECT 5.27 81.09 5.48 81.16 ;
    RECT 5.27 81.45 5.48 81.52 ;
    RECT 1.49 80.73 1.7 80.8 ;
    RECT 1.49 81.09 1.7 81.16 ;
    RECT 1.49 81.45 1.7 81.52 ;
    RECT 1.95 80.73 2.16 80.8 ;
    RECT 1.95 81.09 2.16 81.16 ;
    RECT 1.95 81.45 2.16 81.52 ;
    RECT 64.57 80.73 64.78 80.8 ;
    RECT 64.57 81.09 64.78 81.16 ;
    RECT 64.57 81.45 64.78 81.52 ;
    RECT 65.03 80.73 65.24 80.8 ;
    RECT 65.03 81.09 65.24 81.16 ;
    RECT 65.03 81.45 65.24 81.52 ;
    RECT 61.25 80.01 61.46 80.08 ;
    RECT 61.25 80.37 61.46 80.44 ;
    RECT 61.25 80.73 61.46 80.8 ;
    RECT 61.71 80.01 61.92 80.08 ;
    RECT 61.71 80.37 61.92 80.44 ;
    RECT 61.71 80.73 61.92 80.8 ;
    RECT 57.93 80.01 58.14 80.08 ;
    RECT 57.93 80.37 58.14 80.44 ;
    RECT 57.93 80.73 58.14 80.8 ;
    RECT 58.39 80.01 58.6 80.08 ;
    RECT 58.39 80.37 58.6 80.44 ;
    RECT 58.39 80.73 58.6 80.8 ;
    RECT 54.61 80.01 54.82 80.08 ;
    RECT 54.61 80.37 54.82 80.44 ;
    RECT 54.61 80.73 54.82 80.8 ;
    RECT 55.07 80.01 55.28 80.08 ;
    RECT 55.07 80.37 55.28 80.44 ;
    RECT 55.07 80.73 55.28 80.8 ;
    RECT 51.29 80.01 51.5 80.08 ;
    RECT 51.29 80.37 51.5 80.44 ;
    RECT 51.29 80.73 51.5 80.8 ;
    RECT 51.75 80.01 51.96 80.08 ;
    RECT 51.75 80.37 51.96 80.44 ;
    RECT 51.75 80.73 51.96 80.8 ;
    RECT 47.97 80.01 48.18 80.08 ;
    RECT 47.97 80.37 48.18 80.44 ;
    RECT 47.97 80.73 48.18 80.8 ;
    RECT 48.43 80.01 48.64 80.08 ;
    RECT 48.43 80.37 48.64 80.44 ;
    RECT 48.43 80.73 48.64 80.8 ;
    RECT 44.65 80.01 44.86 80.08 ;
    RECT 44.65 80.37 44.86 80.44 ;
    RECT 44.65 80.73 44.86 80.8 ;
    RECT 45.11 80.01 45.32 80.08 ;
    RECT 45.11 80.37 45.32 80.44 ;
    RECT 45.11 80.73 45.32 80.8 ;
    RECT 41.33 80.01 41.54 80.08 ;
    RECT 41.33 80.37 41.54 80.44 ;
    RECT 41.33 80.73 41.54 80.8 ;
    RECT 41.79 80.01 42.0 80.08 ;
    RECT 41.79 80.37 42.0 80.44 ;
    RECT 41.79 80.73 42.0 80.8 ;
    RECT 38.01 80.01 38.22 80.08 ;
    RECT 38.01 80.37 38.22 80.44 ;
    RECT 38.01 80.73 38.22 80.8 ;
    RECT 38.47 80.01 38.68 80.08 ;
    RECT 38.47 80.37 38.68 80.44 ;
    RECT 38.47 80.73 38.68 80.8 ;
    RECT 0.4 80.37 0.47 80.44 ;
    RECT 34.69 80.01 34.9 80.08 ;
    RECT 34.69 80.37 34.9 80.44 ;
    RECT 34.69 80.73 34.9 80.8 ;
    RECT 35.15 80.01 35.36 80.08 ;
    RECT 35.15 80.37 35.36 80.44 ;
    RECT 35.15 80.73 35.36 80.8 ;
    RECT 117.69 80.01 117.9 80.08 ;
    RECT 117.69 80.37 117.9 80.44 ;
    RECT 117.69 80.73 117.9 80.8 ;
    RECT 118.15 80.01 118.36 80.08 ;
    RECT 118.15 80.37 118.36 80.44 ;
    RECT 118.15 80.73 118.36 80.8 ;
    RECT 114.37 80.01 114.58 80.08 ;
    RECT 114.37 80.37 114.58 80.44 ;
    RECT 114.37 80.73 114.58 80.8 ;
    RECT 114.83 80.01 115.04 80.08 ;
    RECT 114.83 80.37 115.04 80.44 ;
    RECT 114.83 80.73 115.04 80.8 ;
    RECT 111.05 80.01 111.26 80.08 ;
    RECT 111.05 80.37 111.26 80.44 ;
    RECT 111.05 80.73 111.26 80.8 ;
    RECT 111.51 80.01 111.72 80.08 ;
    RECT 111.51 80.37 111.72 80.44 ;
    RECT 111.51 80.73 111.72 80.8 ;
    RECT 107.73 80.01 107.94 80.08 ;
    RECT 107.73 80.37 107.94 80.44 ;
    RECT 107.73 80.73 107.94 80.8 ;
    RECT 108.19 80.01 108.4 80.08 ;
    RECT 108.19 80.37 108.4 80.44 ;
    RECT 108.19 80.73 108.4 80.8 ;
    RECT 104.41 80.01 104.62 80.08 ;
    RECT 104.41 80.37 104.62 80.44 ;
    RECT 104.41 80.73 104.62 80.8 ;
    RECT 104.87 80.01 105.08 80.08 ;
    RECT 104.87 80.37 105.08 80.44 ;
    RECT 104.87 80.73 105.08 80.8 ;
    RECT 101.09 80.01 101.3 80.08 ;
    RECT 101.09 80.37 101.3 80.44 ;
    RECT 101.09 80.73 101.3 80.8 ;
    RECT 101.55 80.01 101.76 80.08 ;
    RECT 101.55 80.37 101.76 80.44 ;
    RECT 101.55 80.73 101.76 80.8 ;
    RECT 97.77 80.01 97.98 80.08 ;
    RECT 97.77 80.37 97.98 80.44 ;
    RECT 97.77 80.73 97.98 80.8 ;
    RECT 98.23 80.01 98.44 80.08 ;
    RECT 98.23 80.37 98.44 80.44 ;
    RECT 98.23 80.73 98.44 80.8 ;
    RECT 94.45 80.01 94.66 80.08 ;
    RECT 94.45 80.37 94.66 80.44 ;
    RECT 94.45 80.73 94.66 80.8 ;
    RECT 94.91 80.01 95.12 80.08 ;
    RECT 94.91 80.37 95.12 80.44 ;
    RECT 94.91 80.73 95.12 80.8 ;
    RECT 91.13 80.01 91.34 80.08 ;
    RECT 91.13 80.37 91.34 80.44 ;
    RECT 91.13 80.73 91.34 80.8 ;
    RECT 91.59 80.01 91.8 80.08 ;
    RECT 91.59 80.37 91.8 80.44 ;
    RECT 91.59 80.73 91.8 80.8 ;
    RECT 87.81 80.01 88.02 80.08 ;
    RECT 87.81 80.37 88.02 80.44 ;
    RECT 87.81 80.73 88.02 80.8 ;
    RECT 88.27 80.01 88.48 80.08 ;
    RECT 88.27 80.37 88.48 80.44 ;
    RECT 88.27 80.73 88.48 80.8 ;
    RECT 84.49 80.01 84.7 80.08 ;
    RECT 84.49 80.37 84.7 80.44 ;
    RECT 84.49 80.73 84.7 80.8 ;
    RECT 84.95 80.01 85.16 80.08 ;
    RECT 84.95 80.37 85.16 80.44 ;
    RECT 84.95 80.73 85.16 80.8 ;
    RECT 81.17 80.01 81.38 80.08 ;
    RECT 81.17 80.37 81.38 80.44 ;
    RECT 81.17 80.73 81.38 80.8 ;
    RECT 81.63 80.01 81.84 80.08 ;
    RECT 81.63 80.37 81.84 80.44 ;
    RECT 81.63 80.73 81.84 80.8 ;
    RECT 77.85 80.01 78.06 80.08 ;
    RECT 77.85 80.37 78.06 80.44 ;
    RECT 77.85 80.73 78.06 80.8 ;
    RECT 78.31 80.01 78.52 80.08 ;
    RECT 78.31 80.37 78.52 80.44 ;
    RECT 78.31 80.73 78.52 80.8 ;
    RECT 74.53 80.01 74.74 80.08 ;
    RECT 74.53 80.37 74.74 80.44 ;
    RECT 74.53 80.73 74.74 80.8 ;
    RECT 74.99 80.01 75.2 80.08 ;
    RECT 74.99 80.37 75.2 80.44 ;
    RECT 74.99 80.73 75.2 80.8 ;
    RECT 71.21 80.01 71.42 80.08 ;
    RECT 71.21 80.37 71.42 80.44 ;
    RECT 71.21 80.73 71.42 80.8 ;
    RECT 71.67 80.01 71.88 80.08 ;
    RECT 71.67 80.37 71.88 80.44 ;
    RECT 71.67 80.73 71.88 80.8 ;
    RECT 31.37 80.01 31.58 80.08 ;
    RECT 31.37 80.37 31.58 80.44 ;
    RECT 31.37 80.73 31.58 80.8 ;
    RECT 31.83 80.01 32.04 80.08 ;
    RECT 31.83 80.37 32.04 80.44 ;
    RECT 31.83 80.73 32.04 80.8 ;
    RECT 67.89 80.01 68.1 80.08 ;
    RECT 67.89 80.37 68.1 80.44 ;
    RECT 67.89 80.73 68.1 80.8 ;
    RECT 68.35 80.01 68.56 80.08 ;
    RECT 68.35 80.37 68.56 80.44 ;
    RECT 68.35 80.73 68.56 80.8 ;
    RECT 28.05 80.01 28.26 80.08 ;
    RECT 28.05 80.37 28.26 80.44 ;
    RECT 28.05 80.73 28.26 80.8 ;
    RECT 28.51 80.01 28.72 80.08 ;
    RECT 28.51 80.37 28.72 80.44 ;
    RECT 28.51 80.73 28.72 80.8 ;
    RECT 24.73 80.01 24.94 80.08 ;
    RECT 24.73 80.37 24.94 80.44 ;
    RECT 24.73 80.73 24.94 80.8 ;
    RECT 25.19 80.01 25.4 80.08 ;
    RECT 25.19 80.37 25.4 80.44 ;
    RECT 25.19 80.73 25.4 80.8 ;
    RECT 21.41 80.01 21.62 80.08 ;
    RECT 21.41 80.37 21.62 80.44 ;
    RECT 21.41 80.73 21.62 80.8 ;
    RECT 21.87 80.01 22.08 80.08 ;
    RECT 21.87 80.37 22.08 80.44 ;
    RECT 21.87 80.73 22.08 80.8 ;
    RECT 18.09 80.01 18.3 80.08 ;
    RECT 18.09 80.37 18.3 80.44 ;
    RECT 18.09 80.73 18.3 80.8 ;
    RECT 18.55 80.01 18.76 80.08 ;
    RECT 18.55 80.37 18.76 80.44 ;
    RECT 18.55 80.73 18.76 80.8 ;
    RECT 120.825 80.37 120.895 80.44 ;
    RECT 14.77 80.01 14.98 80.08 ;
    RECT 14.77 80.37 14.98 80.44 ;
    RECT 14.77 80.73 14.98 80.8 ;
    RECT 15.23 80.01 15.44 80.08 ;
    RECT 15.23 80.37 15.44 80.44 ;
    RECT 15.23 80.73 15.44 80.8 ;
    RECT 11.45 80.01 11.66 80.08 ;
    RECT 11.45 80.37 11.66 80.44 ;
    RECT 11.45 80.73 11.66 80.8 ;
    RECT 11.91 80.01 12.12 80.08 ;
    RECT 11.91 80.37 12.12 80.44 ;
    RECT 11.91 80.73 12.12 80.8 ;
    RECT 8.13 80.01 8.34 80.08 ;
    RECT 8.13 80.37 8.34 80.44 ;
    RECT 8.13 80.73 8.34 80.8 ;
    RECT 8.59 80.01 8.8 80.08 ;
    RECT 8.59 80.37 8.8 80.44 ;
    RECT 8.59 80.73 8.8 80.8 ;
    RECT 4.81 80.01 5.02 80.08 ;
    RECT 4.81 80.37 5.02 80.44 ;
    RECT 4.81 80.73 5.02 80.8 ;
    RECT 5.27 80.01 5.48 80.08 ;
    RECT 5.27 80.37 5.48 80.44 ;
    RECT 5.27 80.73 5.48 80.8 ;
    RECT 1.49 80.01 1.7 80.08 ;
    RECT 1.49 80.37 1.7 80.44 ;
    RECT 1.49 80.73 1.7 80.8 ;
    RECT 1.95 80.01 2.16 80.08 ;
    RECT 1.95 80.37 2.16 80.44 ;
    RECT 1.95 80.73 2.16 80.8 ;
    RECT 64.57 80.01 64.78 80.08 ;
    RECT 64.57 80.37 64.78 80.44 ;
    RECT 64.57 80.73 64.78 80.8 ;
    RECT 65.03 80.01 65.24 80.08 ;
    RECT 65.03 80.37 65.24 80.44 ;
    RECT 65.03 80.73 65.24 80.8 ;
    RECT 61.25 42.55 61.46 42.62 ;
    RECT 61.25 42.91 61.46 42.98 ;
    RECT 61.25 43.27 61.46 43.34 ;
    RECT 61.71 42.55 61.92 42.62 ;
    RECT 61.71 42.91 61.92 42.98 ;
    RECT 61.71 43.27 61.92 43.34 ;
    RECT 57.93 42.55 58.14 42.62 ;
    RECT 57.93 42.91 58.14 42.98 ;
    RECT 57.93 43.27 58.14 43.34 ;
    RECT 58.39 42.55 58.6 42.62 ;
    RECT 58.39 42.91 58.6 42.98 ;
    RECT 58.39 43.27 58.6 43.34 ;
    RECT 54.61 42.55 54.82 42.62 ;
    RECT 54.61 42.91 54.82 42.98 ;
    RECT 54.61 43.27 54.82 43.34 ;
    RECT 55.07 42.55 55.28 42.62 ;
    RECT 55.07 42.91 55.28 42.98 ;
    RECT 55.07 43.27 55.28 43.34 ;
    RECT 51.29 42.55 51.5 42.62 ;
    RECT 51.29 42.91 51.5 42.98 ;
    RECT 51.29 43.27 51.5 43.34 ;
    RECT 51.75 42.55 51.96 42.62 ;
    RECT 51.75 42.91 51.96 42.98 ;
    RECT 51.75 43.27 51.96 43.34 ;
    RECT 47.97 42.55 48.18 42.62 ;
    RECT 47.97 42.91 48.18 42.98 ;
    RECT 47.97 43.27 48.18 43.34 ;
    RECT 48.43 42.55 48.64 42.62 ;
    RECT 48.43 42.91 48.64 42.98 ;
    RECT 48.43 43.27 48.64 43.34 ;
    RECT 44.65 42.55 44.86 42.62 ;
    RECT 44.65 42.91 44.86 42.98 ;
    RECT 44.65 43.27 44.86 43.34 ;
    RECT 45.11 42.55 45.32 42.62 ;
    RECT 45.11 42.91 45.32 42.98 ;
    RECT 45.11 43.27 45.32 43.34 ;
    RECT 41.33 42.55 41.54 42.62 ;
    RECT 41.33 42.91 41.54 42.98 ;
    RECT 41.33 43.27 41.54 43.34 ;
    RECT 41.79 42.55 42.0 42.62 ;
    RECT 41.79 42.91 42.0 42.98 ;
    RECT 41.79 43.27 42.0 43.34 ;
    RECT 38.01 42.55 38.22 42.62 ;
    RECT 38.01 42.91 38.22 42.98 ;
    RECT 38.01 43.27 38.22 43.34 ;
    RECT 38.47 42.55 38.68 42.62 ;
    RECT 38.47 42.91 38.68 42.98 ;
    RECT 38.47 43.27 38.68 43.34 ;
    RECT 0.4 42.91 0.47 42.98 ;
    RECT 34.69 42.55 34.9 42.62 ;
    RECT 34.69 42.91 34.9 42.98 ;
    RECT 34.69 43.27 34.9 43.34 ;
    RECT 35.15 42.55 35.36 42.62 ;
    RECT 35.15 42.91 35.36 42.98 ;
    RECT 35.15 43.27 35.36 43.34 ;
    RECT 117.69 42.55 117.9 42.62 ;
    RECT 117.69 42.91 117.9 42.98 ;
    RECT 117.69 43.27 117.9 43.34 ;
    RECT 118.15 42.55 118.36 42.62 ;
    RECT 118.15 42.91 118.36 42.98 ;
    RECT 118.15 43.27 118.36 43.34 ;
    RECT 114.37 42.55 114.58 42.62 ;
    RECT 114.37 42.91 114.58 42.98 ;
    RECT 114.37 43.27 114.58 43.34 ;
    RECT 114.83 42.55 115.04 42.62 ;
    RECT 114.83 42.91 115.04 42.98 ;
    RECT 114.83 43.27 115.04 43.34 ;
    RECT 111.05 42.55 111.26 42.62 ;
    RECT 111.05 42.91 111.26 42.98 ;
    RECT 111.05 43.27 111.26 43.34 ;
    RECT 111.51 42.55 111.72 42.62 ;
    RECT 111.51 42.91 111.72 42.98 ;
    RECT 111.51 43.27 111.72 43.34 ;
    RECT 107.73 42.55 107.94 42.62 ;
    RECT 107.73 42.91 107.94 42.98 ;
    RECT 107.73 43.27 107.94 43.34 ;
    RECT 108.19 42.55 108.4 42.62 ;
    RECT 108.19 42.91 108.4 42.98 ;
    RECT 108.19 43.27 108.4 43.34 ;
    RECT 104.41 42.55 104.62 42.62 ;
    RECT 104.41 42.91 104.62 42.98 ;
    RECT 104.41 43.27 104.62 43.34 ;
    RECT 104.87 42.55 105.08 42.62 ;
    RECT 104.87 42.91 105.08 42.98 ;
    RECT 104.87 43.27 105.08 43.34 ;
    RECT 101.09 42.55 101.3 42.62 ;
    RECT 101.09 42.91 101.3 42.98 ;
    RECT 101.09 43.27 101.3 43.34 ;
    RECT 101.55 42.55 101.76 42.62 ;
    RECT 101.55 42.91 101.76 42.98 ;
    RECT 101.55 43.27 101.76 43.34 ;
    RECT 97.77 42.55 97.98 42.62 ;
    RECT 97.77 42.91 97.98 42.98 ;
    RECT 97.77 43.27 97.98 43.34 ;
    RECT 98.23 42.55 98.44 42.62 ;
    RECT 98.23 42.91 98.44 42.98 ;
    RECT 98.23 43.27 98.44 43.34 ;
    RECT 94.45 42.55 94.66 42.62 ;
    RECT 94.45 42.91 94.66 42.98 ;
    RECT 94.45 43.27 94.66 43.34 ;
    RECT 94.91 42.55 95.12 42.62 ;
    RECT 94.91 42.91 95.12 42.98 ;
    RECT 94.91 43.27 95.12 43.34 ;
    RECT 91.13 42.55 91.34 42.62 ;
    RECT 91.13 42.91 91.34 42.98 ;
    RECT 91.13 43.27 91.34 43.34 ;
    RECT 91.59 42.55 91.8 42.62 ;
    RECT 91.59 42.91 91.8 42.98 ;
    RECT 91.59 43.27 91.8 43.34 ;
    RECT 87.81 42.55 88.02 42.62 ;
    RECT 87.81 42.91 88.02 42.98 ;
    RECT 87.81 43.27 88.02 43.34 ;
    RECT 88.27 42.55 88.48 42.62 ;
    RECT 88.27 42.91 88.48 42.98 ;
    RECT 88.27 43.27 88.48 43.34 ;
    RECT 84.49 42.55 84.7 42.62 ;
    RECT 84.49 42.91 84.7 42.98 ;
    RECT 84.49 43.27 84.7 43.34 ;
    RECT 84.95 42.55 85.16 42.62 ;
    RECT 84.95 42.91 85.16 42.98 ;
    RECT 84.95 43.27 85.16 43.34 ;
    RECT 81.17 42.55 81.38 42.62 ;
    RECT 81.17 42.91 81.38 42.98 ;
    RECT 81.17 43.27 81.38 43.34 ;
    RECT 81.63 42.55 81.84 42.62 ;
    RECT 81.63 42.91 81.84 42.98 ;
    RECT 81.63 43.27 81.84 43.34 ;
    RECT 77.85 42.55 78.06 42.62 ;
    RECT 77.85 42.91 78.06 42.98 ;
    RECT 77.85 43.27 78.06 43.34 ;
    RECT 78.31 42.55 78.52 42.62 ;
    RECT 78.31 42.91 78.52 42.98 ;
    RECT 78.31 43.27 78.52 43.34 ;
    RECT 74.53 42.55 74.74 42.62 ;
    RECT 74.53 42.91 74.74 42.98 ;
    RECT 74.53 43.27 74.74 43.34 ;
    RECT 74.99 42.55 75.2 42.62 ;
    RECT 74.99 42.91 75.2 42.98 ;
    RECT 74.99 43.27 75.2 43.34 ;
    RECT 71.21 42.55 71.42 42.62 ;
    RECT 71.21 42.91 71.42 42.98 ;
    RECT 71.21 43.27 71.42 43.34 ;
    RECT 71.67 42.55 71.88 42.62 ;
    RECT 71.67 42.91 71.88 42.98 ;
    RECT 71.67 43.27 71.88 43.34 ;
    RECT 31.37 42.55 31.58 42.62 ;
    RECT 31.37 42.91 31.58 42.98 ;
    RECT 31.37 43.27 31.58 43.34 ;
    RECT 31.83 42.55 32.04 42.62 ;
    RECT 31.83 42.91 32.04 42.98 ;
    RECT 31.83 43.27 32.04 43.34 ;
    RECT 67.89 42.55 68.1 42.62 ;
    RECT 67.89 42.91 68.1 42.98 ;
    RECT 67.89 43.27 68.1 43.34 ;
    RECT 68.35 42.55 68.56 42.62 ;
    RECT 68.35 42.91 68.56 42.98 ;
    RECT 68.35 43.27 68.56 43.34 ;
    RECT 28.05 42.55 28.26 42.62 ;
    RECT 28.05 42.91 28.26 42.98 ;
    RECT 28.05 43.27 28.26 43.34 ;
    RECT 28.51 42.55 28.72 42.62 ;
    RECT 28.51 42.91 28.72 42.98 ;
    RECT 28.51 43.27 28.72 43.34 ;
    RECT 24.73 42.55 24.94 42.62 ;
    RECT 24.73 42.91 24.94 42.98 ;
    RECT 24.73 43.27 24.94 43.34 ;
    RECT 25.19 42.55 25.4 42.62 ;
    RECT 25.19 42.91 25.4 42.98 ;
    RECT 25.19 43.27 25.4 43.34 ;
    RECT 21.41 42.55 21.62 42.62 ;
    RECT 21.41 42.91 21.62 42.98 ;
    RECT 21.41 43.27 21.62 43.34 ;
    RECT 21.87 42.55 22.08 42.62 ;
    RECT 21.87 42.91 22.08 42.98 ;
    RECT 21.87 43.27 22.08 43.34 ;
    RECT 18.09 42.55 18.3 42.62 ;
    RECT 18.09 42.91 18.3 42.98 ;
    RECT 18.09 43.27 18.3 43.34 ;
    RECT 18.55 42.55 18.76 42.62 ;
    RECT 18.55 42.91 18.76 42.98 ;
    RECT 18.55 43.27 18.76 43.34 ;
    RECT 120.825 42.91 120.895 42.98 ;
    RECT 14.77 42.55 14.98 42.62 ;
    RECT 14.77 42.91 14.98 42.98 ;
    RECT 14.77 43.27 14.98 43.34 ;
    RECT 15.23 42.55 15.44 42.62 ;
    RECT 15.23 42.91 15.44 42.98 ;
    RECT 15.23 43.27 15.44 43.34 ;
    RECT 11.45 42.55 11.66 42.62 ;
    RECT 11.45 42.91 11.66 42.98 ;
    RECT 11.45 43.27 11.66 43.34 ;
    RECT 11.91 42.55 12.12 42.62 ;
    RECT 11.91 42.91 12.12 42.98 ;
    RECT 11.91 43.27 12.12 43.34 ;
    RECT 8.13 42.55 8.34 42.62 ;
    RECT 8.13 42.91 8.34 42.98 ;
    RECT 8.13 43.27 8.34 43.34 ;
    RECT 8.59 42.55 8.8 42.62 ;
    RECT 8.59 42.91 8.8 42.98 ;
    RECT 8.59 43.27 8.8 43.34 ;
    RECT 4.81 42.55 5.02 42.62 ;
    RECT 4.81 42.91 5.02 42.98 ;
    RECT 4.81 43.27 5.02 43.34 ;
    RECT 5.27 42.55 5.48 42.62 ;
    RECT 5.27 42.91 5.48 42.98 ;
    RECT 5.27 43.27 5.48 43.34 ;
    RECT 1.49 42.55 1.7 42.62 ;
    RECT 1.49 42.91 1.7 42.98 ;
    RECT 1.49 43.27 1.7 43.34 ;
    RECT 1.95 42.55 2.16 42.62 ;
    RECT 1.95 42.91 2.16 42.98 ;
    RECT 1.95 43.27 2.16 43.34 ;
    RECT 64.57 42.55 64.78 42.62 ;
    RECT 64.57 42.91 64.78 42.98 ;
    RECT 64.57 43.27 64.78 43.34 ;
    RECT 65.03 42.55 65.24 42.62 ;
    RECT 65.03 42.91 65.24 42.98 ;
    RECT 65.03 43.27 65.24 43.34 ;
    RECT 61.25 98.01 61.46 98.08 ;
    RECT 61.25 98.37 61.46 98.44 ;
    RECT 61.25 98.73 61.46 98.8 ;
    RECT 61.71 98.01 61.92 98.08 ;
    RECT 61.71 98.37 61.92 98.44 ;
    RECT 61.71 98.73 61.92 98.8 ;
    RECT 57.93 98.01 58.14 98.08 ;
    RECT 57.93 98.37 58.14 98.44 ;
    RECT 57.93 98.73 58.14 98.8 ;
    RECT 58.39 98.01 58.6 98.08 ;
    RECT 58.39 98.37 58.6 98.44 ;
    RECT 58.39 98.73 58.6 98.8 ;
    RECT 54.61 98.01 54.82 98.08 ;
    RECT 54.61 98.37 54.82 98.44 ;
    RECT 54.61 98.73 54.82 98.8 ;
    RECT 55.07 98.01 55.28 98.08 ;
    RECT 55.07 98.37 55.28 98.44 ;
    RECT 55.07 98.73 55.28 98.8 ;
    RECT 117.69 98.01 117.9 98.08 ;
    RECT 117.69 98.37 117.9 98.44 ;
    RECT 117.69 98.73 117.9 98.8 ;
    RECT 118.15 98.01 118.36 98.08 ;
    RECT 118.15 98.37 118.36 98.44 ;
    RECT 118.15 98.73 118.36 98.8 ;
    RECT 51.29 98.01 51.5 98.08 ;
    RECT 51.29 98.37 51.5 98.44 ;
    RECT 51.29 98.73 51.5 98.8 ;
    RECT 51.75 98.01 51.96 98.08 ;
    RECT 51.75 98.37 51.96 98.44 ;
    RECT 51.75 98.73 51.96 98.8 ;
    RECT 47.97 98.01 48.18 98.08 ;
    RECT 47.97 98.37 48.18 98.44 ;
    RECT 47.97 98.73 48.18 98.8 ;
    RECT 48.43 98.01 48.64 98.08 ;
    RECT 48.43 98.37 48.64 98.44 ;
    RECT 48.43 98.73 48.64 98.8 ;
    RECT 44.65 98.01 44.86 98.08 ;
    RECT 44.65 98.37 44.86 98.44 ;
    RECT 44.65 98.73 44.86 98.8 ;
    RECT 45.11 98.01 45.32 98.08 ;
    RECT 45.11 98.37 45.32 98.44 ;
    RECT 45.11 98.73 45.32 98.8 ;
    RECT 41.33 98.01 41.54 98.08 ;
    RECT 41.33 98.37 41.54 98.44 ;
    RECT 41.33 98.73 41.54 98.8 ;
    RECT 41.79 98.01 42.0 98.08 ;
    RECT 41.79 98.37 42.0 98.44 ;
    RECT 41.79 98.73 42.0 98.8 ;
    RECT 38.01 98.01 38.22 98.08 ;
    RECT 38.01 98.37 38.22 98.44 ;
    RECT 38.01 98.73 38.22 98.8 ;
    RECT 38.47 98.01 38.68 98.08 ;
    RECT 38.47 98.37 38.68 98.44 ;
    RECT 38.47 98.73 38.68 98.8 ;
    RECT 34.69 98.01 34.9 98.08 ;
    RECT 34.69 98.37 34.9 98.44 ;
    RECT 34.69 98.73 34.9 98.8 ;
    RECT 35.15 98.01 35.36 98.08 ;
    RECT 35.15 98.37 35.36 98.44 ;
    RECT 35.15 98.73 35.36 98.8 ;
    RECT 1.49 98.01 1.7 98.08 ;
    RECT 1.49 98.37 1.7 98.44 ;
    RECT 1.49 98.73 1.7 98.8 ;
    RECT 1.95 98.01 2.16 98.08 ;
    RECT 1.95 98.37 2.16 98.44 ;
    RECT 1.95 98.73 2.16 98.8 ;
    RECT 0.4 98.37 0.47 98.44 ;
    RECT 114.37 98.01 114.58 98.08 ;
    RECT 114.37 98.37 114.58 98.44 ;
    RECT 114.37 98.73 114.58 98.8 ;
    RECT 114.83 98.01 115.04 98.08 ;
    RECT 114.83 98.37 115.04 98.44 ;
    RECT 114.83 98.73 115.04 98.8 ;
    RECT 111.05 98.01 111.26 98.08 ;
    RECT 111.05 98.37 111.26 98.44 ;
    RECT 111.05 98.73 111.26 98.8 ;
    RECT 111.51 98.01 111.72 98.08 ;
    RECT 111.51 98.37 111.72 98.44 ;
    RECT 111.51 98.73 111.72 98.8 ;
    RECT 107.73 98.01 107.94 98.08 ;
    RECT 107.73 98.37 107.94 98.44 ;
    RECT 107.73 98.73 107.94 98.8 ;
    RECT 108.19 98.01 108.4 98.08 ;
    RECT 108.19 98.37 108.4 98.44 ;
    RECT 108.19 98.73 108.4 98.8 ;
    RECT 104.41 98.01 104.62 98.08 ;
    RECT 104.41 98.37 104.62 98.44 ;
    RECT 104.41 98.73 104.62 98.8 ;
    RECT 104.87 98.01 105.08 98.08 ;
    RECT 104.87 98.37 105.08 98.44 ;
    RECT 104.87 98.73 105.08 98.8 ;
    RECT 101.09 98.01 101.3 98.08 ;
    RECT 101.09 98.37 101.3 98.44 ;
    RECT 101.09 98.73 101.3 98.8 ;
    RECT 101.55 98.01 101.76 98.08 ;
    RECT 101.55 98.37 101.76 98.44 ;
    RECT 101.55 98.73 101.76 98.8 ;
    RECT 97.77 98.01 97.98 98.08 ;
    RECT 97.77 98.37 97.98 98.44 ;
    RECT 97.77 98.73 97.98 98.8 ;
    RECT 98.23 98.01 98.44 98.08 ;
    RECT 98.23 98.37 98.44 98.44 ;
    RECT 98.23 98.73 98.44 98.8 ;
    RECT 94.45 98.01 94.66 98.08 ;
    RECT 94.45 98.37 94.66 98.44 ;
    RECT 94.45 98.73 94.66 98.8 ;
    RECT 94.91 98.01 95.12 98.08 ;
    RECT 94.91 98.37 95.12 98.44 ;
    RECT 94.91 98.73 95.12 98.8 ;
    RECT 91.13 98.01 91.34 98.08 ;
    RECT 91.13 98.37 91.34 98.44 ;
    RECT 91.13 98.73 91.34 98.8 ;
    RECT 91.59 98.01 91.8 98.08 ;
    RECT 91.59 98.37 91.8 98.44 ;
    RECT 91.59 98.73 91.8 98.8 ;
    RECT 87.81 98.01 88.02 98.08 ;
    RECT 87.81 98.37 88.02 98.44 ;
    RECT 87.81 98.73 88.02 98.8 ;
    RECT 88.27 98.01 88.48 98.08 ;
    RECT 88.27 98.37 88.48 98.44 ;
    RECT 88.27 98.73 88.48 98.8 ;
    RECT 84.49 98.01 84.7 98.08 ;
    RECT 84.49 98.37 84.7 98.44 ;
    RECT 84.49 98.73 84.7 98.8 ;
    RECT 84.95 98.01 85.16 98.08 ;
    RECT 84.95 98.37 85.16 98.44 ;
    RECT 84.95 98.73 85.16 98.8 ;
    RECT 81.17 98.01 81.38 98.08 ;
    RECT 81.17 98.37 81.38 98.44 ;
    RECT 81.17 98.73 81.38 98.8 ;
    RECT 81.63 98.01 81.84 98.08 ;
    RECT 81.63 98.37 81.84 98.44 ;
    RECT 81.63 98.73 81.84 98.8 ;
    RECT 77.85 98.01 78.06 98.08 ;
    RECT 77.85 98.37 78.06 98.44 ;
    RECT 77.85 98.73 78.06 98.8 ;
    RECT 78.31 98.01 78.52 98.08 ;
    RECT 78.31 98.37 78.52 98.44 ;
    RECT 78.31 98.73 78.52 98.8 ;
    RECT 74.53 98.01 74.74 98.08 ;
    RECT 74.53 98.37 74.74 98.44 ;
    RECT 74.53 98.73 74.74 98.8 ;
    RECT 74.99 98.01 75.2 98.08 ;
    RECT 74.99 98.37 75.2 98.44 ;
    RECT 74.99 98.73 75.2 98.8 ;
    RECT 71.21 98.01 71.42 98.08 ;
    RECT 71.21 98.37 71.42 98.44 ;
    RECT 71.21 98.73 71.42 98.8 ;
    RECT 71.67 98.01 71.88 98.08 ;
    RECT 71.67 98.37 71.88 98.44 ;
    RECT 71.67 98.73 71.88 98.8 ;
    RECT 31.37 98.01 31.58 98.08 ;
    RECT 31.37 98.37 31.58 98.44 ;
    RECT 31.37 98.73 31.58 98.8 ;
    RECT 31.83 98.01 32.04 98.08 ;
    RECT 31.83 98.37 32.04 98.44 ;
    RECT 31.83 98.73 32.04 98.8 ;
    RECT 67.89 98.01 68.1 98.08 ;
    RECT 67.89 98.37 68.1 98.44 ;
    RECT 67.89 98.73 68.1 98.8 ;
    RECT 68.35 98.01 68.56 98.08 ;
    RECT 68.35 98.37 68.56 98.44 ;
    RECT 68.35 98.73 68.56 98.8 ;
    RECT 28.05 98.01 28.26 98.08 ;
    RECT 28.05 98.37 28.26 98.44 ;
    RECT 28.05 98.73 28.26 98.8 ;
    RECT 28.51 98.01 28.72 98.08 ;
    RECT 28.51 98.37 28.72 98.44 ;
    RECT 28.51 98.73 28.72 98.8 ;
    RECT 24.73 98.01 24.94 98.08 ;
    RECT 24.73 98.37 24.94 98.44 ;
    RECT 24.73 98.73 24.94 98.8 ;
    RECT 25.19 98.01 25.4 98.08 ;
    RECT 25.19 98.37 25.4 98.44 ;
    RECT 25.19 98.73 25.4 98.8 ;
    RECT 21.41 98.01 21.62 98.08 ;
    RECT 21.41 98.37 21.62 98.44 ;
    RECT 21.41 98.73 21.62 98.8 ;
    RECT 21.87 98.01 22.08 98.08 ;
    RECT 21.87 98.37 22.08 98.44 ;
    RECT 21.87 98.73 22.08 98.8 ;
    RECT 18.09 98.01 18.3 98.08 ;
    RECT 18.09 98.37 18.3 98.44 ;
    RECT 18.09 98.73 18.3 98.8 ;
    RECT 18.55 98.01 18.76 98.08 ;
    RECT 18.55 98.37 18.76 98.44 ;
    RECT 18.55 98.73 18.76 98.8 ;
    RECT 14.77 98.01 14.98 98.08 ;
    RECT 14.77 98.37 14.98 98.44 ;
    RECT 14.77 98.73 14.98 98.8 ;
    RECT 15.23 98.01 15.44 98.08 ;
    RECT 15.23 98.37 15.44 98.44 ;
    RECT 15.23 98.73 15.44 98.8 ;
    RECT 11.45 98.01 11.66 98.08 ;
    RECT 11.45 98.37 11.66 98.44 ;
    RECT 11.45 98.73 11.66 98.8 ;
    RECT 11.91 98.01 12.12 98.08 ;
    RECT 11.91 98.37 12.12 98.44 ;
    RECT 11.91 98.73 12.12 98.8 ;
    RECT 120.825 98.37 120.895 98.44 ;
    RECT 8.13 98.01 8.34 98.08 ;
    RECT 8.13 98.37 8.34 98.44 ;
    RECT 8.13 98.73 8.34 98.8 ;
    RECT 8.59 98.01 8.8 98.08 ;
    RECT 8.59 98.37 8.8 98.44 ;
    RECT 8.59 98.73 8.8 98.8 ;
    RECT 4.81 98.01 5.02 98.08 ;
    RECT 4.81 98.37 5.02 98.44 ;
    RECT 4.81 98.73 5.02 98.8 ;
    RECT 5.27 98.01 5.48 98.08 ;
    RECT 5.27 98.37 5.48 98.44 ;
    RECT 5.27 98.73 5.48 98.8 ;
    RECT 64.57 98.01 64.78 98.08 ;
    RECT 64.57 98.37 64.78 98.44 ;
    RECT 64.57 98.73 64.78 98.8 ;
    RECT 65.03 98.01 65.24 98.08 ;
    RECT 65.03 98.37 65.24 98.44 ;
    RECT 65.03 98.73 65.24 98.8 ;
    RECT 61.25 41.83 61.46 41.9 ;
    RECT 61.25 42.19 61.46 42.26 ;
    RECT 61.25 42.55 61.46 42.62 ;
    RECT 61.71 41.83 61.92 41.9 ;
    RECT 61.71 42.19 61.92 42.26 ;
    RECT 61.71 42.55 61.92 42.62 ;
    RECT 57.93 41.83 58.14 41.9 ;
    RECT 57.93 42.19 58.14 42.26 ;
    RECT 57.93 42.55 58.14 42.62 ;
    RECT 58.39 41.83 58.6 41.9 ;
    RECT 58.39 42.19 58.6 42.26 ;
    RECT 58.39 42.55 58.6 42.62 ;
    RECT 54.61 41.83 54.82 41.9 ;
    RECT 54.61 42.19 54.82 42.26 ;
    RECT 54.61 42.55 54.82 42.62 ;
    RECT 55.07 41.83 55.28 41.9 ;
    RECT 55.07 42.19 55.28 42.26 ;
    RECT 55.07 42.55 55.28 42.62 ;
    RECT 51.29 41.83 51.5 41.9 ;
    RECT 51.29 42.19 51.5 42.26 ;
    RECT 51.29 42.55 51.5 42.62 ;
    RECT 51.75 41.83 51.96 41.9 ;
    RECT 51.75 42.19 51.96 42.26 ;
    RECT 51.75 42.55 51.96 42.62 ;
    RECT 47.97 41.83 48.18 41.9 ;
    RECT 47.97 42.19 48.18 42.26 ;
    RECT 47.97 42.55 48.18 42.62 ;
    RECT 48.43 41.83 48.64 41.9 ;
    RECT 48.43 42.19 48.64 42.26 ;
    RECT 48.43 42.55 48.64 42.62 ;
    RECT 44.65 41.83 44.86 41.9 ;
    RECT 44.65 42.19 44.86 42.26 ;
    RECT 44.65 42.55 44.86 42.62 ;
    RECT 45.11 41.83 45.32 41.9 ;
    RECT 45.11 42.19 45.32 42.26 ;
    RECT 45.11 42.55 45.32 42.62 ;
    RECT 41.33 41.83 41.54 41.9 ;
    RECT 41.33 42.19 41.54 42.26 ;
    RECT 41.33 42.55 41.54 42.62 ;
    RECT 41.79 41.83 42.0 41.9 ;
    RECT 41.79 42.19 42.0 42.26 ;
    RECT 41.79 42.55 42.0 42.62 ;
    RECT 38.01 41.83 38.22 41.9 ;
    RECT 38.01 42.19 38.22 42.26 ;
    RECT 38.01 42.55 38.22 42.62 ;
    RECT 38.47 41.83 38.68 41.9 ;
    RECT 38.47 42.19 38.68 42.26 ;
    RECT 38.47 42.55 38.68 42.62 ;
    RECT 0.4 42.19 0.47 42.26 ;
    RECT 34.69 41.83 34.9 41.9 ;
    RECT 34.69 42.19 34.9 42.26 ;
    RECT 34.69 42.55 34.9 42.62 ;
    RECT 35.15 41.83 35.36 41.9 ;
    RECT 35.15 42.19 35.36 42.26 ;
    RECT 35.15 42.55 35.36 42.62 ;
    RECT 117.69 41.83 117.9 41.9 ;
    RECT 117.69 42.19 117.9 42.26 ;
    RECT 117.69 42.55 117.9 42.62 ;
    RECT 118.15 41.83 118.36 41.9 ;
    RECT 118.15 42.19 118.36 42.26 ;
    RECT 118.15 42.55 118.36 42.62 ;
    RECT 114.37 41.83 114.58 41.9 ;
    RECT 114.37 42.19 114.58 42.26 ;
    RECT 114.37 42.55 114.58 42.62 ;
    RECT 114.83 41.83 115.04 41.9 ;
    RECT 114.83 42.19 115.04 42.26 ;
    RECT 114.83 42.55 115.04 42.62 ;
    RECT 111.05 41.83 111.26 41.9 ;
    RECT 111.05 42.19 111.26 42.26 ;
    RECT 111.05 42.55 111.26 42.62 ;
    RECT 111.51 41.83 111.72 41.9 ;
    RECT 111.51 42.19 111.72 42.26 ;
    RECT 111.51 42.55 111.72 42.62 ;
    RECT 107.73 41.83 107.94 41.9 ;
    RECT 107.73 42.19 107.94 42.26 ;
    RECT 107.73 42.55 107.94 42.62 ;
    RECT 108.19 41.83 108.4 41.9 ;
    RECT 108.19 42.19 108.4 42.26 ;
    RECT 108.19 42.55 108.4 42.62 ;
    RECT 104.41 41.83 104.62 41.9 ;
    RECT 104.41 42.19 104.62 42.26 ;
    RECT 104.41 42.55 104.62 42.62 ;
    RECT 104.87 41.83 105.08 41.9 ;
    RECT 104.87 42.19 105.08 42.26 ;
    RECT 104.87 42.55 105.08 42.62 ;
    RECT 101.09 41.83 101.3 41.9 ;
    RECT 101.09 42.19 101.3 42.26 ;
    RECT 101.09 42.55 101.3 42.62 ;
    RECT 101.55 41.83 101.76 41.9 ;
    RECT 101.55 42.19 101.76 42.26 ;
    RECT 101.55 42.55 101.76 42.62 ;
    RECT 97.77 41.83 97.98 41.9 ;
    RECT 97.77 42.19 97.98 42.26 ;
    RECT 97.77 42.55 97.98 42.62 ;
    RECT 98.23 41.83 98.44 41.9 ;
    RECT 98.23 42.19 98.44 42.26 ;
    RECT 98.23 42.55 98.44 42.62 ;
    RECT 94.45 41.83 94.66 41.9 ;
    RECT 94.45 42.19 94.66 42.26 ;
    RECT 94.45 42.55 94.66 42.62 ;
    RECT 94.91 41.83 95.12 41.9 ;
    RECT 94.91 42.19 95.12 42.26 ;
    RECT 94.91 42.55 95.12 42.62 ;
    RECT 91.13 41.83 91.34 41.9 ;
    RECT 91.13 42.19 91.34 42.26 ;
    RECT 91.13 42.55 91.34 42.62 ;
    RECT 91.59 41.83 91.8 41.9 ;
    RECT 91.59 42.19 91.8 42.26 ;
    RECT 91.59 42.55 91.8 42.62 ;
    RECT 87.81 41.83 88.02 41.9 ;
    RECT 87.81 42.19 88.02 42.26 ;
    RECT 87.81 42.55 88.02 42.62 ;
    RECT 88.27 41.83 88.48 41.9 ;
    RECT 88.27 42.19 88.48 42.26 ;
    RECT 88.27 42.55 88.48 42.62 ;
    RECT 84.49 41.83 84.7 41.9 ;
    RECT 84.49 42.19 84.7 42.26 ;
    RECT 84.49 42.55 84.7 42.62 ;
    RECT 84.95 41.83 85.16 41.9 ;
    RECT 84.95 42.19 85.16 42.26 ;
    RECT 84.95 42.55 85.16 42.62 ;
    RECT 81.17 41.83 81.38 41.9 ;
    RECT 81.17 42.19 81.38 42.26 ;
    RECT 81.17 42.55 81.38 42.62 ;
    RECT 81.63 41.83 81.84 41.9 ;
    RECT 81.63 42.19 81.84 42.26 ;
    RECT 81.63 42.55 81.84 42.62 ;
    RECT 77.85 41.83 78.06 41.9 ;
    RECT 77.85 42.19 78.06 42.26 ;
    RECT 77.85 42.55 78.06 42.62 ;
    RECT 78.31 41.83 78.52 41.9 ;
    RECT 78.31 42.19 78.52 42.26 ;
    RECT 78.31 42.55 78.52 42.62 ;
    RECT 74.53 41.83 74.74 41.9 ;
    RECT 74.53 42.19 74.74 42.26 ;
    RECT 74.53 42.55 74.74 42.62 ;
    RECT 74.99 41.83 75.2 41.9 ;
    RECT 74.99 42.19 75.2 42.26 ;
    RECT 74.99 42.55 75.2 42.62 ;
    RECT 71.21 41.83 71.42 41.9 ;
    RECT 71.21 42.19 71.42 42.26 ;
    RECT 71.21 42.55 71.42 42.62 ;
    RECT 71.67 41.83 71.88 41.9 ;
    RECT 71.67 42.19 71.88 42.26 ;
    RECT 71.67 42.55 71.88 42.62 ;
    RECT 31.37 41.83 31.58 41.9 ;
    RECT 31.37 42.19 31.58 42.26 ;
    RECT 31.37 42.55 31.58 42.62 ;
    RECT 31.83 41.83 32.04 41.9 ;
    RECT 31.83 42.19 32.04 42.26 ;
    RECT 31.83 42.55 32.04 42.62 ;
    RECT 67.89 41.83 68.1 41.9 ;
    RECT 67.89 42.19 68.1 42.26 ;
    RECT 67.89 42.55 68.1 42.62 ;
    RECT 68.35 41.83 68.56 41.9 ;
    RECT 68.35 42.19 68.56 42.26 ;
    RECT 68.35 42.55 68.56 42.62 ;
    RECT 28.05 41.83 28.26 41.9 ;
    RECT 28.05 42.19 28.26 42.26 ;
    RECT 28.05 42.55 28.26 42.62 ;
    RECT 28.51 41.83 28.72 41.9 ;
    RECT 28.51 42.19 28.72 42.26 ;
    RECT 28.51 42.55 28.72 42.62 ;
    RECT 24.73 41.83 24.94 41.9 ;
    RECT 24.73 42.19 24.94 42.26 ;
    RECT 24.73 42.55 24.94 42.62 ;
    RECT 25.19 41.83 25.4 41.9 ;
    RECT 25.19 42.19 25.4 42.26 ;
    RECT 25.19 42.55 25.4 42.62 ;
    RECT 21.41 41.83 21.62 41.9 ;
    RECT 21.41 42.19 21.62 42.26 ;
    RECT 21.41 42.55 21.62 42.62 ;
    RECT 21.87 41.83 22.08 41.9 ;
    RECT 21.87 42.19 22.08 42.26 ;
    RECT 21.87 42.55 22.08 42.62 ;
    RECT 18.09 41.83 18.3 41.9 ;
    RECT 18.09 42.19 18.3 42.26 ;
    RECT 18.09 42.55 18.3 42.62 ;
    RECT 18.55 41.83 18.76 41.9 ;
    RECT 18.55 42.19 18.76 42.26 ;
    RECT 18.55 42.55 18.76 42.62 ;
    RECT 120.825 42.19 120.895 42.26 ;
    RECT 14.77 41.83 14.98 41.9 ;
    RECT 14.77 42.19 14.98 42.26 ;
    RECT 14.77 42.55 14.98 42.62 ;
    RECT 15.23 41.83 15.44 41.9 ;
    RECT 15.23 42.19 15.44 42.26 ;
    RECT 15.23 42.55 15.44 42.62 ;
    RECT 11.45 41.83 11.66 41.9 ;
    RECT 11.45 42.19 11.66 42.26 ;
    RECT 11.45 42.55 11.66 42.62 ;
    RECT 11.91 41.83 12.12 41.9 ;
    RECT 11.91 42.19 12.12 42.26 ;
    RECT 11.91 42.55 12.12 42.62 ;
    RECT 8.13 41.83 8.34 41.9 ;
    RECT 8.13 42.19 8.34 42.26 ;
    RECT 8.13 42.55 8.34 42.62 ;
    RECT 8.59 41.83 8.8 41.9 ;
    RECT 8.59 42.19 8.8 42.26 ;
    RECT 8.59 42.55 8.8 42.62 ;
    RECT 4.81 41.83 5.02 41.9 ;
    RECT 4.81 42.19 5.02 42.26 ;
    RECT 4.81 42.55 5.02 42.62 ;
    RECT 5.27 41.83 5.48 41.9 ;
    RECT 5.27 42.19 5.48 42.26 ;
    RECT 5.27 42.55 5.48 42.62 ;
    RECT 1.49 41.83 1.7 41.9 ;
    RECT 1.49 42.19 1.7 42.26 ;
    RECT 1.49 42.55 1.7 42.62 ;
    RECT 1.95 41.83 2.16 41.9 ;
    RECT 1.95 42.19 2.16 42.26 ;
    RECT 1.95 42.55 2.16 42.62 ;
    RECT 64.57 41.83 64.78 41.9 ;
    RECT 64.57 42.19 64.78 42.26 ;
    RECT 64.57 42.55 64.78 42.62 ;
    RECT 65.03 41.83 65.24 41.9 ;
    RECT 65.03 42.19 65.24 42.26 ;
    RECT 65.03 42.55 65.24 42.62 ;
    RECT 61.25 41.11 61.46 41.18 ;
    RECT 61.25 41.47 61.46 41.54 ;
    RECT 61.25 41.83 61.46 41.9 ;
    RECT 61.71 41.11 61.92 41.18 ;
    RECT 61.71 41.47 61.92 41.54 ;
    RECT 61.71 41.83 61.92 41.9 ;
    RECT 57.93 41.11 58.14 41.18 ;
    RECT 57.93 41.47 58.14 41.54 ;
    RECT 57.93 41.83 58.14 41.9 ;
    RECT 58.39 41.11 58.6 41.18 ;
    RECT 58.39 41.47 58.6 41.54 ;
    RECT 58.39 41.83 58.6 41.9 ;
    RECT 54.61 41.11 54.82 41.18 ;
    RECT 54.61 41.47 54.82 41.54 ;
    RECT 54.61 41.83 54.82 41.9 ;
    RECT 55.07 41.11 55.28 41.18 ;
    RECT 55.07 41.47 55.28 41.54 ;
    RECT 55.07 41.83 55.28 41.9 ;
    RECT 51.29 41.11 51.5 41.18 ;
    RECT 51.29 41.47 51.5 41.54 ;
    RECT 51.29 41.83 51.5 41.9 ;
    RECT 51.75 41.11 51.96 41.18 ;
    RECT 51.75 41.47 51.96 41.54 ;
    RECT 51.75 41.83 51.96 41.9 ;
    RECT 47.97 41.11 48.18 41.18 ;
    RECT 47.97 41.47 48.18 41.54 ;
    RECT 47.97 41.83 48.18 41.9 ;
    RECT 48.43 41.11 48.64 41.18 ;
    RECT 48.43 41.47 48.64 41.54 ;
    RECT 48.43 41.83 48.64 41.9 ;
    RECT 44.65 41.11 44.86 41.18 ;
    RECT 44.65 41.47 44.86 41.54 ;
    RECT 44.65 41.83 44.86 41.9 ;
    RECT 45.11 41.11 45.32 41.18 ;
    RECT 45.11 41.47 45.32 41.54 ;
    RECT 45.11 41.83 45.32 41.9 ;
    RECT 41.33 41.11 41.54 41.18 ;
    RECT 41.33 41.47 41.54 41.54 ;
    RECT 41.33 41.83 41.54 41.9 ;
    RECT 41.79 41.11 42.0 41.18 ;
    RECT 41.79 41.47 42.0 41.54 ;
    RECT 41.79 41.83 42.0 41.9 ;
    RECT 38.01 41.11 38.22 41.18 ;
    RECT 38.01 41.47 38.22 41.54 ;
    RECT 38.01 41.83 38.22 41.9 ;
    RECT 38.47 41.11 38.68 41.18 ;
    RECT 38.47 41.47 38.68 41.54 ;
    RECT 38.47 41.83 38.68 41.9 ;
    RECT 0.4 41.47 0.47 41.54 ;
    RECT 34.69 41.11 34.9 41.18 ;
    RECT 34.69 41.47 34.9 41.54 ;
    RECT 34.69 41.83 34.9 41.9 ;
    RECT 35.15 41.11 35.36 41.18 ;
    RECT 35.15 41.47 35.36 41.54 ;
    RECT 35.15 41.83 35.36 41.9 ;
    RECT 117.69 41.11 117.9 41.18 ;
    RECT 117.69 41.47 117.9 41.54 ;
    RECT 117.69 41.83 117.9 41.9 ;
    RECT 118.15 41.11 118.36 41.18 ;
    RECT 118.15 41.47 118.36 41.54 ;
    RECT 118.15 41.83 118.36 41.9 ;
    RECT 114.37 41.11 114.58 41.18 ;
    RECT 114.37 41.47 114.58 41.54 ;
    RECT 114.37 41.83 114.58 41.9 ;
    RECT 114.83 41.11 115.04 41.18 ;
    RECT 114.83 41.47 115.04 41.54 ;
    RECT 114.83 41.83 115.04 41.9 ;
    RECT 111.05 41.11 111.26 41.18 ;
    RECT 111.05 41.47 111.26 41.54 ;
    RECT 111.05 41.83 111.26 41.9 ;
    RECT 111.51 41.11 111.72 41.18 ;
    RECT 111.51 41.47 111.72 41.54 ;
    RECT 111.51 41.83 111.72 41.9 ;
    RECT 107.73 41.11 107.94 41.18 ;
    RECT 107.73 41.47 107.94 41.54 ;
    RECT 107.73 41.83 107.94 41.9 ;
    RECT 108.19 41.11 108.4 41.18 ;
    RECT 108.19 41.47 108.4 41.54 ;
    RECT 108.19 41.83 108.4 41.9 ;
    RECT 104.41 41.11 104.62 41.18 ;
    RECT 104.41 41.47 104.62 41.54 ;
    RECT 104.41 41.83 104.62 41.9 ;
    RECT 104.87 41.11 105.08 41.18 ;
    RECT 104.87 41.47 105.08 41.54 ;
    RECT 104.87 41.83 105.08 41.9 ;
    RECT 101.09 41.11 101.3 41.18 ;
    RECT 101.09 41.47 101.3 41.54 ;
    RECT 101.09 41.83 101.3 41.9 ;
    RECT 101.55 41.11 101.76 41.18 ;
    RECT 101.55 41.47 101.76 41.54 ;
    RECT 101.55 41.83 101.76 41.9 ;
    RECT 97.77 41.11 97.98 41.18 ;
    RECT 97.77 41.47 97.98 41.54 ;
    RECT 97.77 41.83 97.98 41.9 ;
    RECT 98.23 41.11 98.44 41.18 ;
    RECT 98.23 41.47 98.44 41.54 ;
    RECT 98.23 41.83 98.44 41.9 ;
    RECT 94.45 41.11 94.66 41.18 ;
    RECT 94.45 41.47 94.66 41.54 ;
    RECT 94.45 41.83 94.66 41.9 ;
    RECT 94.91 41.11 95.12 41.18 ;
    RECT 94.91 41.47 95.12 41.54 ;
    RECT 94.91 41.83 95.12 41.9 ;
    RECT 91.13 41.11 91.34 41.18 ;
    RECT 91.13 41.47 91.34 41.54 ;
    RECT 91.13 41.83 91.34 41.9 ;
    RECT 91.59 41.11 91.8 41.18 ;
    RECT 91.59 41.47 91.8 41.54 ;
    RECT 91.59 41.83 91.8 41.9 ;
    RECT 87.81 41.11 88.02 41.18 ;
    RECT 87.81 41.47 88.02 41.54 ;
    RECT 87.81 41.83 88.02 41.9 ;
    RECT 88.27 41.11 88.48 41.18 ;
    RECT 88.27 41.47 88.48 41.54 ;
    RECT 88.27 41.83 88.48 41.9 ;
    RECT 84.49 41.11 84.7 41.18 ;
    RECT 84.49 41.47 84.7 41.54 ;
    RECT 84.49 41.83 84.7 41.9 ;
    RECT 84.95 41.11 85.16 41.18 ;
    RECT 84.95 41.47 85.16 41.54 ;
    RECT 84.95 41.83 85.16 41.9 ;
    RECT 81.17 41.11 81.38 41.18 ;
    RECT 81.17 41.47 81.38 41.54 ;
    RECT 81.17 41.83 81.38 41.9 ;
    RECT 81.63 41.11 81.84 41.18 ;
    RECT 81.63 41.47 81.84 41.54 ;
    RECT 81.63 41.83 81.84 41.9 ;
    RECT 77.85 41.11 78.06 41.18 ;
    RECT 77.85 41.47 78.06 41.54 ;
    RECT 77.85 41.83 78.06 41.9 ;
    RECT 78.31 41.11 78.52 41.18 ;
    RECT 78.31 41.47 78.52 41.54 ;
    RECT 78.31 41.83 78.52 41.9 ;
    RECT 74.53 41.11 74.74 41.18 ;
    RECT 74.53 41.47 74.74 41.54 ;
    RECT 74.53 41.83 74.74 41.9 ;
    RECT 74.99 41.11 75.2 41.18 ;
    RECT 74.99 41.47 75.2 41.54 ;
    RECT 74.99 41.83 75.2 41.9 ;
    RECT 71.21 41.11 71.42 41.18 ;
    RECT 71.21 41.47 71.42 41.54 ;
    RECT 71.21 41.83 71.42 41.9 ;
    RECT 71.67 41.11 71.88 41.18 ;
    RECT 71.67 41.47 71.88 41.54 ;
    RECT 71.67 41.83 71.88 41.9 ;
    RECT 31.37 41.11 31.58 41.18 ;
    RECT 31.37 41.47 31.58 41.54 ;
    RECT 31.37 41.83 31.58 41.9 ;
    RECT 31.83 41.11 32.04 41.18 ;
    RECT 31.83 41.47 32.04 41.54 ;
    RECT 31.83 41.83 32.04 41.9 ;
    RECT 67.89 41.11 68.1 41.18 ;
    RECT 67.89 41.47 68.1 41.54 ;
    RECT 67.89 41.83 68.1 41.9 ;
    RECT 68.35 41.11 68.56 41.18 ;
    RECT 68.35 41.47 68.56 41.54 ;
    RECT 68.35 41.83 68.56 41.9 ;
    RECT 28.05 41.11 28.26 41.18 ;
    RECT 28.05 41.47 28.26 41.54 ;
    RECT 28.05 41.83 28.26 41.9 ;
    RECT 28.51 41.11 28.72 41.18 ;
    RECT 28.51 41.47 28.72 41.54 ;
    RECT 28.51 41.83 28.72 41.9 ;
    RECT 24.73 41.11 24.94 41.18 ;
    RECT 24.73 41.47 24.94 41.54 ;
    RECT 24.73 41.83 24.94 41.9 ;
    RECT 25.19 41.11 25.4 41.18 ;
    RECT 25.19 41.47 25.4 41.54 ;
    RECT 25.19 41.83 25.4 41.9 ;
    RECT 21.41 41.11 21.62 41.18 ;
    RECT 21.41 41.47 21.62 41.54 ;
    RECT 21.41 41.83 21.62 41.9 ;
    RECT 21.87 41.11 22.08 41.18 ;
    RECT 21.87 41.47 22.08 41.54 ;
    RECT 21.87 41.83 22.08 41.9 ;
    RECT 18.09 41.11 18.3 41.18 ;
    RECT 18.09 41.47 18.3 41.54 ;
    RECT 18.09 41.83 18.3 41.9 ;
    RECT 18.55 41.11 18.76 41.18 ;
    RECT 18.55 41.47 18.76 41.54 ;
    RECT 18.55 41.83 18.76 41.9 ;
    RECT 120.825 41.47 120.895 41.54 ;
    RECT 14.77 41.11 14.98 41.18 ;
    RECT 14.77 41.47 14.98 41.54 ;
    RECT 14.77 41.83 14.98 41.9 ;
    RECT 15.23 41.11 15.44 41.18 ;
    RECT 15.23 41.47 15.44 41.54 ;
    RECT 15.23 41.83 15.44 41.9 ;
    RECT 11.45 41.11 11.66 41.18 ;
    RECT 11.45 41.47 11.66 41.54 ;
    RECT 11.45 41.83 11.66 41.9 ;
    RECT 11.91 41.11 12.12 41.18 ;
    RECT 11.91 41.47 12.12 41.54 ;
    RECT 11.91 41.83 12.12 41.9 ;
    RECT 8.13 41.11 8.34 41.18 ;
    RECT 8.13 41.47 8.34 41.54 ;
    RECT 8.13 41.83 8.34 41.9 ;
    RECT 8.59 41.11 8.8 41.18 ;
    RECT 8.59 41.47 8.8 41.54 ;
    RECT 8.59 41.83 8.8 41.9 ;
    RECT 4.81 41.11 5.02 41.18 ;
    RECT 4.81 41.47 5.02 41.54 ;
    RECT 4.81 41.83 5.02 41.9 ;
    RECT 5.27 41.11 5.48 41.18 ;
    RECT 5.27 41.47 5.48 41.54 ;
    RECT 5.27 41.83 5.48 41.9 ;
    RECT 1.49 41.11 1.7 41.18 ;
    RECT 1.49 41.47 1.7 41.54 ;
    RECT 1.49 41.83 1.7 41.9 ;
    RECT 1.95 41.11 2.16 41.18 ;
    RECT 1.95 41.47 2.16 41.54 ;
    RECT 1.95 41.83 2.16 41.9 ;
    RECT 64.57 41.11 64.78 41.18 ;
    RECT 64.57 41.47 64.78 41.54 ;
    RECT 64.57 41.83 64.78 41.9 ;
    RECT 65.03 41.11 65.24 41.18 ;
    RECT 65.03 41.47 65.24 41.54 ;
    RECT 65.03 41.83 65.24 41.9 ;
    RECT 61.25 40.39 61.46 40.46 ;
    RECT 61.25 40.75 61.46 40.82 ;
    RECT 61.25 41.11 61.46 41.18 ;
    RECT 61.71 40.39 61.92 40.46 ;
    RECT 61.71 40.75 61.92 40.82 ;
    RECT 61.71 41.11 61.92 41.18 ;
    RECT 57.93 40.39 58.14 40.46 ;
    RECT 57.93 40.75 58.14 40.82 ;
    RECT 57.93 41.11 58.14 41.18 ;
    RECT 58.39 40.39 58.6 40.46 ;
    RECT 58.39 40.75 58.6 40.82 ;
    RECT 58.39 41.11 58.6 41.18 ;
    RECT 54.61 40.39 54.82 40.46 ;
    RECT 54.61 40.75 54.82 40.82 ;
    RECT 54.61 41.11 54.82 41.18 ;
    RECT 55.07 40.39 55.28 40.46 ;
    RECT 55.07 40.75 55.28 40.82 ;
    RECT 55.07 41.11 55.28 41.18 ;
    RECT 51.29 40.39 51.5 40.46 ;
    RECT 51.29 40.75 51.5 40.82 ;
    RECT 51.29 41.11 51.5 41.18 ;
    RECT 51.75 40.39 51.96 40.46 ;
    RECT 51.75 40.75 51.96 40.82 ;
    RECT 51.75 41.11 51.96 41.18 ;
    RECT 47.97 40.39 48.18 40.46 ;
    RECT 47.97 40.75 48.18 40.82 ;
    RECT 47.97 41.11 48.18 41.18 ;
    RECT 48.43 40.39 48.64 40.46 ;
    RECT 48.43 40.75 48.64 40.82 ;
    RECT 48.43 41.11 48.64 41.18 ;
    RECT 44.65 40.39 44.86 40.46 ;
    RECT 44.65 40.75 44.86 40.82 ;
    RECT 44.65 41.11 44.86 41.18 ;
    RECT 45.11 40.39 45.32 40.46 ;
    RECT 45.11 40.75 45.32 40.82 ;
    RECT 45.11 41.11 45.32 41.18 ;
    RECT 41.33 40.39 41.54 40.46 ;
    RECT 41.33 40.75 41.54 40.82 ;
    RECT 41.33 41.11 41.54 41.18 ;
    RECT 41.79 40.39 42.0 40.46 ;
    RECT 41.79 40.75 42.0 40.82 ;
    RECT 41.79 41.11 42.0 41.18 ;
    RECT 38.01 40.39 38.22 40.46 ;
    RECT 38.01 40.75 38.22 40.82 ;
    RECT 38.01 41.11 38.22 41.18 ;
    RECT 38.47 40.39 38.68 40.46 ;
    RECT 38.47 40.75 38.68 40.82 ;
    RECT 38.47 41.11 38.68 41.18 ;
    RECT 0.4 40.75 0.47 40.82 ;
    RECT 34.69 40.39 34.9 40.46 ;
    RECT 34.69 40.75 34.9 40.82 ;
    RECT 34.69 41.11 34.9 41.18 ;
    RECT 35.15 40.39 35.36 40.46 ;
    RECT 35.15 40.75 35.36 40.82 ;
    RECT 35.15 41.11 35.36 41.18 ;
    RECT 117.69 40.39 117.9 40.46 ;
    RECT 117.69 40.75 117.9 40.82 ;
    RECT 117.69 41.11 117.9 41.18 ;
    RECT 118.15 40.39 118.36 40.46 ;
    RECT 118.15 40.75 118.36 40.82 ;
    RECT 118.15 41.11 118.36 41.18 ;
    RECT 114.37 40.39 114.58 40.46 ;
    RECT 114.37 40.75 114.58 40.82 ;
    RECT 114.37 41.11 114.58 41.18 ;
    RECT 114.83 40.39 115.04 40.46 ;
    RECT 114.83 40.75 115.04 40.82 ;
    RECT 114.83 41.11 115.04 41.18 ;
    RECT 111.05 40.39 111.26 40.46 ;
    RECT 111.05 40.75 111.26 40.82 ;
    RECT 111.05 41.11 111.26 41.18 ;
    RECT 111.51 40.39 111.72 40.46 ;
    RECT 111.51 40.75 111.72 40.82 ;
    RECT 111.51 41.11 111.72 41.18 ;
    RECT 107.73 40.39 107.94 40.46 ;
    RECT 107.73 40.75 107.94 40.82 ;
    RECT 107.73 41.11 107.94 41.18 ;
    RECT 108.19 40.39 108.4 40.46 ;
    RECT 108.19 40.75 108.4 40.82 ;
    RECT 108.19 41.11 108.4 41.18 ;
    RECT 104.41 40.39 104.62 40.46 ;
    RECT 104.41 40.75 104.62 40.82 ;
    RECT 104.41 41.11 104.62 41.18 ;
    RECT 104.87 40.39 105.08 40.46 ;
    RECT 104.87 40.75 105.08 40.82 ;
    RECT 104.87 41.11 105.08 41.18 ;
    RECT 101.09 40.39 101.3 40.46 ;
    RECT 101.09 40.75 101.3 40.82 ;
    RECT 101.09 41.11 101.3 41.18 ;
    RECT 101.55 40.39 101.76 40.46 ;
    RECT 101.55 40.75 101.76 40.82 ;
    RECT 101.55 41.11 101.76 41.18 ;
    RECT 97.77 40.39 97.98 40.46 ;
    RECT 97.77 40.75 97.98 40.82 ;
    RECT 97.77 41.11 97.98 41.18 ;
    RECT 98.23 40.39 98.44 40.46 ;
    RECT 98.23 40.75 98.44 40.82 ;
    RECT 98.23 41.11 98.44 41.18 ;
    RECT 94.45 40.39 94.66 40.46 ;
    RECT 94.45 40.75 94.66 40.82 ;
    RECT 94.45 41.11 94.66 41.18 ;
    RECT 94.91 40.39 95.12 40.46 ;
    RECT 94.91 40.75 95.12 40.82 ;
    RECT 94.91 41.11 95.12 41.18 ;
    RECT 91.13 40.39 91.34 40.46 ;
    RECT 91.13 40.75 91.34 40.82 ;
    RECT 91.13 41.11 91.34 41.18 ;
    RECT 91.59 40.39 91.8 40.46 ;
    RECT 91.59 40.75 91.8 40.82 ;
    RECT 91.59 41.11 91.8 41.18 ;
    RECT 87.81 40.39 88.02 40.46 ;
    RECT 87.81 40.75 88.02 40.82 ;
    RECT 87.81 41.11 88.02 41.18 ;
    RECT 88.27 40.39 88.48 40.46 ;
    RECT 88.27 40.75 88.48 40.82 ;
    RECT 88.27 41.11 88.48 41.18 ;
    RECT 84.49 40.39 84.7 40.46 ;
    RECT 84.49 40.75 84.7 40.82 ;
    RECT 84.49 41.11 84.7 41.18 ;
    RECT 84.95 40.39 85.16 40.46 ;
    RECT 84.95 40.75 85.16 40.82 ;
    RECT 84.95 41.11 85.16 41.18 ;
    RECT 81.17 40.39 81.38 40.46 ;
    RECT 81.17 40.75 81.38 40.82 ;
    RECT 81.17 41.11 81.38 41.18 ;
    RECT 81.63 40.39 81.84 40.46 ;
    RECT 81.63 40.75 81.84 40.82 ;
    RECT 81.63 41.11 81.84 41.18 ;
    RECT 77.85 40.39 78.06 40.46 ;
    RECT 77.85 40.75 78.06 40.82 ;
    RECT 77.85 41.11 78.06 41.18 ;
    RECT 78.31 40.39 78.52 40.46 ;
    RECT 78.31 40.75 78.52 40.82 ;
    RECT 78.31 41.11 78.52 41.18 ;
    RECT 74.53 40.39 74.74 40.46 ;
    RECT 74.53 40.75 74.74 40.82 ;
    RECT 74.53 41.11 74.74 41.18 ;
    RECT 74.99 40.39 75.2 40.46 ;
    RECT 74.99 40.75 75.2 40.82 ;
    RECT 74.99 41.11 75.2 41.18 ;
    RECT 71.21 40.39 71.42 40.46 ;
    RECT 71.21 40.75 71.42 40.82 ;
    RECT 71.21 41.11 71.42 41.18 ;
    RECT 71.67 40.39 71.88 40.46 ;
    RECT 71.67 40.75 71.88 40.82 ;
    RECT 71.67 41.11 71.88 41.18 ;
    RECT 31.37 40.39 31.58 40.46 ;
    RECT 31.37 40.75 31.58 40.82 ;
    RECT 31.37 41.11 31.58 41.18 ;
    RECT 31.83 40.39 32.04 40.46 ;
    RECT 31.83 40.75 32.04 40.82 ;
    RECT 31.83 41.11 32.04 41.18 ;
    RECT 67.89 40.39 68.1 40.46 ;
    RECT 67.89 40.75 68.1 40.82 ;
    RECT 67.89 41.11 68.1 41.18 ;
    RECT 68.35 40.39 68.56 40.46 ;
    RECT 68.35 40.75 68.56 40.82 ;
    RECT 68.35 41.11 68.56 41.18 ;
    RECT 28.05 40.39 28.26 40.46 ;
    RECT 28.05 40.75 28.26 40.82 ;
    RECT 28.05 41.11 28.26 41.18 ;
    RECT 28.51 40.39 28.72 40.46 ;
    RECT 28.51 40.75 28.72 40.82 ;
    RECT 28.51 41.11 28.72 41.18 ;
    RECT 24.73 40.39 24.94 40.46 ;
    RECT 24.73 40.75 24.94 40.82 ;
    RECT 24.73 41.11 24.94 41.18 ;
    RECT 25.19 40.39 25.4 40.46 ;
    RECT 25.19 40.75 25.4 40.82 ;
    RECT 25.19 41.11 25.4 41.18 ;
    RECT 21.41 40.39 21.62 40.46 ;
    RECT 21.41 40.75 21.62 40.82 ;
    RECT 21.41 41.11 21.62 41.18 ;
    RECT 21.87 40.39 22.08 40.46 ;
    RECT 21.87 40.75 22.08 40.82 ;
    RECT 21.87 41.11 22.08 41.18 ;
    RECT 18.09 40.39 18.3 40.46 ;
    RECT 18.09 40.75 18.3 40.82 ;
    RECT 18.09 41.11 18.3 41.18 ;
    RECT 18.55 40.39 18.76 40.46 ;
    RECT 18.55 40.75 18.76 40.82 ;
    RECT 18.55 41.11 18.76 41.18 ;
    RECT 120.825 40.75 120.895 40.82 ;
    RECT 14.77 40.39 14.98 40.46 ;
    RECT 14.77 40.75 14.98 40.82 ;
    RECT 14.77 41.11 14.98 41.18 ;
    RECT 15.23 40.39 15.44 40.46 ;
    RECT 15.23 40.75 15.44 40.82 ;
    RECT 15.23 41.11 15.44 41.18 ;
    RECT 11.45 40.39 11.66 40.46 ;
    RECT 11.45 40.75 11.66 40.82 ;
    RECT 11.45 41.11 11.66 41.18 ;
    RECT 11.91 40.39 12.12 40.46 ;
    RECT 11.91 40.75 12.12 40.82 ;
    RECT 11.91 41.11 12.12 41.18 ;
    RECT 8.13 40.39 8.34 40.46 ;
    RECT 8.13 40.75 8.34 40.82 ;
    RECT 8.13 41.11 8.34 41.18 ;
    RECT 8.59 40.39 8.8 40.46 ;
    RECT 8.59 40.75 8.8 40.82 ;
    RECT 8.59 41.11 8.8 41.18 ;
    RECT 4.81 40.39 5.02 40.46 ;
    RECT 4.81 40.75 5.02 40.82 ;
    RECT 4.81 41.11 5.02 41.18 ;
    RECT 5.27 40.39 5.48 40.46 ;
    RECT 5.27 40.75 5.48 40.82 ;
    RECT 5.27 41.11 5.48 41.18 ;
    RECT 1.49 40.39 1.7 40.46 ;
    RECT 1.49 40.75 1.7 40.82 ;
    RECT 1.49 41.11 1.7 41.18 ;
    RECT 1.95 40.39 2.16 40.46 ;
    RECT 1.95 40.75 2.16 40.82 ;
    RECT 1.95 41.11 2.16 41.18 ;
    RECT 64.57 40.39 64.78 40.46 ;
    RECT 64.57 40.75 64.78 40.82 ;
    RECT 64.57 41.11 64.78 41.18 ;
    RECT 65.03 40.39 65.24 40.46 ;
    RECT 65.03 40.75 65.24 40.82 ;
    RECT 65.03 41.11 65.24 41.18 ;
    RECT 61.25 39.67 61.46 39.74 ;
    RECT 61.25 40.03 61.46 40.1 ;
    RECT 61.25 40.39 61.46 40.46 ;
    RECT 61.71 39.67 61.92 39.74 ;
    RECT 61.71 40.03 61.92 40.1 ;
    RECT 61.71 40.39 61.92 40.46 ;
    RECT 57.93 39.67 58.14 39.74 ;
    RECT 57.93 40.03 58.14 40.1 ;
    RECT 57.93 40.39 58.14 40.46 ;
    RECT 58.39 39.67 58.6 39.74 ;
    RECT 58.39 40.03 58.6 40.1 ;
    RECT 58.39 40.39 58.6 40.46 ;
    RECT 54.61 39.67 54.82 39.74 ;
    RECT 54.61 40.03 54.82 40.1 ;
    RECT 54.61 40.39 54.82 40.46 ;
    RECT 55.07 39.67 55.28 39.74 ;
    RECT 55.07 40.03 55.28 40.1 ;
    RECT 55.07 40.39 55.28 40.46 ;
    RECT 51.29 39.67 51.5 39.74 ;
    RECT 51.29 40.03 51.5 40.1 ;
    RECT 51.29 40.39 51.5 40.46 ;
    RECT 51.75 39.67 51.96 39.74 ;
    RECT 51.75 40.03 51.96 40.1 ;
    RECT 51.75 40.39 51.96 40.46 ;
    RECT 47.97 39.67 48.18 39.74 ;
    RECT 47.97 40.03 48.18 40.1 ;
    RECT 47.97 40.39 48.18 40.46 ;
    RECT 48.43 39.67 48.64 39.74 ;
    RECT 48.43 40.03 48.64 40.1 ;
    RECT 48.43 40.39 48.64 40.46 ;
    RECT 44.65 39.67 44.86 39.74 ;
    RECT 44.65 40.03 44.86 40.1 ;
    RECT 44.65 40.39 44.86 40.46 ;
    RECT 45.11 39.67 45.32 39.74 ;
    RECT 45.11 40.03 45.32 40.1 ;
    RECT 45.11 40.39 45.32 40.46 ;
    RECT 41.33 39.67 41.54 39.74 ;
    RECT 41.33 40.03 41.54 40.1 ;
    RECT 41.33 40.39 41.54 40.46 ;
    RECT 41.79 39.67 42.0 39.74 ;
    RECT 41.79 40.03 42.0 40.1 ;
    RECT 41.79 40.39 42.0 40.46 ;
    RECT 38.01 39.67 38.22 39.74 ;
    RECT 38.01 40.03 38.22 40.1 ;
    RECT 38.01 40.39 38.22 40.46 ;
    RECT 38.47 39.67 38.68 39.74 ;
    RECT 38.47 40.03 38.68 40.1 ;
    RECT 38.47 40.39 38.68 40.46 ;
    RECT 0.4 40.03 0.47 40.1 ;
    RECT 34.69 39.67 34.9 39.74 ;
    RECT 34.69 40.03 34.9 40.1 ;
    RECT 34.69 40.39 34.9 40.46 ;
    RECT 35.15 39.67 35.36 39.74 ;
    RECT 35.15 40.03 35.36 40.1 ;
    RECT 35.15 40.39 35.36 40.46 ;
    RECT 117.69 39.67 117.9 39.74 ;
    RECT 117.69 40.03 117.9 40.1 ;
    RECT 117.69 40.39 117.9 40.46 ;
    RECT 118.15 39.67 118.36 39.74 ;
    RECT 118.15 40.03 118.36 40.1 ;
    RECT 118.15 40.39 118.36 40.46 ;
    RECT 114.37 39.67 114.58 39.74 ;
    RECT 114.37 40.03 114.58 40.1 ;
    RECT 114.37 40.39 114.58 40.46 ;
    RECT 114.83 39.67 115.04 39.74 ;
    RECT 114.83 40.03 115.04 40.1 ;
    RECT 114.83 40.39 115.04 40.46 ;
    RECT 111.05 39.67 111.26 39.74 ;
    RECT 111.05 40.03 111.26 40.1 ;
    RECT 111.05 40.39 111.26 40.46 ;
    RECT 111.51 39.67 111.72 39.74 ;
    RECT 111.51 40.03 111.72 40.1 ;
    RECT 111.51 40.39 111.72 40.46 ;
    RECT 107.73 39.67 107.94 39.74 ;
    RECT 107.73 40.03 107.94 40.1 ;
    RECT 107.73 40.39 107.94 40.46 ;
    RECT 108.19 39.67 108.4 39.74 ;
    RECT 108.19 40.03 108.4 40.1 ;
    RECT 108.19 40.39 108.4 40.46 ;
    RECT 104.41 39.67 104.62 39.74 ;
    RECT 104.41 40.03 104.62 40.1 ;
    RECT 104.41 40.39 104.62 40.46 ;
    RECT 104.87 39.67 105.08 39.74 ;
    RECT 104.87 40.03 105.08 40.1 ;
    RECT 104.87 40.39 105.08 40.46 ;
    RECT 101.09 39.67 101.3 39.74 ;
    RECT 101.09 40.03 101.3 40.1 ;
    RECT 101.09 40.39 101.3 40.46 ;
    RECT 101.55 39.67 101.76 39.74 ;
    RECT 101.55 40.03 101.76 40.1 ;
    RECT 101.55 40.39 101.76 40.46 ;
    RECT 97.77 39.67 97.98 39.74 ;
    RECT 97.77 40.03 97.98 40.1 ;
    RECT 97.77 40.39 97.98 40.46 ;
    RECT 98.23 39.67 98.44 39.74 ;
    RECT 98.23 40.03 98.44 40.1 ;
    RECT 98.23 40.39 98.44 40.46 ;
    RECT 94.45 39.67 94.66 39.74 ;
    RECT 94.45 40.03 94.66 40.1 ;
    RECT 94.45 40.39 94.66 40.46 ;
    RECT 94.91 39.67 95.12 39.74 ;
    RECT 94.91 40.03 95.12 40.1 ;
    RECT 94.91 40.39 95.12 40.46 ;
    RECT 91.13 39.67 91.34 39.74 ;
    RECT 91.13 40.03 91.34 40.1 ;
    RECT 91.13 40.39 91.34 40.46 ;
    RECT 91.59 39.67 91.8 39.74 ;
    RECT 91.59 40.03 91.8 40.1 ;
    RECT 91.59 40.39 91.8 40.46 ;
    RECT 87.81 39.67 88.02 39.74 ;
    RECT 87.81 40.03 88.02 40.1 ;
    RECT 87.81 40.39 88.02 40.46 ;
    RECT 88.27 39.67 88.48 39.74 ;
    RECT 88.27 40.03 88.48 40.1 ;
    RECT 88.27 40.39 88.48 40.46 ;
    RECT 84.49 39.67 84.7 39.74 ;
    RECT 84.49 40.03 84.7 40.1 ;
    RECT 84.49 40.39 84.7 40.46 ;
    RECT 84.95 39.67 85.16 39.74 ;
    RECT 84.95 40.03 85.16 40.1 ;
    RECT 84.95 40.39 85.16 40.46 ;
    RECT 81.17 39.67 81.38 39.74 ;
    RECT 81.17 40.03 81.38 40.1 ;
    RECT 81.17 40.39 81.38 40.46 ;
    RECT 81.63 39.67 81.84 39.74 ;
    RECT 81.63 40.03 81.84 40.1 ;
    RECT 81.63 40.39 81.84 40.46 ;
    RECT 77.85 39.67 78.06 39.74 ;
    RECT 77.85 40.03 78.06 40.1 ;
    RECT 77.85 40.39 78.06 40.46 ;
    RECT 78.31 39.67 78.52 39.74 ;
    RECT 78.31 40.03 78.52 40.1 ;
    RECT 78.31 40.39 78.52 40.46 ;
    RECT 74.53 39.67 74.74 39.74 ;
    RECT 74.53 40.03 74.74 40.1 ;
    RECT 74.53 40.39 74.74 40.46 ;
    RECT 74.99 39.67 75.2 39.74 ;
    RECT 74.99 40.03 75.2 40.1 ;
    RECT 74.99 40.39 75.2 40.46 ;
    RECT 71.21 39.67 71.42 39.74 ;
    RECT 71.21 40.03 71.42 40.1 ;
    RECT 71.21 40.39 71.42 40.46 ;
    RECT 71.67 39.67 71.88 39.74 ;
    RECT 71.67 40.03 71.88 40.1 ;
    RECT 71.67 40.39 71.88 40.46 ;
    RECT 31.37 39.67 31.58 39.74 ;
    RECT 31.37 40.03 31.58 40.1 ;
    RECT 31.37 40.39 31.58 40.46 ;
    RECT 31.83 39.67 32.04 39.74 ;
    RECT 31.83 40.03 32.04 40.1 ;
    RECT 31.83 40.39 32.04 40.46 ;
    RECT 67.89 39.67 68.1 39.74 ;
    RECT 67.89 40.03 68.1 40.1 ;
    RECT 67.89 40.39 68.1 40.46 ;
    RECT 68.35 39.67 68.56 39.74 ;
    RECT 68.35 40.03 68.56 40.1 ;
    RECT 68.35 40.39 68.56 40.46 ;
    RECT 28.05 39.67 28.26 39.74 ;
    RECT 28.05 40.03 28.26 40.1 ;
    RECT 28.05 40.39 28.26 40.46 ;
    RECT 28.51 39.67 28.72 39.74 ;
    RECT 28.51 40.03 28.72 40.1 ;
    RECT 28.51 40.39 28.72 40.46 ;
    RECT 24.73 39.67 24.94 39.74 ;
    RECT 24.73 40.03 24.94 40.1 ;
    RECT 24.73 40.39 24.94 40.46 ;
    RECT 25.19 39.67 25.4 39.74 ;
    RECT 25.19 40.03 25.4 40.1 ;
    RECT 25.19 40.39 25.4 40.46 ;
    RECT 21.41 39.67 21.62 39.74 ;
    RECT 21.41 40.03 21.62 40.1 ;
    RECT 21.41 40.39 21.62 40.46 ;
    RECT 21.87 39.67 22.08 39.74 ;
    RECT 21.87 40.03 22.08 40.1 ;
    RECT 21.87 40.39 22.08 40.46 ;
    RECT 18.09 39.67 18.3 39.74 ;
    RECT 18.09 40.03 18.3 40.1 ;
    RECT 18.09 40.39 18.3 40.46 ;
    RECT 18.55 39.67 18.76 39.74 ;
    RECT 18.55 40.03 18.76 40.1 ;
    RECT 18.55 40.39 18.76 40.46 ;
    RECT 120.825 40.03 120.895 40.1 ;
    RECT 14.77 39.67 14.98 39.74 ;
    RECT 14.77 40.03 14.98 40.1 ;
    RECT 14.77 40.39 14.98 40.46 ;
    RECT 15.23 39.67 15.44 39.74 ;
    RECT 15.23 40.03 15.44 40.1 ;
    RECT 15.23 40.39 15.44 40.46 ;
    RECT 11.45 39.67 11.66 39.74 ;
    RECT 11.45 40.03 11.66 40.1 ;
    RECT 11.45 40.39 11.66 40.46 ;
    RECT 11.91 39.67 12.12 39.74 ;
    RECT 11.91 40.03 12.12 40.1 ;
    RECT 11.91 40.39 12.12 40.46 ;
    RECT 8.13 39.67 8.34 39.74 ;
    RECT 8.13 40.03 8.34 40.1 ;
    RECT 8.13 40.39 8.34 40.46 ;
    RECT 8.59 39.67 8.8 39.74 ;
    RECT 8.59 40.03 8.8 40.1 ;
    RECT 8.59 40.39 8.8 40.46 ;
    RECT 4.81 39.67 5.02 39.74 ;
    RECT 4.81 40.03 5.02 40.1 ;
    RECT 4.81 40.39 5.02 40.46 ;
    RECT 5.27 39.67 5.48 39.74 ;
    RECT 5.27 40.03 5.48 40.1 ;
    RECT 5.27 40.39 5.48 40.46 ;
    RECT 1.49 39.67 1.7 39.74 ;
    RECT 1.49 40.03 1.7 40.1 ;
    RECT 1.49 40.39 1.7 40.46 ;
    RECT 1.95 39.67 2.16 39.74 ;
    RECT 1.95 40.03 2.16 40.1 ;
    RECT 1.95 40.39 2.16 40.46 ;
    RECT 64.57 39.67 64.78 39.74 ;
    RECT 64.57 40.03 64.78 40.1 ;
    RECT 64.57 40.39 64.78 40.46 ;
    RECT 65.03 39.67 65.24 39.74 ;
    RECT 65.03 40.03 65.24 40.1 ;
    RECT 65.03 40.39 65.24 40.46 ;
    RECT 61.25 79.29 61.46 79.36 ;
    RECT 61.25 79.65 61.46 79.72 ;
    RECT 61.25 80.01 61.46 80.08 ;
    RECT 61.71 79.29 61.92 79.36 ;
    RECT 61.71 79.65 61.92 79.72 ;
    RECT 61.71 80.01 61.92 80.08 ;
    RECT 57.93 79.29 58.14 79.36 ;
    RECT 57.93 79.65 58.14 79.72 ;
    RECT 57.93 80.01 58.14 80.08 ;
    RECT 58.39 79.29 58.6 79.36 ;
    RECT 58.39 79.65 58.6 79.72 ;
    RECT 58.39 80.01 58.6 80.08 ;
    RECT 54.61 79.29 54.82 79.36 ;
    RECT 54.61 79.65 54.82 79.72 ;
    RECT 54.61 80.01 54.82 80.08 ;
    RECT 55.07 79.29 55.28 79.36 ;
    RECT 55.07 79.65 55.28 79.72 ;
    RECT 55.07 80.01 55.28 80.08 ;
    RECT 51.29 79.29 51.5 79.36 ;
    RECT 51.29 79.65 51.5 79.72 ;
    RECT 51.29 80.01 51.5 80.08 ;
    RECT 51.75 79.29 51.96 79.36 ;
    RECT 51.75 79.65 51.96 79.72 ;
    RECT 51.75 80.01 51.96 80.08 ;
    RECT 47.97 79.29 48.18 79.36 ;
    RECT 47.97 79.65 48.18 79.72 ;
    RECT 47.97 80.01 48.18 80.08 ;
    RECT 48.43 79.29 48.64 79.36 ;
    RECT 48.43 79.65 48.64 79.72 ;
    RECT 48.43 80.01 48.64 80.08 ;
    RECT 44.65 79.29 44.86 79.36 ;
    RECT 44.65 79.65 44.86 79.72 ;
    RECT 44.65 80.01 44.86 80.08 ;
    RECT 45.11 79.29 45.32 79.36 ;
    RECT 45.11 79.65 45.32 79.72 ;
    RECT 45.11 80.01 45.32 80.08 ;
    RECT 41.33 79.29 41.54 79.36 ;
    RECT 41.33 79.65 41.54 79.72 ;
    RECT 41.33 80.01 41.54 80.08 ;
    RECT 41.79 79.29 42.0 79.36 ;
    RECT 41.79 79.65 42.0 79.72 ;
    RECT 41.79 80.01 42.0 80.08 ;
    RECT 38.01 79.29 38.22 79.36 ;
    RECT 38.01 79.65 38.22 79.72 ;
    RECT 38.01 80.01 38.22 80.08 ;
    RECT 38.47 79.29 38.68 79.36 ;
    RECT 38.47 79.65 38.68 79.72 ;
    RECT 38.47 80.01 38.68 80.08 ;
    RECT 0.4 79.65 0.47 79.72 ;
    RECT 34.69 79.29 34.9 79.36 ;
    RECT 34.69 79.65 34.9 79.72 ;
    RECT 34.69 80.01 34.9 80.08 ;
    RECT 35.15 79.29 35.36 79.36 ;
    RECT 35.15 79.65 35.36 79.72 ;
    RECT 35.15 80.01 35.36 80.08 ;
    RECT 117.69 79.29 117.9 79.36 ;
    RECT 117.69 79.65 117.9 79.72 ;
    RECT 117.69 80.01 117.9 80.08 ;
    RECT 118.15 79.29 118.36 79.36 ;
    RECT 118.15 79.65 118.36 79.72 ;
    RECT 118.15 80.01 118.36 80.08 ;
    RECT 114.37 79.29 114.58 79.36 ;
    RECT 114.37 79.65 114.58 79.72 ;
    RECT 114.37 80.01 114.58 80.08 ;
    RECT 114.83 79.29 115.04 79.36 ;
    RECT 114.83 79.65 115.04 79.72 ;
    RECT 114.83 80.01 115.04 80.08 ;
    RECT 111.05 79.29 111.26 79.36 ;
    RECT 111.05 79.65 111.26 79.72 ;
    RECT 111.05 80.01 111.26 80.08 ;
    RECT 111.51 79.29 111.72 79.36 ;
    RECT 111.51 79.65 111.72 79.72 ;
    RECT 111.51 80.01 111.72 80.08 ;
    RECT 107.73 79.29 107.94 79.36 ;
    RECT 107.73 79.65 107.94 79.72 ;
    RECT 107.73 80.01 107.94 80.08 ;
    RECT 108.19 79.29 108.4 79.36 ;
    RECT 108.19 79.65 108.4 79.72 ;
    RECT 108.19 80.01 108.4 80.08 ;
    RECT 104.41 79.29 104.62 79.36 ;
    RECT 104.41 79.65 104.62 79.72 ;
    RECT 104.41 80.01 104.62 80.08 ;
    RECT 104.87 79.29 105.08 79.36 ;
    RECT 104.87 79.65 105.08 79.72 ;
    RECT 104.87 80.01 105.08 80.08 ;
    RECT 101.09 79.29 101.3 79.36 ;
    RECT 101.09 79.65 101.3 79.72 ;
    RECT 101.09 80.01 101.3 80.08 ;
    RECT 101.55 79.29 101.76 79.36 ;
    RECT 101.55 79.65 101.76 79.72 ;
    RECT 101.55 80.01 101.76 80.08 ;
    RECT 97.77 79.29 97.98 79.36 ;
    RECT 97.77 79.65 97.98 79.72 ;
    RECT 97.77 80.01 97.98 80.08 ;
    RECT 98.23 79.29 98.44 79.36 ;
    RECT 98.23 79.65 98.44 79.72 ;
    RECT 98.23 80.01 98.44 80.08 ;
    RECT 94.45 79.29 94.66 79.36 ;
    RECT 94.45 79.65 94.66 79.72 ;
    RECT 94.45 80.01 94.66 80.08 ;
    RECT 94.91 79.29 95.12 79.36 ;
    RECT 94.91 79.65 95.12 79.72 ;
    RECT 94.91 80.01 95.12 80.08 ;
    RECT 91.13 79.29 91.34 79.36 ;
    RECT 91.13 79.65 91.34 79.72 ;
    RECT 91.13 80.01 91.34 80.08 ;
    RECT 91.59 79.29 91.8 79.36 ;
    RECT 91.59 79.65 91.8 79.72 ;
    RECT 91.59 80.01 91.8 80.08 ;
    RECT 87.81 79.29 88.02 79.36 ;
    RECT 87.81 79.65 88.02 79.72 ;
    RECT 87.81 80.01 88.02 80.08 ;
    RECT 88.27 79.29 88.48 79.36 ;
    RECT 88.27 79.65 88.48 79.72 ;
    RECT 88.27 80.01 88.48 80.08 ;
    RECT 84.49 79.29 84.7 79.36 ;
    RECT 84.49 79.65 84.7 79.72 ;
    RECT 84.49 80.01 84.7 80.08 ;
    RECT 84.95 79.29 85.16 79.36 ;
    RECT 84.95 79.65 85.16 79.72 ;
    RECT 84.95 80.01 85.16 80.08 ;
    RECT 81.17 79.29 81.38 79.36 ;
    RECT 81.17 79.65 81.38 79.72 ;
    RECT 81.17 80.01 81.38 80.08 ;
    RECT 81.63 79.29 81.84 79.36 ;
    RECT 81.63 79.65 81.84 79.72 ;
    RECT 81.63 80.01 81.84 80.08 ;
    RECT 77.85 79.29 78.06 79.36 ;
    RECT 77.85 79.65 78.06 79.72 ;
    RECT 77.85 80.01 78.06 80.08 ;
    RECT 78.31 79.29 78.52 79.36 ;
    RECT 78.31 79.65 78.52 79.72 ;
    RECT 78.31 80.01 78.52 80.08 ;
    RECT 74.53 79.29 74.74 79.36 ;
    RECT 74.53 79.65 74.74 79.72 ;
    RECT 74.53 80.01 74.74 80.08 ;
    RECT 74.99 79.29 75.2 79.36 ;
    RECT 74.99 79.65 75.2 79.72 ;
    RECT 74.99 80.01 75.2 80.08 ;
    RECT 71.21 79.29 71.42 79.36 ;
    RECT 71.21 79.65 71.42 79.72 ;
    RECT 71.21 80.01 71.42 80.08 ;
    RECT 71.67 79.29 71.88 79.36 ;
    RECT 71.67 79.65 71.88 79.72 ;
    RECT 71.67 80.01 71.88 80.08 ;
    RECT 31.37 79.29 31.58 79.36 ;
    RECT 31.37 79.65 31.58 79.72 ;
    RECT 31.37 80.01 31.58 80.08 ;
    RECT 31.83 79.29 32.04 79.36 ;
    RECT 31.83 79.65 32.04 79.72 ;
    RECT 31.83 80.01 32.04 80.08 ;
    RECT 67.89 79.29 68.1 79.36 ;
    RECT 67.89 79.65 68.1 79.72 ;
    RECT 67.89 80.01 68.1 80.08 ;
    RECT 68.35 79.29 68.56 79.36 ;
    RECT 68.35 79.65 68.56 79.72 ;
    RECT 68.35 80.01 68.56 80.08 ;
    RECT 28.05 79.29 28.26 79.36 ;
    RECT 28.05 79.65 28.26 79.72 ;
    RECT 28.05 80.01 28.26 80.08 ;
    RECT 28.51 79.29 28.72 79.36 ;
    RECT 28.51 79.65 28.72 79.72 ;
    RECT 28.51 80.01 28.72 80.08 ;
    RECT 24.73 79.29 24.94 79.36 ;
    RECT 24.73 79.65 24.94 79.72 ;
    RECT 24.73 80.01 24.94 80.08 ;
    RECT 25.19 79.29 25.4 79.36 ;
    RECT 25.19 79.65 25.4 79.72 ;
    RECT 25.19 80.01 25.4 80.08 ;
    RECT 21.41 79.29 21.62 79.36 ;
    RECT 21.41 79.65 21.62 79.72 ;
    RECT 21.41 80.01 21.62 80.08 ;
    RECT 21.87 79.29 22.08 79.36 ;
    RECT 21.87 79.65 22.08 79.72 ;
    RECT 21.87 80.01 22.08 80.08 ;
    RECT 18.09 79.29 18.3 79.36 ;
    RECT 18.09 79.65 18.3 79.72 ;
    RECT 18.09 80.01 18.3 80.08 ;
    RECT 18.55 79.29 18.76 79.36 ;
    RECT 18.55 79.65 18.76 79.72 ;
    RECT 18.55 80.01 18.76 80.08 ;
    RECT 120.825 79.65 120.895 79.72 ;
    RECT 14.77 79.29 14.98 79.36 ;
    RECT 14.77 79.65 14.98 79.72 ;
    RECT 14.77 80.01 14.98 80.08 ;
    RECT 15.23 79.29 15.44 79.36 ;
    RECT 15.23 79.65 15.44 79.72 ;
    RECT 15.23 80.01 15.44 80.08 ;
    RECT 11.45 79.29 11.66 79.36 ;
    RECT 11.45 79.65 11.66 79.72 ;
    RECT 11.45 80.01 11.66 80.08 ;
    RECT 11.91 79.29 12.12 79.36 ;
    RECT 11.91 79.65 12.12 79.72 ;
    RECT 11.91 80.01 12.12 80.08 ;
    RECT 8.13 79.29 8.34 79.36 ;
    RECT 8.13 79.65 8.34 79.72 ;
    RECT 8.13 80.01 8.34 80.08 ;
    RECT 8.59 79.29 8.8 79.36 ;
    RECT 8.59 79.65 8.8 79.72 ;
    RECT 8.59 80.01 8.8 80.08 ;
    RECT 4.81 79.29 5.02 79.36 ;
    RECT 4.81 79.65 5.02 79.72 ;
    RECT 4.81 80.01 5.02 80.08 ;
    RECT 5.27 79.29 5.48 79.36 ;
    RECT 5.27 79.65 5.48 79.72 ;
    RECT 5.27 80.01 5.48 80.08 ;
    RECT 1.49 79.29 1.7 79.36 ;
    RECT 1.49 79.65 1.7 79.72 ;
    RECT 1.49 80.01 1.7 80.08 ;
    RECT 1.95 79.29 2.16 79.36 ;
    RECT 1.95 79.65 2.16 79.72 ;
    RECT 1.95 80.01 2.16 80.08 ;
    RECT 64.57 79.29 64.78 79.36 ;
    RECT 64.57 79.65 64.78 79.72 ;
    RECT 64.57 80.01 64.78 80.08 ;
    RECT 65.03 79.29 65.24 79.36 ;
    RECT 65.03 79.65 65.24 79.72 ;
    RECT 65.03 80.01 65.24 80.08 ;
    RECT 61.25 38.95 61.46 39.02 ;
    RECT 61.25 39.31 61.46 39.38 ;
    RECT 61.25 39.67 61.46 39.74 ;
    RECT 61.71 38.95 61.92 39.02 ;
    RECT 61.71 39.31 61.92 39.38 ;
    RECT 61.71 39.67 61.92 39.74 ;
    RECT 57.93 38.95 58.14 39.02 ;
    RECT 57.93 39.31 58.14 39.38 ;
    RECT 57.93 39.67 58.14 39.74 ;
    RECT 58.39 38.95 58.6 39.02 ;
    RECT 58.39 39.31 58.6 39.38 ;
    RECT 58.39 39.67 58.6 39.74 ;
    RECT 54.61 38.95 54.82 39.02 ;
    RECT 54.61 39.31 54.82 39.38 ;
    RECT 54.61 39.67 54.82 39.74 ;
    RECT 55.07 38.95 55.28 39.02 ;
    RECT 55.07 39.31 55.28 39.38 ;
    RECT 55.07 39.67 55.28 39.74 ;
    RECT 51.29 38.95 51.5 39.02 ;
    RECT 51.29 39.31 51.5 39.38 ;
    RECT 51.29 39.67 51.5 39.74 ;
    RECT 51.75 38.95 51.96 39.02 ;
    RECT 51.75 39.31 51.96 39.38 ;
    RECT 51.75 39.67 51.96 39.74 ;
    RECT 47.97 38.95 48.18 39.02 ;
    RECT 47.97 39.31 48.18 39.38 ;
    RECT 47.97 39.67 48.18 39.74 ;
    RECT 48.43 38.95 48.64 39.02 ;
    RECT 48.43 39.31 48.64 39.38 ;
    RECT 48.43 39.67 48.64 39.74 ;
    RECT 44.65 38.95 44.86 39.02 ;
    RECT 44.65 39.31 44.86 39.38 ;
    RECT 44.65 39.67 44.86 39.74 ;
    RECT 45.11 38.95 45.32 39.02 ;
    RECT 45.11 39.31 45.32 39.38 ;
    RECT 45.11 39.67 45.32 39.74 ;
    RECT 41.33 38.95 41.54 39.02 ;
    RECT 41.33 39.31 41.54 39.38 ;
    RECT 41.33 39.67 41.54 39.74 ;
    RECT 41.79 38.95 42.0 39.02 ;
    RECT 41.79 39.31 42.0 39.38 ;
    RECT 41.79 39.67 42.0 39.74 ;
    RECT 38.01 38.95 38.22 39.02 ;
    RECT 38.01 39.31 38.22 39.38 ;
    RECT 38.01 39.67 38.22 39.74 ;
    RECT 38.47 38.95 38.68 39.02 ;
    RECT 38.47 39.31 38.68 39.38 ;
    RECT 38.47 39.67 38.68 39.74 ;
    RECT 0.4 39.31 0.47 39.38 ;
    RECT 34.69 38.95 34.9 39.02 ;
    RECT 34.69 39.31 34.9 39.38 ;
    RECT 34.69 39.67 34.9 39.74 ;
    RECT 35.15 38.95 35.36 39.02 ;
    RECT 35.15 39.31 35.36 39.38 ;
    RECT 35.15 39.67 35.36 39.74 ;
    RECT 117.69 38.95 117.9 39.02 ;
    RECT 117.69 39.31 117.9 39.38 ;
    RECT 117.69 39.67 117.9 39.74 ;
    RECT 118.15 38.95 118.36 39.02 ;
    RECT 118.15 39.31 118.36 39.38 ;
    RECT 118.15 39.67 118.36 39.74 ;
    RECT 114.37 38.95 114.58 39.02 ;
    RECT 114.37 39.31 114.58 39.38 ;
    RECT 114.37 39.67 114.58 39.74 ;
    RECT 114.83 38.95 115.04 39.02 ;
    RECT 114.83 39.31 115.04 39.38 ;
    RECT 114.83 39.67 115.04 39.74 ;
    RECT 111.05 38.95 111.26 39.02 ;
    RECT 111.05 39.31 111.26 39.38 ;
    RECT 111.05 39.67 111.26 39.74 ;
    RECT 111.51 38.95 111.72 39.02 ;
    RECT 111.51 39.31 111.72 39.38 ;
    RECT 111.51 39.67 111.72 39.74 ;
    RECT 107.73 38.95 107.94 39.02 ;
    RECT 107.73 39.31 107.94 39.38 ;
    RECT 107.73 39.67 107.94 39.74 ;
    RECT 108.19 38.95 108.4 39.02 ;
    RECT 108.19 39.31 108.4 39.38 ;
    RECT 108.19 39.67 108.4 39.74 ;
    RECT 104.41 38.95 104.62 39.02 ;
    RECT 104.41 39.31 104.62 39.38 ;
    RECT 104.41 39.67 104.62 39.74 ;
    RECT 104.87 38.95 105.08 39.02 ;
    RECT 104.87 39.31 105.08 39.38 ;
    RECT 104.87 39.67 105.08 39.74 ;
    RECT 101.09 38.95 101.3 39.02 ;
    RECT 101.09 39.31 101.3 39.38 ;
    RECT 101.09 39.67 101.3 39.74 ;
    RECT 101.55 38.95 101.76 39.02 ;
    RECT 101.55 39.31 101.76 39.38 ;
    RECT 101.55 39.67 101.76 39.74 ;
    RECT 97.77 38.95 97.98 39.02 ;
    RECT 97.77 39.31 97.98 39.38 ;
    RECT 97.77 39.67 97.98 39.74 ;
    RECT 98.23 38.95 98.44 39.02 ;
    RECT 98.23 39.31 98.44 39.38 ;
    RECT 98.23 39.67 98.44 39.74 ;
    RECT 94.45 38.95 94.66 39.02 ;
    RECT 94.45 39.31 94.66 39.38 ;
    RECT 94.45 39.67 94.66 39.74 ;
    RECT 94.91 38.95 95.12 39.02 ;
    RECT 94.91 39.31 95.12 39.38 ;
    RECT 94.91 39.67 95.12 39.74 ;
    RECT 91.13 38.95 91.34 39.02 ;
    RECT 91.13 39.31 91.34 39.38 ;
    RECT 91.13 39.67 91.34 39.74 ;
    RECT 91.59 38.95 91.8 39.02 ;
    RECT 91.59 39.31 91.8 39.38 ;
    RECT 91.59 39.67 91.8 39.74 ;
    RECT 87.81 38.95 88.02 39.02 ;
    RECT 87.81 39.31 88.02 39.38 ;
    RECT 87.81 39.67 88.02 39.74 ;
    RECT 88.27 38.95 88.48 39.02 ;
    RECT 88.27 39.31 88.48 39.38 ;
    RECT 88.27 39.67 88.48 39.74 ;
    RECT 84.49 38.95 84.7 39.02 ;
    RECT 84.49 39.31 84.7 39.38 ;
    RECT 84.49 39.67 84.7 39.74 ;
    RECT 84.95 38.95 85.16 39.02 ;
    RECT 84.95 39.31 85.16 39.38 ;
    RECT 84.95 39.67 85.16 39.74 ;
    RECT 81.17 38.95 81.38 39.02 ;
    RECT 81.17 39.31 81.38 39.38 ;
    RECT 81.17 39.67 81.38 39.74 ;
    RECT 81.63 38.95 81.84 39.02 ;
    RECT 81.63 39.31 81.84 39.38 ;
    RECT 81.63 39.67 81.84 39.74 ;
    RECT 77.85 38.95 78.06 39.02 ;
    RECT 77.85 39.31 78.06 39.38 ;
    RECT 77.85 39.67 78.06 39.74 ;
    RECT 78.31 38.95 78.52 39.02 ;
    RECT 78.31 39.31 78.52 39.38 ;
    RECT 78.31 39.67 78.52 39.74 ;
    RECT 74.53 38.95 74.74 39.02 ;
    RECT 74.53 39.31 74.74 39.38 ;
    RECT 74.53 39.67 74.74 39.74 ;
    RECT 74.99 38.95 75.2 39.02 ;
    RECT 74.99 39.31 75.2 39.38 ;
    RECT 74.99 39.67 75.2 39.74 ;
    RECT 71.21 38.95 71.42 39.02 ;
    RECT 71.21 39.31 71.42 39.38 ;
    RECT 71.21 39.67 71.42 39.74 ;
    RECT 71.67 38.95 71.88 39.02 ;
    RECT 71.67 39.31 71.88 39.38 ;
    RECT 71.67 39.67 71.88 39.74 ;
    RECT 31.37 38.95 31.58 39.02 ;
    RECT 31.37 39.31 31.58 39.38 ;
    RECT 31.37 39.67 31.58 39.74 ;
    RECT 31.83 38.95 32.04 39.02 ;
    RECT 31.83 39.31 32.04 39.38 ;
    RECT 31.83 39.67 32.04 39.74 ;
    RECT 67.89 38.95 68.1 39.02 ;
    RECT 67.89 39.31 68.1 39.38 ;
    RECT 67.89 39.67 68.1 39.74 ;
    RECT 68.35 38.95 68.56 39.02 ;
    RECT 68.35 39.31 68.56 39.38 ;
    RECT 68.35 39.67 68.56 39.74 ;
    RECT 28.05 38.95 28.26 39.02 ;
    RECT 28.05 39.31 28.26 39.38 ;
    RECT 28.05 39.67 28.26 39.74 ;
    RECT 28.51 38.95 28.72 39.02 ;
    RECT 28.51 39.31 28.72 39.38 ;
    RECT 28.51 39.67 28.72 39.74 ;
    RECT 24.73 38.95 24.94 39.02 ;
    RECT 24.73 39.31 24.94 39.38 ;
    RECT 24.73 39.67 24.94 39.74 ;
    RECT 25.19 38.95 25.4 39.02 ;
    RECT 25.19 39.31 25.4 39.38 ;
    RECT 25.19 39.67 25.4 39.74 ;
    RECT 21.41 38.95 21.62 39.02 ;
    RECT 21.41 39.31 21.62 39.38 ;
    RECT 21.41 39.67 21.62 39.74 ;
    RECT 21.87 38.95 22.08 39.02 ;
    RECT 21.87 39.31 22.08 39.38 ;
    RECT 21.87 39.67 22.08 39.74 ;
    RECT 18.09 38.95 18.3 39.02 ;
    RECT 18.09 39.31 18.3 39.38 ;
    RECT 18.09 39.67 18.3 39.74 ;
    RECT 18.55 38.95 18.76 39.02 ;
    RECT 18.55 39.31 18.76 39.38 ;
    RECT 18.55 39.67 18.76 39.74 ;
    RECT 120.825 39.31 120.895 39.38 ;
    RECT 14.77 38.95 14.98 39.02 ;
    RECT 14.77 39.31 14.98 39.38 ;
    RECT 14.77 39.67 14.98 39.74 ;
    RECT 15.23 38.95 15.44 39.02 ;
    RECT 15.23 39.31 15.44 39.38 ;
    RECT 15.23 39.67 15.44 39.74 ;
    RECT 11.45 38.95 11.66 39.02 ;
    RECT 11.45 39.31 11.66 39.38 ;
    RECT 11.45 39.67 11.66 39.74 ;
    RECT 11.91 38.95 12.12 39.02 ;
    RECT 11.91 39.31 12.12 39.38 ;
    RECT 11.91 39.67 12.12 39.74 ;
    RECT 8.13 38.95 8.34 39.02 ;
    RECT 8.13 39.31 8.34 39.38 ;
    RECT 8.13 39.67 8.34 39.74 ;
    RECT 8.59 38.95 8.8 39.02 ;
    RECT 8.59 39.31 8.8 39.38 ;
    RECT 8.59 39.67 8.8 39.74 ;
    RECT 4.81 38.95 5.02 39.02 ;
    RECT 4.81 39.31 5.02 39.38 ;
    RECT 4.81 39.67 5.02 39.74 ;
    RECT 5.27 38.95 5.48 39.02 ;
    RECT 5.27 39.31 5.48 39.38 ;
    RECT 5.27 39.67 5.48 39.74 ;
    RECT 1.49 38.95 1.7 39.02 ;
    RECT 1.49 39.31 1.7 39.38 ;
    RECT 1.49 39.67 1.7 39.74 ;
    RECT 1.95 38.95 2.16 39.02 ;
    RECT 1.95 39.31 2.16 39.38 ;
    RECT 1.95 39.67 2.16 39.74 ;
    RECT 64.57 38.95 64.78 39.02 ;
    RECT 64.57 39.31 64.78 39.38 ;
    RECT 64.57 39.67 64.78 39.74 ;
    RECT 65.03 38.95 65.24 39.02 ;
    RECT 65.03 39.31 65.24 39.38 ;
    RECT 65.03 39.67 65.24 39.74 ;
    RECT 61.25 78.57 61.46 78.64 ;
    RECT 61.25 78.93 61.46 79.0 ;
    RECT 61.25 79.29 61.46 79.36 ;
    RECT 61.71 78.57 61.92 78.64 ;
    RECT 61.71 78.93 61.92 79.0 ;
    RECT 61.71 79.29 61.92 79.36 ;
    RECT 57.93 78.57 58.14 78.64 ;
    RECT 57.93 78.93 58.14 79.0 ;
    RECT 57.93 79.29 58.14 79.36 ;
    RECT 58.39 78.57 58.6 78.64 ;
    RECT 58.39 78.93 58.6 79.0 ;
    RECT 58.39 79.29 58.6 79.36 ;
    RECT 54.61 78.57 54.82 78.64 ;
    RECT 54.61 78.93 54.82 79.0 ;
    RECT 54.61 79.29 54.82 79.36 ;
    RECT 55.07 78.57 55.28 78.64 ;
    RECT 55.07 78.93 55.28 79.0 ;
    RECT 55.07 79.29 55.28 79.36 ;
    RECT 51.29 78.57 51.5 78.64 ;
    RECT 51.29 78.93 51.5 79.0 ;
    RECT 51.29 79.29 51.5 79.36 ;
    RECT 51.75 78.57 51.96 78.64 ;
    RECT 51.75 78.93 51.96 79.0 ;
    RECT 51.75 79.29 51.96 79.36 ;
    RECT 47.97 78.57 48.18 78.64 ;
    RECT 47.97 78.93 48.18 79.0 ;
    RECT 47.97 79.29 48.18 79.36 ;
    RECT 48.43 78.57 48.64 78.64 ;
    RECT 48.43 78.93 48.64 79.0 ;
    RECT 48.43 79.29 48.64 79.36 ;
    RECT 44.65 78.57 44.86 78.64 ;
    RECT 44.65 78.93 44.86 79.0 ;
    RECT 44.65 79.29 44.86 79.36 ;
    RECT 45.11 78.57 45.32 78.64 ;
    RECT 45.11 78.93 45.32 79.0 ;
    RECT 45.11 79.29 45.32 79.36 ;
    RECT 41.33 78.57 41.54 78.64 ;
    RECT 41.33 78.93 41.54 79.0 ;
    RECT 41.33 79.29 41.54 79.36 ;
    RECT 41.79 78.57 42.0 78.64 ;
    RECT 41.79 78.93 42.0 79.0 ;
    RECT 41.79 79.29 42.0 79.36 ;
    RECT 38.01 78.57 38.22 78.64 ;
    RECT 38.01 78.93 38.22 79.0 ;
    RECT 38.01 79.29 38.22 79.36 ;
    RECT 38.47 78.57 38.68 78.64 ;
    RECT 38.47 78.93 38.68 79.0 ;
    RECT 38.47 79.29 38.68 79.36 ;
    RECT 0.4 78.93 0.47 79.0 ;
    RECT 34.69 78.57 34.9 78.64 ;
    RECT 34.69 78.93 34.9 79.0 ;
    RECT 34.69 79.29 34.9 79.36 ;
    RECT 35.15 78.57 35.36 78.64 ;
    RECT 35.15 78.93 35.36 79.0 ;
    RECT 35.15 79.29 35.36 79.36 ;
    RECT 117.69 78.57 117.9 78.64 ;
    RECT 117.69 78.93 117.9 79.0 ;
    RECT 117.69 79.29 117.9 79.36 ;
    RECT 118.15 78.57 118.36 78.64 ;
    RECT 118.15 78.93 118.36 79.0 ;
    RECT 118.15 79.29 118.36 79.36 ;
    RECT 114.37 78.57 114.58 78.64 ;
    RECT 114.37 78.93 114.58 79.0 ;
    RECT 114.37 79.29 114.58 79.36 ;
    RECT 114.83 78.57 115.04 78.64 ;
    RECT 114.83 78.93 115.04 79.0 ;
    RECT 114.83 79.29 115.04 79.36 ;
    RECT 111.05 78.57 111.26 78.64 ;
    RECT 111.05 78.93 111.26 79.0 ;
    RECT 111.05 79.29 111.26 79.36 ;
    RECT 111.51 78.57 111.72 78.64 ;
    RECT 111.51 78.93 111.72 79.0 ;
    RECT 111.51 79.29 111.72 79.36 ;
    RECT 107.73 78.57 107.94 78.64 ;
    RECT 107.73 78.93 107.94 79.0 ;
    RECT 107.73 79.29 107.94 79.36 ;
    RECT 108.19 78.57 108.4 78.64 ;
    RECT 108.19 78.93 108.4 79.0 ;
    RECT 108.19 79.29 108.4 79.36 ;
    RECT 104.41 78.57 104.62 78.64 ;
    RECT 104.41 78.93 104.62 79.0 ;
    RECT 104.41 79.29 104.62 79.36 ;
    RECT 104.87 78.57 105.08 78.64 ;
    RECT 104.87 78.93 105.08 79.0 ;
    RECT 104.87 79.29 105.08 79.36 ;
    RECT 101.09 78.57 101.3 78.64 ;
    RECT 101.09 78.93 101.3 79.0 ;
    RECT 101.09 79.29 101.3 79.36 ;
    RECT 101.55 78.57 101.76 78.64 ;
    RECT 101.55 78.93 101.76 79.0 ;
    RECT 101.55 79.29 101.76 79.36 ;
    RECT 97.77 78.57 97.98 78.64 ;
    RECT 97.77 78.93 97.98 79.0 ;
    RECT 97.77 79.29 97.98 79.36 ;
    RECT 98.23 78.57 98.44 78.64 ;
    RECT 98.23 78.93 98.44 79.0 ;
    RECT 98.23 79.29 98.44 79.36 ;
    RECT 94.45 78.57 94.66 78.64 ;
    RECT 94.45 78.93 94.66 79.0 ;
    RECT 94.45 79.29 94.66 79.36 ;
    RECT 94.91 78.57 95.12 78.64 ;
    RECT 94.91 78.93 95.12 79.0 ;
    RECT 94.91 79.29 95.12 79.36 ;
    RECT 91.13 78.57 91.34 78.64 ;
    RECT 91.13 78.93 91.34 79.0 ;
    RECT 91.13 79.29 91.34 79.36 ;
    RECT 91.59 78.57 91.8 78.64 ;
    RECT 91.59 78.93 91.8 79.0 ;
    RECT 91.59 79.29 91.8 79.36 ;
    RECT 87.81 78.57 88.02 78.64 ;
    RECT 87.81 78.93 88.02 79.0 ;
    RECT 87.81 79.29 88.02 79.36 ;
    RECT 88.27 78.57 88.48 78.64 ;
    RECT 88.27 78.93 88.48 79.0 ;
    RECT 88.27 79.29 88.48 79.36 ;
    RECT 84.49 78.57 84.7 78.64 ;
    RECT 84.49 78.93 84.7 79.0 ;
    RECT 84.49 79.29 84.7 79.36 ;
    RECT 84.95 78.57 85.16 78.64 ;
    RECT 84.95 78.93 85.16 79.0 ;
    RECT 84.95 79.29 85.16 79.36 ;
    RECT 81.17 78.57 81.38 78.64 ;
    RECT 81.17 78.93 81.38 79.0 ;
    RECT 81.17 79.29 81.38 79.36 ;
    RECT 81.63 78.57 81.84 78.64 ;
    RECT 81.63 78.93 81.84 79.0 ;
    RECT 81.63 79.29 81.84 79.36 ;
    RECT 77.85 78.57 78.06 78.64 ;
    RECT 77.85 78.93 78.06 79.0 ;
    RECT 77.85 79.29 78.06 79.36 ;
    RECT 78.31 78.57 78.52 78.64 ;
    RECT 78.31 78.93 78.52 79.0 ;
    RECT 78.31 79.29 78.52 79.36 ;
    RECT 74.53 78.57 74.74 78.64 ;
    RECT 74.53 78.93 74.74 79.0 ;
    RECT 74.53 79.29 74.74 79.36 ;
    RECT 74.99 78.57 75.2 78.64 ;
    RECT 74.99 78.93 75.2 79.0 ;
    RECT 74.99 79.29 75.2 79.36 ;
    RECT 71.21 78.57 71.42 78.64 ;
    RECT 71.21 78.93 71.42 79.0 ;
    RECT 71.21 79.29 71.42 79.36 ;
    RECT 71.67 78.57 71.88 78.64 ;
    RECT 71.67 78.93 71.88 79.0 ;
    RECT 71.67 79.29 71.88 79.36 ;
    RECT 31.37 78.57 31.58 78.64 ;
    RECT 31.37 78.93 31.58 79.0 ;
    RECT 31.37 79.29 31.58 79.36 ;
    RECT 31.83 78.57 32.04 78.64 ;
    RECT 31.83 78.93 32.04 79.0 ;
    RECT 31.83 79.29 32.04 79.36 ;
    RECT 67.89 78.57 68.1 78.64 ;
    RECT 67.89 78.93 68.1 79.0 ;
    RECT 67.89 79.29 68.1 79.36 ;
    RECT 68.35 78.57 68.56 78.64 ;
    RECT 68.35 78.93 68.56 79.0 ;
    RECT 68.35 79.29 68.56 79.36 ;
    RECT 28.05 78.57 28.26 78.64 ;
    RECT 28.05 78.93 28.26 79.0 ;
    RECT 28.05 79.29 28.26 79.36 ;
    RECT 28.51 78.57 28.72 78.64 ;
    RECT 28.51 78.93 28.72 79.0 ;
    RECT 28.51 79.29 28.72 79.36 ;
    RECT 24.73 78.57 24.94 78.64 ;
    RECT 24.73 78.93 24.94 79.0 ;
    RECT 24.73 79.29 24.94 79.36 ;
    RECT 25.19 78.57 25.4 78.64 ;
    RECT 25.19 78.93 25.4 79.0 ;
    RECT 25.19 79.29 25.4 79.36 ;
    RECT 21.41 78.57 21.62 78.64 ;
    RECT 21.41 78.93 21.62 79.0 ;
    RECT 21.41 79.29 21.62 79.36 ;
    RECT 21.87 78.57 22.08 78.64 ;
    RECT 21.87 78.93 22.08 79.0 ;
    RECT 21.87 79.29 22.08 79.36 ;
    RECT 18.09 78.57 18.3 78.64 ;
    RECT 18.09 78.93 18.3 79.0 ;
    RECT 18.09 79.29 18.3 79.36 ;
    RECT 18.55 78.57 18.76 78.64 ;
    RECT 18.55 78.93 18.76 79.0 ;
    RECT 18.55 79.29 18.76 79.36 ;
    RECT 120.825 78.93 120.895 79.0 ;
    RECT 14.77 78.57 14.98 78.64 ;
    RECT 14.77 78.93 14.98 79.0 ;
    RECT 14.77 79.29 14.98 79.36 ;
    RECT 15.23 78.57 15.44 78.64 ;
    RECT 15.23 78.93 15.44 79.0 ;
    RECT 15.23 79.29 15.44 79.36 ;
    RECT 11.45 78.57 11.66 78.64 ;
    RECT 11.45 78.93 11.66 79.0 ;
    RECT 11.45 79.29 11.66 79.36 ;
    RECT 11.91 78.57 12.12 78.64 ;
    RECT 11.91 78.93 12.12 79.0 ;
    RECT 11.91 79.29 12.12 79.36 ;
    RECT 8.13 78.57 8.34 78.64 ;
    RECT 8.13 78.93 8.34 79.0 ;
    RECT 8.13 79.29 8.34 79.36 ;
    RECT 8.59 78.57 8.8 78.64 ;
    RECT 8.59 78.93 8.8 79.0 ;
    RECT 8.59 79.29 8.8 79.36 ;
    RECT 4.81 78.57 5.02 78.64 ;
    RECT 4.81 78.93 5.02 79.0 ;
    RECT 4.81 79.29 5.02 79.36 ;
    RECT 5.27 78.57 5.48 78.64 ;
    RECT 5.27 78.93 5.48 79.0 ;
    RECT 5.27 79.29 5.48 79.36 ;
    RECT 1.49 78.57 1.7 78.64 ;
    RECT 1.49 78.93 1.7 79.0 ;
    RECT 1.49 79.29 1.7 79.36 ;
    RECT 1.95 78.57 2.16 78.64 ;
    RECT 1.95 78.93 2.16 79.0 ;
    RECT 1.95 79.29 2.16 79.36 ;
    RECT 64.57 78.57 64.78 78.64 ;
    RECT 64.57 78.93 64.78 79.0 ;
    RECT 64.57 79.29 64.78 79.36 ;
    RECT 65.03 78.57 65.24 78.64 ;
    RECT 65.03 78.93 65.24 79.0 ;
    RECT 65.03 79.29 65.24 79.36 ;
    RECT 61.25 38.23 61.46 38.3 ;
    RECT 61.25 38.59 61.46 38.66 ;
    RECT 61.25 38.95 61.46 39.02 ;
    RECT 61.71 38.23 61.92 38.3 ;
    RECT 61.71 38.59 61.92 38.66 ;
    RECT 61.71 38.95 61.92 39.02 ;
    RECT 57.93 38.23 58.14 38.3 ;
    RECT 57.93 38.59 58.14 38.66 ;
    RECT 57.93 38.95 58.14 39.02 ;
    RECT 58.39 38.23 58.6 38.3 ;
    RECT 58.39 38.59 58.6 38.66 ;
    RECT 58.39 38.95 58.6 39.02 ;
    RECT 54.61 38.23 54.82 38.3 ;
    RECT 54.61 38.59 54.82 38.66 ;
    RECT 54.61 38.95 54.82 39.02 ;
    RECT 55.07 38.23 55.28 38.3 ;
    RECT 55.07 38.59 55.28 38.66 ;
    RECT 55.07 38.95 55.28 39.02 ;
    RECT 51.29 38.23 51.5 38.3 ;
    RECT 51.29 38.59 51.5 38.66 ;
    RECT 51.29 38.95 51.5 39.02 ;
    RECT 51.75 38.23 51.96 38.3 ;
    RECT 51.75 38.59 51.96 38.66 ;
    RECT 51.75 38.95 51.96 39.02 ;
    RECT 47.97 38.23 48.18 38.3 ;
    RECT 47.97 38.59 48.18 38.66 ;
    RECT 47.97 38.95 48.18 39.02 ;
    RECT 48.43 38.23 48.64 38.3 ;
    RECT 48.43 38.59 48.64 38.66 ;
    RECT 48.43 38.95 48.64 39.02 ;
    RECT 44.65 38.23 44.86 38.3 ;
    RECT 44.65 38.59 44.86 38.66 ;
    RECT 44.65 38.95 44.86 39.02 ;
    RECT 45.11 38.23 45.32 38.3 ;
    RECT 45.11 38.59 45.32 38.66 ;
    RECT 45.11 38.95 45.32 39.02 ;
    RECT 41.33 38.23 41.54 38.3 ;
    RECT 41.33 38.59 41.54 38.66 ;
    RECT 41.33 38.95 41.54 39.02 ;
    RECT 41.79 38.23 42.0 38.3 ;
    RECT 41.79 38.59 42.0 38.66 ;
    RECT 41.79 38.95 42.0 39.02 ;
    RECT 38.01 38.23 38.22 38.3 ;
    RECT 38.01 38.59 38.22 38.66 ;
    RECT 38.01 38.95 38.22 39.02 ;
    RECT 38.47 38.23 38.68 38.3 ;
    RECT 38.47 38.59 38.68 38.66 ;
    RECT 38.47 38.95 38.68 39.02 ;
    RECT 0.4 38.59 0.47 38.66 ;
    RECT 34.69 38.23 34.9 38.3 ;
    RECT 34.69 38.59 34.9 38.66 ;
    RECT 34.69 38.95 34.9 39.02 ;
    RECT 35.15 38.23 35.36 38.3 ;
    RECT 35.15 38.59 35.36 38.66 ;
    RECT 35.15 38.95 35.36 39.02 ;
    RECT 117.69 38.23 117.9 38.3 ;
    RECT 117.69 38.59 117.9 38.66 ;
    RECT 117.69 38.95 117.9 39.02 ;
    RECT 118.15 38.23 118.36 38.3 ;
    RECT 118.15 38.59 118.36 38.66 ;
    RECT 118.15 38.95 118.36 39.02 ;
    RECT 114.37 38.23 114.58 38.3 ;
    RECT 114.37 38.59 114.58 38.66 ;
    RECT 114.37 38.95 114.58 39.02 ;
    RECT 114.83 38.23 115.04 38.3 ;
    RECT 114.83 38.59 115.04 38.66 ;
    RECT 114.83 38.95 115.04 39.02 ;
    RECT 111.05 38.23 111.26 38.3 ;
    RECT 111.05 38.59 111.26 38.66 ;
    RECT 111.05 38.95 111.26 39.02 ;
    RECT 111.51 38.23 111.72 38.3 ;
    RECT 111.51 38.59 111.72 38.66 ;
    RECT 111.51 38.95 111.72 39.02 ;
    RECT 107.73 38.23 107.94 38.3 ;
    RECT 107.73 38.59 107.94 38.66 ;
    RECT 107.73 38.95 107.94 39.02 ;
    RECT 108.19 38.23 108.4 38.3 ;
    RECT 108.19 38.59 108.4 38.66 ;
    RECT 108.19 38.95 108.4 39.02 ;
    RECT 104.41 38.23 104.62 38.3 ;
    RECT 104.41 38.59 104.62 38.66 ;
    RECT 104.41 38.95 104.62 39.02 ;
    RECT 104.87 38.23 105.08 38.3 ;
    RECT 104.87 38.59 105.08 38.66 ;
    RECT 104.87 38.95 105.08 39.02 ;
    RECT 101.09 38.23 101.3 38.3 ;
    RECT 101.09 38.59 101.3 38.66 ;
    RECT 101.09 38.95 101.3 39.02 ;
    RECT 101.55 38.23 101.76 38.3 ;
    RECT 101.55 38.59 101.76 38.66 ;
    RECT 101.55 38.95 101.76 39.02 ;
    RECT 97.77 38.23 97.98 38.3 ;
    RECT 97.77 38.59 97.98 38.66 ;
    RECT 97.77 38.95 97.98 39.02 ;
    RECT 98.23 38.23 98.44 38.3 ;
    RECT 98.23 38.59 98.44 38.66 ;
    RECT 98.23 38.95 98.44 39.02 ;
    RECT 94.45 38.23 94.66 38.3 ;
    RECT 94.45 38.59 94.66 38.66 ;
    RECT 94.45 38.95 94.66 39.02 ;
    RECT 94.91 38.23 95.12 38.3 ;
    RECT 94.91 38.59 95.12 38.66 ;
    RECT 94.91 38.95 95.12 39.02 ;
    RECT 91.13 38.23 91.34 38.3 ;
    RECT 91.13 38.59 91.34 38.66 ;
    RECT 91.13 38.95 91.34 39.02 ;
    RECT 91.59 38.23 91.8 38.3 ;
    RECT 91.59 38.59 91.8 38.66 ;
    RECT 91.59 38.95 91.8 39.02 ;
    RECT 87.81 38.23 88.02 38.3 ;
    RECT 87.81 38.59 88.02 38.66 ;
    RECT 87.81 38.95 88.02 39.02 ;
    RECT 88.27 38.23 88.48 38.3 ;
    RECT 88.27 38.59 88.48 38.66 ;
    RECT 88.27 38.95 88.48 39.02 ;
    RECT 84.49 38.23 84.7 38.3 ;
    RECT 84.49 38.59 84.7 38.66 ;
    RECT 84.49 38.95 84.7 39.02 ;
    RECT 84.95 38.23 85.16 38.3 ;
    RECT 84.95 38.59 85.16 38.66 ;
    RECT 84.95 38.95 85.16 39.02 ;
    RECT 81.17 38.23 81.38 38.3 ;
    RECT 81.17 38.59 81.38 38.66 ;
    RECT 81.17 38.95 81.38 39.02 ;
    RECT 81.63 38.23 81.84 38.3 ;
    RECT 81.63 38.59 81.84 38.66 ;
    RECT 81.63 38.95 81.84 39.02 ;
    RECT 77.85 38.23 78.06 38.3 ;
    RECT 77.85 38.59 78.06 38.66 ;
    RECT 77.85 38.95 78.06 39.02 ;
    RECT 78.31 38.23 78.52 38.3 ;
    RECT 78.31 38.59 78.52 38.66 ;
    RECT 78.31 38.95 78.52 39.02 ;
    RECT 74.53 38.23 74.74 38.3 ;
    RECT 74.53 38.59 74.74 38.66 ;
    RECT 74.53 38.95 74.74 39.02 ;
    RECT 74.99 38.23 75.2 38.3 ;
    RECT 74.99 38.59 75.2 38.66 ;
    RECT 74.99 38.95 75.2 39.02 ;
    RECT 71.21 38.23 71.42 38.3 ;
    RECT 71.21 38.59 71.42 38.66 ;
    RECT 71.21 38.95 71.42 39.02 ;
    RECT 71.67 38.23 71.88 38.3 ;
    RECT 71.67 38.59 71.88 38.66 ;
    RECT 71.67 38.95 71.88 39.02 ;
    RECT 31.37 38.23 31.58 38.3 ;
    RECT 31.37 38.59 31.58 38.66 ;
    RECT 31.37 38.95 31.58 39.02 ;
    RECT 31.83 38.23 32.04 38.3 ;
    RECT 31.83 38.59 32.04 38.66 ;
    RECT 31.83 38.95 32.04 39.02 ;
    RECT 67.89 38.23 68.1 38.3 ;
    RECT 67.89 38.59 68.1 38.66 ;
    RECT 67.89 38.95 68.1 39.02 ;
    RECT 68.35 38.23 68.56 38.3 ;
    RECT 68.35 38.59 68.56 38.66 ;
    RECT 68.35 38.95 68.56 39.02 ;
    RECT 28.05 38.23 28.26 38.3 ;
    RECT 28.05 38.59 28.26 38.66 ;
    RECT 28.05 38.95 28.26 39.02 ;
    RECT 28.51 38.23 28.72 38.3 ;
    RECT 28.51 38.59 28.72 38.66 ;
    RECT 28.51 38.95 28.72 39.02 ;
    RECT 24.73 38.23 24.94 38.3 ;
    RECT 24.73 38.59 24.94 38.66 ;
    RECT 24.73 38.95 24.94 39.02 ;
    RECT 25.19 38.23 25.4 38.3 ;
    RECT 25.19 38.59 25.4 38.66 ;
    RECT 25.19 38.95 25.4 39.02 ;
    RECT 21.41 38.23 21.62 38.3 ;
    RECT 21.41 38.59 21.62 38.66 ;
    RECT 21.41 38.95 21.62 39.02 ;
    RECT 21.87 38.23 22.08 38.3 ;
    RECT 21.87 38.59 22.08 38.66 ;
    RECT 21.87 38.95 22.08 39.02 ;
    RECT 18.09 38.23 18.3 38.3 ;
    RECT 18.09 38.59 18.3 38.66 ;
    RECT 18.09 38.95 18.3 39.02 ;
    RECT 18.55 38.23 18.76 38.3 ;
    RECT 18.55 38.59 18.76 38.66 ;
    RECT 18.55 38.95 18.76 39.02 ;
    RECT 120.825 38.59 120.895 38.66 ;
    RECT 14.77 38.23 14.98 38.3 ;
    RECT 14.77 38.59 14.98 38.66 ;
    RECT 14.77 38.95 14.98 39.02 ;
    RECT 15.23 38.23 15.44 38.3 ;
    RECT 15.23 38.59 15.44 38.66 ;
    RECT 15.23 38.95 15.44 39.02 ;
    RECT 11.45 38.23 11.66 38.3 ;
    RECT 11.45 38.59 11.66 38.66 ;
    RECT 11.45 38.95 11.66 39.02 ;
    RECT 11.91 38.23 12.12 38.3 ;
    RECT 11.91 38.59 12.12 38.66 ;
    RECT 11.91 38.95 12.12 39.02 ;
    RECT 8.13 38.23 8.34 38.3 ;
    RECT 8.13 38.59 8.34 38.66 ;
    RECT 8.13 38.95 8.34 39.02 ;
    RECT 8.59 38.23 8.8 38.3 ;
    RECT 8.59 38.59 8.8 38.66 ;
    RECT 8.59 38.95 8.8 39.02 ;
    RECT 4.81 38.23 5.02 38.3 ;
    RECT 4.81 38.59 5.02 38.66 ;
    RECT 4.81 38.95 5.02 39.02 ;
    RECT 5.27 38.23 5.48 38.3 ;
    RECT 5.27 38.59 5.48 38.66 ;
    RECT 5.27 38.95 5.48 39.02 ;
    RECT 1.49 38.23 1.7 38.3 ;
    RECT 1.49 38.59 1.7 38.66 ;
    RECT 1.49 38.95 1.7 39.02 ;
    RECT 1.95 38.23 2.16 38.3 ;
    RECT 1.95 38.59 2.16 38.66 ;
    RECT 1.95 38.95 2.16 39.02 ;
    RECT 64.57 38.23 64.78 38.3 ;
    RECT 64.57 38.59 64.78 38.66 ;
    RECT 64.57 38.95 64.78 39.02 ;
    RECT 65.03 38.23 65.24 38.3 ;
    RECT 65.03 38.59 65.24 38.66 ;
    RECT 65.03 38.95 65.24 39.02 ;
    RECT 61.25 77.85 61.46 77.92 ;
    RECT 61.25 78.21 61.46 78.28 ;
    RECT 61.25 78.57 61.46 78.64 ;
    RECT 61.71 77.85 61.92 77.92 ;
    RECT 61.71 78.21 61.92 78.28 ;
    RECT 61.71 78.57 61.92 78.64 ;
    RECT 57.93 77.85 58.14 77.92 ;
    RECT 57.93 78.21 58.14 78.28 ;
    RECT 57.93 78.57 58.14 78.64 ;
    RECT 58.39 77.85 58.6 77.92 ;
    RECT 58.39 78.21 58.6 78.28 ;
    RECT 58.39 78.57 58.6 78.64 ;
    RECT 54.61 77.85 54.82 77.92 ;
    RECT 54.61 78.21 54.82 78.28 ;
    RECT 54.61 78.57 54.82 78.64 ;
    RECT 55.07 77.85 55.28 77.92 ;
    RECT 55.07 78.21 55.28 78.28 ;
    RECT 55.07 78.57 55.28 78.64 ;
    RECT 51.29 77.85 51.5 77.92 ;
    RECT 51.29 78.21 51.5 78.28 ;
    RECT 51.29 78.57 51.5 78.64 ;
    RECT 51.75 77.85 51.96 77.92 ;
    RECT 51.75 78.21 51.96 78.28 ;
    RECT 51.75 78.57 51.96 78.64 ;
    RECT 47.97 77.85 48.18 77.92 ;
    RECT 47.97 78.21 48.18 78.28 ;
    RECT 47.97 78.57 48.18 78.64 ;
    RECT 48.43 77.85 48.64 77.92 ;
    RECT 48.43 78.21 48.64 78.28 ;
    RECT 48.43 78.57 48.64 78.64 ;
    RECT 44.65 77.85 44.86 77.92 ;
    RECT 44.65 78.21 44.86 78.28 ;
    RECT 44.65 78.57 44.86 78.64 ;
    RECT 45.11 77.85 45.32 77.92 ;
    RECT 45.11 78.21 45.32 78.28 ;
    RECT 45.11 78.57 45.32 78.64 ;
    RECT 41.33 77.85 41.54 77.92 ;
    RECT 41.33 78.21 41.54 78.28 ;
    RECT 41.33 78.57 41.54 78.64 ;
    RECT 41.79 77.85 42.0 77.92 ;
    RECT 41.79 78.21 42.0 78.28 ;
    RECT 41.79 78.57 42.0 78.64 ;
    RECT 38.01 77.85 38.22 77.92 ;
    RECT 38.01 78.21 38.22 78.28 ;
    RECT 38.01 78.57 38.22 78.64 ;
    RECT 38.47 77.85 38.68 77.92 ;
    RECT 38.47 78.21 38.68 78.28 ;
    RECT 38.47 78.57 38.68 78.64 ;
    RECT 0.4 78.21 0.47 78.28 ;
    RECT 34.69 77.85 34.9 77.92 ;
    RECT 34.69 78.21 34.9 78.28 ;
    RECT 34.69 78.57 34.9 78.64 ;
    RECT 35.15 77.85 35.36 77.92 ;
    RECT 35.15 78.21 35.36 78.28 ;
    RECT 35.15 78.57 35.36 78.64 ;
    RECT 117.69 77.85 117.9 77.92 ;
    RECT 117.69 78.21 117.9 78.28 ;
    RECT 117.69 78.57 117.9 78.64 ;
    RECT 118.15 77.85 118.36 77.92 ;
    RECT 118.15 78.21 118.36 78.28 ;
    RECT 118.15 78.57 118.36 78.64 ;
    RECT 114.37 77.85 114.58 77.92 ;
    RECT 114.37 78.21 114.58 78.28 ;
    RECT 114.37 78.57 114.58 78.64 ;
    RECT 114.83 77.85 115.04 77.92 ;
    RECT 114.83 78.21 115.04 78.28 ;
    RECT 114.83 78.57 115.04 78.64 ;
    RECT 111.05 77.85 111.26 77.92 ;
    RECT 111.05 78.21 111.26 78.28 ;
    RECT 111.05 78.57 111.26 78.64 ;
    RECT 111.51 77.85 111.72 77.92 ;
    RECT 111.51 78.21 111.72 78.28 ;
    RECT 111.51 78.57 111.72 78.64 ;
    RECT 107.73 77.85 107.94 77.92 ;
    RECT 107.73 78.21 107.94 78.28 ;
    RECT 107.73 78.57 107.94 78.64 ;
    RECT 108.19 77.85 108.4 77.92 ;
    RECT 108.19 78.21 108.4 78.28 ;
    RECT 108.19 78.57 108.4 78.64 ;
    RECT 104.41 77.85 104.62 77.92 ;
    RECT 104.41 78.21 104.62 78.28 ;
    RECT 104.41 78.57 104.62 78.64 ;
    RECT 104.87 77.85 105.08 77.92 ;
    RECT 104.87 78.21 105.08 78.28 ;
    RECT 104.87 78.57 105.08 78.64 ;
    RECT 101.09 77.85 101.3 77.92 ;
    RECT 101.09 78.21 101.3 78.28 ;
    RECT 101.09 78.57 101.3 78.64 ;
    RECT 101.55 77.85 101.76 77.92 ;
    RECT 101.55 78.21 101.76 78.28 ;
    RECT 101.55 78.57 101.76 78.64 ;
    RECT 97.77 77.85 97.98 77.92 ;
    RECT 97.77 78.21 97.98 78.28 ;
    RECT 97.77 78.57 97.98 78.64 ;
    RECT 98.23 77.85 98.44 77.92 ;
    RECT 98.23 78.21 98.44 78.28 ;
    RECT 98.23 78.57 98.44 78.64 ;
    RECT 94.45 77.85 94.66 77.92 ;
    RECT 94.45 78.21 94.66 78.28 ;
    RECT 94.45 78.57 94.66 78.64 ;
    RECT 94.91 77.85 95.12 77.92 ;
    RECT 94.91 78.21 95.12 78.28 ;
    RECT 94.91 78.57 95.12 78.64 ;
    RECT 91.13 77.85 91.34 77.92 ;
    RECT 91.13 78.21 91.34 78.28 ;
    RECT 91.13 78.57 91.34 78.64 ;
    RECT 91.59 77.85 91.8 77.92 ;
    RECT 91.59 78.21 91.8 78.28 ;
    RECT 91.59 78.57 91.8 78.64 ;
    RECT 87.81 77.85 88.02 77.92 ;
    RECT 87.81 78.21 88.02 78.28 ;
    RECT 87.81 78.57 88.02 78.64 ;
    RECT 88.27 77.85 88.48 77.92 ;
    RECT 88.27 78.21 88.48 78.28 ;
    RECT 88.27 78.57 88.48 78.64 ;
    RECT 84.49 77.85 84.7 77.92 ;
    RECT 84.49 78.21 84.7 78.28 ;
    RECT 84.49 78.57 84.7 78.64 ;
    RECT 84.95 77.85 85.16 77.92 ;
    RECT 84.95 78.21 85.16 78.28 ;
    RECT 84.95 78.57 85.16 78.64 ;
    RECT 81.17 77.85 81.38 77.92 ;
    RECT 81.17 78.21 81.38 78.28 ;
    RECT 81.17 78.57 81.38 78.64 ;
    RECT 81.63 77.85 81.84 77.92 ;
    RECT 81.63 78.21 81.84 78.28 ;
    RECT 81.63 78.57 81.84 78.64 ;
    RECT 77.85 77.85 78.06 77.92 ;
    RECT 77.85 78.21 78.06 78.28 ;
    RECT 77.85 78.57 78.06 78.64 ;
    RECT 78.31 77.85 78.52 77.92 ;
    RECT 78.31 78.21 78.52 78.28 ;
    RECT 78.31 78.57 78.52 78.64 ;
    RECT 74.53 77.85 74.74 77.92 ;
    RECT 74.53 78.21 74.74 78.28 ;
    RECT 74.53 78.57 74.74 78.64 ;
    RECT 74.99 77.85 75.2 77.92 ;
    RECT 74.99 78.21 75.2 78.28 ;
    RECT 74.99 78.57 75.2 78.64 ;
    RECT 71.21 77.85 71.42 77.92 ;
    RECT 71.21 78.21 71.42 78.28 ;
    RECT 71.21 78.57 71.42 78.64 ;
    RECT 71.67 77.85 71.88 77.92 ;
    RECT 71.67 78.21 71.88 78.28 ;
    RECT 71.67 78.57 71.88 78.64 ;
    RECT 31.37 77.85 31.58 77.92 ;
    RECT 31.37 78.21 31.58 78.28 ;
    RECT 31.37 78.57 31.58 78.64 ;
    RECT 31.83 77.85 32.04 77.92 ;
    RECT 31.83 78.21 32.04 78.28 ;
    RECT 31.83 78.57 32.04 78.64 ;
    RECT 67.89 77.85 68.1 77.92 ;
    RECT 67.89 78.21 68.1 78.28 ;
    RECT 67.89 78.57 68.1 78.64 ;
    RECT 68.35 77.85 68.56 77.92 ;
    RECT 68.35 78.21 68.56 78.28 ;
    RECT 68.35 78.57 68.56 78.64 ;
    RECT 28.05 77.85 28.26 77.92 ;
    RECT 28.05 78.21 28.26 78.28 ;
    RECT 28.05 78.57 28.26 78.64 ;
    RECT 28.51 77.85 28.72 77.92 ;
    RECT 28.51 78.21 28.72 78.28 ;
    RECT 28.51 78.57 28.72 78.64 ;
    RECT 24.73 77.85 24.94 77.92 ;
    RECT 24.73 78.21 24.94 78.28 ;
    RECT 24.73 78.57 24.94 78.64 ;
    RECT 25.19 77.85 25.4 77.92 ;
    RECT 25.19 78.21 25.4 78.28 ;
    RECT 25.19 78.57 25.4 78.64 ;
    RECT 21.41 77.85 21.62 77.92 ;
    RECT 21.41 78.21 21.62 78.28 ;
    RECT 21.41 78.57 21.62 78.64 ;
    RECT 21.87 77.85 22.08 77.92 ;
    RECT 21.87 78.21 22.08 78.28 ;
    RECT 21.87 78.57 22.08 78.64 ;
    RECT 18.09 77.85 18.3 77.92 ;
    RECT 18.09 78.21 18.3 78.28 ;
    RECT 18.09 78.57 18.3 78.64 ;
    RECT 18.55 77.85 18.76 77.92 ;
    RECT 18.55 78.21 18.76 78.28 ;
    RECT 18.55 78.57 18.76 78.64 ;
    RECT 120.825 78.21 120.895 78.28 ;
    RECT 14.77 77.85 14.98 77.92 ;
    RECT 14.77 78.21 14.98 78.28 ;
    RECT 14.77 78.57 14.98 78.64 ;
    RECT 15.23 77.85 15.44 77.92 ;
    RECT 15.23 78.21 15.44 78.28 ;
    RECT 15.23 78.57 15.44 78.64 ;
    RECT 11.45 77.85 11.66 77.92 ;
    RECT 11.45 78.21 11.66 78.28 ;
    RECT 11.45 78.57 11.66 78.64 ;
    RECT 11.91 77.85 12.12 77.92 ;
    RECT 11.91 78.21 12.12 78.28 ;
    RECT 11.91 78.57 12.12 78.64 ;
    RECT 8.13 77.85 8.34 77.92 ;
    RECT 8.13 78.21 8.34 78.28 ;
    RECT 8.13 78.57 8.34 78.64 ;
    RECT 8.59 77.85 8.8 77.92 ;
    RECT 8.59 78.21 8.8 78.28 ;
    RECT 8.59 78.57 8.8 78.64 ;
    RECT 4.81 77.85 5.02 77.92 ;
    RECT 4.81 78.21 5.02 78.28 ;
    RECT 4.81 78.57 5.02 78.64 ;
    RECT 5.27 77.85 5.48 77.92 ;
    RECT 5.27 78.21 5.48 78.28 ;
    RECT 5.27 78.57 5.48 78.64 ;
    RECT 1.49 77.85 1.7 77.92 ;
    RECT 1.49 78.21 1.7 78.28 ;
    RECT 1.49 78.57 1.7 78.64 ;
    RECT 1.95 77.85 2.16 77.92 ;
    RECT 1.95 78.21 2.16 78.28 ;
    RECT 1.95 78.57 2.16 78.64 ;
    RECT 64.57 77.85 64.78 77.92 ;
    RECT 64.57 78.21 64.78 78.28 ;
    RECT 64.57 78.57 64.78 78.64 ;
    RECT 65.03 77.85 65.24 77.92 ;
    RECT 65.03 78.21 65.24 78.28 ;
    RECT 65.03 78.57 65.24 78.64 ;
    RECT 61.25 37.51 61.46 37.58 ;
    RECT 61.25 37.87 61.46 37.94 ;
    RECT 61.25 38.23 61.46 38.3 ;
    RECT 61.71 37.51 61.92 37.58 ;
    RECT 61.71 37.87 61.92 37.94 ;
    RECT 61.71 38.23 61.92 38.3 ;
    RECT 57.93 37.51 58.14 37.58 ;
    RECT 57.93 37.87 58.14 37.94 ;
    RECT 57.93 38.23 58.14 38.3 ;
    RECT 58.39 37.51 58.6 37.58 ;
    RECT 58.39 37.87 58.6 37.94 ;
    RECT 58.39 38.23 58.6 38.3 ;
    RECT 54.61 37.51 54.82 37.58 ;
    RECT 54.61 37.87 54.82 37.94 ;
    RECT 54.61 38.23 54.82 38.3 ;
    RECT 55.07 37.51 55.28 37.58 ;
    RECT 55.07 37.87 55.28 37.94 ;
    RECT 55.07 38.23 55.28 38.3 ;
    RECT 51.29 37.51 51.5 37.58 ;
    RECT 51.29 37.87 51.5 37.94 ;
    RECT 51.29 38.23 51.5 38.3 ;
    RECT 51.75 37.51 51.96 37.58 ;
    RECT 51.75 37.87 51.96 37.94 ;
    RECT 51.75 38.23 51.96 38.3 ;
    RECT 47.97 37.51 48.18 37.58 ;
    RECT 47.97 37.87 48.18 37.94 ;
    RECT 47.97 38.23 48.18 38.3 ;
    RECT 48.43 37.51 48.64 37.58 ;
    RECT 48.43 37.87 48.64 37.94 ;
    RECT 48.43 38.23 48.64 38.3 ;
    RECT 44.65 37.51 44.86 37.58 ;
    RECT 44.65 37.87 44.86 37.94 ;
    RECT 44.65 38.23 44.86 38.3 ;
    RECT 45.11 37.51 45.32 37.58 ;
    RECT 45.11 37.87 45.32 37.94 ;
    RECT 45.11 38.23 45.32 38.3 ;
    RECT 41.33 37.51 41.54 37.58 ;
    RECT 41.33 37.87 41.54 37.94 ;
    RECT 41.33 38.23 41.54 38.3 ;
    RECT 41.79 37.51 42.0 37.58 ;
    RECT 41.79 37.87 42.0 37.94 ;
    RECT 41.79 38.23 42.0 38.3 ;
    RECT 38.01 37.51 38.22 37.58 ;
    RECT 38.01 37.87 38.22 37.94 ;
    RECT 38.01 38.23 38.22 38.3 ;
    RECT 38.47 37.51 38.68 37.58 ;
    RECT 38.47 37.87 38.68 37.94 ;
    RECT 38.47 38.23 38.68 38.3 ;
    RECT 0.4 37.87 0.47 37.94 ;
    RECT 34.69 37.51 34.9 37.58 ;
    RECT 34.69 37.87 34.9 37.94 ;
    RECT 34.69 38.23 34.9 38.3 ;
    RECT 35.15 37.51 35.36 37.58 ;
    RECT 35.15 37.87 35.36 37.94 ;
    RECT 35.15 38.23 35.36 38.3 ;
    RECT 117.69 37.51 117.9 37.58 ;
    RECT 117.69 37.87 117.9 37.94 ;
    RECT 117.69 38.23 117.9 38.3 ;
    RECT 118.15 37.51 118.36 37.58 ;
    RECT 118.15 37.87 118.36 37.94 ;
    RECT 118.15 38.23 118.36 38.3 ;
    RECT 114.37 37.51 114.58 37.58 ;
    RECT 114.37 37.87 114.58 37.94 ;
    RECT 114.37 38.23 114.58 38.3 ;
    RECT 114.83 37.51 115.04 37.58 ;
    RECT 114.83 37.87 115.04 37.94 ;
    RECT 114.83 38.23 115.04 38.3 ;
    RECT 111.05 37.51 111.26 37.58 ;
    RECT 111.05 37.87 111.26 37.94 ;
    RECT 111.05 38.23 111.26 38.3 ;
    RECT 111.51 37.51 111.72 37.58 ;
    RECT 111.51 37.87 111.72 37.94 ;
    RECT 111.51 38.23 111.72 38.3 ;
    RECT 107.73 37.51 107.94 37.58 ;
    RECT 107.73 37.87 107.94 37.94 ;
    RECT 107.73 38.23 107.94 38.3 ;
    RECT 108.19 37.51 108.4 37.58 ;
    RECT 108.19 37.87 108.4 37.94 ;
    RECT 108.19 38.23 108.4 38.3 ;
    RECT 104.41 37.51 104.62 37.58 ;
    RECT 104.41 37.87 104.62 37.94 ;
    RECT 104.41 38.23 104.62 38.3 ;
    RECT 104.87 37.51 105.08 37.58 ;
    RECT 104.87 37.87 105.08 37.94 ;
    RECT 104.87 38.23 105.08 38.3 ;
    RECT 101.09 37.51 101.3 37.58 ;
    RECT 101.09 37.87 101.3 37.94 ;
    RECT 101.09 38.23 101.3 38.3 ;
    RECT 101.55 37.51 101.76 37.58 ;
    RECT 101.55 37.87 101.76 37.94 ;
    RECT 101.55 38.23 101.76 38.3 ;
    RECT 97.77 37.51 97.98 37.58 ;
    RECT 97.77 37.87 97.98 37.94 ;
    RECT 97.77 38.23 97.98 38.3 ;
    RECT 98.23 37.51 98.44 37.58 ;
    RECT 98.23 37.87 98.44 37.94 ;
    RECT 98.23 38.23 98.44 38.3 ;
    RECT 94.45 37.51 94.66 37.58 ;
    RECT 94.45 37.87 94.66 37.94 ;
    RECT 94.45 38.23 94.66 38.3 ;
    RECT 94.91 37.51 95.12 37.58 ;
    RECT 94.91 37.87 95.12 37.94 ;
    RECT 94.91 38.23 95.12 38.3 ;
    RECT 91.13 37.51 91.34 37.58 ;
    RECT 91.13 37.87 91.34 37.94 ;
    RECT 91.13 38.23 91.34 38.3 ;
    RECT 91.59 37.51 91.8 37.58 ;
    RECT 91.59 37.87 91.8 37.94 ;
    RECT 91.59 38.23 91.8 38.3 ;
    RECT 87.81 37.51 88.02 37.58 ;
    RECT 87.81 37.87 88.02 37.94 ;
    RECT 87.81 38.23 88.02 38.3 ;
    RECT 88.27 37.51 88.48 37.58 ;
    RECT 88.27 37.87 88.48 37.94 ;
    RECT 88.27 38.23 88.48 38.3 ;
    RECT 84.49 37.51 84.7 37.58 ;
    RECT 84.49 37.87 84.7 37.94 ;
    RECT 84.49 38.23 84.7 38.3 ;
    RECT 84.95 37.51 85.16 37.58 ;
    RECT 84.95 37.87 85.16 37.94 ;
    RECT 84.95 38.23 85.16 38.3 ;
    RECT 81.17 37.51 81.38 37.58 ;
    RECT 81.17 37.87 81.38 37.94 ;
    RECT 81.17 38.23 81.38 38.3 ;
    RECT 81.63 37.51 81.84 37.58 ;
    RECT 81.63 37.87 81.84 37.94 ;
    RECT 81.63 38.23 81.84 38.3 ;
    RECT 77.85 37.51 78.06 37.58 ;
    RECT 77.85 37.87 78.06 37.94 ;
    RECT 77.85 38.23 78.06 38.3 ;
    RECT 78.31 37.51 78.52 37.58 ;
    RECT 78.31 37.87 78.52 37.94 ;
    RECT 78.31 38.23 78.52 38.3 ;
    RECT 74.53 37.51 74.74 37.58 ;
    RECT 74.53 37.87 74.74 37.94 ;
    RECT 74.53 38.23 74.74 38.3 ;
    RECT 74.99 37.51 75.2 37.58 ;
    RECT 74.99 37.87 75.2 37.94 ;
    RECT 74.99 38.23 75.2 38.3 ;
    RECT 71.21 37.51 71.42 37.58 ;
    RECT 71.21 37.87 71.42 37.94 ;
    RECT 71.21 38.23 71.42 38.3 ;
    RECT 71.67 37.51 71.88 37.58 ;
    RECT 71.67 37.87 71.88 37.94 ;
    RECT 71.67 38.23 71.88 38.3 ;
    RECT 31.37 37.51 31.58 37.58 ;
    RECT 31.37 37.87 31.58 37.94 ;
    RECT 31.37 38.23 31.58 38.3 ;
    RECT 31.83 37.51 32.04 37.58 ;
    RECT 31.83 37.87 32.04 37.94 ;
    RECT 31.83 38.23 32.04 38.3 ;
    RECT 67.89 37.51 68.1 37.58 ;
    RECT 67.89 37.87 68.1 37.94 ;
    RECT 67.89 38.23 68.1 38.3 ;
    RECT 68.35 37.51 68.56 37.58 ;
    RECT 68.35 37.87 68.56 37.94 ;
    RECT 68.35 38.23 68.56 38.3 ;
    RECT 28.05 37.51 28.26 37.58 ;
    RECT 28.05 37.87 28.26 37.94 ;
    RECT 28.05 38.23 28.26 38.3 ;
    RECT 28.51 37.51 28.72 37.58 ;
    RECT 28.51 37.87 28.72 37.94 ;
    RECT 28.51 38.23 28.72 38.3 ;
    RECT 24.73 37.51 24.94 37.58 ;
    RECT 24.73 37.87 24.94 37.94 ;
    RECT 24.73 38.23 24.94 38.3 ;
    RECT 25.19 37.51 25.4 37.58 ;
    RECT 25.19 37.87 25.4 37.94 ;
    RECT 25.19 38.23 25.4 38.3 ;
    RECT 21.41 37.51 21.62 37.58 ;
    RECT 21.41 37.87 21.62 37.94 ;
    RECT 21.41 38.23 21.62 38.3 ;
    RECT 21.87 37.51 22.08 37.58 ;
    RECT 21.87 37.87 22.08 37.94 ;
    RECT 21.87 38.23 22.08 38.3 ;
    RECT 18.09 37.51 18.3 37.58 ;
    RECT 18.09 37.87 18.3 37.94 ;
    RECT 18.09 38.23 18.3 38.3 ;
    RECT 18.55 37.51 18.76 37.58 ;
    RECT 18.55 37.87 18.76 37.94 ;
    RECT 18.55 38.23 18.76 38.3 ;
    RECT 120.825 37.87 120.895 37.94 ;
    RECT 14.77 37.51 14.98 37.58 ;
    RECT 14.77 37.87 14.98 37.94 ;
    RECT 14.77 38.23 14.98 38.3 ;
    RECT 15.23 37.51 15.44 37.58 ;
    RECT 15.23 37.87 15.44 37.94 ;
    RECT 15.23 38.23 15.44 38.3 ;
    RECT 11.45 37.51 11.66 37.58 ;
    RECT 11.45 37.87 11.66 37.94 ;
    RECT 11.45 38.23 11.66 38.3 ;
    RECT 11.91 37.51 12.12 37.58 ;
    RECT 11.91 37.87 12.12 37.94 ;
    RECT 11.91 38.23 12.12 38.3 ;
    RECT 8.13 37.51 8.34 37.58 ;
    RECT 8.13 37.87 8.34 37.94 ;
    RECT 8.13 38.23 8.34 38.3 ;
    RECT 8.59 37.51 8.8 37.58 ;
    RECT 8.59 37.87 8.8 37.94 ;
    RECT 8.59 38.23 8.8 38.3 ;
    RECT 4.81 37.51 5.02 37.58 ;
    RECT 4.81 37.87 5.02 37.94 ;
    RECT 4.81 38.23 5.02 38.3 ;
    RECT 5.27 37.51 5.48 37.58 ;
    RECT 5.27 37.87 5.48 37.94 ;
    RECT 5.27 38.23 5.48 38.3 ;
    RECT 1.49 37.51 1.7 37.58 ;
    RECT 1.49 37.87 1.7 37.94 ;
    RECT 1.49 38.23 1.7 38.3 ;
    RECT 1.95 37.51 2.16 37.58 ;
    RECT 1.95 37.87 2.16 37.94 ;
    RECT 1.95 38.23 2.16 38.3 ;
    RECT 64.57 37.51 64.78 37.58 ;
    RECT 64.57 37.87 64.78 37.94 ;
    RECT 64.57 38.23 64.78 38.3 ;
    RECT 65.03 37.51 65.24 37.58 ;
    RECT 65.03 37.87 65.24 37.94 ;
    RECT 65.03 38.23 65.24 38.3 ;
    RECT 61.25 77.13 61.46 77.2 ;
    RECT 61.25 77.49 61.46 77.56 ;
    RECT 61.25 77.85 61.46 77.92 ;
    RECT 61.71 77.13 61.92 77.2 ;
    RECT 61.71 77.49 61.92 77.56 ;
    RECT 61.71 77.85 61.92 77.92 ;
    RECT 57.93 77.13 58.14 77.2 ;
    RECT 57.93 77.49 58.14 77.56 ;
    RECT 57.93 77.85 58.14 77.92 ;
    RECT 58.39 77.13 58.6 77.2 ;
    RECT 58.39 77.49 58.6 77.56 ;
    RECT 58.39 77.85 58.6 77.92 ;
    RECT 54.61 77.13 54.82 77.2 ;
    RECT 54.61 77.49 54.82 77.56 ;
    RECT 54.61 77.85 54.82 77.92 ;
    RECT 55.07 77.13 55.28 77.2 ;
    RECT 55.07 77.49 55.28 77.56 ;
    RECT 55.07 77.85 55.28 77.92 ;
    RECT 51.29 77.13 51.5 77.2 ;
    RECT 51.29 77.49 51.5 77.56 ;
    RECT 51.29 77.85 51.5 77.92 ;
    RECT 51.75 77.13 51.96 77.2 ;
    RECT 51.75 77.49 51.96 77.56 ;
    RECT 51.75 77.85 51.96 77.92 ;
    RECT 47.97 77.13 48.18 77.2 ;
    RECT 47.97 77.49 48.18 77.56 ;
    RECT 47.97 77.85 48.18 77.92 ;
    RECT 48.43 77.13 48.64 77.2 ;
    RECT 48.43 77.49 48.64 77.56 ;
    RECT 48.43 77.85 48.64 77.92 ;
    RECT 44.65 77.13 44.86 77.2 ;
    RECT 44.65 77.49 44.86 77.56 ;
    RECT 44.65 77.85 44.86 77.92 ;
    RECT 45.11 77.13 45.32 77.2 ;
    RECT 45.11 77.49 45.32 77.56 ;
    RECT 45.11 77.85 45.32 77.92 ;
    RECT 41.33 77.13 41.54 77.2 ;
    RECT 41.33 77.49 41.54 77.56 ;
    RECT 41.33 77.85 41.54 77.92 ;
    RECT 41.79 77.13 42.0 77.2 ;
    RECT 41.79 77.49 42.0 77.56 ;
    RECT 41.79 77.85 42.0 77.92 ;
    RECT 38.01 77.13 38.22 77.2 ;
    RECT 38.01 77.49 38.22 77.56 ;
    RECT 38.01 77.85 38.22 77.92 ;
    RECT 38.47 77.13 38.68 77.2 ;
    RECT 38.47 77.49 38.68 77.56 ;
    RECT 38.47 77.85 38.68 77.92 ;
    RECT 0.4 77.49 0.47 77.56 ;
    RECT 34.69 77.13 34.9 77.2 ;
    RECT 34.69 77.49 34.9 77.56 ;
    RECT 34.69 77.85 34.9 77.92 ;
    RECT 35.15 77.13 35.36 77.2 ;
    RECT 35.15 77.49 35.36 77.56 ;
    RECT 35.15 77.85 35.36 77.92 ;
    RECT 117.69 77.13 117.9 77.2 ;
    RECT 117.69 77.49 117.9 77.56 ;
    RECT 117.69 77.85 117.9 77.92 ;
    RECT 118.15 77.13 118.36 77.2 ;
    RECT 118.15 77.49 118.36 77.56 ;
    RECT 118.15 77.85 118.36 77.92 ;
    RECT 114.37 77.13 114.58 77.2 ;
    RECT 114.37 77.49 114.58 77.56 ;
    RECT 114.37 77.85 114.58 77.92 ;
    RECT 114.83 77.13 115.04 77.2 ;
    RECT 114.83 77.49 115.04 77.56 ;
    RECT 114.83 77.85 115.04 77.92 ;
    RECT 111.05 77.13 111.26 77.2 ;
    RECT 111.05 77.49 111.26 77.56 ;
    RECT 111.05 77.85 111.26 77.92 ;
    RECT 111.51 77.13 111.72 77.2 ;
    RECT 111.51 77.49 111.72 77.56 ;
    RECT 111.51 77.85 111.72 77.92 ;
    RECT 107.73 77.13 107.94 77.2 ;
    RECT 107.73 77.49 107.94 77.56 ;
    RECT 107.73 77.85 107.94 77.92 ;
    RECT 108.19 77.13 108.4 77.2 ;
    RECT 108.19 77.49 108.4 77.56 ;
    RECT 108.19 77.85 108.4 77.92 ;
    RECT 104.41 77.13 104.62 77.2 ;
    RECT 104.41 77.49 104.62 77.56 ;
    RECT 104.41 77.85 104.62 77.92 ;
    RECT 104.87 77.13 105.08 77.2 ;
    RECT 104.87 77.49 105.08 77.56 ;
    RECT 104.87 77.85 105.08 77.92 ;
    RECT 101.09 77.13 101.3 77.2 ;
    RECT 101.09 77.49 101.3 77.56 ;
    RECT 101.09 77.85 101.3 77.92 ;
    RECT 101.55 77.13 101.76 77.2 ;
    RECT 101.55 77.49 101.76 77.56 ;
    RECT 101.55 77.85 101.76 77.92 ;
    RECT 97.77 77.13 97.98 77.2 ;
    RECT 97.77 77.49 97.98 77.56 ;
    RECT 97.77 77.85 97.98 77.92 ;
    RECT 98.23 77.13 98.44 77.2 ;
    RECT 98.23 77.49 98.44 77.56 ;
    RECT 98.23 77.85 98.44 77.92 ;
    RECT 94.45 77.13 94.66 77.2 ;
    RECT 94.45 77.49 94.66 77.56 ;
    RECT 94.45 77.85 94.66 77.92 ;
    RECT 94.91 77.13 95.12 77.2 ;
    RECT 94.91 77.49 95.12 77.56 ;
    RECT 94.91 77.85 95.12 77.92 ;
    RECT 91.13 77.13 91.34 77.2 ;
    RECT 91.13 77.49 91.34 77.56 ;
    RECT 91.13 77.85 91.34 77.92 ;
    RECT 91.59 77.13 91.8 77.2 ;
    RECT 91.59 77.49 91.8 77.56 ;
    RECT 91.59 77.85 91.8 77.92 ;
    RECT 87.81 77.13 88.02 77.2 ;
    RECT 87.81 77.49 88.02 77.56 ;
    RECT 87.81 77.85 88.02 77.92 ;
    RECT 88.27 77.13 88.48 77.2 ;
    RECT 88.27 77.49 88.48 77.56 ;
    RECT 88.27 77.85 88.48 77.92 ;
    RECT 84.49 77.13 84.7 77.2 ;
    RECT 84.49 77.49 84.7 77.56 ;
    RECT 84.49 77.85 84.7 77.92 ;
    RECT 84.95 77.13 85.16 77.2 ;
    RECT 84.95 77.49 85.16 77.56 ;
    RECT 84.95 77.85 85.16 77.92 ;
    RECT 81.17 77.13 81.38 77.2 ;
    RECT 81.17 77.49 81.38 77.56 ;
    RECT 81.17 77.85 81.38 77.92 ;
    RECT 81.63 77.13 81.84 77.2 ;
    RECT 81.63 77.49 81.84 77.56 ;
    RECT 81.63 77.85 81.84 77.92 ;
    RECT 77.85 77.13 78.06 77.2 ;
    RECT 77.85 77.49 78.06 77.56 ;
    RECT 77.85 77.85 78.06 77.92 ;
    RECT 78.31 77.13 78.52 77.2 ;
    RECT 78.31 77.49 78.52 77.56 ;
    RECT 78.31 77.85 78.52 77.92 ;
    RECT 74.53 77.13 74.74 77.2 ;
    RECT 74.53 77.49 74.74 77.56 ;
    RECT 74.53 77.85 74.74 77.92 ;
    RECT 74.99 77.13 75.2 77.2 ;
    RECT 74.99 77.49 75.2 77.56 ;
    RECT 74.99 77.85 75.2 77.92 ;
    RECT 71.21 77.13 71.42 77.2 ;
    RECT 71.21 77.49 71.42 77.56 ;
    RECT 71.21 77.85 71.42 77.92 ;
    RECT 71.67 77.13 71.88 77.2 ;
    RECT 71.67 77.49 71.88 77.56 ;
    RECT 71.67 77.85 71.88 77.92 ;
    RECT 31.37 77.13 31.58 77.2 ;
    RECT 31.37 77.49 31.58 77.56 ;
    RECT 31.37 77.85 31.58 77.92 ;
    RECT 31.83 77.13 32.04 77.2 ;
    RECT 31.83 77.49 32.04 77.56 ;
    RECT 31.83 77.85 32.04 77.92 ;
    RECT 67.89 77.13 68.1 77.2 ;
    RECT 67.89 77.49 68.1 77.56 ;
    RECT 67.89 77.85 68.1 77.92 ;
    RECT 68.35 77.13 68.56 77.2 ;
    RECT 68.35 77.49 68.56 77.56 ;
    RECT 68.35 77.85 68.56 77.92 ;
    RECT 28.05 77.13 28.26 77.2 ;
    RECT 28.05 77.49 28.26 77.56 ;
    RECT 28.05 77.85 28.26 77.92 ;
    RECT 28.51 77.13 28.72 77.2 ;
    RECT 28.51 77.49 28.72 77.56 ;
    RECT 28.51 77.85 28.72 77.92 ;
    RECT 24.73 77.13 24.94 77.2 ;
    RECT 24.73 77.49 24.94 77.56 ;
    RECT 24.73 77.85 24.94 77.92 ;
    RECT 25.19 77.13 25.4 77.2 ;
    RECT 25.19 77.49 25.4 77.56 ;
    RECT 25.19 77.85 25.4 77.92 ;
    RECT 21.41 77.13 21.62 77.2 ;
    RECT 21.41 77.49 21.62 77.56 ;
    RECT 21.41 77.85 21.62 77.92 ;
    RECT 21.87 77.13 22.08 77.2 ;
    RECT 21.87 77.49 22.08 77.56 ;
    RECT 21.87 77.85 22.08 77.92 ;
    RECT 18.09 77.13 18.3 77.2 ;
    RECT 18.09 77.49 18.3 77.56 ;
    RECT 18.09 77.85 18.3 77.92 ;
    RECT 18.55 77.13 18.76 77.2 ;
    RECT 18.55 77.49 18.76 77.56 ;
    RECT 18.55 77.85 18.76 77.92 ;
    RECT 120.825 77.49 120.895 77.56 ;
    RECT 14.77 77.13 14.98 77.2 ;
    RECT 14.77 77.49 14.98 77.56 ;
    RECT 14.77 77.85 14.98 77.92 ;
    RECT 15.23 77.13 15.44 77.2 ;
    RECT 15.23 77.49 15.44 77.56 ;
    RECT 15.23 77.85 15.44 77.92 ;
    RECT 11.45 77.13 11.66 77.2 ;
    RECT 11.45 77.49 11.66 77.56 ;
    RECT 11.45 77.85 11.66 77.92 ;
    RECT 11.91 77.13 12.12 77.2 ;
    RECT 11.91 77.49 12.12 77.56 ;
    RECT 11.91 77.85 12.12 77.92 ;
    RECT 8.13 77.13 8.34 77.2 ;
    RECT 8.13 77.49 8.34 77.56 ;
    RECT 8.13 77.85 8.34 77.92 ;
    RECT 8.59 77.13 8.8 77.2 ;
    RECT 8.59 77.49 8.8 77.56 ;
    RECT 8.59 77.85 8.8 77.92 ;
    RECT 4.81 77.13 5.02 77.2 ;
    RECT 4.81 77.49 5.02 77.56 ;
    RECT 4.81 77.85 5.02 77.92 ;
    RECT 5.27 77.13 5.48 77.2 ;
    RECT 5.27 77.49 5.48 77.56 ;
    RECT 5.27 77.85 5.48 77.92 ;
    RECT 1.49 77.13 1.7 77.2 ;
    RECT 1.49 77.49 1.7 77.56 ;
    RECT 1.49 77.85 1.7 77.92 ;
    RECT 1.95 77.13 2.16 77.2 ;
    RECT 1.95 77.49 2.16 77.56 ;
    RECT 1.95 77.85 2.16 77.92 ;
    RECT 64.57 77.13 64.78 77.2 ;
    RECT 64.57 77.49 64.78 77.56 ;
    RECT 64.57 77.85 64.78 77.92 ;
    RECT 65.03 77.13 65.24 77.2 ;
    RECT 65.03 77.49 65.24 77.56 ;
    RECT 65.03 77.85 65.24 77.92 ;
    RECT 61.25 36.79 61.46 36.86 ;
    RECT 61.25 37.15 61.46 37.22 ;
    RECT 61.25 37.51 61.46 37.58 ;
    RECT 61.71 36.79 61.92 36.86 ;
    RECT 61.71 37.15 61.92 37.22 ;
    RECT 61.71 37.51 61.92 37.58 ;
    RECT 57.93 36.79 58.14 36.86 ;
    RECT 57.93 37.15 58.14 37.22 ;
    RECT 57.93 37.51 58.14 37.58 ;
    RECT 58.39 36.79 58.6 36.86 ;
    RECT 58.39 37.15 58.6 37.22 ;
    RECT 58.39 37.51 58.6 37.58 ;
    RECT 54.61 36.79 54.82 36.86 ;
    RECT 54.61 37.15 54.82 37.22 ;
    RECT 54.61 37.51 54.82 37.58 ;
    RECT 55.07 36.79 55.28 36.86 ;
    RECT 55.07 37.15 55.28 37.22 ;
    RECT 55.07 37.51 55.28 37.58 ;
    RECT 51.29 36.79 51.5 36.86 ;
    RECT 51.29 37.15 51.5 37.22 ;
    RECT 51.29 37.51 51.5 37.58 ;
    RECT 51.75 36.79 51.96 36.86 ;
    RECT 51.75 37.15 51.96 37.22 ;
    RECT 51.75 37.51 51.96 37.58 ;
    RECT 47.97 36.79 48.18 36.86 ;
    RECT 47.97 37.15 48.18 37.22 ;
    RECT 47.97 37.51 48.18 37.58 ;
    RECT 48.43 36.79 48.64 36.86 ;
    RECT 48.43 37.15 48.64 37.22 ;
    RECT 48.43 37.51 48.64 37.58 ;
    RECT 44.65 36.79 44.86 36.86 ;
    RECT 44.65 37.15 44.86 37.22 ;
    RECT 44.65 37.51 44.86 37.58 ;
    RECT 45.11 36.79 45.32 36.86 ;
    RECT 45.11 37.15 45.32 37.22 ;
    RECT 45.11 37.51 45.32 37.58 ;
    RECT 41.33 36.79 41.54 36.86 ;
    RECT 41.33 37.15 41.54 37.22 ;
    RECT 41.33 37.51 41.54 37.58 ;
    RECT 41.79 36.79 42.0 36.86 ;
    RECT 41.79 37.15 42.0 37.22 ;
    RECT 41.79 37.51 42.0 37.58 ;
    RECT 38.01 36.79 38.22 36.86 ;
    RECT 38.01 37.15 38.22 37.22 ;
    RECT 38.01 37.51 38.22 37.58 ;
    RECT 38.47 36.79 38.68 36.86 ;
    RECT 38.47 37.15 38.68 37.22 ;
    RECT 38.47 37.51 38.68 37.58 ;
    RECT 0.4 37.15 0.47 37.22 ;
    RECT 34.69 36.79 34.9 36.86 ;
    RECT 34.69 37.15 34.9 37.22 ;
    RECT 34.69 37.51 34.9 37.58 ;
    RECT 35.15 36.79 35.36 36.86 ;
    RECT 35.15 37.15 35.36 37.22 ;
    RECT 35.15 37.51 35.36 37.58 ;
    RECT 117.69 36.79 117.9 36.86 ;
    RECT 117.69 37.15 117.9 37.22 ;
    RECT 117.69 37.51 117.9 37.58 ;
    RECT 118.15 36.79 118.36 36.86 ;
    RECT 118.15 37.15 118.36 37.22 ;
    RECT 118.15 37.51 118.36 37.58 ;
    RECT 114.37 36.79 114.58 36.86 ;
    RECT 114.37 37.15 114.58 37.22 ;
    RECT 114.37 37.51 114.58 37.58 ;
    RECT 114.83 36.79 115.04 36.86 ;
    RECT 114.83 37.15 115.04 37.22 ;
    RECT 114.83 37.51 115.04 37.58 ;
    RECT 111.05 36.79 111.26 36.86 ;
    RECT 111.05 37.15 111.26 37.22 ;
    RECT 111.05 37.51 111.26 37.58 ;
    RECT 111.51 36.79 111.72 36.86 ;
    RECT 111.51 37.15 111.72 37.22 ;
    RECT 111.51 37.51 111.72 37.58 ;
    RECT 107.73 36.79 107.94 36.86 ;
    RECT 107.73 37.15 107.94 37.22 ;
    RECT 107.73 37.51 107.94 37.58 ;
    RECT 108.19 36.79 108.4 36.86 ;
    RECT 108.19 37.15 108.4 37.22 ;
    RECT 108.19 37.51 108.4 37.58 ;
    RECT 104.41 36.79 104.62 36.86 ;
    RECT 104.41 37.15 104.62 37.22 ;
    RECT 104.41 37.51 104.62 37.58 ;
    RECT 104.87 36.79 105.08 36.86 ;
    RECT 104.87 37.15 105.08 37.22 ;
    RECT 104.87 37.51 105.08 37.58 ;
    RECT 101.09 36.79 101.3 36.86 ;
    RECT 101.09 37.15 101.3 37.22 ;
    RECT 101.09 37.51 101.3 37.58 ;
    RECT 101.55 36.79 101.76 36.86 ;
    RECT 101.55 37.15 101.76 37.22 ;
    RECT 101.55 37.51 101.76 37.58 ;
    RECT 97.77 36.79 97.98 36.86 ;
    RECT 97.77 37.15 97.98 37.22 ;
    RECT 97.77 37.51 97.98 37.58 ;
    RECT 98.23 36.79 98.44 36.86 ;
    RECT 98.23 37.15 98.44 37.22 ;
    RECT 98.23 37.51 98.44 37.58 ;
    RECT 94.45 36.79 94.66 36.86 ;
    RECT 94.45 37.15 94.66 37.22 ;
    RECT 94.45 37.51 94.66 37.58 ;
    RECT 94.91 36.79 95.12 36.86 ;
    RECT 94.91 37.15 95.12 37.22 ;
    RECT 94.91 37.51 95.12 37.58 ;
    RECT 91.13 36.79 91.34 36.86 ;
    RECT 91.13 37.15 91.34 37.22 ;
    RECT 91.13 37.51 91.34 37.58 ;
    RECT 91.59 36.79 91.8 36.86 ;
    RECT 91.59 37.15 91.8 37.22 ;
    RECT 91.59 37.51 91.8 37.58 ;
    RECT 87.81 36.79 88.02 36.86 ;
    RECT 87.81 37.15 88.02 37.22 ;
    RECT 87.81 37.51 88.02 37.58 ;
    RECT 88.27 36.79 88.48 36.86 ;
    RECT 88.27 37.15 88.48 37.22 ;
    RECT 88.27 37.51 88.48 37.58 ;
    RECT 84.49 36.79 84.7 36.86 ;
    RECT 84.49 37.15 84.7 37.22 ;
    RECT 84.49 37.51 84.7 37.58 ;
    RECT 84.95 36.79 85.16 36.86 ;
    RECT 84.95 37.15 85.16 37.22 ;
    RECT 84.95 37.51 85.16 37.58 ;
    RECT 81.17 36.79 81.38 36.86 ;
    RECT 81.17 37.15 81.38 37.22 ;
    RECT 81.17 37.51 81.38 37.58 ;
    RECT 81.63 36.79 81.84 36.86 ;
    RECT 81.63 37.15 81.84 37.22 ;
    RECT 81.63 37.51 81.84 37.58 ;
    RECT 77.85 36.79 78.06 36.86 ;
    RECT 77.85 37.15 78.06 37.22 ;
    RECT 77.85 37.51 78.06 37.58 ;
    RECT 78.31 36.79 78.52 36.86 ;
    RECT 78.31 37.15 78.52 37.22 ;
    RECT 78.31 37.51 78.52 37.58 ;
    RECT 74.53 36.79 74.74 36.86 ;
    RECT 74.53 37.15 74.74 37.22 ;
    RECT 74.53 37.51 74.74 37.58 ;
    RECT 74.99 36.79 75.2 36.86 ;
    RECT 74.99 37.15 75.2 37.22 ;
    RECT 74.99 37.51 75.2 37.58 ;
    RECT 71.21 36.79 71.42 36.86 ;
    RECT 71.21 37.15 71.42 37.22 ;
    RECT 71.21 37.51 71.42 37.58 ;
    RECT 71.67 36.79 71.88 36.86 ;
    RECT 71.67 37.15 71.88 37.22 ;
    RECT 71.67 37.51 71.88 37.58 ;
    RECT 31.37 36.79 31.58 36.86 ;
    RECT 31.37 37.15 31.58 37.22 ;
    RECT 31.37 37.51 31.58 37.58 ;
    RECT 31.83 36.79 32.04 36.86 ;
    RECT 31.83 37.15 32.04 37.22 ;
    RECT 31.83 37.51 32.04 37.58 ;
    RECT 67.89 36.79 68.1 36.86 ;
    RECT 67.89 37.15 68.1 37.22 ;
    RECT 67.89 37.51 68.1 37.58 ;
    RECT 68.35 36.79 68.56 36.86 ;
    RECT 68.35 37.15 68.56 37.22 ;
    RECT 68.35 37.51 68.56 37.58 ;
    RECT 28.05 36.79 28.26 36.86 ;
    RECT 28.05 37.15 28.26 37.22 ;
    RECT 28.05 37.51 28.26 37.58 ;
    RECT 28.51 36.79 28.72 36.86 ;
    RECT 28.51 37.15 28.72 37.22 ;
    RECT 28.51 37.51 28.72 37.58 ;
    RECT 24.73 36.79 24.94 36.86 ;
    RECT 24.73 37.15 24.94 37.22 ;
    RECT 24.73 37.51 24.94 37.58 ;
    RECT 25.19 36.79 25.4 36.86 ;
    RECT 25.19 37.15 25.4 37.22 ;
    RECT 25.19 37.51 25.4 37.58 ;
    RECT 21.41 36.79 21.62 36.86 ;
    RECT 21.41 37.15 21.62 37.22 ;
    RECT 21.41 37.51 21.62 37.58 ;
    RECT 21.87 36.79 22.08 36.86 ;
    RECT 21.87 37.15 22.08 37.22 ;
    RECT 21.87 37.51 22.08 37.58 ;
    RECT 18.09 36.79 18.3 36.86 ;
    RECT 18.09 37.15 18.3 37.22 ;
    RECT 18.09 37.51 18.3 37.58 ;
    RECT 18.55 36.79 18.76 36.86 ;
    RECT 18.55 37.15 18.76 37.22 ;
    RECT 18.55 37.51 18.76 37.58 ;
    RECT 120.825 37.15 120.895 37.22 ;
    RECT 14.77 36.79 14.98 36.86 ;
    RECT 14.77 37.15 14.98 37.22 ;
    RECT 14.77 37.51 14.98 37.58 ;
    RECT 15.23 36.79 15.44 36.86 ;
    RECT 15.23 37.15 15.44 37.22 ;
    RECT 15.23 37.51 15.44 37.58 ;
    RECT 11.45 36.79 11.66 36.86 ;
    RECT 11.45 37.15 11.66 37.22 ;
    RECT 11.45 37.51 11.66 37.58 ;
    RECT 11.91 36.79 12.12 36.86 ;
    RECT 11.91 37.15 12.12 37.22 ;
    RECT 11.91 37.51 12.12 37.58 ;
    RECT 8.13 36.79 8.34 36.86 ;
    RECT 8.13 37.15 8.34 37.22 ;
    RECT 8.13 37.51 8.34 37.58 ;
    RECT 8.59 36.79 8.8 36.86 ;
    RECT 8.59 37.15 8.8 37.22 ;
    RECT 8.59 37.51 8.8 37.58 ;
    RECT 4.81 36.79 5.02 36.86 ;
    RECT 4.81 37.15 5.02 37.22 ;
    RECT 4.81 37.51 5.02 37.58 ;
    RECT 5.27 36.79 5.48 36.86 ;
    RECT 5.27 37.15 5.48 37.22 ;
    RECT 5.27 37.51 5.48 37.58 ;
    RECT 1.49 36.79 1.7 36.86 ;
    RECT 1.49 37.15 1.7 37.22 ;
    RECT 1.49 37.51 1.7 37.58 ;
    RECT 1.95 36.79 2.16 36.86 ;
    RECT 1.95 37.15 2.16 37.22 ;
    RECT 1.95 37.51 2.16 37.58 ;
    RECT 64.57 36.79 64.78 36.86 ;
    RECT 64.57 37.15 64.78 37.22 ;
    RECT 64.57 37.51 64.78 37.58 ;
    RECT 65.03 36.79 65.24 36.86 ;
    RECT 65.03 37.15 65.24 37.22 ;
    RECT 65.03 37.51 65.24 37.58 ;
    RECT 61.25 76.41 61.46 76.48 ;
    RECT 61.25 76.77 61.46 76.84 ;
    RECT 61.25 77.13 61.46 77.2 ;
    RECT 61.71 76.41 61.92 76.48 ;
    RECT 61.71 76.77 61.92 76.84 ;
    RECT 61.71 77.13 61.92 77.2 ;
    RECT 57.93 76.41 58.14 76.48 ;
    RECT 57.93 76.77 58.14 76.84 ;
    RECT 57.93 77.13 58.14 77.2 ;
    RECT 58.39 76.41 58.6 76.48 ;
    RECT 58.39 76.77 58.6 76.84 ;
    RECT 58.39 77.13 58.6 77.2 ;
    RECT 54.61 76.41 54.82 76.48 ;
    RECT 54.61 76.77 54.82 76.84 ;
    RECT 54.61 77.13 54.82 77.2 ;
    RECT 55.07 76.41 55.28 76.48 ;
    RECT 55.07 76.77 55.28 76.84 ;
    RECT 55.07 77.13 55.28 77.2 ;
    RECT 51.29 76.41 51.5 76.48 ;
    RECT 51.29 76.77 51.5 76.84 ;
    RECT 51.29 77.13 51.5 77.2 ;
    RECT 51.75 76.41 51.96 76.48 ;
    RECT 51.75 76.77 51.96 76.84 ;
    RECT 51.75 77.13 51.96 77.2 ;
    RECT 47.97 76.41 48.18 76.48 ;
    RECT 47.97 76.77 48.18 76.84 ;
    RECT 47.97 77.13 48.18 77.2 ;
    RECT 48.43 76.41 48.64 76.48 ;
    RECT 48.43 76.77 48.64 76.84 ;
    RECT 48.43 77.13 48.64 77.2 ;
    RECT 44.65 76.41 44.86 76.48 ;
    RECT 44.65 76.77 44.86 76.84 ;
    RECT 44.65 77.13 44.86 77.2 ;
    RECT 45.11 76.41 45.32 76.48 ;
    RECT 45.11 76.77 45.32 76.84 ;
    RECT 45.11 77.13 45.32 77.2 ;
    RECT 41.33 76.41 41.54 76.48 ;
    RECT 41.33 76.77 41.54 76.84 ;
    RECT 41.33 77.13 41.54 77.2 ;
    RECT 41.79 76.41 42.0 76.48 ;
    RECT 41.79 76.77 42.0 76.84 ;
    RECT 41.79 77.13 42.0 77.2 ;
    RECT 38.01 76.41 38.22 76.48 ;
    RECT 38.01 76.77 38.22 76.84 ;
    RECT 38.01 77.13 38.22 77.2 ;
    RECT 38.47 76.41 38.68 76.48 ;
    RECT 38.47 76.77 38.68 76.84 ;
    RECT 38.47 77.13 38.68 77.2 ;
    RECT 0.4 76.77 0.47 76.84 ;
    RECT 34.69 76.41 34.9 76.48 ;
    RECT 34.69 76.77 34.9 76.84 ;
    RECT 34.69 77.13 34.9 77.2 ;
    RECT 35.15 76.41 35.36 76.48 ;
    RECT 35.15 76.77 35.36 76.84 ;
    RECT 35.15 77.13 35.36 77.2 ;
    RECT 117.69 76.41 117.9 76.48 ;
    RECT 117.69 76.77 117.9 76.84 ;
    RECT 117.69 77.13 117.9 77.2 ;
    RECT 118.15 76.41 118.36 76.48 ;
    RECT 118.15 76.77 118.36 76.84 ;
    RECT 118.15 77.13 118.36 77.2 ;
    RECT 114.37 76.41 114.58 76.48 ;
    RECT 114.37 76.77 114.58 76.84 ;
    RECT 114.37 77.13 114.58 77.2 ;
    RECT 114.83 76.41 115.04 76.48 ;
    RECT 114.83 76.77 115.04 76.84 ;
    RECT 114.83 77.13 115.04 77.2 ;
    RECT 111.05 76.41 111.26 76.48 ;
    RECT 111.05 76.77 111.26 76.84 ;
    RECT 111.05 77.13 111.26 77.2 ;
    RECT 111.51 76.41 111.72 76.48 ;
    RECT 111.51 76.77 111.72 76.84 ;
    RECT 111.51 77.13 111.72 77.2 ;
    RECT 107.73 76.41 107.94 76.48 ;
    RECT 107.73 76.77 107.94 76.84 ;
    RECT 107.73 77.13 107.94 77.2 ;
    RECT 108.19 76.41 108.4 76.48 ;
    RECT 108.19 76.77 108.4 76.84 ;
    RECT 108.19 77.13 108.4 77.2 ;
    RECT 104.41 76.41 104.62 76.48 ;
    RECT 104.41 76.77 104.62 76.84 ;
    RECT 104.41 77.13 104.62 77.2 ;
    RECT 104.87 76.41 105.08 76.48 ;
    RECT 104.87 76.77 105.08 76.84 ;
    RECT 104.87 77.13 105.08 77.2 ;
    RECT 101.09 76.41 101.3 76.48 ;
    RECT 101.09 76.77 101.3 76.84 ;
    RECT 101.09 77.13 101.3 77.2 ;
    RECT 101.55 76.41 101.76 76.48 ;
    RECT 101.55 76.77 101.76 76.84 ;
    RECT 101.55 77.13 101.76 77.2 ;
    RECT 97.77 76.41 97.98 76.48 ;
    RECT 97.77 76.77 97.98 76.84 ;
    RECT 97.77 77.13 97.98 77.2 ;
    RECT 98.23 76.41 98.44 76.48 ;
    RECT 98.23 76.77 98.44 76.84 ;
    RECT 98.23 77.13 98.44 77.2 ;
    RECT 94.45 76.41 94.66 76.48 ;
    RECT 94.45 76.77 94.66 76.84 ;
    RECT 94.45 77.13 94.66 77.2 ;
    RECT 94.91 76.41 95.12 76.48 ;
    RECT 94.91 76.77 95.12 76.84 ;
    RECT 94.91 77.13 95.12 77.2 ;
    RECT 91.13 76.41 91.34 76.48 ;
    RECT 91.13 76.77 91.34 76.84 ;
    RECT 91.13 77.13 91.34 77.2 ;
    RECT 91.59 76.41 91.8 76.48 ;
    RECT 91.59 76.77 91.8 76.84 ;
    RECT 91.59 77.13 91.8 77.2 ;
    RECT 87.81 76.41 88.02 76.48 ;
    RECT 87.81 76.77 88.02 76.84 ;
    RECT 87.81 77.13 88.02 77.2 ;
    RECT 88.27 76.41 88.48 76.48 ;
    RECT 88.27 76.77 88.48 76.84 ;
    RECT 88.27 77.13 88.48 77.2 ;
    RECT 84.49 76.41 84.7 76.48 ;
    RECT 84.49 76.77 84.7 76.84 ;
    RECT 84.49 77.13 84.7 77.2 ;
    RECT 84.95 76.41 85.16 76.48 ;
    RECT 84.95 76.77 85.16 76.84 ;
    RECT 84.95 77.13 85.16 77.2 ;
    RECT 81.17 76.41 81.38 76.48 ;
    RECT 81.17 76.77 81.38 76.84 ;
    RECT 81.17 77.13 81.38 77.2 ;
    RECT 81.63 76.41 81.84 76.48 ;
    RECT 81.63 76.77 81.84 76.84 ;
    RECT 81.63 77.13 81.84 77.2 ;
    RECT 77.85 76.41 78.06 76.48 ;
    RECT 77.85 76.77 78.06 76.84 ;
    RECT 77.85 77.13 78.06 77.2 ;
    RECT 78.31 76.41 78.52 76.48 ;
    RECT 78.31 76.77 78.52 76.84 ;
    RECT 78.31 77.13 78.52 77.2 ;
    RECT 74.53 76.41 74.74 76.48 ;
    RECT 74.53 76.77 74.74 76.84 ;
    RECT 74.53 77.13 74.74 77.2 ;
    RECT 74.99 76.41 75.2 76.48 ;
    RECT 74.99 76.77 75.2 76.84 ;
    RECT 74.99 77.13 75.2 77.2 ;
    RECT 71.21 76.41 71.42 76.48 ;
    RECT 71.21 76.77 71.42 76.84 ;
    RECT 71.21 77.13 71.42 77.2 ;
    RECT 71.67 76.41 71.88 76.48 ;
    RECT 71.67 76.77 71.88 76.84 ;
    RECT 71.67 77.13 71.88 77.2 ;
    RECT 31.37 76.41 31.58 76.48 ;
    RECT 31.37 76.77 31.58 76.84 ;
    RECT 31.37 77.13 31.58 77.2 ;
    RECT 31.83 76.41 32.04 76.48 ;
    RECT 31.83 76.77 32.04 76.84 ;
    RECT 31.83 77.13 32.04 77.2 ;
    RECT 67.89 76.41 68.1 76.48 ;
    RECT 67.89 76.77 68.1 76.84 ;
    RECT 67.89 77.13 68.1 77.2 ;
    RECT 68.35 76.41 68.56 76.48 ;
    RECT 68.35 76.77 68.56 76.84 ;
    RECT 68.35 77.13 68.56 77.2 ;
    RECT 28.05 76.41 28.26 76.48 ;
    RECT 28.05 76.77 28.26 76.84 ;
    RECT 28.05 77.13 28.26 77.2 ;
    RECT 28.51 76.41 28.72 76.48 ;
    RECT 28.51 76.77 28.72 76.84 ;
    RECT 28.51 77.13 28.72 77.2 ;
    RECT 24.73 76.41 24.94 76.48 ;
    RECT 24.73 76.77 24.94 76.84 ;
    RECT 24.73 77.13 24.94 77.2 ;
    RECT 25.19 76.41 25.4 76.48 ;
    RECT 25.19 76.77 25.4 76.84 ;
    RECT 25.19 77.13 25.4 77.2 ;
    RECT 21.41 76.41 21.62 76.48 ;
    RECT 21.41 76.77 21.62 76.84 ;
    RECT 21.41 77.13 21.62 77.2 ;
    RECT 21.87 76.41 22.08 76.48 ;
    RECT 21.87 76.77 22.08 76.84 ;
    RECT 21.87 77.13 22.08 77.2 ;
    RECT 18.09 76.41 18.3 76.48 ;
    RECT 18.09 76.77 18.3 76.84 ;
    RECT 18.09 77.13 18.3 77.2 ;
    RECT 18.55 76.41 18.76 76.48 ;
    RECT 18.55 76.77 18.76 76.84 ;
    RECT 18.55 77.13 18.76 77.2 ;
    RECT 120.825 76.77 120.895 76.84 ;
    RECT 14.77 76.41 14.98 76.48 ;
    RECT 14.77 76.77 14.98 76.84 ;
    RECT 14.77 77.13 14.98 77.2 ;
    RECT 15.23 76.41 15.44 76.48 ;
    RECT 15.23 76.77 15.44 76.84 ;
    RECT 15.23 77.13 15.44 77.2 ;
    RECT 11.45 76.41 11.66 76.48 ;
    RECT 11.45 76.77 11.66 76.84 ;
    RECT 11.45 77.13 11.66 77.2 ;
    RECT 11.91 76.41 12.12 76.48 ;
    RECT 11.91 76.77 12.12 76.84 ;
    RECT 11.91 77.13 12.12 77.2 ;
    RECT 8.13 76.41 8.34 76.48 ;
    RECT 8.13 76.77 8.34 76.84 ;
    RECT 8.13 77.13 8.34 77.2 ;
    RECT 8.59 76.41 8.8 76.48 ;
    RECT 8.59 76.77 8.8 76.84 ;
    RECT 8.59 77.13 8.8 77.2 ;
    RECT 4.81 76.41 5.02 76.48 ;
    RECT 4.81 76.77 5.02 76.84 ;
    RECT 4.81 77.13 5.02 77.2 ;
    RECT 5.27 76.41 5.48 76.48 ;
    RECT 5.27 76.77 5.48 76.84 ;
    RECT 5.27 77.13 5.48 77.2 ;
    RECT 1.49 76.41 1.7 76.48 ;
    RECT 1.49 76.77 1.7 76.84 ;
    RECT 1.49 77.13 1.7 77.2 ;
    RECT 1.95 76.41 2.16 76.48 ;
    RECT 1.95 76.77 2.16 76.84 ;
    RECT 1.95 77.13 2.16 77.2 ;
    RECT 64.57 76.41 64.78 76.48 ;
    RECT 64.57 76.77 64.78 76.84 ;
    RECT 64.57 77.13 64.78 77.2 ;
    RECT 65.03 76.41 65.24 76.48 ;
    RECT 65.03 76.77 65.24 76.84 ;
    RECT 65.03 77.13 65.24 77.2 ;
    RECT 61.25 36.07 61.46 36.14 ;
    RECT 61.25 36.43 61.46 36.5 ;
    RECT 61.25 36.79 61.46 36.86 ;
    RECT 61.71 36.07 61.92 36.14 ;
    RECT 61.71 36.43 61.92 36.5 ;
    RECT 61.71 36.79 61.92 36.86 ;
    RECT 57.93 36.07 58.14 36.14 ;
    RECT 57.93 36.43 58.14 36.5 ;
    RECT 57.93 36.79 58.14 36.86 ;
    RECT 58.39 36.07 58.6 36.14 ;
    RECT 58.39 36.43 58.6 36.5 ;
    RECT 58.39 36.79 58.6 36.86 ;
    RECT 54.61 36.07 54.82 36.14 ;
    RECT 54.61 36.43 54.82 36.5 ;
    RECT 54.61 36.79 54.82 36.86 ;
    RECT 55.07 36.07 55.28 36.14 ;
    RECT 55.07 36.43 55.28 36.5 ;
    RECT 55.07 36.79 55.28 36.86 ;
    RECT 51.29 36.07 51.5 36.14 ;
    RECT 51.29 36.43 51.5 36.5 ;
    RECT 51.29 36.79 51.5 36.86 ;
    RECT 51.75 36.07 51.96 36.14 ;
    RECT 51.75 36.43 51.96 36.5 ;
    RECT 51.75 36.79 51.96 36.86 ;
    RECT 47.97 36.07 48.18 36.14 ;
    RECT 47.97 36.43 48.18 36.5 ;
    RECT 47.97 36.79 48.18 36.86 ;
    RECT 48.43 36.07 48.64 36.14 ;
    RECT 48.43 36.43 48.64 36.5 ;
    RECT 48.43 36.79 48.64 36.86 ;
    RECT 44.65 36.07 44.86 36.14 ;
    RECT 44.65 36.43 44.86 36.5 ;
    RECT 44.65 36.79 44.86 36.86 ;
    RECT 45.11 36.07 45.32 36.14 ;
    RECT 45.11 36.43 45.32 36.5 ;
    RECT 45.11 36.79 45.32 36.86 ;
    RECT 41.33 36.07 41.54 36.14 ;
    RECT 41.33 36.43 41.54 36.5 ;
    RECT 41.33 36.79 41.54 36.86 ;
    RECT 41.79 36.07 42.0 36.14 ;
    RECT 41.79 36.43 42.0 36.5 ;
    RECT 41.79 36.79 42.0 36.86 ;
    RECT 38.01 36.07 38.22 36.14 ;
    RECT 38.01 36.43 38.22 36.5 ;
    RECT 38.01 36.79 38.22 36.86 ;
    RECT 38.47 36.07 38.68 36.14 ;
    RECT 38.47 36.43 38.68 36.5 ;
    RECT 38.47 36.79 38.68 36.86 ;
    RECT 0.4 36.43 0.47 36.5 ;
    RECT 34.69 36.07 34.9 36.14 ;
    RECT 34.69 36.43 34.9 36.5 ;
    RECT 34.69 36.79 34.9 36.86 ;
    RECT 35.15 36.07 35.36 36.14 ;
    RECT 35.15 36.43 35.36 36.5 ;
    RECT 35.15 36.79 35.36 36.86 ;
    RECT 117.69 36.07 117.9 36.14 ;
    RECT 117.69 36.43 117.9 36.5 ;
    RECT 117.69 36.79 117.9 36.86 ;
    RECT 118.15 36.07 118.36 36.14 ;
    RECT 118.15 36.43 118.36 36.5 ;
    RECT 118.15 36.79 118.36 36.86 ;
    RECT 114.37 36.07 114.58 36.14 ;
    RECT 114.37 36.43 114.58 36.5 ;
    RECT 114.37 36.79 114.58 36.86 ;
    RECT 114.83 36.07 115.04 36.14 ;
    RECT 114.83 36.43 115.04 36.5 ;
    RECT 114.83 36.79 115.04 36.86 ;
    RECT 111.05 36.07 111.26 36.14 ;
    RECT 111.05 36.43 111.26 36.5 ;
    RECT 111.05 36.79 111.26 36.86 ;
    RECT 111.51 36.07 111.72 36.14 ;
    RECT 111.51 36.43 111.72 36.5 ;
    RECT 111.51 36.79 111.72 36.86 ;
    RECT 107.73 36.07 107.94 36.14 ;
    RECT 107.73 36.43 107.94 36.5 ;
    RECT 107.73 36.79 107.94 36.86 ;
    RECT 108.19 36.07 108.4 36.14 ;
    RECT 108.19 36.43 108.4 36.5 ;
    RECT 108.19 36.79 108.4 36.86 ;
    RECT 104.41 36.07 104.62 36.14 ;
    RECT 104.41 36.43 104.62 36.5 ;
    RECT 104.41 36.79 104.62 36.86 ;
    RECT 104.87 36.07 105.08 36.14 ;
    RECT 104.87 36.43 105.08 36.5 ;
    RECT 104.87 36.79 105.08 36.86 ;
    RECT 101.09 36.07 101.3 36.14 ;
    RECT 101.09 36.43 101.3 36.5 ;
    RECT 101.09 36.79 101.3 36.86 ;
    RECT 101.55 36.07 101.76 36.14 ;
    RECT 101.55 36.43 101.76 36.5 ;
    RECT 101.55 36.79 101.76 36.86 ;
    RECT 97.77 36.07 97.98 36.14 ;
    RECT 97.77 36.43 97.98 36.5 ;
    RECT 97.77 36.79 97.98 36.86 ;
    RECT 98.23 36.07 98.44 36.14 ;
    RECT 98.23 36.43 98.44 36.5 ;
    RECT 98.23 36.79 98.44 36.86 ;
    RECT 94.45 36.07 94.66 36.14 ;
    RECT 94.45 36.43 94.66 36.5 ;
    RECT 94.45 36.79 94.66 36.86 ;
    RECT 94.91 36.07 95.12 36.14 ;
    RECT 94.91 36.43 95.12 36.5 ;
    RECT 94.91 36.79 95.12 36.86 ;
    RECT 91.13 36.07 91.34 36.14 ;
    RECT 91.13 36.43 91.34 36.5 ;
    RECT 91.13 36.79 91.34 36.86 ;
    RECT 91.59 36.07 91.8 36.14 ;
    RECT 91.59 36.43 91.8 36.5 ;
    RECT 91.59 36.79 91.8 36.86 ;
    RECT 87.81 36.07 88.02 36.14 ;
    RECT 87.81 36.43 88.02 36.5 ;
    RECT 87.81 36.79 88.02 36.86 ;
    RECT 88.27 36.07 88.48 36.14 ;
    RECT 88.27 36.43 88.48 36.5 ;
    RECT 88.27 36.79 88.48 36.86 ;
    RECT 84.49 36.07 84.7 36.14 ;
    RECT 84.49 36.43 84.7 36.5 ;
    RECT 84.49 36.79 84.7 36.86 ;
    RECT 84.95 36.07 85.16 36.14 ;
    RECT 84.95 36.43 85.16 36.5 ;
    RECT 84.95 36.79 85.16 36.86 ;
    RECT 81.17 36.07 81.38 36.14 ;
    RECT 81.17 36.43 81.38 36.5 ;
    RECT 81.17 36.79 81.38 36.86 ;
    RECT 81.63 36.07 81.84 36.14 ;
    RECT 81.63 36.43 81.84 36.5 ;
    RECT 81.63 36.79 81.84 36.86 ;
    RECT 77.85 36.07 78.06 36.14 ;
    RECT 77.85 36.43 78.06 36.5 ;
    RECT 77.85 36.79 78.06 36.86 ;
    RECT 78.31 36.07 78.52 36.14 ;
    RECT 78.31 36.43 78.52 36.5 ;
    RECT 78.31 36.79 78.52 36.86 ;
    RECT 74.53 36.07 74.74 36.14 ;
    RECT 74.53 36.43 74.74 36.5 ;
    RECT 74.53 36.79 74.74 36.86 ;
    RECT 74.99 36.07 75.2 36.14 ;
    RECT 74.99 36.43 75.2 36.5 ;
    RECT 74.99 36.79 75.2 36.86 ;
    RECT 71.21 36.07 71.42 36.14 ;
    RECT 71.21 36.43 71.42 36.5 ;
    RECT 71.21 36.79 71.42 36.86 ;
    RECT 71.67 36.07 71.88 36.14 ;
    RECT 71.67 36.43 71.88 36.5 ;
    RECT 71.67 36.79 71.88 36.86 ;
    RECT 31.37 36.07 31.58 36.14 ;
    RECT 31.37 36.43 31.58 36.5 ;
    RECT 31.37 36.79 31.58 36.86 ;
    RECT 31.83 36.07 32.04 36.14 ;
    RECT 31.83 36.43 32.04 36.5 ;
    RECT 31.83 36.79 32.04 36.86 ;
    RECT 67.89 36.07 68.1 36.14 ;
    RECT 67.89 36.43 68.1 36.5 ;
    RECT 67.89 36.79 68.1 36.86 ;
    RECT 68.35 36.07 68.56 36.14 ;
    RECT 68.35 36.43 68.56 36.5 ;
    RECT 68.35 36.79 68.56 36.86 ;
    RECT 28.05 36.07 28.26 36.14 ;
    RECT 28.05 36.43 28.26 36.5 ;
    RECT 28.05 36.79 28.26 36.86 ;
    RECT 28.51 36.07 28.72 36.14 ;
    RECT 28.51 36.43 28.72 36.5 ;
    RECT 28.51 36.79 28.72 36.86 ;
    RECT 24.73 36.07 24.94 36.14 ;
    RECT 24.73 36.43 24.94 36.5 ;
    RECT 24.73 36.79 24.94 36.86 ;
    RECT 25.19 36.07 25.4 36.14 ;
    RECT 25.19 36.43 25.4 36.5 ;
    RECT 25.19 36.79 25.4 36.86 ;
    RECT 21.41 36.07 21.62 36.14 ;
    RECT 21.41 36.43 21.62 36.5 ;
    RECT 21.41 36.79 21.62 36.86 ;
    RECT 21.87 36.07 22.08 36.14 ;
    RECT 21.87 36.43 22.08 36.5 ;
    RECT 21.87 36.79 22.08 36.86 ;
    RECT 18.09 36.07 18.3 36.14 ;
    RECT 18.09 36.43 18.3 36.5 ;
    RECT 18.09 36.79 18.3 36.86 ;
    RECT 18.55 36.07 18.76 36.14 ;
    RECT 18.55 36.43 18.76 36.5 ;
    RECT 18.55 36.79 18.76 36.86 ;
    RECT 120.825 36.43 120.895 36.5 ;
    RECT 14.77 36.07 14.98 36.14 ;
    RECT 14.77 36.43 14.98 36.5 ;
    RECT 14.77 36.79 14.98 36.86 ;
    RECT 15.23 36.07 15.44 36.14 ;
    RECT 15.23 36.43 15.44 36.5 ;
    RECT 15.23 36.79 15.44 36.86 ;
    RECT 11.45 36.07 11.66 36.14 ;
    RECT 11.45 36.43 11.66 36.5 ;
    RECT 11.45 36.79 11.66 36.86 ;
    RECT 11.91 36.07 12.12 36.14 ;
    RECT 11.91 36.43 12.12 36.5 ;
    RECT 11.91 36.79 12.12 36.86 ;
    RECT 8.13 36.07 8.34 36.14 ;
    RECT 8.13 36.43 8.34 36.5 ;
    RECT 8.13 36.79 8.34 36.86 ;
    RECT 8.59 36.07 8.8 36.14 ;
    RECT 8.59 36.43 8.8 36.5 ;
    RECT 8.59 36.79 8.8 36.86 ;
    RECT 4.81 36.07 5.02 36.14 ;
    RECT 4.81 36.43 5.02 36.5 ;
    RECT 4.81 36.79 5.02 36.86 ;
    RECT 5.27 36.07 5.48 36.14 ;
    RECT 5.27 36.43 5.48 36.5 ;
    RECT 5.27 36.79 5.48 36.86 ;
    RECT 1.49 36.07 1.7 36.14 ;
    RECT 1.49 36.43 1.7 36.5 ;
    RECT 1.49 36.79 1.7 36.86 ;
    RECT 1.95 36.07 2.16 36.14 ;
    RECT 1.95 36.43 2.16 36.5 ;
    RECT 1.95 36.79 2.16 36.86 ;
    RECT 64.57 36.07 64.78 36.14 ;
    RECT 64.57 36.43 64.78 36.5 ;
    RECT 64.57 36.79 64.78 36.86 ;
    RECT 65.03 36.07 65.24 36.14 ;
    RECT 65.03 36.43 65.24 36.5 ;
    RECT 65.03 36.79 65.24 36.86 ;
    RECT 61.25 75.69 61.46 75.76 ;
    RECT 61.25 76.05 61.46 76.12 ;
    RECT 61.25 76.41 61.46 76.48 ;
    RECT 61.71 75.69 61.92 75.76 ;
    RECT 61.71 76.05 61.92 76.12 ;
    RECT 61.71 76.41 61.92 76.48 ;
    RECT 57.93 75.69 58.14 75.76 ;
    RECT 57.93 76.05 58.14 76.12 ;
    RECT 57.93 76.41 58.14 76.48 ;
    RECT 58.39 75.69 58.6 75.76 ;
    RECT 58.39 76.05 58.6 76.12 ;
    RECT 58.39 76.41 58.6 76.48 ;
    RECT 54.61 75.69 54.82 75.76 ;
    RECT 54.61 76.05 54.82 76.12 ;
    RECT 54.61 76.41 54.82 76.48 ;
    RECT 55.07 75.69 55.28 75.76 ;
    RECT 55.07 76.05 55.28 76.12 ;
    RECT 55.07 76.41 55.28 76.48 ;
    RECT 51.29 75.69 51.5 75.76 ;
    RECT 51.29 76.05 51.5 76.12 ;
    RECT 51.29 76.41 51.5 76.48 ;
    RECT 51.75 75.69 51.96 75.76 ;
    RECT 51.75 76.05 51.96 76.12 ;
    RECT 51.75 76.41 51.96 76.48 ;
    RECT 47.97 75.69 48.18 75.76 ;
    RECT 47.97 76.05 48.18 76.12 ;
    RECT 47.97 76.41 48.18 76.48 ;
    RECT 48.43 75.69 48.64 75.76 ;
    RECT 48.43 76.05 48.64 76.12 ;
    RECT 48.43 76.41 48.64 76.48 ;
    RECT 44.65 75.69 44.86 75.76 ;
    RECT 44.65 76.05 44.86 76.12 ;
    RECT 44.65 76.41 44.86 76.48 ;
    RECT 45.11 75.69 45.32 75.76 ;
    RECT 45.11 76.05 45.32 76.12 ;
    RECT 45.11 76.41 45.32 76.48 ;
    RECT 41.33 75.69 41.54 75.76 ;
    RECT 41.33 76.05 41.54 76.12 ;
    RECT 41.33 76.41 41.54 76.48 ;
    RECT 41.79 75.69 42.0 75.76 ;
    RECT 41.79 76.05 42.0 76.12 ;
    RECT 41.79 76.41 42.0 76.48 ;
    RECT 38.01 75.69 38.22 75.76 ;
    RECT 38.01 76.05 38.22 76.12 ;
    RECT 38.01 76.41 38.22 76.48 ;
    RECT 38.47 75.69 38.68 75.76 ;
    RECT 38.47 76.05 38.68 76.12 ;
    RECT 38.47 76.41 38.68 76.48 ;
    RECT 0.4 76.05 0.47 76.12 ;
    RECT 34.69 75.69 34.9 75.76 ;
    RECT 34.69 76.05 34.9 76.12 ;
    RECT 34.69 76.41 34.9 76.48 ;
    RECT 35.15 75.69 35.36 75.76 ;
    RECT 35.15 76.05 35.36 76.12 ;
    RECT 35.15 76.41 35.36 76.48 ;
    RECT 117.69 75.69 117.9 75.76 ;
    RECT 117.69 76.05 117.9 76.12 ;
    RECT 117.69 76.41 117.9 76.48 ;
    RECT 118.15 75.69 118.36 75.76 ;
    RECT 118.15 76.05 118.36 76.12 ;
    RECT 118.15 76.41 118.36 76.48 ;
    RECT 114.37 75.69 114.58 75.76 ;
    RECT 114.37 76.05 114.58 76.12 ;
    RECT 114.37 76.41 114.58 76.48 ;
    RECT 114.83 75.69 115.04 75.76 ;
    RECT 114.83 76.05 115.04 76.12 ;
    RECT 114.83 76.41 115.04 76.48 ;
    RECT 111.05 75.69 111.26 75.76 ;
    RECT 111.05 76.05 111.26 76.12 ;
    RECT 111.05 76.41 111.26 76.48 ;
    RECT 111.51 75.69 111.72 75.76 ;
    RECT 111.51 76.05 111.72 76.12 ;
    RECT 111.51 76.41 111.72 76.48 ;
    RECT 107.73 75.69 107.94 75.76 ;
    RECT 107.73 76.05 107.94 76.12 ;
    RECT 107.73 76.41 107.94 76.48 ;
    RECT 108.19 75.69 108.4 75.76 ;
    RECT 108.19 76.05 108.4 76.12 ;
    RECT 108.19 76.41 108.4 76.48 ;
    RECT 104.41 75.69 104.62 75.76 ;
    RECT 104.41 76.05 104.62 76.12 ;
    RECT 104.41 76.41 104.62 76.48 ;
    RECT 104.87 75.69 105.08 75.76 ;
    RECT 104.87 76.05 105.08 76.12 ;
    RECT 104.87 76.41 105.08 76.48 ;
    RECT 101.09 75.69 101.3 75.76 ;
    RECT 101.09 76.05 101.3 76.12 ;
    RECT 101.09 76.41 101.3 76.48 ;
    RECT 101.55 75.69 101.76 75.76 ;
    RECT 101.55 76.05 101.76 76.12 ;
    RECT 101.55 76.41 101.76 76.48 ;
    RECT 97.77 75.69 97.98 75.76 ;
    RECT 97.77 76.05 97.98 76.12 ;
    RECT 97.77 76.41 97.98 76.48 ;
    RECT 98.23 75.69 98.44 75.76 ;
    RECT 98.23 76.05 98.44 76.12 ;
    RECT 98.23 76.41 98.44 76.48 ;
    RECT 94.45 75.69 94.66 75.76 ;
    RECT 94.45 76.05 94.66 76.12 ;
    RECT 94.45 76.41 94.66 76.48 ;
    RECT 94.91 75.69 95.12 75.76 ;
    RECT 94.91 76.05 95.12 76.12 ;
    RECT 94.91 76.41 95.12 76.48 ;
    RECT 91.13 75.69 91.34 75.76 ;
    RECT 91.13 76.05 91.34 76.12 ;
    RECT 91.13 76.41 91.34 76.48 ;
    RECT 91.59 75.69 91.8 75.76 ;
    RECT 91.59 76.05 91.8 76.12 ;
    RECT 91.59 76.41 91.8 76.48 ;
    RECT 87.81 75.69 88.02 75.76 ;
    RECT 87.81 76.05 88.02 76.12 ;
    RECT 87.81 76.41 88.02 76.48 ;
    RECT 88.27 75.69 88.48 75.76 ;
    RECT 88.27 76.05 88.48 76.12 ;
    RECT 88.27 76.41 88.48 76.48 ;
    RECT 84.49 75.69 84.7 75.76 ;
    RECT 84.49 76.05 84.7 76.12 ;
    RECT 84.49 76.41 84.7 76.48 ;
    RECT 84.95 75.69 85.16 75.76 ;
    RECT 84.95 76.05 85.16 76.12 ;
    RECT 84.95 76.41 85.16 76.48 ;
    RECT 81.17 75.69 81.38 75.76 ;
    RECT 81.17 76.05 81.38 76.12 ;
    RECT 81.17 76.41 81.38 76.48 ;
    RECT 81.63 75.69 81.84 75.76 ;
    RECT 81.63 76.05 81.84 76.12 ;
    RECT 81.63 76.41 81.84 76.48 ;
    RECT 77.85 75.69 78.06 75.76 ;
    RECT 77.85 76.05 78.06 76.12 ;
    RECT 77.85 76.41 78.06 76.48 ;
    RECT 78.31 75.69 78.52 75.76 ;
    RECT 78.31 76.05 78.52 76.12 ;
    RECT 78.31 76.41 78.52 76.48 ;
    RECT 74.53 75.69 74.74 75.76 ;
    RECT 74.53 76.05 74.74 76.12 ;
    RECT 74.53 76.41 74.74 76.48 ;
    RECT 74.99 75.69 75.2 75.76 ;
    RECT 74.99 76.05 75.2 76.12 ;
    RECT 74.99 76.41 75.2 76.48 ;
    RECT 71.21 75.69 71.42 75.76 ;
    RECT 71.21 76.05 71.42 76.12 ;
    RECT 71.21 76.41 71.42 76.48 ;
    RECT 71.67 75.69 71.88 75.76 ;
    RECT 71.67 76.05 71.88 76.12 ;
    RECT 71.67 76.41 71.88 76.48 ;
    RECT 31.37 75.69 31.58 75.76 ;
    RECT 31.37 76.05 31.58 76.12 ;
    RECT 31.37 76.41 31.58 76.48 ;
    RECT 31.83 75.69 32.04 75.76 ;
    RECT 31.83 76.05 32.04 76.12 ;
    RECT 31.83 76.41 32.04 76.48 ;
    RECT 67.89 75.69 68.1 75.76 ;
    RECT 67.89 76.05 68.1 76.12 ;
    RECT 67.89 76.41 68.1 76.48 ;
    RECT 68.35 75.69 68.56 75.76 ;
    RECT 68.35 76.05 68.56 76.12 ;
    RECT 68.35 76.41 68.56 76.48 ;
    RECT 28.05 75.69 28.26 75.76 ;
    RECT 28.05 76.05 28.26 76.12 ;
    RECT 28.05 76.41 28.26 76.48 ;
    RECT 28.51 75.69 28.72 75.76 ;
    RECT 28.51 76.05 28.72 76.12 ;
    RECT 28.51 76.41 28.72 76.48 ;
    RECT 24.73 75.69 24.94 75.76 ;
    RECT 24.73 76.05 24.94 76.12 ;
    RECT 24.73 76.41 24.94 76.48 ;
    RECT 25.19 75.69 25.4 75.76 ;
    RECT 25.19 76.05 25.4 76.12 ;
    RECT 25.19 76.41 25.4 76.48 ;
    RECT 21.41 75.69 21.62 75.76 ;
    RECT 21.41 76.05 21.62 76.12 ;
    RECT 21.41 76.41 21.62 76.48 ;
    RECT 21.87 75.69 22.08 75.76 ;
    RECT 21.87 76.05 22.08 76.12 ;
    RECT 21.87 76.41 22.08 76.48 ;
    RECT 18.09 75.69 18.3 75.76 ;
    RECT 18.09 76.05 18.3 76.12 ;
    RECT 18.09 76.41 18.3 76.48 ;
    RECT 18.55 75.69 18.76 75.76 ;
    RECT 18.55 76.05 18.76 76.12 ;
    RECT 18.55 76.41 18.76 76.48 ;
    RECT 120.825 76.05 120.895 76.12 ;
    RECT 14.77 75.69 14.98 75.76 ;
    RECT 14.77 76.05 14.98 76.12 ;
    RECT 14.77 76.41 14.98 76.48 ;
    RECT 15.23 75.69 15.44 75.76 ;
    RECT 15.23 76.05 15.44 76.12 ;
    RECT 15.23 76.41 15.44 76.48 ;
    RECT 11.45 75.69 11.66 75.76 ;
    RECT 11.45 76.05 11.66 76.12 ;
    RECT 11.45 76.41 11.66 76.48 ;
    RECT 11.91 75.69 12.12 75.76 ;
    RECT 11.91 76.05 12.12 76.12 ;
    RECT 11.91 76.41 12.12 76.48 ;
    RECT 8.13 75.69 8.34 75.76 ;
    RECT 8.13 76.05 8.34 76.12 ;
    RECT 8.13 76.41 8.34 76.48 ;
    RECT 8.59 75.69 8.8 75.76 ;
    RECT 8.59 76.05 8.8 76.12 ;
    RECT 8.59 76.41 8.8 76.48 ;
    RECT 4.81 75.69 5.02 75.76 ;
    RECT 4.81 76.05 5.02 76.12 ;
    RECT 4.81 76.41 5.02 76.48 ;
    RECT 5.27 75.69 5.48 75.76 ;
    RECT 5.27 76.05 5.48 76.12 ;
    RECT 5.27 76.41 5.48 76.48 ;
    RECT 1.49 75.69 1.7 75.76 ;
    RECT 1.49 76.05 1.7 76.12 ;
    RECT 1.49 76.41 1.7 76.48 ;
    RECT 1.95 75.69 2.16 75.76 ;
    RECT 1.95 76.05 2.16 76.12 ;
    RECT 1.95 76.41 2.16 76.48 ;
    RECT 64.57 75.69 64.78 75.76 ;
    RECT 64.57 76.05 64.78 76.12 ;
    RECT 64.57 76.41 64.78 76.48 ;
    RECT 65.03 75.69 65.24 75.76 ;
    RECT 65.03 76.05 65.24 76.12 ;
    RECT 65.03 76.41 65.24 76.48 ;
    RECT 61.25 74.97 61.46 75.04 ;
    RECT 61.25 75.33 61.46 75.4 ;
    RECT 61.25 75.69 61.46 75.76 ;
    RECT 61.71 74.97 61.92 75.04 ;
    RECT 61.71 75.33 61.92 75.4 ;
    RECT 61.71 75.69 61.92 75.76 ;
    RECT 57.93 74.97 58.14 75.04 ;
    RECT 57.93 75.33 58.14 75.4 ;
    RECT 57.93 75.69 58.14 75.76 ;
    RECT 58.39 74.97 58.6 75.04 ;
    RECT 58.39 75.33 58.6 75.4 ;
    RECT 58.39 75.69 58.6 75.76 ;
    RECT 54.61 74.97 54.82 75.04 ;
    RECT 54.61 75.33 54.82 75.4 ;
    RECT 54.61 75.69 54.82 75.76 ;
    RECT 55.07 74.97 55.28 75.04 ;
    RECT 55.07 75.33 55.28 75.4 ;
    RECT 55.07 75.69 55.28 75.76 ;
    RECT 51.29 74.97 51.5 75.04 ;
    RECT 51.29 75.33 51.5 75.4 ;
    RECT 51.29 75.69 51.5 75.76 ;
    RECT 51.75 74.97 51.96 75.04 ;
    RECT 51.75 75.33 51.96 75.4 ;
    RECT 51.75 75.69 51.96 75.76 ;
    RECT 47.97 74.97 48.18 75.04 ;
    RECT 47.97 75.33 48.18 75.4 ;
    RECT 47.97 75.69 48.18 75.76 ;
    RECT 48.43 74.97 48.64 75.04 ;
    RECT 48.43 75.33 48.64 75.4 ;
    RECT 48.43 75.69 48.64 75.76 ;
    RECT 44.65 74.97 44.86 75.04 ;
    RECT 44.65 75.33 44.86 75.4 ;
    RECT 44.65 75.69 44.86 75.76 ;
    RECT 45.11 74.97 45.32 75.04 ;
    RECT 45.11 75.33 45.32 75.4 ;
    RECT 45.11 75.69 45.32 75.76 ;
    RECT 41.33 74.97 41.54 75.04 ;
    RECT 41.33 75.33 41.54 75.4 ;
    RECT 41.33 75.69 41.54 75.76 ;
    RECT 41.79 74.97 42.0 75.04 ;
    RECT 41.79 75.33 42.0 75.4 ;
    RECT 41.79 75.69 42.0 75.76 ;
    RECT 38.01 74.97 38.22 75.04 ;
    RECT 38.01 75.33 38.22 75.4 ;
    RECT 38.01 75.69 38.22 75.76 ;
    RECT 38.47 74.97 38.68 75.04 ;
    RECT 38.47 75.33 38.68 75.4 ;
    RECT 38.47 75.69 38.68 75.76 ;
    RECT 0.4 75.33 0.47 75.4 ;
    RECT 34.69 74.97 34.9 75.04 ;
    RECT 34.69 75.33 34.9 75.4 ;
    RECT 34.69 75.69 34.9 75.76 ;
    RECT 35.15 74.97 35.36 75.04 ;
    RECT 35.15 75.33 35.36 75.4 ;
    RECT 35.15 75.69 35.36 75.76 ;
    RECT 117.69 74.97 117.9 75.04 ;
    RECT 117.69 75.33 117.9 75.4 ;
    RECT 117.69 75.69 117.9 75.76 ;
    RECT 118.15 74.97 118.36 75.04 ;
    RECT 118.15 75.33 118.36 75.4 ;
    RECT 118.15 75.69 118.36 75.76 ;
    RECT 114.37 74.97 114.58 75.04 ;
    RECT 114.37 75.33 114.58 75.4 ;
    RECT 114.37 75.69 114.58 75.76 ;
    RECT 114.83 74.97 115.04 75.04 ;
    RECT 114.83 75.33 115.04 75.4 ;
    RECT 114.83 75.69 115.04 75.76 ;
    RECT 111.05 74.97 111.26 75.04 ;
    RECT 111.05 75.33 111.26 75.4 ;
    RECT 111.05 75.69 111.26 75.76 ;
    RECT 111.51 74.97 111.72 75.04 ;
    RECT 111.51 75.33 111.72 75.4 ;
    RECT 111.51 75.69 111.72 75.76 ;
    RECT 107.73 74.97 107.94 75.04 ;
    RECT 107.73 75.33 107.94 75.4 ;
    RECT 107.73 75.69 107.94 75.76 ;
    RECT 108.19 74.97 108.4 75.04 ;
    RECT 108.19 75.33 108.4 75.4 ;
    RECT 108.19 75.69 108.4 75.76 ;
    RECT 104.41 74.97 104.62 75.04 ;
    RECT 104.41 75.33 104.62 75.4 ;
    RECT 104.41 75.69 104.62 75.76 ;
    RECT 104.87 74.97 105.08 75.04 ;
    RECT 104.87 75.33 105.08 75.4 ;
    RECT 104.87 75.69 105.08 75.76 ;
    RECT 101.09 74.97 101.3 75.04 ;
    RECT 101.09 75.33 101.3 75.4 ;
    RECT 101.09 75.69 101.3 75.76 ;
    RECT 101.55 74.97 101.76 75.04 ;
    RECT 101.55 75.33 101.76 75.4 ;
    RECT 101.55 75.69 101.76 75.76 ;
    RECT 97.77 74.97 97.98 75.04 ;
    RECT 97.77 75.33 97.98 75.4 ;
    RECT 97.77 75.69 97.98 75.76 ;
    RECT 98.23 74.97 98.44 75.04 ;
    RECT 98.23 75.33 98.44 75.4 ;
    RECT 98.23 75.69 98.44 75.76 ;
    RECT 94.45 74.97 94.66 75.04 ;
    RECT 94.45 75.33 94.66 75.4 ;
    RECT 94.45 75.69 94.66 75.76 ;
    RECT 94.91 74.97 95.12 75.04 ;
    RECT 94.91 75.33 95.12 75.4 ;
    RECT 94.91 75.69 95.12 75.76 ;
    RECT 91.13 74.97 91.34 75.04 ;
    RECT 91.13 75.33 91.34 75.4 ;
    RECT 91.13 75.69 91.34 75.76 ;
    RECT 91.59 74.97 91.8 75.04 ;
    RECT 91.59 75.33 91.8 75.4 ;
    RECT 91.59 75.69 91.8 75.76 ;
    RECT 87.81 74.97 88.02 75.04 ;
    RECT 87.81 75.33 88.02 75.4 ;
    RECT 87.81 75.69 88.02 75.76 ;
    RECT 88.27 74.97 88.48 75.04 ;
    RECT 88.27 75.33 88.48 75.4 ;
    RECT 88.27 75.69 88.48 75.76 ;
    RECT 84.49 74.97 84.7 75.04 ;
    RECT 84.49 75.33 84.7 75.4 ;
    RECT 84.49 75.69 84.7 75.76 ;
    RECT 84.95 74.97 85.16 75.04 ;
    RECT 84.95 75.33 85.16 75.4 ;
    RECT 84.95 75.69 85.16 75.76 ;
    RECT 81.17 74.97 81.38 75.04 ;
    RECT 81.17 75.33 81.38 75.4 ;
    RECT 81.17 75.69 81.38 75.76 ;
    RECT 81.63 74.97 81.84 75.04 ;
    RECT 81.63 75.33 81.84 75.4 ;
    RECT 81.63 75.69 81.84 75.76 ;
    RECT 77.85 74.97 78.06 75.04 ;
    RECT 77.85 75.33 78.06 75.4 ;
    RECT 77.85 75.69 78.06 75.76 ;
    RECT 78.31 74.97 78.52 75.04 ;
    RECT 78.31 75.33 78.52 75.4 ;
    RECT 78.31 75.69 78.52 75.76 ;
    RECT 74.53 74.97 74.74 75.04 ;
    RECT 74.53 75.33 74.74 75.4 ;
    RECT 74.53 75.69 74.74 75.76 ;
    RECT 74.99 74.97 75.2 75.04 ;
    RECT 74.99 75.33 75.2 75.4 ;
    RECT 74.99 75.69 75.2 75.76 ;
    RECT 71.21 74.97 71.42 75.04 ;
    RECT 71.21 75.33 71.42 75.4 ;
    RECT 71.21 75.69 71.42 75.76 ;
    RECT 71.67 74.97 71.88 75.04 ;
    RECT 71.67 75.33 71.88 75.4 ;
    RECT 71.67 75.69 71.88 75.76 ;
    RECT 31.37 74.97 31.58 75.04 ;
    RECT 31.37 75.33 31.58 75.4 ;
    RECT 31.37 75.69 31.58 75.76 ;
    RECT 31.83 74.97 32.04 75.04 ;
    RECT 31.83 75.33 32.04 75.4 ;
    RECT 31.83 75.69 32.04 75.76 ;
    RECT 67.89 74.97 68.1 75.04 ;
    RECT 67.89 75.33 68.1 75.4 ;
    RECT 67.89 75.69 68.1 75.76 ;
    RECT 68.35 74.97 68.56 75.04 ;
    RECT 68.35 75.33 68.56 75.4 ;
    RECT 68.35 75.69 68.56 75.76 ;
    RECT 28.05 74.97 28.26 75.04 ;
    RECT 28.05 75.33 28.26 75.4 ;
    RECT 28.05 75.69 28.26 75.76 ;
    RECT 28.51 74.97 28.72 75.04 ;
    RECT 28.51 75.33 28.72 75.4 ;
    RECT 28.51 75.69 28.72 75.76 ;
    RECT 24.73 74.97 24.94 75.04 ;
    RECT 24.73 75.33 24.94 75.4 ;
    RECT 24.73 75.69 24.94 75.76 ;
    RECT 25.19 74.97 25.4 75.04 ;
    RECT 25.19 75.33 25.4 75.4 ;
    RECT 25.19 75.69 25.4 75.76 ;
    RECT 21.41 74.97 21.62 75.04 ;
    RECT 21.41 75.33 21.62 75.4 ;
    RECT 21.41 75.69 21.62 75.76 ;
    RECT 21.87 74.97 22.08 75.04 ;
    RECT 21.87 75.33 22.08 75.4 ;
    RECT 21.87 75.69 22.08 75.76 ;
    RECT 18.09 74.97 18.3 75.04 ;
    RECT 18.09 75.33 18.3 75.4 ;
    RECT 18.09 75.69 18.3 75.76 ;
    RECT 18.55 74.97 18.76 75.04 ;
    RECT 18.55 75.33 18.76 75.4 ;
    RECT 18.55 75.69 18.76 75.76 ;
    RECT 120.825 75.33 120.895 75.4 ;
    RECT 14.77 74.97 14.98 75.04 ;
    RECT 14.77 75.33 14.98 75.4 ;
    RECT 14.77 75.69 14.98 75.76 ;
    RECT 15.23 74.97 15.44 75.04 ;
    RECT 15.23 75.33 15.44 75.4 ;
    RECT 15.23 75.69 15.44 75.76 ;
    RECT 11.45 74.97 11.66 75.04 ;
    RECT 11.45 75.33 11.66 75.4 ;
    RECT 11.45 75.69 11.66 75.76 ;
    RECT 11.91 74.97 12.12 75.04 ;
    RECT 11.91 75.33 12.12 75.4 ;
    RECT 11.91 75.69 12.12 75.76 ;
    RECT 8.13 74.97 8.34 75.04 ;
    RECT 8.13 75.33 8.34 75.4 ;
    RECT 8.13 75.69 8.34 75.76 ;
    RECT 8.59 74.97 8.8 75.04 ;
    RECT 8.59 75.33 8.8 75.4 ;
    RECT 8.59 75.69 8.8 75.76 ;
    RECT 4.81 74.97 5.02 75.04 ;
    RECT 4.81 75.33 5.02 75.4 ;
    RECT 4.81 75.69 5.02 75.76 ;
    RECT 5.27 74.97 5.48 75.04 ;
    RECT 5.27 75.33 5.48 75.4 ;
    RECT 5.27 75.69 5.48 75.76 ;
    RECT 1.49 74.97 1.7 75.04 ;
    RECT 1.49 75.33 1.7 75.4 ;
    RECT 1.49 75.69 1.7 75.76 ;
    RECT 1.95 74.97 2.16 75.04 ;
    RECT 1.95 75.33 2.16 75.4 ;
    RECT 1.95 75.69 2.16 75.76 ;
    RECT 64.57 74.97 64.78 75.04 ;
    RECT 64.57 75.33 64.78 75.4 ;
    RECT 64.57 75.69 64.78 75.76 ;
    RECT 65.03 74.97 65.24 75.04 ;
    RECT 65.03 75.33 65.24 75.4 ;
    RECT 65.03 75.69 65.24 75.76 ;
    RECT 61.25 74.25 61.46 74.32 ;
    RECT 61.25 74.61 61.46 74.68 ;
    RECT 61.25 74.97 61.46 75.04 ;
    RECT 61.71 74.25 61.92 74.32 ;
    RECT 61.71 74.61 61.92 74.68 ;
    RECT 61.71 74.97 61.92 75.04 ;
    RECT 57.93 74.25 58.14 74.32 ;
    RECT 57.93 74.61 58.14 74.68 ;
    RECT 57.93 74.97 58.14 75.04 ;
    RECT 58.39 74.25 58.6 74.32 ;
    RECT 58.39 74.61 58.6 74.68 ;
    RECT 58.39 74.97 58.6 75.04 ;
    RECT 54.61 74.25 54.82 74.32 ;
    RECT 54.61 74.61 54.82 74.68 ;
    RECT 54.61 74.97 54.82 75.04 ;
    RECT 55.07 74.25 55.28 74.32 ;
    RECT 55.07 74.61 55.28 74.68 ;
    RECT 55.07 74.97 55.28 75.04 ;
    RECT 51.29 74.25 51.5 74.32 ;
    RECT 51.29 74.61 51.5 74.68 ;
    RECT 51.29 74.97 51.5 75.04 ;
    RECT 51.75 74.25 51.96 74.32 ;
    RECT 51.75 74.61 51.96 74.68 ;
    RECT 51.75 74.97 51.96 75.04 ;
    RECT 47.97 74.25 48.18 74.32 ;
    RECT 47.97 74.61 48.18 74.68 ;
    RECT 47.97 74.97 48.18 75.04 ;
    RECT 48.43 74.25 48.64 74.32 ;
    RECT 48.43 74.61 48.64 74.68 ;
    RECT 48.43 74.97 48.64 75.04 ;
    RECT 44.65 74.25 44.86 74.32 ;
    RECT 44.65 74.61 44.86 74.68 ;
    RECT 44.65 74.97 44.86 75.04 ;
    RECT 45.11 74.25 45.32 74.32 ;
    RECT 45.11 74.61 45.32 74.68 ;
    RECT 45.11 74.97 45.32 75.04 ;
    RECT 41.33 74.25 41.54 74.32 ;
    RECT 41.33 74.61 41.54 74.68 ;
    RECT 41.33 74.97 41.54 75.04 ;
    RECT 41.79 74.25 42.0 74.32 ;
    RECT 41.79 74.61 42.0 74.68 ;
    RECT 41.79 74.97 42.0 75.04 ;
    RECT 38.01 74.25 38.22 74.32 ;
    RECT 38.01 74.61 38.22 74.68 ;
    RECT 38.01 74.97 38.22 75.04 ;
    RECT 38.47 74.25 38.68 74.32 ;
    RECT 38.47 74.61 38.68 74.68 ;
    RECT 38.47 74.97 38.68 75.04 ;
    RECT 0.4 74.61 0.47 74.68 ;
    RECT 34.69 74.25 34.9 74.32 ;
    RECT 34.69 74.61 34.9 74.68 ;
    RECT 34.69 74.97 34.9 75.04 ;
    RECT 35.15 74.25 35.36 74.32 ;
    RECT 35.15 74.61 35.36 74.68 ;
    RECT 35.15 74.97 35.36 75.04 ;
    RECT 117.69 74.25 117.9 74.32 ;
    RECT 117.69 74.61 117.9 74.68 ;
    RECT 117.69 74.97 117.9 75.04 ;
    RECT 118.15 74.25 118.36 74.32 ;
    RECT 118.15 74.61 118.36 74.68 ;
    RECT 118.15 74.97 118.36 75.04 ;
    RECT 114.37 74.25 114.58 74.32 ;
    RECT 114.37 74.61 114.58 74.68 ;
    RECT 114.37 74.97 114.58 75.04 ;
    RECT 114.83 74.25 115.04 74.32 ;
    RECT 114.83 74.61 115.04 74.68 ;
    RECT 114.83 74.97 115.04 75.04 ;
    RECT 111.05 74.25 111.26 74.32 ;
    RECT 111.05 74.61 111.26 74.68 ;
    RECT 111.05 74.97 111.26 75.04 ;
    RECT 111.51 74.25 111.72 74.32 ;
    RECT 111.51 74.61 111.72 74.68 ;
    RECT 111.51 74.97 111.72 75.04 ;
    RECT 107.73 74.25 107.94 74.32 ;
    RECT 107.73 74.61 107.94 74.68 ;
    RECT 107.73 74.97 107.94 75.04 ;
    RECT 108.19 74.25 108.4 74.32 ;
    RECT 108.19 74.61 108.4 74.68 ;
    RECT 108.19 74.97 108.4 75.04 ;
    RECT 104.41 74.25 104.62 74.32 ;
    RECT 104.41 74.61 104.62 74.68 ;
    RECT 104.41 74.97 104.62 75.04 ;
    RECT 104.87 74.25 105.08 74.32 ;
    RECT 104.87 74.61 105.08 74.68 ;
    RECT 104.87 74.97 105.08 75.04 ;
    RECT 101.09 74.25 101.3 74.32 ;
    RECT 101.09 74.61 101.3 74.68 ;
    RECT 101.09 74.97 101.3 75.04 ;
    RECT 101.55 74.25 101.76 74.32 ;
    RECT 101.55 74.61 101.76 74.68 ;
    RECT 101.55 74.97 101.76 75.04 ;
    RECT 97.77 74.25 97.98 74.32 ;
    RECT 97.77 74.61 97.98 74.68 ;
    RECT 97.77 74.97 97.98 75.04 ;
    RECT 98.23 74.25 98.44 74.32 ;
    RECT 98.23 74.61 98.44 74.68 ;
    RECT 98.23 74.97 98.44 75.04 ;
    RECT 94.45 74.25 94.66 74.32 ;
    RECT 94.45 74.61 94.66 74.68 ;
    RECT 94.45 74.97 94.66 75.04 ;
    RECT 94.91 74.25 95.12 74.32 ;
    RECT 94.91 74.61 95.12 74.68 ;
    RECT 94.91 74.97 95.12 75.04 ;
    RECT 91.13 74.25 91.34 74.32 ;
    RECT 91.13 74.61 91.34 74.68 ;
    RECT 91.13 74.97 91.34 75.04 ;
    RECT 91.59 74.25 91.8 74.32 ;
    RECT 91.59 74.61 91.8 74.68 ;
    RECT 91.59 74.97 91.8 75.04 ;
    RECT 87.81 74.25 88.02 74.32 ;
    RECT 87.81 74.61 88.02 74.68 ;
    RECT 87.81 74.97 88.02 75.04 ;
    RECT 88.27 74.25 88.48 74.32 ;
    RECT 88.27 74.61 88.48 74.68 ;
    RECT 88.27 74.97 88.48 75.04 ;
    RECT 84.49 74.25 84.7 74.32 ;
    RECT 84.49 74.61 84.7 74.68 ;
    RECT 84.49 74.97 84.7 75.04 ;
    RECT 84.95 74.25 85.16 74.32 ;
    RECT 84.95 74.61 85.16 74.68 ;
    RECT 84.95 74.97 85.16 75.04 ;
    RECT 81.17 74.25 81.38 74.32 ;
    RECT 81.17 74.61 81.38 74.68 ;
    RECT 81.17 74.97 81.38 75.04 ;
    RECT 81.63 74.25 81.84 74.32 ;
    RECT 81.63 74.61 81.84 74.68 ;
    RECT 81.63 74.97 81.84 75.04 ;
    RECT 77.85 74.25 78.06 74.32 ;
    RECT 77.85 74.61 78.06 74.68 ;
    RECT 77.85 74.97 78.06 75.04 ;
    RECT 78.31 74.25 78.52 74.32 ;
    RECT 78.31 74.61 78.52 74.68 ;
    RECT 78.31 74.97 78.52 75.04 ;
    RECT 74.53 74.25 74.74 74.32 ;
    RECT 74.53 74.61 74.74 74.68 ;
    RECT 74.53 74.97 74.74 75.04 ;
    RECT 74.99 74.25 75.2 74.32 ;
    RECT 74.99 74.61 75.2 74.68 ;
    RECT 74.99 74.97 75.2 75.04 ;
    RECT 71.21 74.25 71.42 74.32 ;
    RECT 71.21 74.61 71.42 74.68 ;
    RECT 71.21 74.97 71.42 75.04 ;
    RECT 71.67 74.25 71.88 74.32 ;
    RECT 71.67 74.61 71.88 74.68 ;
    RECT 71.67 74.97 71.88 75.04 ;
    RECT 31.37 74.25 31.58 74.32 ;
    RECT 31.37 74.61 31.58 74.68 ;
    RECT 31.37 74.97 31.58 75.04 ;
    RECT 31.83 74.25 32.04 74.32 ;
    RECT 31.83 74.61 32.04 74.68 ;
    RECT 31.83 74.97 32.04 75.04 ;
    RECT 67.89 74.25 68.1 74.32 ;
    RECT 67.89 74.61 68.1 74.68 ;
    RECT 67.89 74.97 68.1 75.04 ;
    RECT 68.35 74.25 68.56 74.32 ;
    RECT 68.35 74.61 68.56 74.68 ;
    RECT 68.35 74.97 68.56 75.04 ;
    RECT 28.05 74.25 28.26 74.32 ;
    RECT 28.05 74.61 28.26 74.68 ;
    RECT 28.05 74.97 28.26 75.04 ;
    RECT 28.51 74.25 28.72 74.32 ;
    RECT 28.51 74.61 28.72 74.68 ;
    RECT 28.51 74.97 28.72 75.04 ;
    RECT 24.73 74.25 24.94 74.32 ;
    RECT 24.73 74.61 24.94 74.68 ;
    RECT 24.73 74.97 24.94 75.04 ;
    RECT 25.19 74.25 25.4 74.32 ;
    RECT 25.19 74.61 25.4 74.68 ;
    RECT 25.19 74.97 25.4 75.04 ;
    RECT 21.41 74.25 21.62 74.32 ;
    RECT 21.41 74.61 21.62 74.68 ;
    RECT 21.41 74.97 21.62 75.04 ;
    RECT 21.87 74.25 22.08 74.32 ;
    RECT 21.87 74.61 22.08 74.68 ;
    RECT 21.87 74.97 22.08 75.04 ;
    RECT 18.09 74.25 18.3 74.32 ;
    RECT 18.09 74.61 18.3 74.68 ;
    RECT 18.09 74.97 18.3 75.04 ;
    RECT 18.55 74.25 18.76 74.32 ;
    RECT 18.55 74.61 18.76 74.68 ;
    RECT 18.55 74.97 18.76 75.04 ;
    RECT 120.825 74.61 120.895 74.68 ;
    RECT 14.77 74.25 14.98 74.32 ;
    RECT 14.77 74.61 14.98 74.68 ;
    RECT 14.77 74.97 14.98 75.04 ;
    RECT 15.23 74.25 15.44 74.32 ;
    RECT 15.23 74.61 15.44 74.68 ;
    RECT 15.23 74.97 15.44 75.04 ;
    RECT 11.45 74.25 11.66 74.32 ;
    RECT 11.45 74.61 11.66 74.68 ;
    RECT 11.45 74.97 11.66 75.04 ;
    RECT 11.91 74.25 12.12 74.32 ;
    RECT 11.91 74.61 12.12 74.68 ;
    RECT 11.91 74.97 12.12 75.04 ;
    RECT 8.13 74.25 8.34 74.32 ;
    RECT 8.13 74.61 8.34 74.68 ;
    RECT 8.13 74.97 8.34 75.04 ;
    RECT 8.59 74.25 8.8 74.32 ;
    RECT 8.59 74.61 8.8 74.68 ;
    RECT 8.59 74.97 8.8 75.04 ;
    RECT 4.81 74.25 5.02 74.32 ;
    RECT 4.81 74.61 5.02 74.68 ;
    RECT 4.81 74.97 5.02 75.04 ;
    RECT 5.27 74.25 5.48 74.32 ;
    RECT 5.27 74.61 5.48 74.68 ;
    RECT 5.27 74.97 5.48 75.04 ;
    RECT 1.49 74.25 1.7 74.32 ;
    RECT 1.49 74.61 1.7 74.68 ;
    RECT 1.49 74.97 1.7 75.04 ;
    RECT 1.95 74.25 2.16 74.32 ;
    RECT 1.95 74.61 2.16 74.68 ;
    RECT 1.95 74.97 2.16 75.04 ;
    RECT 64.57 74.25 64.78 74.32 ;
    RECT 64.57 74.61 64.78 74.68 ;
    RECT 64.57 74.97 64.78 75.04 ;
    RECT 65.03 74.25 65.24 74.32 ;
    RECT 65.03 74.61 65.24 74.68 ;
    RECT 65.03 74.97 65.24 75.04 ;
    RECT 61.25 73.53 61.46 73.6 ;
    RECT 61.25 73.89 61.46 73.96 ;
    RECT 61.25 74.25 61.46 74.32 ;
    RECT 61.71 73.53 61.92 73.6 ;
    RECT 61.71 73.89 61.92 73.96 ;
    RECT 61.71 74.25 61.92 74.32 ;
    RECT 57.93 73.53 58.14 73.6 ;
    RECT 57.93 73.89 58.14 73.96 ;
    RECT 57.93 74.25 58.14 74.32 ;
    RECT 58.39 73.53 58.6 73.6 ;
    RECT 58.39 73.89 58.6 73.96 ;
    RECT 58.39 74.25 58.6 74.32 ;
    RECT 54.61 73.53 54.82 73.6 ;
    RECT 54.61 73.89 54.82 73.96 ;
    RECT 54.61 74.25 54.82 74.32 ;
    RECT 55.07 73.53 55.28 73.6 ;
    RECT 55.07 73.89 55.28 73.96 ;
    RECT 55.07 74.25 55.28 74.32 ;
    RECT 51.29 73.53 51.5 73.6 ;
    RECT 51.29 73.89 51.5 73.96 ;
    RECT 51.29 74.25 51.5 74.32 ;
    RECT 51.75 73.53 51.96 73.6 ;
    RECT 51.75 73.89 51.96 73.96 ;
    RECT 51.75 74.25 51.96 74.32 ;
    RECT 47.97 73.53 48.18 73.6 ;
    RECT 47.97 73.89 48.18 73.96 ;
    RECT 47.97 74.25 48.18 74.32 ;
    RECT 48.43 73.53 48.64 73.6 ;
    RECT 48.43 73.89 48.64 73.96 ;
    RECT 48.43 74.25 48.64 74.32 ;
    RECT 44.65 73.53 44.86 73.6 ;
    RECT 44.65 73.89 44.86 73.96 ;
    RECT 44.65 74.25 44.86 74.32 ;
    RECT 45.11 73.53 45.32 73.6 ;
    RECT 45.11 73.89 45.32 73.96 ;
    RECT 45.11 74.25 45.32 74.32 ;
    RECT 41.33 73.53 41.54 73.6 ;
    RECT 41.33 73.89 41.54 73.96 ;
    RECT 41.33 74.25 41.54 74.32 ;
    RECT 41.79 73.53 42.0 73.6 ;
    RECT 41.79 73.89 42.0 73.96 ;
    RECT 41.79 74.25 42.0 74.32 ;
    RECT 38.01 73.53 38.22 73.6 ;
    RECT 38.01 73.89 38.22 73.96 ;
    RECT 38.01 74.25 38.22 74.32 ;
    RECT 38.47 73.53 38.68 73.6 ;
    RECT 38.47 73.89 38.68 73.96 ;
    RECT 38.47 74.25 38.68 74.32 ;
    RECT 0.4 73.89 0.47 73.96 ;
    RECT 34.69 73.53 34.9 73.6 ;
    RECT 34.69 73.89 34.9 73.96 ;
    RECT 34.69 74.25 34.9 74.32 ;
    RECT 35.15 73.53 35.36 73.6 ;
    RECT 35.15 73.89 35.36 73.96 ;
    RECT 35.15 74.25 35.36 74.32 ;
    RECT 117.69 73.53 117.9 73.6 ;
    RECT 117.69 73.89 117.9 73.96 ;
    RECT 117.69 74.25 117.9 74.32 ;
    RECT 118.15 73.53 118.36 73.6 ;
    RECT 118.15 73.89 118.36 73.96 ;
    RECT 118.15 74.25 118.36 74.32 ;
    RECT 114.37 73.53 114.58 73.6 ;
    RECT 114.37 73.89 114.58 73.96 ;
    RECT 114.37 74.25 114.58 74.32 ;
    RECT 114.83 73.53 115.04 73.6 ;
    RECT 114.83 73.89 115.04 73.96 ;
    RECT 114.83 74.25 115.04 74.32 ;
    RECT 111.05 73.53 111.26 73.6 ;
    RECT 111.05 73.89 111.26 73.96 ;
    RECT 111.05 74.25 111.26 74.32 ;
    RECT 111.51 73.53 111.72 73.6 ;
    RECT 111.51 73.89 111.72 73.96 ;
    RECT 111.51 74.25 111.72 74.32 ;
    RECT 107.73 73.53 107.94 73.6 ;
    RECT 107.73 73.89 107.94 73.96 ;
    RECT 107.73 74.25 107.94 74.32 ;
    RECT 108.19 73.53 108.4 73.6 ;
    RECT 108.19 73.89 108.4 73.96 ;
    RECT 108.19 74.25 108.4 74.32 ;
    RECT 104.41 73.53 104.62 73.6 ;
    RECT 104.41 73.89 104.62 73.96 ;
    RECT 104.41 74.25 104.62 74.32 ;
    RECT 104.87 73.53 105.08 73.6 ;
    RECT 104.87 73.89 105.08 73.96 ;
    RECT 104.87 74.25 105.08 74.32 ;
    RECT 101.09 73.53 101.3 73.6 ;
    RECT 101.09 73.89 101.3 73.96 ;
    RECT 101.09 74.25 101.3 74.32 ;
    RECT 101.55 73.53 101.76 73.6 ;
    RECT 101.55 73.89 101.76 73.96 ;
    RECT 101.55 74.25 101.76 74.32 ;
    RECT 97.77 73.53 97.98 73.6 ;
    RECT 97.77 73.89 97.98 73.96 ;
    RECT 97.77 74.25 97.98 74.32 ;
    RECT 98.23 73.53 98.44 73.6 ;
    RECT 98.23 73.89 98.44 73.96 ;
    RECT 98.23 74.25 98.44 74.32 ;
    RECT 94.45 73.53 94.66 73.6 ;
    RECT 94.45 73.89 94.66 73.96 ;
    RECT 94.45 74.25 94.66 74.32 ;
    RECT 94.91 73.53 95.12 73.6 ;
    RECT 94.91 73.89 95.12 73.96 ;
    RECT 94.91 74.25 95.12 74.32 ;
    RECT 91.13 73.53 91.34 73.6 ;
    RECT 91.13 73.89 91.34 73.96 ;
    RECT 91.13 74.25 91.34 74.32 ;
    RECT 91.59 73.53 91.8 73.6 ;
    RECT 91.59 73.89 91.8 73.96 ;
    RECT 91.59 74.25 91.8 74.32 ;
    RECT 87.81 73.53 88.02 73.6 ;
    RECT 87.81 73.89 88.02 73.96 ;
    RECT 87.81 74.25 88.02 74.32 ;
    RECT 88.27 73.53 88.48 73.6 ;
    RECT 88.27 73.89 88.48 73.96 ;
    RECT 88.27 74.25 88.48 74.32 ;
    RECT 84.49 73.53 84.7 73.6 ;
    RECT 84.49 73.89 84.7 73.96 ;
    RECT 84.49 74.25 84.7 74.32 ;
    RECT 84.95 73.53 85.16 73.6 ;
    RECT 84.95 73.89 85.16 73.96 ;
    RECT 84.95 74.25 85.16 74.32 ;
    RECT 81.17 73.53 81.38 73.6 ;
    RECT 81.17 73.89 81.38 73.96 ;
    RECT 81.17 74.25 81.38 74.32 ;
    RECT 81.63 73.53 81.84 73.6 ;
    RECT 81.63 73.89 81.84 73.96 ;
    RECT 81.63 74.25 81.84 74.32 ;
    RECT 77.85 73.53 78.06 73.6 ;
    RECT 77.85 73.89 78.06 73.96 ;
    RECT 77.85 74.25 78.06 74.32 ;
    RECT 78.31 73.53 78.52 73.6 ;
    RECT 78.31 73.89 78.52 73.96 ;
    RECT 78.31 74.25 78.52 74.32 ;
    RECT 74.53 73.53 74.74 73.6 ;
    RECT 74.53 73.89 74.74 73.96 ;
    RECT 74.53 74.25 74.74 74.32 ;
    RECT 74.99 73.53 75.2 73.6 ;
    RECT 74.99 73.89 75.2 73.96 ;
    RECT 74.99 74.25 75.2 74.32 ;
    RECT 71.21 73.53 71.42 73.6 ;
    RECT 71.21 73.89 71.42 73.96 ;
    RECT 71.21 74.25 71.42 74.32 ;
    RECT 71.67 73.53 71.88 73.6 ;
    RECT 71.67 73.89 71.88 73.96 ;
    RECT 71.67 74.25 71.88 74.32 ;
    RECT 31.37 73.53 31.58 73.6 ;
    RECT 31.37 73.89 31.58 73.96 ;
    RECT 31.37 74.25 31.58 74.32 ;
    RECT 31.83 73.53 32.04 73.6 ;
    RECT 31.83 73.89 32.04 73.96 ;
    RECT 31.83 74.25 32.04 74.32 ;
    RECT 67.89 73.53 68.1 73.6 ;
    RECT 67.89 73.89 68.1 73.96 ;
    RECT 67.89 74.25 68.1 74.32 ;
    RECT 68.35 73.53 68.56 73.6 ;
    RECT 68.35 73.89 68.56 73.96 ;
    RECT 68.35 74.25 68.56 74.32 ;
    RECT 28.05 73.53 28.26 73.6 ;
    RECT 28.05 73.89 28.26 73.96 ;
    RECT 28.05 74.25 28.26 74.32 ;
    RECT 28.51 73.53 28.72 73.6 ;
    RECT 28.51 73.89 28.72 73.96 ;
    RECT 28.51 74.25 28.72 74.32 ;
    RECT 24.73 73.53 24.94 73.6 ;
    RECT 24.73 73.89 24.94 73.96 ;
    RECT 24.73 74.25 24.94 74.32 ;
    RECT 25.19 73.53 25.4 73.6 ;
    RECT 25.19 73.89 25.4 73.96 ;
    RECT 25.19 74.25 25.4 74.32 ;
    RECT 21.41 73.53 21.62 73.6 ;
    RECT 21.41 73.89 21.62 73.96 ;
    RECT 21.41 74.25 21.62 74.32 ;
    RECT 21.87 73.53 22.08 73.6 ;
    RECT 21.87 73.89 22.08 73.96 ;
    RECT 21.87 74.25 22.08 74.32 ;
    RECT 18.09 73.53 18.3 73.6 ;
    RECT 18.09 73.89 18.3 73.96 ;
    RECT 18.09 74.25 18.3 74.32 ;
    RECT 18.55 73.53 18.76 73.6 ;
    RECT 18.55 73.89 18.76 73.96 ;
    RECT 18.55 74.25 18.76 74.32 ;
    RECT 120.825 73.89 120.895 73.96 ;
    RECT 14.77 73.53 14.98 73.6 ;
    RECT 14.77 73.89 14.98 73.96 ;
    RECT 14.77 74.25 14.98 74.32 ;
    RECT 15.23 73.53 15.44 73.6 ;
    RECT 15.23 73.89 15.44 73.96 ;
    RECT 15.23 74.25 15.44 74.32 ;
    RECT 11.45 73.53 11.66 73.6 ;
    RECT 11.45 73.89 11.66 73.96 ;
    RECT 11.45 74.25 11.66 74.32 ;
    RECT 11.91 73.53 12.12 73.6 ;
    RECT 11.91 73.89 12.12 73.96 ;
    RECT 11.91 74.25 12.12 74.32 ;
    RECT 8.13 73.53 8.34 73.6 ;
    RECT 8.13 73.89 8.34 73.96 ;
    RECT 8.13 74.25 8.34 74.32 ;
    RECT 8.59 73.53 8.8 73.6 ;
    RECT 8.59 73.89 8.8 73.96 ;
    RECT 8.59 74.25 8.8 74.32 ;
    RECT 4.81 73.53 5.02 73.6 ;
    RECT 4.81 73.89 5.02 73.96 ;
    RECT 4.81 74.25 5.02 74.32 ;
    RECT 5.27 73.53 5.48 73.6 ;
    RECT 5.27 73.89 5.48 73.96 ;
    RECT 5.27 74.25 5.48 74.32 ;
    RECT 1.49 73.53 1.7 73.6 ;
    RECT 1.49 73.89 1.7 73.96 ;
    RECT 1.49 74.25 1.7 74.32 ;
    RECT 1.95 73.53 2.16 73.6 ;
    RECT 1.95 73.89 2.16 73.96 ;
    RECT 1.95 74.25 2.16 74.32 ;
    RECT 64.57 73.53 64.78 73.6 ;
    RECT 64.57 73.89 64.78 73.96 ;
    RECT 64.57 74.25 64.78 74.32 ;
    RECT 65.03 73.53 65.24 73.6 ;
    RECT 65.03 73.89 65.24 73.96 ;
    RECT 65.03 74.25 65.24 74.32 ;
    RECT 61.25 72.81 61.46 72.88 ;
    RECT 61.25 73.17 61.46 73.24 ;
    RECT 61.25 73.53 61.46 73.6 ;
    RECT 61.71 72.81 61.92 72.88 ;
    RECT 61.71 73.17 61.92 73.24 ;
    RECT 61.71 73.53 61.92 73.6 ;
    RECT 57.93 72.81 58.14 72.88 ;
    RECT 57.93 73.17 58.14 73.24 ;
    RECT 57.93 73.53 58.14 73.6 ;
    RECT 58.39 72.81 58.6 72.88 ;
    RECT 58.39 73.17 58.6 73.24 ;
    RECT 58.39 73.53 58.6 73.6 ;
    RECT 54.61 72.81 54.82 72.88 ;
    RECT 54.61 73.17 54.82 73.24 ;
    RECT 54.61 73.53 54.82 73.6 ;
    RECT 55.07 72.81 55.28 72.88 ;
    RECT 55.07 73.17 55.28 73.24 ;
    RECT 55.07 73.53 55.28 73.6 ;
    RECT 51.29 72.81 51.5 72.88 ;
    RECT 51.29 73.17 51.5 73.24 ;
    RECT 51.29 73.53 51.5 73.6 ;
    RECT 51.75 72.81 51.96 72.88 ;
    RECT 51.75 73.17 51.96 73.24 ;
    RECT 51.75 73.53 51.96 73.6 ;
    RECT 47.97 72.81 48.18 72.88 ;
    RECT 47.97 73.17 48.18 73.24 ;
    RECT 47.97 73.53 48.18 73.6 ;
    RECT 48.43 72.81 48.64 72.88 ;
    RECT 48.43 73.17 48.64 73.24 ;
    RECT 48.43 73.53 48.64 73.6 ;
    RECT 44.65 72.81 44.86 72.88 ;
    RECT 44.65 73.17 44.86 73.24 ;
    RECT 44.65 73.53 44.86 73.6 ;
    RECT 45.11 72.81 45.32 72.88 ;
    RECT 45.11 73.17 45.32 73.24 ;
    RECT 45.11 73.53 45.32 73.6 ;
    RECT 41.33 72.81 41.54 72.88 ;
    RECT 41.33 73.17 41.54 73.24 ;
    RECT 41.33 73.53 41.54 73.6 ;
    RECT 41.79 72.81 42.0 72.88 ;
    RECT 41.79 73.17 42.0 73.24 ;
    RECT 41.79 73.53 42.0 73.6 ;
    RECT 38.01 72.81 38.22 72.88 ;
    RECT 38.01 73.17 38.22 73.24 ;
    RECT 38.01 73.53 38.22 73.6 ;
    RECT 38.47 72.81 38.68 72.88 ;
    RECT 38.47 73.17 38.68 73.24 ;
    RECT 38.47 73.53 38.68 73.6 ;
    RECT 0.4 73.17 0.47 73.24 ;
    RECT 34.69 72.81 34.9 72.88 ;
    RECT 34.69 73.17 34.9 73.24 ;
    RECT 34.69 73.53 34.9 73.6 ;
    RECT 35.15 72.81 35.36 72.88 ;
    RECT 35.15 73.17 35.36 73.24 ;
    RECT 35.15 73.53 35.36 73.6 ;
    RECT 117.69 72.81 117.9 72.88 ;
    RECT 117.69 73.17 117.9 73.24 ;
    RECT 117.69 73.53 117.9 73.6 ;
    RECT 118.15 72.81 118.36 72.88 ;
    RECT 118.15 73.17 118.36 73.24 ;
    RECT 118.15 73.53 118.36 73.6 ;
    RECT 114.37 72.81 114.58 72.88 ;
    RECT 114.37 73.17 114.58 73.24 ;
    RECT 114.37 73.53 114.58 73.6 ;
    RECT 114.83 72.81 115.04 72.88 ;
    RECT 114.83 73.17 115.04 73.24 ;
    RECT 114.83 73.53 115.04 73.6 ;
    RECT 111.05 72.81 111.26 72.88 ;
    RECT 111.05 73.17 111.26 73.24 ;
    RECT 111.05 73.53 111.26 73.6 ;
    RECT 111.51 72.81 111.72 72.88 ;
    RECT 111.51 73.17 111.72 73.24 ;
    RECT 111.51 73.53 111.72 73.6 ;
    RECT 107.73 72.81 107.94 72.88 ;
    RECT 107.73 73.17 107.94 73.24 ;
    RECT 107.73 73.53 107.94 73.6 ;
    RECT 108.19 72.81 108.4 72.88 ;
    RECT 108.19 73.17 108.4 73.24 ;
    RECT 108.19 73.53 108.4 73.6 ;
    RECT 104.41 72.81 104.62 72.88 ;
    RECT 104.41 73.17 104.62 73.24 ;
    RECT 104.41 73.53 104.62 73.6 ;
    RECT 104.87 72.81 105.08 72.88 ;
    RECT 104.87 73.17 105.08 73.24 ;
    RECT 104.87 73.53 105.08 73.6 ;
    RECT 101.09 72.81 101.3 72.88 ;
    RECT 101.09 73.17 101.3 73.24 ;
    RECT 101.09 73.53 101.3 73.6 ;
    RECT 101.55 72.81 101.76 72.88 ;
    RECT 101.55 73.17 101.76 73.24 ;
    RECT 101.55 73.53 101.76 73.6 ;
    RECT 97.77 72.81 97.98 72.88 ;
    RECT 97.77 73.17 97.98 73.24 ;
    RECT 97.77 73.53 97.98 73.6 ;
    RECT 98.23 72.81 98.44 72.88 ;
    RECT 98.23 73.17 98.44 73.24 ;
    RECT 98.23 73.53 98.44 73.6 ;
    RECT 94.45 72.81 94.66 72.88 ;
    RECT 94.45 73.17 94.66 73.24 ;
    RECT 94.45 73.53 94.66 73.6 ;
    RECT 94.91 72.81 95.12 72.88 ;
    RECT 94.91 73.17 95.12 73.24 ;
    RECT 94.91 73.53 95.12 73.6 ;
    RECT 91.13 72.81 91.34 72.88 ;
    RECT 91.13 73.17 91.34 73.24 ;
    RECT 91.13 73.53 91.34 73.6 ;
    RECT 91.59 72.81 91.8 72.88 ;
    RECT 91.59 73.17 91.8 73.24 ;
    RECT 91.59 73.53 91.8 73.6 ;
    RECT 87.81 72.81 88.02 72.88 ;
    RECT 87.81 73.17 88.02 73.24 ;
    RECT 87.81 73.53 88.02 73.6 ;
    RECT 88.27 72.81 88.48 72.88 ;
    RECT 88.27 73.17 88.48 73.24 ;
    RECT 88.27 73.53 88.48 73.6 ;
    RECT 84.49 72.81 84.7 72.88 ;
    RECT 84.49 73.17 84.7 73.24 ;
    RECT 84.49 73.53 84.7 73.6 ;
    RECT 84.95 72.81 85.16 72.88 ;
    RECT 84.95 73.17 85.16 73.24 ;
    RECT 84.95 73.53 85.16 73.6 ;
    RECT 81.17 72.81 81.38 72.88 ;
    RECT 81.17 73.17 81.38 73.24 ;
    RECT 81.17 73.53 81.38 73.6 ;
    RECT 81.63 72.81 81.84 72.88 ;
    RECT 81.63 73.17 81.84 73.24 ;
    RECT 81.63 73.53 81.84 73.6 ;
    RECT 77.85 72.81 78.06 72.88 ;
    RECT 77.85 73.17 78.06 73.24 ;
    RECT 77.85 73.53 78.06 73.6 ;
    RECT 78.31 72.81 78.52 72.88 ;
    RECT 78.31 73.17 78.52 73.24 ;
    RECT 78.31 73.53 78.52 73.6 ;
    RECT 74.53 72.81 74.74 72.88 ;
    RECT 74.53 73.17 74.74 73.24 ;
    RECT 74.53 73.53 74.74 73.6 ;
    RECT 74.99 72.81 75.2 72.88 ;
    RECT 74.99 73.17 75.2 73.24 ;
    RECT 74.99 73.53 75.2 73.6 ;
    RECT 71.21 72.81 71.42 72.88 ;
    RECT 71.21 73.17 71.42 73.24 ;
    RECT 71.21 73.53 71.42 73.6 ;
    RECT 71.67 72.81 71.88 72.88 ;
    RECT 71.67 73.17 71.88 73.24 ;
    RECT 71.67 73.53 71.88 73.6 ;
    RECT 31.37 72.81 31.58 72.88 ;
    RECT 31.37 73.17 31.58 73.24 ;
    RECT 31.37 73.53 31.58 73.6 ;
    RECT 31.83 72.81 32.04 72.88 ;
    RECT 31.83 73.17 32.04 73.24 ;
    RECT 31.83 73.53 32.04 73.6 ;
    RECT 67.89 72.81 68.1 72.88 ;
    RECT 67.89 73.17 68.1 73.24 ;
    RECT 67.89 73.53 68.1 73.6 ;
    RECT 68.35 72.81 68.56 72.88 ;
    RECT 68.35 73.17 68.56 73.24 ;
    RECT 68.35 73.53 68.56 73.6 ;
    RECT 28.05 72.81 28.26 72.88 ;
    RECT 28.05 73.17 28.26 73.24 ;
    RECT 28.05 73.53 28.26 73.6 ;
    RECT 28.51 72.81 28.72 72.88 ;
    RECT 28.51 73.17 28.72 73.24 ;
    RECT 28.51 73.53 28.72 73.6 ;
    RECT 24.73 72.81 24.94 72.88 ;
    RECT 24.73 73.17 24.94 73.24 ;
    RECT 24.73 73.53 24.94 73.6 ;
    RECT 25.19 72.81 25.4 72.88 ;
    RECT 25.19 73.17 25.4 73.24 ;
    RECT 25.19 73.53 25.4 73.6 ;
    RECT 21.41 72.81 21.62 72.88 ;
    RECT 21.41 73.17 21.62 73.24 ;
    RECT 21.41 73.53 21.62 73.6 ;
    RECT 21.87 72.81 22.08 72.88 ;
    RECT 21.87 73.17 22.08 73.24 ;
    RECT 21.87 73.53 22.08 73.6 ;
    RECT 18.09 72.81 18.3 72.88 ;
    RECT 18.09 73.17 18.3 73.24 ;
    RECT 18.09 73.53 18.3 73.6 ;
    RECT 18.55 72.81 18.76 72.88 ;
    RECT 18.55 73.17 18.76 73.24 ;
    RECT 18.55 73.53 18.76 73.6 ;
    RECT 120.825 73.17 120.895 73.24 ;
    RECT 14.77 72.81 14.98 72.88 ;
    RECT 14.77 73.17 14.98 73.24 ;
    RECT 14.77 73.53 14.98 73.6 ;
    RECT 15.23 72.81 15.44 72.88 ;
    RECT 15.23 73.17 15.44 73.24 ;
    RECT 15.23 73.53 15.44 73.6 ;
    RECT 11.45 72.81 11.66 72.88 ;
    RECT 11.45 73.17 11.66 73.24 ;
    RECT 11.45 73.53 11.66 73.6 ;
    RECT 11.91 72.81 12.12 72.88 ;
    RECT 11.91 73.17 12.12 73.24 ;
    RECT 11.91 73.53 12.12 73.6 ;
    RECT 8.13 72.81 8.34 72.88 ;
    RECT 8.13 73.17 8.34 73.24 ;
    RECT 8.13 73.53 8.34 73.6 ;
    RECT 8.59 72.81 8.8 72.88 ;
    RECT 8.59 73.17 8.8 73.24 ;
    RECT 8.59 73.53 8.8 73.6 ;
    RECT 4.81 72.81 5.02 72.88 ;
    RECT 4.81 73.17 5.02 73.24 ;
    RECT 4.81 73.53 5.02 73.6 ;
    RECT 5.27 72.81 5.48 72.88 ;
    RECT 5.27 73.17 5.48 73.24 ;
    RECT 5.27 73.53 5.48 73.6 ;
    RECT 1.49 72.81 1.7 72.88 ;
    RECT 1.49 73.17 1.7 73.24 ;
    RECT 1.49 73.53 1.7 73.6 ;
    RECT 1.95 72.81 2.16 72.88 ;
    RECT 1.95 73.17 2.16 73.24 ;
    RECT 1.95 73.53 2.16 73.6 ;
    RECT 64.57 72.81 64.78 72.88 ;
    RECT 64.57 73.17 64.78 73.24 ;
    RECT 64.57 73.53 64.78 73.6 ;
    RECT 65.03 72.81 65.24 72.88 ;
    RECT 65.03 73.17 65.24 73.24 ;
    RECT 65.03 73.53 65.24 73.6 ;
    RECT 61.25 35.35 61.46 35.42 ;
    RECT 61.25 35.71 61.46 35.78 ;
    RECT 61.25 36.07 61.46 36.14 ;
    RECT 61.71 35.35 61.92 35.42 ;
    RECT 61.71 35.71 61.92 35.78 ;
    RECT 61.71 36.07 61.92 36.14 ;
    RECT 57.93 35.35 58.14 35.42 ;
    RECT 57.93 35.71 58.14 35.78 ;
    RECT 57.93 36.07 58.14 36.14 ;
    RECT 58.39 35.35 58.6 35.42 ;
    RECT 58.39 35.71 58.6 35.78 ;
    RECT 58.39 36.07 58.6 36.14 ;
    RECT 54.61 35.35 54.82 35.42 ;
    RECT 54.61 35.71 54.82 35.78 ;
    RECT 54.61 36.07 54.82 36.14 ;
    RECT 55.07 35.35 55.28 35.42 ;
    RECT 55.07 35.71 55.28 35.78 ;
    RECT 55.07 36.07 55.28 36.14 ;
    RECT 51.29 35.35 51.5 35.42 ;
    RECT 51.29 35.71 51.5 35.78 ;
    RECT 51.29 36.07 51.5 36.14 ;
    RECT 51.75 35.35 51.96 35.42 ;
    RECT 51.75 35.71 51.96 35.78 ;
    RECT 51.75 36.07 51.96 36.14 ;
    RECT 47.97 35.35 48.18 35.42 ;
    RECT 47.97 35.71 48.18 35.78 ;
    RECT 47.97 36.07 48.18 36.14 ;
    RECT 48.43 35.35 48.64 35.42 ;
    RECT 48.43 35.71 48.64 35.78 ;
    RECT 48.43 36.07 48.64 36.14 ;
    RECT 44.65 35.35 44.86 35.42 ;
    RECT 44.65 35.71 44.86 35.78 ;
    RECT 44.65 36.07 44.86 36.14 ;
    RECT 45.11 35.35 45.32 35.42 ;
    RECT 45.11 35.71 45.32 35.78 ;
    RECT 45.11 36.07 45.32 36.14 ;
    RECT 41.33 35.35 41.54 35.42 ;
    RECT 41.33 35.71 41.54 35.78 ;
    RECT 41.33 36.07 41.54 36.14 ;
    RECT 41.79 35.35 42.0 35.42 ;
    RECT 41.79 35.71 42.0 35.78 ;
    RECT 41.79 36.07 42.0 36.14 ;
    RECT 38.01 35.35 38.22 35.42 ;
    RECT 38.01 35.71 38.22 35.78 ;
    RECT 38.01 36.07 38.22 36.14 ;
    RECT 38.47 35.35 38.68 35.42 ;
    RECT 38.47 35.71 38.68 35.78 ;
    RECT 38.47 36.07 38.68 36.14 ;
    RECT 0.4 35.71 0.47 35.78 ;
    RECT 34.69 35.35 34.9 35.42 ;
    RECT 34.69 35.71 34.9 35.78 ;
    RECT 34.69 36.07 34.9 36.14 ;
    RECT 35.15 35.35 35.36 35.42 ;
    RECT 35.15 35.71 35.36 35.78 ;
    RECT 35.15 36.07 35.36 36.14 ;
    RECT 117.69 35.35 117.9 35.42 ;
    RECT 117.69 35.71 117.9 35.78 ;
    RECT 117.69 36.07 117.9 36.14 ;
    RECT 118.15 35.35 118.36 35.42 ;
    RECT 118.15 35.71 118.36 35.78 ;
    RECT 118.15 36.07 118.36 36.14 ;
    RECT 114.37 35.35 114.58 35.42 ;
    RECT 114.37 35.71 114.58 35.78 ;
    RECT 114.37 36.07 114.58 36.14 ;
    RECT 114.83 35.35 115.04 35.42 ;
    RECT 114.83 35.71 115.04 35.78 ;
    RECT 114.83 36.07 115.04 36.14 ;
    RECT 111.05 35.35 111.26 35.42 ;
    RECT 111.05 35.71 111.26 35.78 ;
    RECT 111.05 36.07 111.26 36.14 ;
    RECT 111.51 35.35 111.72 35.42 ;
    RECT 111.51 35.71 111.72 35.78 ;
    RECT 111.51 36.07 111.72 36.14 ;
    RECT 107.73 35.35 107.94 35.42 ;
    RECT 107.73 35.71 107.94 35.78 ;
    RECT 107.73 36.07 107.94 36.14 ;
    RECT 108.19 35.35 108.4 35.42 ;
    RECT 108.19 35.71 108.4 35.78 ;
    RECT 108.19 36.07 108.4 36.14 ;
    RECT 104.41 35.35 104.62 35.42 ;
    RECT 104.41 35.71 104.62 35.78 ;
    RECT 104.41 36.07 104.62 36.14 ;
    RECT 104.87 35.35 105.08 35.42 ;
    RECT 104.87 35.71 105.08 35.78 ;
    RECT 104.87 36.07 105.08 36.14 ;
    RECT 101.09 35.35 101.3 35.42 ;
    RECT 101.09 35.71 101.3 35.78 ;
    RECT 101.09 36.07 101.3 36.14 ;
    RECT 101.55 35.35 101.76 35.42 ;
    RECT 101.55 35.71 101.76 35.78 ;
    RECT 101.55 36.07 101.76 36.14 ;
    RECT 97.77 35.35 97.98 35.42 ;
    RECT 97.77 35.71 97.98 35.78 ;
    RECT 97.77 36.07 97.98 36.14 ;
    RECT 98.23 35.35 98.44 35.42 ;
    RECT 98.23 35.71 98.44 35.78 ;
    RECT 98.23 36.07 98.44 36.14 ;
    RECT 94.45 35.35 94.66 35.42 ;
    RECT 94.45 35.71 94.66 35.78 ;
    RECT 94.45 36.07 94.66 36.14 ;
    RECT 94.91 35.35 95.12 35.42 ;
    RECT 94.91 35.71 95.12 35.78 ;
    RECT 94.91 36.07 95.12 36.14 ;
    RECT 91.13 35.35 91.34 35.42 ;
    RECT 91.13 35.71 91.34 35.78 ;
    RECT 91.13 36.07 91.34 36.14 ;
    RECT 91.59 35.35 91.8 35.42 ;
    RECT 91.59 35.71 91.8 35.78 ;
    RECT 91.59 36.07 91.8 36.14 ;
    RECT 87.81 35.35 88.02 35.42 ;
    RECT 87.81 35.71 88.02 35.78 ;
    RECT 87.81 36.07 88.02 36.14 ;
    RECT 88.27 35.35 88.48 35.42 ;
    RECT 88.27 35.71 88.48 35.78 ;
    RECT 88.27 36.07 88.48 36.14 ;
    RECT 84.49 35.35 84.7 35.42 ;
    RECT 84.49 35.71 84.7 35.78 ;
    RECT 84.49 36.07 84.7 36.14 ;
    RECT 84.95 35.35 85.16 35.42 ;
    RECT 84.95 35.71 85.16 35.78 ;
    RECT 84.95 36.07 85.16 36.14 ;
    RECT 81.17 35.35 81.38 35.42 ;
    RECT 81.17 35.71 81.38 35.78 ;
    RECT 81.17 36.07 81.38 36.14 ;
    RECT 81.63 35.35 81.84 35.42 ;
    RECT 81.63 35.71 81.84 35.78 ;
    RECT 81.63 36.07 81.84 36.14 ;
    RECT 77.85 35.35 78.06 35.42 ;
    RECT 77.85 35.71 78.06 35.78 ;
    RECT 77.85 36.07 78.06 36.14 ;
    RECT 78.31 35.35 78.52 35.42 ;
    RECT 78.31 35.71 78.52 35.78 ;
    RECT 78.31 36.07 78.52 36.14 ;
    RECT 74.53 35.35 74.74 35.42 ;
    RECT 74.53 35.71 74.74 35.78 ;
    RECT 74.53 36.07 74.74 36.14 ;
    RECT 74.99 35.35 75.2 35.42 ;
    RECT 74.99 35.71 75.2 35.78 ;
    RECT 74.99 36.07 75.2 36.14 ;
    RECT 71.21 35.35 71.42 35.42 ;
    RECT 71.21 35.71 71.42 35.78 ;
    RECT 71.21 36.07 71.42 36.14 ;
    RECT 71.67 35.35 71.88 35.42 ;
    RECT 71.67 35.71 71.88 35.78 ;
    RECT 71.67 36.07 71.88 36.14 ;
    RECT 31.37 35.35 31.58 35.42 ;
    RECT 31.37 35.71 31.58 35.78 ;
    RECT 31.37 36.07 31.58 36.14 ;
    RECT 31.83 35.35 32.04 35.42 ;
    RECT 31.83 35.71 32.04 35.78 ;
    RECT 31.83 36.07 32.04 36.14 ;
    RECT 67.89 35.35 68.1 35.42 ;
    RECT 67.89 35.71 68.1 35.78 ;
    RECT 67.89 36.07 68.1 36.14 ;
    RECT 68.35 35.35 68.56 35.42 ;
    RECT 68.35 35.71 68.56 35.78 ;
    RECT 68.35 36.07 68.56 36.14 ;
    RECT 28.05 35.35 28.26 35.42 ;
    RECT 28.05 35.71 28.26 35.78 ;
    RECT 28.05 36.07 28.26 36.14 ;
    RECT 28.51 35.35 28.72 35.42 ;
    RECT 28.51 35.71 28.72 35.78 ;
    RECT 28.51 36.07 28.72 36.14 ;
    RECT 24.73 35.35 24.94 35.42 ;
    RECT 24.73 35.71 24.94 35.78 ;
    RECT 24.73 36.07 24.94 36.14 ;
    RECT 25.19 35.35 25.4 35.42 ;
    RECT 25.19 35.71 25.4 35.78 ;
    RECT 25.19 36.07 25.4 36.14 ;
    RECT 21.41 35.35 21.62 35.42 ;
    RECT 21.41 35.71 21.62 35.78 ;
    RECT 21.41 36.07 21.62 36.14 ;
    RECT 21.87 35.35 22.08 35.42 ;
    RECT 21.87 35.71 22.08 35.78 ;
    RECT 21.87 36.07 22.08 36.14 ;
    RECT 18.09 35.35 18.3 35.42 ;
    RECT 18.09 35.71 18.3 35.78 ;
    RECT 18.09 36.07 18.3 36.14 ;
    RECT 18.55 35.35 18.76 35.42 ;
    RECT 18.55 35.71 18.76 35.78 ;
    RECT 18.55 36.07 18.76 36.14 ;
    RECT 120.825 35.71 120.895 35.78 ;
    RECT 14.77 35.35 14.98 35.42 ;
    RECT 14.77 35.71 14.98 35.78 ;
    RECT 14.77 36.07 14.98 36.14 ;
    RECT 15.23 35.35 15.44 35.42 ;
    RECT 15.23 35.71 15.44 35.78 ;
    RECT 15.23 36.07 15.44 36.14 ;
    RECT 11.45 35.35 11.66 35.42 ;
    RECT 11.45 35.71 11.66 35.78 ;
    RECT 11.45 36.07 11.66 36.14 ;
    RECT 11.91 35.35 12.12 35.42 ;
    RECT 11.91 35.71 12.12 35.78 ;
    RECT 11.91 36.07 12.12 36.14 ;
    RECT 8.13 35.35 8.34 35.42 ;
    RECT 8.13 35.71 8.34 35.78 ;
    RECT 8.13 36.07 8.34 36.14 ;
    RECT 8.59 35.35 8.8 35.42 ;
    RECT 8.59 35.71 8.8 35.78 ;
    RECT 8.59 36.07 8.8 36.14 ;
    RECT 4.81 35.35 5.02 35.42 ;
    RECT 4.81 35.71 5.02 35.78 ;
    RECT 4.81 36.07 5.02 36.14 ;
    RECT 5.27 35.35 5.48 35.42 ;
    RECT 5.27 35.71 5.48 35.78 ;
    RECT 5.27 36.07 5.48 36.14 ;
    RECT 1.49 35.35 1.7 35.42 ;
    RECT 1.49 35.71 1.7 35.78 ;
    RECT 1.49 36.07 1.7 36.14 ;
    RECT 1.95 35.35 2.16 35.42 ;
    RECT 1.95 35.71 2.16 35.78 ;
    RECT 1.95 36.07 2.16 36.14 ;
    RECT 64.57 35.35 64.78 35.42 ;
    RECT 64.57 35.71 64.78 35.78 ;
    RECT 64.57 36.07 64.78 36.14 ;
    RECT 65.03 35.35 65.24 35.42 ;
    RECT 65.03 35.71 65.24 35.78 ;
    RECT 65.03 36.07 65.24 36.14 ;
    RECT 61.25 34.63 61.46 34.7 ;
    RECT 61.25 34.99 61.46 35.06 ;
    RECT 61.25 35.35 61.46 35.42 ;
    RECT 61.71 34.63 61.92 34.7 ;
    RECT 61.71 34.99 61.92 35.06 ;
    RECT 61.71 35.35 61.92 35.42 ;
    RECT 57.93 34.63 58.14 34.7 ;
    RECT 57.93 34.99 58.14 35.06 ;
    RECT 57.93 35.35 58.14 35.42 ;
    RECT 58.39 34.63 58.6 34.7 ;
    RECT 58.39 34.99 58.6 35.06 ;
    RECT 58.39 35.35 58.6 35.42 ;
    RECT 54.61 34.63 54.82 34.7 ;
    RECT 54.61 34.99 54.82 35.06 ;
    RECT 54.61 35.35 54.82 35.42 ;
    RECT 55.07 34.63 55.28 34.7 ;
    RECT 55.07 34.99 55.28 35.06 ;
    RECT 55.07 35.35 55.28 35.42 ;
    RECT 51.29 34.63 51.5 34.7 ;
    RECT 51.29 34.99 51.5 35.06 ;
    RECT 51.29 35.35 51.5 35.42 ;
    RECT 51.75 34.63 51.96 34.7 ;
    RECT 51.75 34.99 51.96 35.06 ;
    RECT 51.75 35.35 51.96 35.42 ;
    RECT 47.97 34.63 48.18 34.7 ;
    RECT 47.97 34.99 48.18 35.06 ;
    RECT 47.97 35.35 48.18 35.42 ;
    RECT 48.43 34.63 48.64 34.7 ;
    RECT 48.43 34.99 48.64 35.06 ;
    RECT 48.43 35.35 48.64 35.42 ;
    RECT 44.65 34.63 44.86 34.7 ;
    RECT 44.65 34.99 44.86 35.06 ;
    RECT 44.65 35.35 44.86 35.42 ;
    RECT 45.11 34.63 45.32 34.7 ;
    RECT 45.11 34.99 45.32 35.06 ;
    RECT 45.11 35.35 45.32 35.42 ;
    RECT 41.33 34.63 41.54 34.7 ;
    RECT 41.33 34.99 41.54 35.06 ;
    RECT 41.33 35.35 41.54 35.42 ;
    RECT 41.79 34.63 42.0 34.7 ;
    RECT 41.79 34.99 42.0 35.06 ;
    RECT 41.79 35.35 42.0 35.42 ;
    RECT 38.01 34.63 38.22 34.7 ;
    RECT 38.01 34.99 38.22 35.06 ;
    RECT 38.01 35.35 38.22 35.42 ;
    RECT 38.47 34.63 38.68 34.7 ;
    RECT 38.47 34.99 38.68 35.06 ;
    RECT 38.47 35.35 38.68 35.42 ;
    RECT 0.4 34.99 0.47 35.06 ;
    RECT 34.69 34.63 34.9 34.7 ;
    RECT 34.69 34.99 34.9 35.06 ;
    RECT 34.69 35.35 34.9 35.42 ;
    RECT 35.15 34.63 35.36 34.7 ;
    RECT 35.15 34.99 35.36 35.06 ;
    RECT 35.15 35.35 35.36 35.42 ;
    RECT 117.69 34.63 117.9 34.7 ;
    RECT 117.69 34.99 117.9 35.06 ;
    RECT 117.69 35.35 117.9 35.42 ;
    RECT 118.15 34.63 118.36 34.7 ;
    RECT 118.15 34.99 118.36 35.06 ;
    RECT 118.15 35.35 118.36 35.42 ;
    RECT 114.37 34.63 114.58 34.7 ;
    RECT 114.37 34.99 114.58 35.06 ;
    RECT 114.37 35.35 114.58 35.42 ;
    RECT 114.83 34.63 115.04 34.7 ;
    RECT 114.83 34.99 115.04 35.06 ;
    RECT 114.83 35.35 115.04 35.42 ;
    RECT 111.05 34.63 111.26 34.7 ;
    RECT 111.05 34.99 111.26 35.06 ;
    RECT 111.05 35.35 111.26 35.42 ;
    RECT 111.51 34.63 111.72 34.7 ;
    RECT 111.51 34.99 111.72 35.06 ;
    RECT 111.51 35.35 111.72 35.42 ;
    RECT 107.73 34.63 107.94 34.7 ;
    RECT 107.73 34.99 107.94 35.06 ;
    RECT 107.73 35.35 107.94 35.42 ;
    RECT 108.19 34.63 108.4 34.7 ;
    RECT 108.19 34.99 108.4 35.06 ;
    RECT 108.19 35.35 108.4 35.42 ;
    RECT 104.41 34.63 104.62 34.7 ;
    RECT 104.41 34.99 104.62 35.06 ;
    RECT 104.41 35.35 104.62 35.42 ;
    RECT 104.87 34.63 105.08 34.7 ;
    RECT 104.87 34.99 105.08 35.06 ;
    RECT 104.87 35.35 105.08 35.42 ;
    RECT 101.09 34.63 101.3 34.7 ;
    RECT 101.09 34.99 101.3 35.06 ;
    RECT 101.09 35.35 101.3 35.42 ;
    RECT 101.55 34.63 101.76 34.7 ;
    RECT 101.55 34.99 101.76 35.06 ;
    RECT 101.55 35.35 101.76 35.42 ;
    RECT 97.77 34.63 97.98 34.7 ;
    RECT 97.77 34.99 97.98 35.06 ;
    RECT 97.77 35.35 97.98 35.42 ;
    RECT 98.23 34.63 98.44 34.7 ;
    RECT 98.23 34.99 98.44 35.06 ;
    RECT 98.23 35.35 98.44 35.42 ;
    RECT 94.45 34.63 94.66 34.7 ;
    RECT 94.45 34.99 94.66 35.06 ;
    RECT 94.45 35.35 94.66 35.42 ;
    RECT 94.91 34.63 95.12 34.7 ;
    RECT 94.91 34.99 95.12 35.06 ;
    RECT 94.91 35.35 95.12 35.42 ;
    RECT 91.13 34.63 91.34 34.7 ;
    RECT 91.13 34.99 91.34 35.06 ;
    RECT 91.13 35.35 91.34 35.42 ;
    RECT 91.59 34.63 91.8 34.7 ;
    RECT 91.59 34.99 91.8 35.06 ;
    RECT 91.59 35.35 91.8 35.42 ;
    RECT 87.81 34.63 88.02 34.7 ;
    RECT 87.81 34.99 88.02 35.06 ;
    RECT 87.81 35.35 88.02 35.42 ;
    RECT 88.27 34.63 88.48 34.7 ;
    RECT 88.27 34.99 88.48 35.06 ;
    RECT 88.27 35.35 88.48 35.42 ;
    RECT 84.49 34.63 84.7 34.7 ;
    RECT 84.49 34.99 84.7 35.06 ;
    RECT 84.49 35.35 84.7 35.42 ;
    RECT 84.95 34.63 85.16 34.7 ;
    RECT 84.95 34.99 85.16 35.06 ;
    RECT 84.95 35.35 85.16 35.42 ;
    RECT 81.17 34.63 81.38 34.7 ;
    RECT 81.17 34.99 81.38 35.06 ;
    RECT 81.17 35.35 81.38 35.42 ;
    RECT 81.63 34.63 81.84 34.7 ;
    RECT 81.63 34.99 81.84 35.06 ;
    RECT 81.63 35.35 81.84 35.42 ;
    RECT 77.85 34.63 78.06 34.7 ;
    RECT 77.85 34.99 78.06 35.06 ;
    RECT 77.85 35.35 78.06 35.42 ;
    RECT 78.31 34.63 78.52 34.7 ;
    RECT 78.31 34.99 78.52 35.06 ;
    RECT 78.31 35.35 78.52 35.42 ;
    RECT 74.53 34.63 74.74 34.7 ;
    RECT 74.53 34.99 74.74 35.06 ;
    RECT 74.53 35.35 74.74 35.42 ;
    RECT 74.99 34.63 75.2 34.7 ;
    RECT 74.99 34.99 75.2 35.06 ;
    RECT 74.99 35.35 75.2 35.42 ;
    RECT 71.21 34.63 71.42 34.7 ;
    RECT 71.21 34.99 71.42 35.06 ;
    RECT 71.21 35.35 71.42 35.42 ;
    RECT 71.67 34.63 71.88 34.7 ;
    RECT 71.67 34.99 71.88 35.06 ;
    RECT 71.67 35.35 71.88 35.42 ;
    RECT 31.37 34.63 31.58 34.7 ;
    RECT 31.37 34.99 31.58 35.06 ;
    RECT 31.37 35.35 31.58 35.42 ;
    RECT 31.83 34.63 32.04 34.7 ;
    RECT 31.83 34.99 32.04 35.06 ;
    RECT 31.83 35.35 32.04 35.42 ;
    RECT 67.89 34.63 68.1 34.7 ;
    RECT 67.89 34.99 68.1 35.06 ;
    RECT 67.89 35.35 68.1 35.42 ;
    RECT 68.35 34.63 68.56 34.7 ;
    RECT 68.35 34.99 68.56 35.06 ;
    RECT 68.35 35.35 68.56 35.42 ;
    RECT 28.05 34.63 28.26 34.7 ;
    RECT 28.05 34.99 28.26 35.06 ;
    RECT 28.05 35.35 28.26 35.42 ;
    RECT 28.51 34.63 28.72 34.7 ;
    RECT 28.51 34.99 28.72 35.06 ;
    RECT 28.51 35.35 28.72 35.42 ;
    RECT 24.73 34.63 24.94 34.7 ;
    RECT 24.73 34.99 24.94 35.06 ;
    RECT 24.73 35.35 24.94 35.42 ;
    RECT 25.19 34.63 25.4 34.7 ;
    RECT 25.19 34.99 25.4 35.06 ;
    RECT 25.19 35.35 25.4 35.42 ;
    RECT 21.41 34.63 21.62 34.7 ;
    RECT 21.41 34.99 21.62 35.06 ;
    RECT 21.41 35.35 21.62 35.42 ;
    RECT 21.87 34.63 22.08 34.7 ;
    RECT 21.87 34.99 22.08 35.06 ;
    RECT 21.87 35.35 22.08 35.42 ;
    RECT 18.09 34.63 18.3 34.7 ;
    RECT 18.09 34.99 18.3 35.06 ;
    RECT 18.09 35.35 18.3 35.42 ;
    RECT 18.55 34.63 18.76 34.7 ;
    RECT 18.55 34.99 18.76 35.06 ;
    RECT 18.55 35.35 18.76 35.42 ;
    RECT 120.825 34.99 120.895 35.06 ;
    RECT 14.77 34.63 14.98 34.7 ;
    RECT 14.77 34.99 14.98 35.06 ;
    RECT 14.77 35.35 14.98 35.42 ;
    RECT 15.23 34.63 15.44 34.7 ;
    RECT 15.23 34.99 15.44 35.06 ;
    RECT 15.23 35.35 15.44 35.42 ;
    RECT 11.45 34.63 11.66 34.7 ;
    RECT 11.45 34.99 11.66 35.06 ;
    RECT 11.45 35.35 11.66 35.42 ;
    RECT 11.91 34.63 12.12 34.7 ;
    RECT 11.91 34.99 12.12 35.06 ;
    RECT 11.91 35.35 12.12 35.42 ;
    RECT 8.13 34.63 8.34 34.7 ;
    RECT 8.13 34.99 8.34 35.06 ;
    RECT 8.13 35.35 8.34 35.42 ;
    RECT 8.59 34.63 8.8 34.7 ;
    RECT 8.59 34.99 8.8 35.06 ;
    RECT 8.59 35.35 8.8 35.42 ;
    RECT 4.81 34.63 5.02 34.7 ;
    RECT 4.81 34.99 5.02 35.06 ;
    RECT 4.81 35.35 5.02 35.42 ;
    RECT 5.27 34.63 5.48 34.7 ;
    RECT 5.27 34.99 5.48 35.06 ;
    RECT 5.27 35.35 5.48 35.42 ;
    RECT 1.49 34.63 1.7 34.7 ;
    RECT 1.49 34.99 1.7 35.06 ;
    RECT 1.49 35.35 1.7 35.42 ;
    RECT 1.95 34.63 2.16 34.7 ;
    RECT 1.95 34.99 2.16 35.06 ;
    RECT 1.95 35.35 2.16 35.42 ;
    RECT 64.57 34.63 64.78 34.7 ;
    RECT 64.57 34.99 64.78 35.06 ;
    RECT 64.57 35.35 64.78 35.42 ;
    RECT 65.03 34.63 65.24 34.7 ;
    RECT 65.03 34.99 65.24 35.06 ;
    RECT 65.03 35.35 65.24 35.42 ;
    RECT 61.25 33.91 61.46 33.98 ;
    RECT 61.25 34.27 61.46 34.34 ;
    RECT 61.25 34.63 61.46 34.7 ;
    RECT 61.71 33.91 61.92 33.98 ;
    RECT 61.71 34.27 61.92 34.34 ;
    RECT 61.71 34.63 61.92 34.7 ;
    RECT 57.93 33.91 58.14 33.98 ;
    RECT 57.93 34.27 58.14 34.34 ;
    RECT 57.93 34.63 58.14 34.7 ;
    RECT 58.39 33.91 58.6 33.98 ;
    RECT 58.39 34.27 58.6 34.34 ;
    RECT 58.39 34.63 58.6 34.7 ;
    RECT 54.61 33.91 54.82 33.98 ;
    RECT 54.61 34.27 54.82 34.34 ;
    RECT 54.61 34.63 54.82 34.7 ;
    RECT 55.07 33.91 55.28 33.98 ;
    RECT 55.07 34.27 55.28 34.34 ;
    RECT 55.07 34.63 55.28 34.7 ;
    RECT 51.29 33.91 51.5 33.98 ;
    RECT 51.29 34.27 51.5 34.34 ;
    RECT 51.29 34.63 51.5 34.7 ;
    RECT 51.75 33.91 51.96 33.98 ;
    RECT 51.75 34.27 51.96 34.34 ;
    RECT 51.75 34.63 51.96 34.7 ;
    RECT 47.97 33.91 48.18 33.98 ;
    RECT 47.97 34.27 48.18 34.34 ;
    RECT 47.97 34.63 48.18 34.7 ;
    RECT 48.43 33.91 48.64 33.98 ;
    RECT 48.43 34.27 48.64 34.34 ;
    RECT 48.43 34.63 48.64 34.7 ;
    RECT 44.65 33.91 44.86 33.98 ;
    RECT 44.65 34.27 44.86 34.34 ;
    RECT 44.65 34.63 44.86 34.7 ;
    RECT 45.11 33.91 45.32 33.98 ;
    RECT 45.11 34.27 45.32 34.34 ;
    RECT 45.11 34.63 45.32 34.7 ;
    RECT 41.33 33.91 41.54 33.98 ;
    RECT 41.33 34.27 41.54 34.34 ;
    RECT 41.33 34.63 41.54 34.7 ;
    RECT 41.79 33.91 42.0 33.98 ;
    RECT 41.79 34.27 42.0 34.34 ;
    RECT 41.79 34.63 42.0 34.7 ;
    RECT 38.01 33.91 38.22 33.98 ;
    RECT 38.01 34.27 38.22 34.34 ;
    RECT 38.01 34.63 38.22 34.7 ;
    RECT 38.47 33.91 38.68 33.98 ;
    RECT 38.47 34.27 38.68 34.34 ;
    RECT 38.47 34.63 38.68 34.7 ;
    RECT 0.4 34.27 0.47 34.34 ;
    RECT 34.69 33.91 34.9 33.98 ;
    RECT 34.69 34.27 34.9 34.34 ;
    RECT 34.69 34.63 34.9 34.7 ;
    RECT 35.15 33.91 35.36 33.98 ;
    RECT 35.15 34.27 35.36 34.34 ;
    RECT 35.15 34.63 35.36 34.7 ;
    RECT 117.69 33.91 117.9 33.98 ;
    RECT 117.69 34.27 117.9 34.34 ;
    RECT 117.69 34.63 117.9 34.7 ;
    RECT 118.15 33.91 118.36 33.98 ;
    RECT 118.15 34.27 118.36 34.34 ;
    RECT 118.15 34.63 118.36 34.7 ;
    RECT 114.37 33.91 114.58 33.98 ;
    RECT 114.37 34.27 114.58 34.34 ;
    RECT 114.37 34.63 114.58 34.7 ;
    RECT 114.83 33.91 115.04 33.98 ;
    RECT 114.83 34.27 115.04 34.34 ;
    RECT 114.83 34.63 115.04 34.7 ;
    RECT 111.05 33.91 111.26 33.98 ;
    RECT 111.05 34.27 111.26 34.34 ;
    RECT 111.05 34.63 111.26 34.7 ;
    RECT 111.51 33.91 111.72 33.98 ;
    RECT 111.51 34.27 111.72 34.34 ;
    RECT 111.51 34.63 111.72 34.7 ;
    RECT 107.73 33.91 107.94 33.98 ;
    RECT 107.73 34.27 107.94 34.34 ;
    RECT 107.73 34.63 107.94 34.7 ;
    RECT 108.19 33.91 108.4 33.98 ;
    RECT 108.19 34.27 108.4 34.34 ;
    RECT 108.19 34.63 108.4 34.7 ;
    RECT 104.41 33.91 104.62 33.98 ;
    RECT 104.41 34.27 104.62 34.34 ;
    RECT 104.41 34.63 104.62 34.7 ;
    RECT 104.87 33.91 105.08 33.98 ;
    RECT 104.87 34.27 105.08 34.34 ;
    RECT 104.87 34.63 105.08 34.7 ;
    RECT 101.09 33.91 101.3 33.98 ;
    RECT 101.09 34.27 101.3 34.34 ;
    RECT 101.09 34.63 101.3 34.7 ;
    RECT 101.55 33.91 101.76 33.98 ;
    RECT 101.55 34.27 101.76 34.34 ;
    RECT 101.55 34.63 101.76 34.7 ;
    RECT 97.77 33.91 97.98 33.98 ;
    RECT 97.77 34.27 97.98 34.34 ;
    RECT 97.77 34.63 97.98 34.7 ;
    RECT 98.23 33.91 98.44 33.98 ;
    RECT 98.23 34.27 98.44 34.34 ;
    RECT 98.23 34.63 98.44 34.7 ;
    RECT 94.45 33.91 94.66 33.98 ;
    RECT 94.45 34.27 94.66 34.34 ;
    RECT 94.45 34.63 94.66 34.7 ;
    RECT 94.91 33.91 95.12 33.98 ;
    RECT 94.91 34.27 95.12 34.34 ;
    RECT 94.91 34.63 95.12 34.7 ;
    RECT 91.13 33.91 91.34 33.98 ;
    RECT 91.13 34.27 91.34 34.34 ;
    RECT 91.13 34.63 91.34 34.7 ;
    RECT 91.59 33.91 91.8 33.98 ;
    RECT 91.59 34.27 91.8 34.34 ;
    RECT 91.59 34.63 91.8 34.7 ;
    RECT 87.81 33.91 88.02 33.98 ;
    RECT 87.81 34.27 88.02 34.34 ;
    RECT 87.81 34.63 88.02 34.7 ;
    RECT 88.27 33.91 88.48 33.98 ;
    RECT 88.27 34.27 88.48 34.34 ;
    RECT 88.27 34.63 88.48 34.7 ;
    RECT 84.49 33.91 84.7 33.98 ;
    RECT 84.49 34.27 84.7 34.34 ;
    RECT 84.49 34.63 84.7 34.7 ;
    RECT 84.95 33.91 85.16 33.98 ;
    RECT 84.95 34.27 85.16 34.34 ;
    RECT 84.95 34.63 85.16 34.7 ;
    RECT 81.17 33.91 81.38 33.98 ;
    RECT 81.17 34.27 81.38 34.34 ;
    RECT 81.17 34.63 81.38 34.7 ;
    RECT 81.63 33.91 81.84 33.98 ;
    RECT 81.63 34.27 81.84 34.34 ;
    RECT 81.63 34.63 81.84 34.7 ;
    RECT 77.85 33.91 78.06 33.98 ;
    RECT 77.85 34.27 78.06 34.34 ;
    RECT 77.85 34.63 78.06 34.7 ;
    RECT 78.31 33.91 78.52 33.98 ;
    RECT 78.31 34.27 78.52 34.34 ;
    RECT 78.31 34.63 78.52 34.7 ;
    RECT 74.53 33.91 74.74 33.98 ;
    RECT 74.53 34.27 74.74 34.34 ;
    RECT 74.53 34.63 74.74 34.7 ;
    RECT 74.99 33.91 75.2 33.98 ;
    RECT 74.99 34.27 75.2 34.34 ;
    RECT 74.99 34.63 75.2 34.7 ;
    RECT 71.21 33.91 71.42 33.98 ;
    RECT 71.21 34.27 71.42 34.34 ;
    RECT 71.21 34.63 71.42 34.7 ;
    RECT 71.67 33.91 71.88 33.98 ;
    RECT 71.67 34.27 71.88 34.34 ;
    RECT 71.67 34.63 71.88 34.7 ;
    RECT 31.37 33.91 31.58 33.98 ;
    RECT 31.37 34.27 31.58 34.34 ;
    RECT 31.37 34.63 31.58 34.7 ;
    RECT 31.83 33.91 32.04 33.98 ;
    RECT 31.83 34.27 32.04 34.34 ;
    RECT 31.83 34.63 32.04 34.7 ;
    RECT 67.89 33.91 68.1 33.98 ;
    RECT 67.89 34.27 68.1 34.34 ;
    RECT 67.89 34.63 68.1 34.7 ;
    RECT 68.35 33.91 68.56 33.98 ;
    RECT 68.35 34.27 68.56 34.34 ;
    RECT 68.35 34.63 68.56 34.7 ;
    RECT 28.05 33.91 28.26 33.98 ;
    RECT 28.05 34.27 28.26 34.34 ;
    RECT 28.05 34.63 28.26 34.7 ;
    RECT 28.51 33.91 28.72 33.98 ;
    RECT 28.51 34.27 28.72 34.34 ;
    RECT 28.51 34.63 28.72 34.7 ;
    RECT 24.73 33.91 24.94 33.98 ;
    RECT 24.73 34.27 24.94 34.34 ;
    RECT 24.73 34.63 24.94 34.7 ;
    RECT 25.19 33.91 25.4 33.98 ;
    RECT 25.19 34.27 25.4 34.34 ;
    RECT 25.19 34.63 25.4 34.7 ;
    RECT 21.41 33.91 21.62 33.98 ;
    RECT 21.41 34.27 21.62 34.34 ;
    RECT 21.41 34.63 21.62 34.7 ;
    RECT 21.87 33.91 22.08 33.98 ;
    RECT 21.87 34.27 22.08 34.34 ;
    RECT 21.87 34.63 22.08 34.7 ;
    RECT 18.09 33.91 18.3 33.98 ;
    RECT 18.09 34.27 18.3 34.34 ;
    RECT 18.09 34.63 18.3 34.7 ;
    RECT 18.55 33.91 18.76 33.98 ;
    RECT 18.55 34.27 18.76 34.34 ;
    RECT 18.55 34.63 18.76 34.7 ;
    RECT 120.825 34.27 120.895 34.34 ;
    RECT 14.77 33.91 14.98 33.98 ;
    RECT 14.77 34.27 14.98 34.34 ;
    RECT 14.77 34.63 14.98 34.7 ;
    RECT 15.23 33.91 15.44 33.98 ;
    RECT 15.23 34.27 15.44 34.34 ;
    RECT 15.23 34.63 15.44 34.7 ;
    RECT 11.45 33.91 11.66 33.98 ;
    RECT 11.45 34.27 11.66 34.34 ;
    RECT 11.45 34.63 11.66 34.7 ;
    RECT 11.91 33.91 12.12 33.98 ;
    RECT 11.91 34.27 12.12 34.34 ;
    RECT 11.91 34.63 12.12 34.7 ;
    RECT 8.13 33.91 8.34 33.98 ;
    RECT 8.13 34.27 8.34 34.34 ;
    RECT 8.13 34.63 8.34 34.7 ;
    RECT 8.59 33.91 8.8 33.98 ;
    RECT 8.59 34.27 8.8 34.34 ;
    RECT 8.59 34.63 8.8 34.7 ;
    RECT 4.81 33.91 5.02 33.98 ;
    RECT 4.81 34.27 5.02 34.34 ;
    RECT 4.81 34.63 5.02 34.7 ;
    RECT 5.27 33.91 5.48 33.98 ;
    RECT 5.27 34.27 5.48 34.34 ;
    RECT 5.27 34.63 5.48 34.7 ;
    RECT 1.49 33.91 1.7 33.98 ;
    RECT 1.49 34.27 1.7 34.34 ;
    RECT 1.49 34.63 1.7 34.7 ;
    RECT 1.95 33.91 2.16 33.98 ;
    RECT 1.95 34.27 2.16 34.34 ;
    RECT 1.95 34.63 2.16 34.7 ;
    RECT 64.57 33.91 64.78 33.98 ;
    RECT 64.57 34.27 64.78 34.34 ;
    RECT 64.57 34.63 64.78 34.7 ;
    RECT 65.03 33.91 65.24 33.98 ;
    RECT 65.03 34.27 65.24 34.34 ;
    RECT 65.03 34.63 65.24 34.7 ;
    RECT 61.25 33.19 61.46 33.26 ;
    RECT 61.25 33.55 61.46 33.62 ;
    RECT 61.25 33.91 61.46 33.98 ;
    RECT 61.71 33.19 61.92 33.26 ;
    RECT 61.71 33.55 61.92 33.62 ;
    RECT 61.71 33.91 61.92 33.98 ;
    RECT 57.93 33.19 58.14 33.26 ;
    RECT 57.93 33.55 58.14 33.62 ;
    RECT 57.93 33.91 58.14 33.98 ;
    RECT 58.39 33.19 58.6 33.26 ;
    RECT 58.39 33.55 58.6 33.62 ;
    RECT 58.39 33.91 58.6 33.98 ;
    RECT 54.61 33.19 54.82 33.26 ;
    RECT 54.61 33.55 54.82 33.62 ;
    RECT 54.61 33.91 54.82 33.98 ;
    RECT 55.07 33.19 55.28 33.26 ;
    RECT 55.07 33.55 55.28 33.62 ;
    RECT 55.07 33.91 55.28 33.98 ;
    RECT 51.29 33.19 51.5 33.26 ;
    RECT 51.29 33.55 51.5 33.62 ;
    RECT 51.29 33.91 51.5 33.98 ;
    RECT 51.75 33.19 51.96 33.26 ;
    RECT 51.75 33.55 51.96 33.62 ;
    RECT 51.75 33.91 51.96 33.98 ;
    RECT 47.97 33.19 48.18 33.26 ;
    RECT 47.97 33.55 48.18 33.62 ;
    RECT 47.97 33.91 48.18 33.98 ;
    RECT 48.43 33.19 48.64 33.26 ;
    RECT 48.43 33.55 48.64 33.62 ;
    RECT 48.43 33.91 48.64 33.98 ;
    RECT 44.65 33.19 44.86 33.26 ;
    RECT 44.65 33.55 44.86 33.62 ;
    RECT 44.65 33.91 44.86 33.98 ;
    RECT 45.11 33.19 45.32 33.26 ;
    RECT 45.11 33.55 45.32 33.62 ;
    RECT 45.11 33.91 45.32 33.98 ;
    RECT 41.33 33.19 41.54 33.26 ;
    RECT 41.33 33.55 41.54 33.62 ;
    RECT 41.33 33.91 41.54 33.98 ;
    RECT 41.79 33.19 42.0 33.26 ;
    RECT 41.79 33.55 42.0 33.62 ;
    RECT 41.79 33.91 42.0 33.98 ;
    RECT 38.01 33.19 38.22 33.26 ;
    RECT 38.01 33.55 38.22 33.62 ;
    RECT 38.01 33.91 38.22 33.98 ;
    RECT 38.47 33.19 38.68 33.26 ;
    RECT 38.47 33.55 38.68 33.62 ;
    RECT 38.47 33.91 38.68 33.98 ;
    RECT 0.4 33.55 0.47 33.62 ;
    RECT 34.69 33.19 34.9 33.26 ;
    RECT 34.69 33.55 34.9 33.62 ;
    RECT 34.69 33.91 34.9 33.98 ;
    RECT 35.15 33.19 35.36 33.26 ;
    RECT 35.15 33.55 35.36 33.62 ;
    RECT 35.15 33.91 35.36 33.98 ;
    RECT 117.69 33.19 117.9 33.26 ;
    RECT 117.69 33.55 117.9 33.62 ;
    RECT 117.69 33.91 117.9 33.98 ;
    RECT 118.15 33.19 118.36 33.26 ;
    RECT 118.15 33.55 118.36 33.62 ;
    RECT 118.15 33.91 118.36 33.98 ;
    RECT 114.37 33.19 114.58 33.26 ;
    RECT 114.37 33.55 114.58 33.62 ;
    RECT 114.37 33.91 114.58 33.98 ;
    RECT 114.83 33.19 115.04 33.26 ;
    RECT 114.83 33.55 115.04 33.62 ;
    RECT 114.83 33.91 115.04 33.98 ;
    RECT 111.05 33.19 111.26 33.26 ;
    RECT 111.05 33.55 111.26 33.62 ;
    RECT 111.05 33.91 111.26 33.98 ;
    RECT 111.51 33.19 111.72 33.26 ;
    RECT 111.51 33.55 111.72 33.62 ;
    RECT 111.51 33.91 111.72 33.98 ;
    RECT 107.73 33.19 107.94 33.26 ;
    RECT 107.73 33.55 107.94 33.62 ;
    RECT 107.73 33.91 107.94 33.98 ;
    RECT 108.19 33.19 108.4 33.26 ;
    RECT 108.19 33.55 108.4 33.62 ;
    RECT 108.19 33.91 108.4 33.98 ;
    RECT 104.41 33.19 104.62 33.26 ;
    RECT 104.41 33.55 104.62 33.62 ;
    RECT 104.41 33.91 104.62 33.98 ;
    RECT 104.87 33.19 105.08 33.26 ;
    RECT 104.87 33.55 105.08 33.62 ;
    RECT 104.87 33.91 105.08 33.98 ;
    RECT 101.09 33.19 101.3 33.26 ;
    RECT 101.09 33.55 101.3 33.62 ;
    RECT 101.09 33.91 101.3 33.98 ;
    RECT 101.55 33.19 101.76 33.26 ;
    RECT 101.55 33.55 101.76 33.62 ;
    RECT 101.55 33.91 101.76 33.98 ;
    RECT 97.77 33.19 97.98 33.26 ;
    RECT 97.77 33.55 97.98 33.62 ;
    RECT 97.77 33.91 97.98 33.98 ;
    RECT 98.23 33.19 98.44 33.26 ;
    RECT 98.23 33.55 98.44 33.62 ;
    RECT 98.23 33.91 98.44 33.98 ;
    RECT 94.45 33.19 94.66 33.26 ;
    RECT 94.45 33.55 94.66 33.62 ;
    RECT 94.45 33.91 94.66 33.98 ;
    RECT 94.91 33.19 95.12 33.26 ;
    RECT 94.91 33.55 95.12 33.62 ;
    RECT 94.91 33.91 95.12 33.98 ;
    RECT 91.13 33.19 91.34 33.26 ;
    RECT 91.13 33.55 91.34 33.62 ;
    RECT 91.13 33.91 91.34 33.98 ;
    RECT 91.59 33.19 91.8 33.26 ;
    RECT 91.59 33.55 91.8 33.62 ;
    RECT 91.59 33.91 91.8 33.98 ;
    RECT 87.81 33.19 88.02 33.26 ;
    RECT 87.81 33.55 88.02 33.62 ;
    RECT 87.81 33.91 88.02 33.98 ;
    RECT 88.27 33.19 88.48 33.26 ;
    RECT 88.27 33.55 88.48 33.62 ;
    RECT 88.27 33.91 88.48 33.98 ;
    RECT 84.49 33.19 84.7 33.26 ;
    RECT 84.49 33.55 84.7 33.62 ;
    RECT 84.49 33.91 84.7 33.98 ;
    RECT 84.95 33.19 85.16 33.26 ;
    RECT 84.95 33.55 85.16 33.62 ;
    RECT 84.95 33.91 85.16 33.98 ;
    RECT 81.17 33.19 81.38 33.26 ;
    RECT 81.17 33.55 81.38 33.62 ;
    RECT 81.17 33.91 81.38 33.98 ;
    RECT 81.63 33.19 81.84 33.26 ;
    RECT 81.63 33.55 81.84 33.62 ;
    RECT 81.63 33.91 81.84 33.98 ;
    RECT 77.85 33.19 78.06 33.26 ;
    RECT 77.85 33.55 78.06 33.62 ;
    RECT 77.85 33.91 78.06 33.98 ;
    RECT 78.31 33.19 78.52 33.26 ;
    RECT 78.31 33.55 78.52 33.62 ;
    RECT 78.31 33.91 78.52 33.98 ;
    RECT 74.53 33.19 74.74 33.26 ;
    RECT 74.53 33.55 74.74 33.62 ;
    RECT 74.53 33.91 74.74 33.98 ;
    RECT 74.99 33.19 75.2 33.26 ;
    RECT 74.99 33.55 75.2 33.62 ;
    RECT 74.99 33.91 75.2 33.98 ;
    RECT 71.21 33.19 71.42 33.26 ;
    RECT 71.21 33.55 71.42 33.62 ;
    RECT 71.21 33.91 71.42 33.98 ;
    RECT 71.67 33.19 71.88 33.26 ;
    RECT 71.67 33.55 71.88 33.62 ;
    RECT 71.67 33.91 71.88 33.98 ;
    RECT 31.37 33.19 31.58 33.26 ;
    RECT 31.37 33.55 31.58 33.62 ;
    RECT 31.37 33.91 31.58 33.98 ;
    RECT 31.83 33.19 32.04 33.26 ;
    RECT 31.83 33.55 32.04 33.62 ;
    RECT 31.83 33.91 32.04 33.98 ;
    RECT 67.89 33.19 68.1 33.26 ;
    RECT 67.89 33.55 68.1 33.62 ;
    RECT 67.89 33.91 68.1 33.98 ;
    RECT 68.35 33.19 68.56 33.26 ;
    RECT 68.35 33.55 68.56 33.62 ;
    RECT 68.35 33.91 68.56 33.98 ;
    RECT 28.05 33.19 28.26 33.26 ;
    RECT 28.05 33.55 28.26 33.62 ;
    RECT 28.05 33.91 28.26 33.98 ;
    RECT 28.51 33.19 28.72 33.26 ;
    RECT 28.51 33.55 28.72 33.62 ;
    RECT 28.51 33.91 28.72 33.98 ;
    RECT 24.73 33.19 24.94 33.26 ;
    RECT 24.73 33.55 24.94 33.62 ;
    RECT 24.73 33.91 24.94 33.98 ;
    RECT 25.19 33.19 25.4 33.26 ;
    RECT 25.19 33.55 25.4 33.62 ;
    RECT 25.19 33.91 25.4 33.98 ;
    RECT 21.41 33.19 21.62 33.26 ;
    RECT 21.41 33.55 21.62 33.62 ;
    RECT 21.41 33.91 21.62 33.98 ;
    RECT 21.87 33.19 22.08 33.26 ;
    RECT 21.87 33.55 22.08 33.62 ;
    RECT 21.87 33.91 22.08 33.98 ;
    RECT 18.09 33.19 18.3 33.26 ;
    RECT 18.09 33.55 18.3 33.62 ;
    RECT 18.09 33.91 18.3 33.98 ;
    RECT 18.55 33.19 18.76 33.26 ;
    RECT 18.55 33.55 18.76 33.62 ;
    RECT 18.55 33.91 18.76 33.98 ;
    RECT 120.825 33.55 120.895 33.62 ;
    RECT 14.77 33.19 14.98 33.26 ;
    RECT 14.77 33.55 14.98 33.62 ;
    RECT 14.77 33.91 14.98 33.98 ;
    RECT 15.23 33.19 15.44 33.26 ;
    RECT 15.23 33.55 15.44 33.62 ;
    RECT 15.23 33.91 15.44 33.98 ;
    RECT 11.45 33.19 11.66 33.26 ;
    RECT 11.45 33.55 11.66 33.62 ;
    RECT 11.45 33.91 11.66 33.98 ;
    RECT 11.91 33.19 12.12 33.26 ;
    RECT 11.91 33.55 12.12 33.62 ;
    RECT 11.91 33.91 12.12 33.98 ;
    RECT 8.13 33.19 8.34 33.26 ;
    RECT 8.13 33.55 8.34 33.62 ;
    RECT 8.13 33.91 8.34 33.98 ;
    RECT 8.59 33.19 8.8 33.26 ;
    RECT 8.59 33.55 8.8 33.62 ;
    RECT 8.59 33.91 8.8 33.98 ;
    RECT 4.81 33.19 5.02 33.26 ;
    RECT 4.81 33.55 5.02 33.62 ;
    RECT 4.81 33.91 5.02 33.98 ;
    RECT 5.27 33.19 5.48 33.26 ;
    RECT 5.27 33.55 5.48 33.62 ;
    RECT 5.27 33.91 5.48 33.98 ;
    RECT 1.49 33.19 1.7 33.26 ;
    RECT 1.49 33.55 1.7 33.62 ;
    RECT 1.49 33.91 1.7 33.98 ;
    RECT 1.95 33.19 2.16 33.26 ;
    RECT 1.95 33.55 2.16 33.62 ;
    RECT 1.95 33.91 2.16 33.98 ;
    RECT 64.57 33.19 64.78 33.26 ;
    RECT 64.57 33.55 64.78 33.62 ;
    RECT 64.57 33.91 64.78 33.98 ;
    RECT 65.03 33.19 65.24 33.26 ;
    RECT 65.03 33.55 65.24 33.62 ;
    RECT 65.03 33.91 65.24 33.98 ;
    RECT 61.25 32.47 61.46 32.54 ;
    RECT 61.25 32.83 61.46 32.9 ;
    RECT 61.25 33.19 61.46 33.26 ;
    RECT 61.71 32.47 61.92 32.54 ;
    RECT 61.71 32.83 61.92 32.9 ;
    RECT 61.71 33.19 61.92 33.26 ;
    RECT 57.93 32.47 58.14 32.54 ;
    RECT 57.93 32.83 58.14 32.9 ;
    RECT 57.93 33.19 58.14 33.26 ;
    RECT 58.39 32.47 58.6 32.54 ;
    RECT 58.39 32.83 58.6 32.9 ;
    RECT 58.39 33.19 58.6 33.26 ;
    RECT 54.61 32.47 54.82 32.54 ;
    RECT 54.61 32.83 54.82 32.9 ;
    RECT 54.61 33.19 54.82 33.26 ;
    RECT 55.07 32.47 55.28 32.54 ;
    RECT 55.07 32.83 55.28 32.9 ;
    RECT 55.07 33.19 55.28 33.26 ;
    RECT 51.29 32.47 51.5 32.54 ;
    RECT 51.29 32.83 51.5 32.9 ;
    RECT 51.29 33.19 51.5 33.26 ;
    RECT 51.75 32.47 51.96 32.54 ;
    RECT 51.75 32.83 51.96 32.9 ;
    RECT 51.75 33.19 51.96 33.26 ;
    RECT 47.97 32.47 48.18 32.54 ;
    RECT 47.97 32.83 48.18 32.9 ;
    RECT 47.97 33.19 48.18 33.26 ;
    RECT 48.43 32.47 48.64 32.54 ;
    RECT 48.43 32.83 48.64 32.9 ;
    RECT 48.43 33.19 48.64 33.26 ;
    RECT 44.65 32.47 44.86 32.54 ;
    RECT 44.65 32.83 44.86 32.9 ;
    RECT 44.65 33.19 44.86 33.26 ;
    RECT 45.11 32.47 45.32 32.54 ;
    RECT 45.11 32.83 45.32 32.9 ;
    RECT 45.11 33.19 45.32 33.26 ;
    RECT 41.33 32.47 41.54 32.54 ;
    RECT 41.33 32.83 41.54 32.9 ;
    RECT 41.33 33.19 41.54 33.26 ;
    RECT 41.79 32.47 42.0 32.54 ;
    RECT 41.79 32.83 42.0 32.9 ;
    RECT 41.79 33.19 42.0 33.26 ;
    RECT 38.01 32.47 38.22 32.54 ;
    RECT 38.01 32.83 38.22 32.9 ;
    RECT 38.01 33.19 38.22 33.26 ;
    RECT 38.47 32.47 38.68 32.54 ;
    RECT 38.47 32.83 38.68 32.9 ;
    RECT 38.47 33.19 38.68 33.26 ;
    RECT 0.4 32.83 0.47 32.9 ;
    RECT 34.69 32.47 34.9 32.54 ;
    RECT 34.69 32.83 34.9 32.9 ;
    RECT 34.69 33.19 34.9 33.26 ;
    RECT 35.15 32.47 35.36 32.54 ;
    RECT 35.15 32.83 35.36 32.9 ;
    RECT 35.15 33.19 35.36 33.26 ;
    RECT 117.69 32.47 117.9 32.54 ;
    RECT 117.69 32.83 117.9 32.9 ;
    RECT 117.69 33.19 117.9 33.26 ;
    RECT 118.15 32.47 118.36 32.54 ;
    RECT 118.15 32.83 118.36 32.9 ;
    RECT 118.15 33.19 118.36 33.26 ;
    RECT 114.37 32.47 114.58 32.54 ;
    RECT 114.37 32.83 114.58 32.9 ;
    RECT 114.37 33.19 114.58 33.26 ;
    RECT 114.83 32.47 115.04 32.54 ;
    RECT 114.83 32.83 115.04 32.9 ;
    RECT 114.83 33.19 115.04 33.26 ;
    RECT 111.05 32.47 111.26 32.54 ;
    RECT 111.05 32.83 111.26 32.9 ;
    RECT 111.05 33.19 111.26 33.26 ;
    RECT 111.51 32.47 111.72 32.54 ;
    RECT 111.51 32.83 111.72 32.9 ;
    RECT 111.51 33.19 111.72 33.26 ;
    RECT 107.73 32.47 107.94 32.54 ;
    RECT 107.73 32.83 107.94 32.9 ;
    RECT 107.73 33.19 107.94 33.26 ;
    RECT 108.19 32.47 108.4 32.54 ;
    RECT 108.19 32.83 108.4 32.9 ;
    RECT 108.19 33.19 108.4 33.26 ;
    RECT 104.41 32.47 104.62 32.54 ;
    RECT 104.41 32.83 104.62 32.9 ;
    RECT 104.41 33.19 104.62 33.26 ;
    RECT 104.87 32.47 105.08 32.54 ;
    RECT 104.87 32.83 105.08 32.9 ;
    RECT 104.87 33.19 105.08 33.26 ;
    RECT 101.09 32.47 101.3 32.54 ;
    RECT 101.09 32.83 101.3 32.9 ;
    RECT 101.09 33.19 101.3 33.26 ;
    RECT 101.55 32.47 101.76 32.54 ;
    RECT 101.55 32.83 101.76 32.9 ;
    RECT 101.55 33.19 101.76 33.26 ;
    RECT 97.77 32.47 97.98 32.54 ;
    RECT 97.77 32.83 97.98 32.9 ;
    RECT 97.77 33.19 97.98 33.26 ;
    RECT 98.23 32.47 98.44 32.54 ;
    RECT 98.23 32.83 98.44 32.9 ;
    RECT 98.23 33.19 98.44 33.26 ;
    RECT 94.45 32.47 94.66 32.54 ;
    RECT 94.45 32.83 94.66 32.9 ;
    RECT 94.45 33.19 94.66 33.26 ;
    RECT 94.91 32.47 95.12 32.54 ;
    RECT 94.91 32.83 95.12 32.9 ;
    RECT 94.91 33.19 95.12 33.26 ;
    RECT 91.13 32.47 91.34 32.54 ;
    RECT 91.13 32.83 91.34 32.9 ;
    RECT 91.13 33.19 91.34 33.26 ;
    RECT 91.59 32.47 91.8 32.54 ;
    RECT 91.59 32.83 91.8 32.9 ;
    RECT 91.59 33.19 91.8 33.26 ;
    RECT 87.81 32.47 88.02 32.54 ;
    RECT 87.81 32.83 88.02 32.9 ;
    RECT 87.81 33.19 88.02 33.26 ;
    RECT 88.27 32.47 88.48 32.54 ;
    RECT 88.27 32.83 88.48 32.9 ;
    RECT 88.27 33.19 88.48 33.26 ;
    RECT 84.49 32.47 84.7 32.54 ;
    RECT 84.49 32.83 84.7 32.9 ;
    RECT 84.49 33.19 84.7 33.26 ;
    RECT 84.95 32.47 85.16 32.54 ;
    RECT 84.95 32.83 85.16 32.9 ;
    RECT 84.95 33.19 85.16 33.26 ;
    RECT 81.17 32.47 81.38 32.54 ;
    RECT 81.17 32.83 81.38 32.9 ;
    RECT 81.17 33.19 81.38 33.26 ;
    RECT 81.63 32.47 81.84 32.54 ;
    RECT 81.63 32.83 81.84 32.9 ;
    RECT 81.63 33.19 81.84 33.26 ;
    RECT 77.85 32.47 78.06 32.54 ;
    RECT 77.85 32.83 78.06 32.9 ;
    RECT 77.85 33.19 78.06 33.26 ;
    RECT 78.31 32.47 78.52 32.54 ;
    RECT 78.31 32.83 78.52 32.9 ;
    RECT 78.31 33.19 78.52 33.26 ;
    RECT 74.53 32.47 74.74 32.54 ;
    RECT 74.53 32.83 74.74 32.9 ;
    RECT 74.53 33.19 74.74 33.26 ;
    RECT 74.99 32.47 75.2 32.54 ;
    RECT 74.99 32.83 75.2 32.9 ;
    RECT 74.99 33.19 75.2 33.26 ;
    RECT 71.21 32.47 71.42 32.54 ;
    RECT 71.21 32.83 71.42 32.9 ;
    RECT 71.21 33.19 71.42 33.26 ;
    RECT 71.67 32.47 71.88 32.54 ;
    RECT 71.67 32.83 71.88 32.9 ;
    RECT 71.67 33.19 71.88 33.26 ;
    RECT 31.37 32.47 31.58 32.54 ;
    RECT 31.37 32.83 31.58 32.9 ;
    RECT 31.37 33.19 31.58 33.26 ;
    RECT 31.83 32.47 32.04 32.54 ;
    RECT 31.83 32.83 32.04 32.9 ;
    RECT 31.83 33.19 32.04 33.26 ;
    RECT 67.89 32.47 68.1 32.54 ;
    RECT 67.89 32.83 68.1 32.9 ;
    RECT 67.89 33.19 68.1 33.26 ;
    RECT 68.35 32.47 68.56 32.54 ;
    RECT 68.35 32.83 68.56 32.9 ;
    RECT 68.35 33.19 68.56 33.26 ;
    RECT 28.05 32.47 28.26 32.54 ;
    RECT 28.05 32.83 28.26 32.9 ;
    RECT 28.05 33.19 28.26 33.26 ;
    RECT 28.51 32.47 28.72 32.54 ;
    RECT 28.51 32.83 28.72 32.9 ;
    RECT 28.51 33.19 28.72 33.26 ;
    RECT 24.73 32.47 24.94 32.54 ;
    RECT 24.73 32.83 24.94 32.9 ;
    RECT 24.73 33.19 24.94 33.26 ;
    RECT 25.19 32.47 25.4 32.54 ;
    RECT 25.19 32.83 25.4 32.9 ;
    RECT 25.19 33.19 25.4 33.26 ;
    RECT 21.41 32.47 21.62 32.54 ;
    RECT 21.41 32.83 21.62 32.9 ;
    RECT 21.41 33.19 21.62 33.26 ;
    RECT 21.87 32.47 22.08 32.54 ;
    RECT 21.87 32.83 22.08 32.9 ;
    RECT 21.87 33.19 22.08 33.26 ;
    RECT 18.09 32.47 18.3 32.54 ;
    RECT 18.09 32.83 18.3 32.9 ;
    RECT 18.09 33.19 18.3 33.26 ;
    RECT 18.55 32.47 18.76 32.54 ;
    RECT 18.55 32.83 18.76 32.9 ;
    RECT 18.55 33.19 18.76 33.26 ;
    RECT 120.825 32.83 120.895 32.9 ;
    RECT 14.77 32.47 14.98 32.54 ;
    RECT 14.77 32.83 14.98 32.9 ;
    RECT 14.77 33.19 14.98 33.26 ;
    RECT 15.23 32.47 15.44 32.54 ;
    RECT 15.23 32.83 15.44 32.9 ;
    RECT 15.23 33.19 15.44 33.26 ;
    RECT 11.45 32.47 11.66 32.54 ;
    RECT 11.45 32.83 11.66 32.9 ;
    RECT 11.45 33.19 11.66 33.26 ;
    RECT 11.91 32.47 12.12 32.54 ;
    RECT 11.91 32.83 12.12 32.9 ;
    RECT 11.91 33.19 12.12 33.26 ;
    RECT 8.13 32.47 8.34 32.54 ;
    RECT 8.13 32.83 8.34 32.9 ;
    RECT 8.13 33.19 8.34 33.26 ;
    RECT 8.59 32.47 8.8 32.54 ;
    RECT 8.59 32.83 8.8 32.9 ;
    RECT 8.59 33.19 8.8 33.26 ;
    RECT 4.81 32.47 5.02 32.54 ;
    RECT 4.81 32.83 5.02 32.9 ;
    RECT 4.81 33.19 5.02 33.26 ;
    RECT 5.27 32.47 5.48 32.54 ;
    RECT 5.27 32.83 5.48 32.9 ;
    RECT 5.27 33.19 5.48 33.26 ;
    RECT 1.49 32.47 1.7 32.54 ;
    RECT 1.49 32.83 1.7 32.9 ;
    RECT 1.49 33.19 1.7 33.26 ;
    RECT 1.95 32.47 2.16 32.54 ;
    RECT 1.95 32.83 2.16 32.9 ;
    RECT 1.95 33.19 2.16 33.26 ;
    RECT 64.57 32.47 64.78 32.54 ;
    RECT 64.57 32.83 64.78 32.9 ;
    RECT 64.57 33.19 64.78 33.26 ;
    RECT 65.03 32.47 65.24 32.54 ;
    RECT 65.03 32.83 65.24 32.9 ;
    RECT 65.03 33.19 65.24 33.26 ;
    RECT 61.25 72.09 61.46 72.16 ;
    RECT 61.25 72.45 61.46 72.52 ;
    RECT 61.25 72.81 61.46 72.88 ;
    RECT 61.71 72.09 61.92 72.16 ;
    RECT 61.71 72.45 61.92 72.52 ;
    RECT 61.71 72.81 61.92 72.88 ;
    RECT 57.93 72.09 58.14 72.16 ;
    RECT 57.93 72.45 58.14 72.52 ;
    RECT 57.93 72.81 58.14 72.88 ;
    RECT 58.39 72.09 58.6 72.16 ;
    RECT 58.39 72.45 58.6 72.52 ;
    RECT 58.39 72.81 58.6 72.88 ;
    RECT 54.61 72.09 54.82 72.16 ;
    RECT 54.61 72.45 54.82 72.52 ;
    RECT 54.61 72.81 54.82 72.88 ;
    RECT 55.07 72.09 55.28 72.16 ;
    RECT 55.07 72.45 55.28 72.52 ;
    RECT 55.07 72.81 55.28 72.88 ;
    RECT 51.29 72.09 51.5 72.16 ;
    RECT 51.29 72.45 51.5 72.52 ;
    RECT 51.29 72.81 51.5 72.88 ;
    RECT 51.75 72.09 51.96 72.16 ;
    RECT 51.75 72.45 51.96 72.52 ;
    RECT 51.75 72.81 51.96 72.88 ;
    RECT 47.97 72.09 48.18 72.16 ;
    RECT 47.97 72.45 48.18 72.52 ;
    RECT 47.97 72.81 48.18 72.88 ;
    RECT 48.43 72.09 48.64 72.16 ;
    RECT 48.43 72.45 48.64 72.52 ;
    RECT 48.43 72.81 48.64 72.88 ;
    RECT 44.65 72.09 44.86 72.16 ;
    RECT 44.65 72.45 44.86 72.52 ;
    RECT 44.65 72.81 44.86 72.88 ;
    RECT 45.11 72.09 45.32 72.16 ;
    RECT 45.11 72.45 45.32 72.52 ;
    RECT 45.11 72.81 45.32 72.88 ;
    RECT 41.33 72.09 41.54 72.16 ;
    RECT 41.33 72.45 41.54 72.52 ;
    RECT 41.33 72.81 41.54 72.88 ;
    RECT 41.79 72.09 42.0 72.16 ;
    RECT 41.79 72.45 42.0 72.52 ;
    RECT 41.79 72.81 42.0 72.88 ;
    RECT 38.01 72.09 38.22 72.16 ;
    RECT 38.01 72.45 38.22 72.52 ;
    RECT 38.01 72.81 38.22 72.88 ;
    RECT 38.47 72.09 38.68 72.16 ;
    RECT 38.47 72.45 38.68 72.52 ;
    RECT 38.47 72.81 38.68 72.88 ;
    RECT 0.4 72.45 0.47 72.52 ;
    RECT 34.69 72.09 34.9 72.16 ;
    RECT 34.69 72.45 34.9 72.52 ;
    RECT 34.69 72.81 34.9 72.88 ;
    RECT 35.15 72.09 35.36 72.16 ;
    RECT 35.15 72.45 35.36 72.52 ;
    RECT 35.15 72.81 35.36 72.88 ;
    RECT 117.69 72.09 117.9 72.16 ;
    RECT 117.69 72.45 117.9 72.52 ;
    RECT 117.69 72.81 117.9 72.88 ;
    RECT 118.15 72.09 118.36 72.16 ;
    RECT 118.15 72.45 118.36 72.52 ;
    RECT 118.15 72.81 118.36 72.88 ;
    RECT 114.37 72.09 114.58 72.16 ;
    RECT 114.37 72.45 114.58 72.52 ;
    RECT 114.37 72.81 114.58 72.88 ;
    RECT 114.83 72.09 115.04 72.16 ;
    RECT 114.83 72.45 115.04 72.52 ;
    RECT 114.83 72.81 115.04 72.88 ;
    RECT 111.05 72.09 111.26 72.16 ;
    RECT 111.05 72.45 111.26 72.52 ;
    RECT 111.05 72.81 111.26 72.88 ;
    RECT 111.51 72.09 111.72 72.16 ;
    RECT 111.51 72.45 111.72 72.52 ;
    RECT 111.51 72.81 111.72 72.88 ;
    RECT 107.73 72.09 107.94 72.16 ;
    RECT 107.73 72.45 107.94 72.52 ;
    RECT 107.73 72.81 107.94 72.88 ;
    RECT 108.19 72.09 108.4 72.16 ;
    RECT 108.19 72.45 108.4 72.52 ;
    RECT 108.19 72.81 108.4 72.88 ;
    RECT 104.41 72.09 104.62 72.16 ;
    RECT 104.41 72.45 104.62 72.52 ;
    RECT 104.41 72.81 104.62 72.88 ;
    RECT 104.87 72.09 105.08 72.16 ;
    RECT 104.87 72.45 105.08 72.52 ;
    RECT 104.87 72.81 105.08 72.88 ;
    RECT 101.09 72.09 101.3 72.16 ;
    RECT 101.09 72.45 101.3 72.52 ;
    RECT 101.09 72.81 101.3 72.88 ;
    RECT 101.55 72.09 101.76 72.16 ;
    RECT 101.55 72.45 101.76 72.52 ;
    RECT 101.55 72.81 101.76 72.88 ;
    RECT 97.77 72.09 97.98 72.16 ;
    RECT 97.77 72.45 97.98 72.52 ;
    RECT 97.77 72.81 97.98 72.88 ;
    RECT 98.23 72.09 98.44 72.16 ;
    RECT 98.23 72.45 98.44 72.52 ;
    RECT 98.23 72.81 98.44 72.88 ;
    RECT 94.45 72.09 94.66 72.16 ;
    RECT 94.45 72.45 94.66 72.52 ;
    RECT 94.45 72.81 94.66 72.88 ;
    RECT 94.91 72.09 95.12 72.16 ;
    RECT 94.91 72.45 95.12 72.52 ;
    RECT 94.91 72.81 95.12 72.88 ;
    RECT 91.13 72.09 91.34 72.16 ;
    RECT 91.13 72.45 91.34 72.52 ;
    RECT 91.13 72.81 91.34 72.88 ;
    RECT 91.59 72.09 91.8 72.16 ;
    RECT 91.59 72.45 91.8 72.52 ;
    RECT 91.59 72.81 91.8 72.88 ;
    RECT 87.81 72.09 88.02 72.16 ;
    RECT 87.81 72.45 88.02 72.52 ;
    RECT 87.81 72.81 88.02 72.88 ;
    RECT 88.27 72.09 88.48 72.16 ;
    RECT 88.27 72.45 88.48 72.52 ;
    RECT 88.27 72.81 88.48 72.88 ;
    RECT 84.49 72.09 84.7 72.16 ;
    RECT 84.49 72.45 84.7 72.52 ;
    RECT 84.49 72.81 84.7 72.88 ;
    RECT 84.95 72.09 85.16 72.16 ;
    RECT 84.95 72.45 85.16 72.52 ;
    RECT 84.95 72.81 85.16 72.88 ;
    RECT 81.17 72.09 81.38 72.16 ;
    RECT 81.17 72.45 81.38 72.52 ;
    RECT 81.17 72.81 81.38 72.88 ;
    RECT 81.63 72.09 81.84 72.16 ;
    RECT 81.63 72.45 81.84 72.52 ;
    RECT 81.63 72.81 81.84 72.88 ;
    RECT 77.85 72.09 78.06 72.16 ;
    RECT 77.85 72.45 78.06 72.52 ;
    RECT 77.85 72.81 78.06 72.88 ;
    RECT 78.31 72.09 78.52 72.16 ;
    RECT 78.31 72.45 78.52 72.52 ;
    RECT 78.31 72.81 78.52 72.88 ;
    RECT 74.53 72.09 74.74 72.16 ;
    RECT 74.53 72.45 74.74 72.52 ;
    RECT 74.53 72.81 74.74 72.88 ;
    RECT 74.99 72.09 75.2 72.16 ;
    RECT 74.99 72.45 75.2 72.52 ;
    RECT 74.99 72.81 75.2 72.88 ;
    RECT 71.21 72.09 71.42 72.16 ;
    RECT 71.21 72.45 71.42 72.52 ;
    RECT 71.21 72.81 71.42 72.88 ;
    RECT 71.67 72.09 71.88 72.16 ;
    RECT 71.67 72.45 71.88 72.52 ;
    RECT 71.67 72.81 71.88 72.88 ;
    RECT 31.37 72.09 31.58 72.16 ;
    RECT 31.37 72.45 31.58 72.52 ;
    RECT 31.37 72.81 31.58 72.88 ;
    RECT 31.83 72.09 32.04 72.16 ;
    RECT 31.83 72.45 32.04 72.52 ;
    RECT 31.83 72.81 32.04 72.88 ;
    RECT 67.89 72.09 68.1 72.16 ;
    RECT 67.89 72.45 68.1 72.52 ;
    RECT 67.89 72.81 68.1 72.88 ;
    RECT 68.35 72.09 68.56 72.16 ;
    RECT 68.35 72.45 68.56 72.52 ;
    RECT 68.35 72.81 68.56 72.88 ;
    RECT 28.05 72.09 28.26 72.16 ;
    RECT 28.05 72.45 28.26 72.52 ;
    RECT 28.05 72.81 28.26 72.88 ;
    RECT 28.51 72.09 28.72 72.16 ;
    RECT 28.51 72.45 28.72 72.52 ;
    RECT 28.51 72.81 28.72 72.88 ;
    RECT 24.73 72.09 24.94 72.16 ;
    RECT 24.73 72.45 24.94 72.52 ;
    RECT 24.73 72.81 24.94 72.88 ;
    RECT 25.19 72.09 25.4 72.16 ;
    RECT 25.19 72.45 25.4 72.52 ;
    RECT 25.19 72.81 25.4 72.88 ;
    RECT 21.41 72.09 21.62 72.16 ;
    RECT 21.41 72.45 21.62 72.52 ;
    RECT 21.41 72.81 21.62 72.88 ;
    RECT 21.87 72.09 22.08 72.16 ;
    RECT 21.87 72.45 22.08 72.52 ;
    RECT 21.87 72.81 22.08 72.88 ;
    RECT 18.09 72.09 18.3 72.16 ;
    RECT 18.09 72.45 18.3 72.52 ;
    RECT 18.09 72.81 18.3 72.88 ;
    RECT 18.55 72.09 18.76 72.16 ;
    RECT 18.55 72.45 18.76 72.52 ;
    RECT 18.55 72.81 18.76 72.88 ;
    RECT 120.825 72.45 120.895 72.52 ;
    RECT 14.77 72.09 14.98 72.16 ;
    RECT 14.77 72.45 14.98 72.52 ;
    RECT 14.77 72.81 14.98 72.88 ;
    RECT 15.23 72.09 15.44 72.16 ;
    RECT 15.23 72.45 15.44 72.52 ;
    RECT 15.23 72.81 15.44 72.88 ;
    RECT 11.45 72.09 11.66 72.16 ;
    RECT 11.45 72.45 11.66 72.52 ;
    RECT 11.45 72.81 11.66 72.88 ;
    RECT 11.91 72.09 12.12 72.16 ;
    RECT 11.91 72.45 12.12 72.52 ;
    RECT 11.91 72.81 12.12 72.88 ;
    RECT 8.13 72.09 8.34 72.16 ;
    RECT 8.13 72.45 8.34 72.52 ;
    RECT 8.13 72.81 8.34 72.88 ;
    RECT 8.59 72.09 8.8 72.16 ;
    RECT 8.59 72.45 8.8 72.52 ;
    RECT 8.59 72.81 8.8 72.88 ;
    RECT 4.81 72.09 5.02 72.16 ;
    RECT 4.81 72.45 5.02 72.52 ;
    RECT 4.81 72.81 5.02 72.88 ;
    RECT 5.27 72.09 5.48 72.16 ;
    RECT 5.27 72.45 5.48 72.52 ;
    RECT 5.27 72.81 5.48 72.88 ;
    RECT 1.49 72.09 1.7 72.16 ;
    RECT 1.49 72.45 1.7 72.52 ;
    RECT 1.49 72.81 1.7 72.88 ;
    RECT 1.95 72.09 2.16 72.16 ;
    RECT 1.95 72.45 2.16 72.52 ;
    RECT 1.95 72.81 2.16 72.88 ;
    RECT 64.57 72.09 64.78 72.16 ;
    RECT 64.57 72.45 64.78 72.52 ;
    RECT 64.57 72.81 64.78 72.88 ;
    RECT 65.03 72.09 65.24 72.16 ;
    RECT 65.03 72.45 65.24 72.52 ;
    RECT 65.03 72.81 65.24 72.88 ;
    RECT 61.25 31.75 61.46 31.82 ;
    RECT 61.25 32.11 61.46 32.18 ;
    RECT 61.25 32.47 61.46 32.54 ;
    RECT 61.71 31.75 61.92 31.82 ;
    RECT 61.71 32.11 61.92 32.18 ;
    RECT 61.71 32.47 61.92 32.54 ;
    RECT 57.93 31.75 58.14 31.82 ;
    RECT 57.93 32.11 58.14 32.18 ;
    RECT 57.93 32.47 58.14 32.54 ;
    RECT 58.39 31.75 58.6 31.82 ;
    RECT 58.39 32.11 58.6 32.18 ;
    RECT 58.39 32.47 58.6 32.54 ;
    RECT 54.61 31.75 54.82 31.82 ;
    RECT 54.61 32.11 54.82 32.18 ;
    RECT 54.61 32.47 54.82 32.54 ;
    RECT 55.07 31.75 55.28 31.82 ;
    RECT 55.07 32.11 55.28 32.18 ;
    RECT 55.07 32.47 55.28 32.54 ;
    RECT 51.29 31.75 51.5 31.82 ;
    RECT 51.29 32.11 51.5 32.18 ;
    RECT 51.29 32.47 51.5 32.54 ;
    RECT 51.75 31.75 51.96 31.82 ;
    RECT 51.75 32.11 51.96 32.18 ;
    RECT 51.75 32.47 51.96 32.54 ;
    RECT 47.97 31.75 48.18 31.82 ;
    RECT 47.97 32.11 48.18 32.18 ;
    RECT 47.97 32.47 48.18 32.54 ;
    RECT 48.43 31.75 48.64 31.82 ;
    RECT 48.43 32.11 48.64 32.18 ;
    RECT 48.43 32.47 48.64 32.54 ;
    RECT 44.65 31.75 44.86 31.82 ;
    RECT 44.65 32.11 44.86 32.18 ;
    RECT 44.65 32.47 44.86 32.54 ;
    RECT 45.11 31.75 45.32 31.82 ;
    RECT 45.11 32.11 45.32 32.18 ;
    RECT 45.11 32.47 45.32 32.54 ;
    RECT 41.33 31.75 41.54 31.82 ;
    RECT 41.33 32.11 41.54 32.18 ;
    RECT 41.33 32.47 41.54 32.54 ;
    RECT 41.79 31.75 42.0 31.82 ;
    RECT 41.79 32.11 42.0 32.18 ;
    RECT 41.79 32.47 42.0 32.54 ;
    RECT 38.01 31.75 38.22 31.82 ;
    RECT 38.01 32.11 38.22 32.18 ;
    RECT 38.01 32.47 38.22 32.54 ;
    RECT 38.47 31.75 38.68 31.82 ;
    RECT 38.47 32.11 38.68 32.18 ;
    RECT 38.47 32.47 38.68 32.54 ;
    RECT 0.4 32.11 0.47 32.18 ;
    RECT 34.69 31.75 34.9 31.82 ;
    RECT 34.69 32.11 34.9 32.18 ;
    RECT 34.69 32.47 34.9 32.54 ;
    RECT 35.15 31.75 35.36 31.82 ;
    RECT 35.15 32.11 35.36 32.18 ;
    RECT 35.15 32.47 35.36 32.54 ;
    RECT 117.69 31.75 117.9 31.82 ;
    RECT 117.69 32.11 117.9 32.18 ;
    RECT 117.69 32.47 117.9 32.54 ;
    RECT 118.15 31.75 118.36 31.82 ;
    RECT 118.15 32.11 118.36 32.18 ;
    RECT 118.15 32.47 118.36 32.54 ;
    RECT 114.37 31.75 114.58 31.82 ;
    RECT 114.37 32.11 114.58 32.18 ;
    RECT 114.37 32.47 114.58 32.54 ;
    RECT 114.83 31.75 115.04 31.82 ;
    RECT 114.83 32.11 115.04 32.18 ;
    RECT 114.83 32.47 115.04 32.54 ;
    RECT 111.05 31.75 111.26 31.82 ;
    RECT 111.05 32.11 111.26 32.18 ;
    RECT 111.05 32.47 111.26 32.54 ;
    RECT 111.51 31.75 111.72 31.82 ;
    RECT 111.51 32.11 111.72 32.18 ;
    RECT 111.51 32.47 111.72 32.54 ;
    RECT 107.73 31.75 107.94 31.82 ;
    RECT 107.73 32.11 107.94 32.18 ;
    RECT 107.73 32.47 107.94 32.54 ;
    RECT 108.19 31.75 108.4 31.82 ;
    RECT 108.19 32.11 108.4 32.18 ;
    RECT 108.19 32.47 108.4 32.54 ;
    RECT 104.41 31.75 104.62 31.82 ;
    RECT 104.41 32.11 104.62 32.18 ;
    RECT 104.41 32.47 104.62 32.54 ;
    RECT 104.87 31.75 105.08 31.82 ;
    RECT 104.87 32.11 105.08 32.18 ;
    RECT 104.87 32.47 105.08 32.54 ;
    RECT 101.09 31.75 101.3 31.82 ;
    RECT 101.09 32.11 101.3 32.18 ;
    RECT 101.09 32.47 101.3 32.54 ;
    RECT 101.55 31.75 101.76 31.82 ;
    RECT 101.55 32.11 101.76 32.18 ;
    RECT 101.55 32.47 101.76 32.54 ;
    RECT 97.77 31.75 97.98 31.82 ;
    RECT 97.77 32.11 97.98 32.18 ;
    RECT 97.77 32.47 97.98 32.54 ;
    RECT 98.23 31.75 98.44 31.82 ;
    RECT 98.23 32.11 98.44 32.18 ;
    RECT 98.23 32.47 98.44 32.54 ;
    RECT 94.45 31.75 94.66 31.82 ;
    RECT 94.45 32.11 94.66 32.18 ;
    RECT 94.45 32.47 94.66 32.54 ;
    RECT 94.91 31.75 95.12 31.82 ;
    RECT 94.91 32.11 95.12 32.18 ;
    RECT 94.91 32.47 95.12 32.54 ;
    RECT 91.13 31.75 91.34 31.82 ;
    RECT 91.13 32.11 91.34 32.18 ;
    RECT 91.13 32.47 91.34 32.54 ;
    RECT 91.59 31.75 91.8 31.82 ;
    RECT 91.59 32.11 91.8 32.18 ;
    RECT 91.59 32.47 91.8 32.54 ;
    RECT 87.81 31.75 88.02 31.82 ;
    RECT 87.81 32.11 88.02 32.18 ;
    RECT 87.81 32.47 88.02 32.54 ;
    RECT 88.27 31.75 88.48 31.82 ;
    RECT 88.27 32.11 88.48 32.18 ;
    RECT 88.27 32.47 88.48 32.54 ;
    RECT 84.49 31.75 84.7 31.82 ;
    RECT 84.49 32.11 84.7 32.18 ;
    RECT 84.49 32.47 84.7 32.54 ;
    RECT 84.95 31.75 85.16 31.82 ;
    RECT 84.95 32.11 85.16 32.18 ;
    RECT 84.95 32.47 85.16 32.54 ;
    RECT 81.17 31.75 81.38 31.82 ;
    RECT 81.17 32.11 81.38 32.18 ;
    RECT 81.17 32.47 81.38 32.54 ;
    RECT 81.63 31.75 81.84 31.82 ;
    RECT 81.63 32.11 81.84 32.18 ;
    RECT 81.63 32.47 81.84 32.54 ;
    RECT 77.85 31.75 78.06 31.82 ;
    RECT 77.85 32.11 78.06 32.18 ;
    RECT 77.85 32.47 78.06 32.54 ;
    RECT 78.31 31.75 78.52 31.82 ;
    RECT 78.31 32.11 78.52 32.18 ;
    RECT 78.31 32.47 78.52 32.54 ;
    RECT 74.53 31.75 74.74 31.82 ;
    RECT 74.53 32.11 74.74 32.18 ;
    RECT 74.53 32.47 74.74 32.54 ;
    RECT 74.99 31.75 75.2 31.82 ;
    RECT 74.99 32.11 75.2 32.18 ;
    RECT 74.99 32.47 75.2 32.54 ;
    RECT 71.21 31.75 71.42 31.82 ;
    RECT 71.21 32.11 71.42 32.18 ;
    RECT 71.21 32.47 71.42 32.54 ;
    RECT 71.67 31.75 71.88 31.82 ;
    RECT 71.67 32.11 71.88 32.18 ;
    RECT 71.67 32.47 71.88 32.54 ;
    RECT 31.37 31.75 31.58 31.82 ;
    RECT 31.37 32.11 31.58 32.18 ;
    RECT 31.37 32.47 31.58 32.54 ;
    RECT 31.83 31.75 32.04 31.82 ;
    RECT 31.83 32.11 32.04 32.18 ;
    RECT 31.83 32.47 32.04 32.54 ;
    RECT 67.89 31.75 68.1 31.82 ;
    RECT 67.89 32.11 68.1 32.18 ;
    RECT 67.89 32.47 68.1 32.54 ;
    RECT 68.35 31.75 68.56 31.82 ;
    RECT 68.35 32.11 68.56 32.18 ;
    RECT 68.35 32.47 68.56 32.54 ;
    RECT 28.05 31.75 28.26 31.82 ;
    RECT 28.05 32.11 28.26 32.18 ;
    RECT 28.05 32.47 28.26 32.54 ;
    RECT 28.51 31.75 28.72 31.82 ;
    RECT 28.51 32.11 28.72 32.18 ;
    RECT 28.51 32.47 28.72 32.54 ;
    RECT 24.73 31.75 24.94 31.82 ;
    RECT 24.73 32.11 24.94 32.18 ;
    RECT 24.73 32.47 24.94 32.54 ;
    RECT 25.19 31.75 25.4 31.82 ;
    RECT 25.19 32.11 25.4 32.18 ;
    RECT 25.19 32.47 25.4 32.54 ;
    RECT 21.41 31.75 21.62 31.82 ;
    RECT 21.41 32.11 21.62 32.18 ;
    RECT 21.41 32.47 21.62 32.54 ;
    RECT 21.87 31.75 22.08 31.82 ;
    RECT 21.87 32.11 22.08 32.18 ;
    RECT 21.87 32.47 22.08 32.54 ;
    RECT 18.09 31.75 18.3 31.82 ;
    RECT 18.09 32.11 18.3 32.18 ;
    RECT 18.09 32.47 18.3 32.54 ;
    RECT 18.55 31.75 18.76 31.82 ;
    RECT 18.55 32.11 18.76 32.18 ;
    RECT 18.55 32.47 18.76 32.54 ;
    RECT 120.825 32.11 120.895 32.18 ;
    RECT 14.77 31.75 14.98 31.82 ;
    RECT 14.77 32.11 14.98 32.18 ;
    RECT 14.77 32.47 14.98 32.54 ;
    RECT 15.23 31.75 15.44 31.82 ;
    RECT 15.23 32.11 15.44 32.18 ;
    RECT 15.23 32.47 15.44 32.54 ;
    RECT 11.45 31.75 11.66 31.82 ;
    RECT 11.45 32.11 11.66 32.18 ;
    RECT 11.45 32.47 11.66 32.54 ;
    RECT 11.91 31.75 12.12 31.82 ;
    RECT 11.91 32.11 12.12 32.18 ;
    RECT 11.91 32.47 12.12 32.54 ;
    RECT 8.13 31.75 8.34 31.82 ;
    RECT 8.13 32.11 8.34 32.18 ;
    RECT 8.13 32.47 8.34 32.54 ;
    RECT 8.59 31.75 8.8 31.82 ;
    RECT 8.59 32.11 8.8 32.18 ;
    RECT 8.59 32.47 8.8 32.54 ;
    RECT 4.81 31.75 5.02 31.82 ;
    RECT 4.81 32.11 5.02 32.18 ;
    RECT 4.81 32.47 5.02 32.54 ;
    RECT 5.27 31.75 5.48 31.82 ;
    RECT 5.27 32.11 5.48 32.18 ;
    RECT 5.27 32.47 5.48 32.54 ;
    RECT 1.49 31.75 1.7 31.82 ;
    RECT 1.49 32.11 1.7 32.18 ;
    RECT 1.49 32.47 1.7 32.54 ;
    RECT 1.95 31.75 2.16 31.82 ;
    RECT 1.95 32.11 2.16 32.18 ;
    RECT 1.95 32.47 2.16 32.54 ;
    RECT 64.57 31.75 64.78 31.82 ;
    RECT 64.57 32.11 64.78 32.18 ;
    RECT 64.57 32.47 64.78 32.54 ;
    RECT 65.03 31.75 65.24 31.82 ;
    RECT 65.03 32.11 65.24 32.18 ;
    RECT 65.03 32.47 65.24 32.54 ;
    RECT 61.25 71.37 61.46 71.44 ;
    RECT 61.25 71.73 61.46 71.8 ;
    RECT 61.25 72.09 61.46 72.16 ;
    RECT 61.71 71.37 61.92 71.44 ;
    RECT 61.71 71.73 61.92 71.8 ;
    RECT 61.71 72.09 61.92 72.16 ;
    RECT 57.93 71.37 58.14 71.44 ;
    RECT 57.93 71.73 58.14 71.8 ;
    RECT 57.93 72.09 58.14 72.16 ;
    RECT 58.39 71.37 58.6 71.44 ;
    RECT 58.39 71.73 58.6 71.8 ;
    RECT 58.39 72.09 58.6 72.16 ;
    RECT 54.61 71.37 54.82 71.44 ;
    RECT 54.61 71.73 54.82 71.8 ;
    RECT 54.61 72.09 54.82 72.16 ;
    RECT 55.07 71.37 55.28 71.44 ;
    RECT 55.07 71.73 55.28 71.8 ;
    RECT 55.07 72.09 55.28 72.16 ;
    RECT 51.29 71.37 51.5 71.44 ;
    RECT 51.29 71.73 51.5 71.8 ;
    RECT 51.29 72.09 51.5 72.16 ;
    RECT 51.75 71.37 51.96 71.44 ;
    RECT 51.75 71.73 51.96 71.8 ;
    RECT 51.75 72.09 51.96 72.16 ;
    RECT 47.97 71.37 48.18 71.44 ;
    RECT 47.97 71.73 48.18 71.8 ;
    RECT 47.97 72.09 48.18 72.16 ;
    RECT 48.43 71.37 48.64 71.44 ;
    RECT 48.43 71.73 48.64 71.8 ;
    RECT 48.43 72.09 48.64 72.16 ;
    RECT 44.65 71.37 44.86 71.44 ;
    RECT 44.65 71.73 44.86 71.8 ;
    RECT 44.65 72.09 44.86 72.16 ;
    RECT 45.11 71.37 45.32 71.44 ;
    RECT 45.11 71.73 45.32 71.8 ;
    RECT 45.11 72.09 45.32 72.16 ;
    RECT 41.33 71.37 41.54 71.44 ;
    RECT 41.33 71.73 41.54 71.8 ;
    RECT 41.33 72.09 41.54 72.16 ;
    RECT 41.79 71.37 42.0 71.44 ;
    RECT 41.79 71.73 42.0 71.8 ;
    RECT 41.79 72.09 42.0 72.16 ;
    RECT 38.01 71.37 38.22 71.44 ;
    RECT 38.01 71.73 38.22 71.8 ;
    RECT 38.01 72.09 38.22 72.16 ;
    RECT 38.47 71.37 38.68 71.44 ;
    RECT 38.47 71.73 38.68 71.8 ;
    RECT 38.47 72.09 38.68 72.16 ;
    RECT 0.4 71.73 0.47 71.8 ;
    RECT 34.69 71.37 34.9 71.44 ;
    RECT 34.69 71.73 34.9 71.8 ;
    RECT 34.69 72.09 34.9 72.16 ;
    RECT 35.15 71.37 35.36 71.44 ;
    RECT 35.15 71.73 35.36 71.8 ;
    RECT 35.15 72.09 35.36 72.16 ;
    RECT 117.69 71.37 117.9 71.44 ;
    RECT 117.69 71.73 117.9 71.8 ;
    RECT 117.69 72.09 117.9 72.16 ;
    RECT 118.15 71.37 118.36 71.44 ;
    RECT 118.15 71.73 118.36 71.8 ;
    RECT 118.15 72.09 118.36 72.16 ;
    RECT 114.37 71.37 114.58 71.44 ;
    RECT 114.37 71.73 114.58 71.8 ;
    RECT 114.37 72.09 114.58 72.16 ;
    RECT 114.83 71.37 115.04 71.44 ;
    RECT 114.83 71.73 115.04 71.8 ;
    RECT 114.83 72.09 115.04 72.16 ;
    RECT 111.05 71.37 111.26 71.44 ;
    RECT 111.05 71.73 111.26 71.8 ;
    RECT 111.05 72.09 111.26 72.16 ;
    RECT 111.51 71.37 111.72 71.44 ;
    RECT 111.51 71.73 111.72 71.8 ;
    RECT 111.51 72.09 111.72 72.16 ;
    RECT 107.73 71.37 107.94 71.44 ;
    RECT 107.73 71.73 107.94 71.8 ;
    RECT 107.73 72.09 107.94 72.16 ;
    RECT 108.19 71.37 108.4 71.44 ;
    RECT 108.19 71.73 108.4 71.8 ;
    RECT 108.19 72.09 108.4 72.16 ;
    RECT 104.41 71.37 104.62 71.44 ;
    RECT 104.41 71.73 104.62 71.8 ;
    RECT 104.41 72.09 104.62 72.16 ;
    RECT 104.87 71.37 105.08 71.44 ;
    RECT 104.87 71.73 105.08 71.8 ;
    RECT 104.87 72.09 105.08 72.16 ;
    RECT 101.09 71.37 101.3 71.44 ;
    RECT 101.09 71.73 101.3 71.8 ;
    RECT 101.09 72.09 101.3 72.16 ;
    RECT 101.55 71.37 101.76 71.44 ;
    RECT 101.55 71.73 101.76 71.8 ;
    RECT 101.55 72.09 101.76 72.16 ;
    RECT 97.77 71.37 97.98 71.44 ;
    RECT 97.77 71.73 97.98 71.8 ;
    RECT 97.77 72.09 97.98 72.16 ;
    RECT 98.23 71.37 98.44 71.44 ;
    RECT 98.23 71.73 98.44 71.8 ;
    RECT 98.23 72.09 98.44 72.16 ;
    RECT 94.45 71.37 94.66 71.44 ;
    RECT 94.45 71.73 94.66 71.8 ;
    RECT 94.45 72.09 94.66 72.16 ;
    RECT 94.91 71.37 95.12 71.44 ;
    RECT 94.91 71.73 95.12 71.8 ;
    RECT 94.91 72.09 95.12 72.16 ;
    RECT 91.13 71.37 91.34 71.44 ;
    RECT 91.13 71.73 91.34 71.8 ;
    RECT 91.13 72.09 91.34 72.16 ;
    RECT 91.59 71.37 91.8 71.44 ;
    RECT 91.59 71.73 91.8 71.8 ;
    RECT 91.59 72.09 91.8 72.16 ;
    RECT 87.81 71.37 88.02 71.44 ;
    RECT 87.81 71.73 88.02 71.8 ;
    RECT 87.81 72.09 88.02 72.16 ;
    RECT 88.27 71.37 88.48 71.44 ;
    RECT 88.27 71.73 88.48 71.8 ;
    RECT 88.27 72.09 88.48 72.16 ;
    RECT 84.49 71.37 84.7 71.44 ;
    RECT 84.49 71.73 84.7 71.8 ;
    RECT 84.49 72.09 84.7 72.16 ;
    RECT 84.95 71.37 85.16 71.44 ;
    RECT 84.95 71.73 85.16 71.8 ;
    RECT 84.95 72.09 85.16 72.16 ;
    RECT 81.17 71.37 81.38 71.44 ;
    RECT 81.17 71.73 81.38 71.8 ;
    RECT 81.17 72.09 81.38 72.16 ;
    RECT 81.63 71.37 81.84 71.44 ;
    RECT 81.63 71.73 81.84 71.8 ;
    RECT 81.63 72.09 81.84 72.16 ;
    RECT 77.85 71.37 78.06 71.44 ;
    RECT 77.85 71.73 78.06 71.8 ;
    RECT 77.85 72.09 78.06 72.16 ;
    RECT 78.31 71.37 78.52 71.44 ;
    RECT 78.31 71.73 78.52 71.8 ;
    RECT 78.31 72.09 78.52 72.16 ;
    RECT 74.53 71.37 74.74 71.44 ;
    RECT 74.53 71.73 74.74 71.8 ;
    RECT 74.53 72.09 74.74 72.16 ;
    RECT 74.99 71.37 75.2 71.44 ;
    RECT 74.99 71.73 75.2 71.8 ;
    RECT 74.99 72.09 75.2 72.16 ;
    RECT 71.21 71.37 71.42 71.44 ;
    RECT 71.21 71.73 71.42 71.8 ;
    RECT 71.21 72.09 71.42 72.16 ;
    RECT 71.67 71.37 71.88 71.44 ;
    RECT 71.67 71.73 71.88 71.8 ;
    RECT 71.67 72.09 71.88 72.16 ;
    RECT 31.37 71.37 31.58 71.44 ;
    RECT 31.37 71.73 31.58 71.8 ;
    RECT 31.37 72.09 31.58 72.16 ;
    RECT 31.83 71.37 32.04 71.44 ;
    RECT 31.83 71.73 32.04 71.8 ;
    RECT 31.83 72.09 32.04 72.16 ;
    RECT 67.89 71.37 68.1 71.44 ;
    RECT 67.89 71.73 68.1 71.8 ;
    RECT 67.89 72.09 68.1 72.16 ;
    RECT 68.35 71.37 68.56 71.44 ;
    RECT 68.35 71.73 68.56 71.8 ;
    RECT 68.35 72.09 68.56 72.16 ;
    RECT 28.05 71.37 28.26 71.44 ;
    RECT 28.05 71.73 28.26 71.8 ;
    RECT 28.05 72.09 28.26 72.16 ;
    RECT 28.51 71.37 28.72 71.44 ;
    RECT 28.51 71.73 28.72 71.8 ;
    RECT 28.51 72.09 28.72 72.16 ;
    RECT 24.73 71.37 24.94 71.44 ;
    RECT 24.73 71.73 24.94 71.8 ;
    RECT 24.73 72.09 24.94 72.16 ;
    RECT 25.19 71.37 25.4 71.44 ;
    RECT 25.19 71.73 25.4 71.8 ;
    RECT 25.19 72.09 25.4 72.16 ;
    RECT 21.41 71.37 21.62 71.44 ;
    RECT 21.41 71.73 21.62 71.8 ;
    RECT 21.41 72.09 21.62 72.16 ;
    RECT 21.87 71.37 22.08 71.44 ;
    RECT 21.87 71.73 22.08 71.8 ;
    RECT 21.87 72.09 22.08 72.16 ;
    RECT 18.09 71.37 18.3 71.44 ;
    RECT 18.09 71.73 18.3 71.8 ;
    RECT 18.09 72.09 18.3 72.16 ;
    RECT 18.55 71.37 18.76 71.44 ;
    RECT 18.55 71.73 18.76 71.8 ;
    RECT 18.55 72.09 18.76 72.16 ;
    RECT 120.825 71.73 120.895 71.8 ;
    RECT 14.77 71.37 14.98 71.44 ;
    RECT 14.77 71.73 14.98 71.8 ;
    RECT 14.77 72.09 14.98 72.16 ;
    RECT 15.23 71.37 15.44 71.44 ;
    RECT 15.23 71.73 15.44 71.8 ;
    RECT 15.23 72.09 15.44 72.16 ;
    RECT 11.45 71.37 11.66 71.44 ;
    RECT 11.45 71.73 11.66 71.8 ;
    RECT 11.45 72.09 11.66 72.16 ;
    RECT 11.91 71.37 12.12 71.44 ;
    RECT 11.91 71.73 12.12 71.8 ;
    RECT 11.91 72.09 12.12 72.16 ;
    RECT 8.13 71.37 8.34 71.44 ;
    RECT 8.13 71.73 8.34 71.8 ;
    RECT 8.13 72.09 8.34 72.16 ;
    RECT 8.59 71.37 8.8 71.44 ;
    RECT 8.59 71.73 8.8 71.8 ;
    RECT 8.59 72.09 8.8 72.16 ;
    RECT 4.81 71.37 5.02 71.44 ;
    RECT 4.81 71.73 5.02 71.8 ;
    RECT 4.81 72.09 5.02 72.16 ;
    RECT 5.27 71.37 5.48 71.44 ;
    RECT 5.27 71.73 5.48 71.8 ;
    RECT 5.27 72.09 5.48 72.16 ;
    RECT 1.49 71.37 1.7 71.44 ;
    RECT 1.49 71.73 1.7 71.8 ;
    RECT 1.49 72.09 1.7 72.16 ;
    RECT 1.95 71.37 2.16 71.44 ;
    RECT 1.95 71.73 2.16 71.8 ;
    RECT 1.95 72.09 2.16 72.16 ;
    RECT 64.57 71.37 64.78 71.44 ;
    RECT 64.57 71.73 64.78 71.8 ;
    RECT 64.57 72.09 64.78 72.16 ;
    RECT 65.03 71.37 65.24 71.44 ;
    RECT 65.03 71.73 65.24 71.8 ;
    RECT 65.03 72.09 65.24 72.16 ;
    RECT 61.25 31.03 61.46 31.1 ;
    RECT 61.25 31.39 61.46 31.46 ;
    RECT 61.25 31.75 61.46 31.82 ;
    RECT 61.71 31.03 61.92 31.1 ;
    RECT 61.71 31.39 61.92 31.46 ;
    RECT 61.71 31.75 61.92 31.82 ;
    RECT 57.93 31.03 58.14 31.1 ;
    RECT 57.93 31.39 58.14 31.46 ;
    RECT 57.93 31.75 58.14 31.82 ;
    RECT 58.39 31.03 58.6 31.1 ;
    RECT 58.39 31.39 58.6 31.46 ;
    RECT 58.39 31.75 58.6 31.82 ;
    RECT 54.61 31.03 54.82 31.1 ;
    RECT 54.61 31.39 54.82 31.46 ;
    RECT 54.61 31.75 54.82 31.82 ;
    RECT 55.07 31.03 55.28 31.1 ;
    RECT 55.07 31.39 55.28 31.46 ;
    RECT 55.07 31.75 55.28 31.82 ;
    RECT 51.29 31.03 51.5 31.1 ;
    RECT 51.29 31.39 51.5 31.46 ;
    RECT 51.29 31.75 51.5 31.82 ;
    RECT 51.75 31.03 51.96 31.1 ;
    RECT 51.75 31.39 51.96 31.46 ;
    RECT 51.75 31.75 51.96 31.82 ;
    RECT 47.97 31.03 48.18 31.1 ;
    RECT 47.97 31.39 48.18 31.46 ;
    RECT 47.97 31.75 48.18 31.82 ;
    RECT 48.43 31.03 48.64 31.1 ;
    RECT 48.43 31.39 48.64 31.46 ;
    RECT 48.43 31.75 48.64 31.82 ;
    RECT 44.65 31.03 44.86 31.1 ;
    RECT 44.65 31.39 44.86 31.46 ;
    RECT 44.65 31.75 44.86 31.82 ;
    RECT 45.11 31.03 45.32 31.1 ;
    RECT 45.11 31.39 45.32 31.46 ;
    RECT 45.11 31.75 45.32 31.82 ;
    RECT 41.33 31.03 41.54 31.1 ;
    RECT 41.33 31.39 41.54 31.46 ;
    RECT 41.33 31.75 41.54 31.82 ;
    RECT 41.79 31.03 42.0 31.1 ;
    RECT 41.79 31.39 42.0 31.46 ;
    RECT 41.79 31.75 42.0 31.82 ;
    RECT 38.01 31.03 38.22 31.1 ;
    RECT 38.01 31.39 38.22 31.46 ;
    RECT 38.01 31.75 38.22 31.82 ;
    RECT 38.47 31.03 38.68 31.1 ;
    RECT 38.47 31.39 38.68 31.46 ;
    RECT 38.47 31.75 38.68 31.82 ;
    RECT 0.4 31.39 0.47 31.46 ;
    RECT 34.69 31.03 34.9 31.1 ;
    RECT 34.69 31.39 34.9 31.46 ;
    RECT 34.69 31.75 34.9 31.82 ;
    RECT 35.15 31.03 35.36 31.1 ;
    RECT 35.15 31.39 35.36 31.46 ;
    RECT 35.15 31.75 35.36 31.82 ;
    RECT 117.69 31.03 117.9 31.1 ;
    RECT 117.69 31.39 117.9 31.46 ;
    RECT 117.69 31.75 117.9 31.82 ;
    RECT 118.15 31.03 118.36 31.1 ;
    RECT 118.15 31.39 118.36 31.46 ;
    RECT 118.15 31.75 118.36 31.82 ;
    RECT 114.37 31.03 114.58 31.1 ;
    RECT 114.37 31.39 114.58 31.46 ;
    RECT 114.37 31.75 114.58 31.82 ;
    RECT 114.83 31.03 115.04 31.1 ;
    RECT 114.83 31.39 115.04 31.46 ;
    RECT 114.83 31.75 115.04 31.82 ;
    RECT 111.05 31.03 111.26 31.1 ;
    RECT 111.05 31.39 111.26 31.46 ;
    RECT 111.05 31.75 111.26 31.82 ;
    RECT 111.51 31.03 111.72 31.1 ;
    RECT 111.51 31.39 111.72 31.46 ;
    RECT 111.51 31.75 111.72 31.82 ;
    RECT 107.73 31.03 107.94 31.1 ;
    RECT 107.73 31.39 107.94 31.46 ;
    RECT 107.73 31.75 107.94 31.82 ;
    RECT 108.19 31.03 108.4 31.1 ;
    RECT 108.19 31.39 108.4 31.46 ;
    RECT 108.19 31.75 108.4 31.82 ;
    RECT 104.41 31.03 104.62 31.1 ;
    RECT 104.41 31.39 104.62 31.46 ;
    RECT 104.41 31.75 104.62 31.82 ;
    RECT 104.87 31.03 105.08 31.1 ;
    RECT 104.87 31.39 105.08 31.46 ;
    RECT 104.87 31.75 105.08 31.82 ;
    RECT 101.09 31.03 101.3 31.1 ;
    RECT 101.09 31.39 101.3 31.46 ;
    RECT 101.09 31.75 101.3 31.82 ;
    RECT 101.55 31.03 101.76 31.1 ;
    RECT 101.55 31.39 101.76 31.46 ;
    RECT 101.55 31.75 101.76 31.82 ;
    RECT 97.77 31.03 97.98 31.1 ;
    RECT 97.77 31.39 97.98 31.46 ;
    RECT 97.77 31.75 97.98 31.82 ;
    RECT 98.23 31.03 98.44 31.1 ;
    RECT 98.23 31.39 98.44 31.46 ;
    RECT 98.23 31.75 98.44 31.82 ;
    RECT 94.45 31.03 94.66 31.1 ;
    RECT 94.45 31.39 94.66 31.46 ;
    RECT 94.45 31.75 94.66 31.82 ;
    RECT 94.91 31.03 95.12 31.1 ;
    RECT 94.91 31.39 95.12 31.46 ;
    RECT 94.91 31.75 95.12 31.82 ;
    RECT 91.13 31.03 91.34 31.1 ;
    RECT 91.13 31.39 91.34 31.46 ;
    RECT 91.13 31.75 91.34 31.82 ;
    RECT 91.59 31.03 91.8 31.1 ;
    RECT 91.59 31.39 91.8 31.46 ;
    RECT 91.59 31.75 91.8 31.82 ;
    RECT 87.81 31.03 88.02 31.1 ;
    RECT 87.81 31.39 88.02 31.46 ;
    RECT 87.81 31.75 88.02 31.82 ;
    RECT 88.27 31.03 88.48 31.1 ;
    RECT 88.27 31.39 88.48 31.46 ;
    RECT 88.27 31.75 88.48 31.82 ;
    RECT 84.49 31.03 84.7 31.1 ;
    RECT 84.49 31.39 84.7 31.46 ;
    RECT 84.49 31.75 84.7 31.82 ;
    RECT 84.95 31.03 85.16 31.1 ;
    RECT 84.95 31.39 85.16 31.46 ;
    RECT 84.95 31.75 85.16 31.82 ;
    RECT 81.17 31.03 81.38 31.1 ;
    RECT 81.17 31.39 81.38 31.46 ;
    RECT 81.17 31.75 81.38 31.82 ;
    RECT 81.63 31.03 81.84 31.1 ;
    RECT 81.63 31.39 81.84 31.46 ;
    RECT 81.63 31.75 81.84 31.82 ;
    RECT 77.85 31.03 78.06 31.1 ;
    RECT 77.85 31.39 78.06 31.46 ;
    RECT 77.85 31.75 78.06 31.82 ;
    RECT 78.31 31.03 78.52 31.1 ;
    RECT 78.31 31.39 78.52 31.46 ;
    RECT 78.31 31.75 78.52 31.82 ;
    RECT 74.53 31.03 74.74 31.1 ;
    RECT 74.53 31.39 74.74 31.46 ;
    RECT 74.53 31.75 74.74 31.82 ;
    RECT 74.99 31.03 75.2 31.1 ;
    RECT 74.99 31.39 75.2 31.46 ;
    RECT 74.99 31.75 75.2 31.82 ;
    RECT 71.21 31.03 71.42 31.1 ;
    RECT 71.21 31.39 71.42 31.46 ;
    RECT 71.21 31.75 71.42 31.82 ;
    RECT 71.67 31.03 71.88 31.1 ;
    RECT 71.67 31.39 71.88 31.46 ;
    RECT 71.67 31.75 71.88 31.82 ;
    RECT 31.37 31.03 31.58 31.1 ;
    RECT 31.37 31.39 31.58 31.46 ;
    RECT 31.37 31.75 31.58 31.82 ;
    RECT 31.83 31.03 32.04 31.1 ;
    RECT 31.83 31.39 32.04 31.46 ;
    RECT 31.83 31.75 32.04 31.82 ;
    RECT 67.89 31.03 68.1 31.1 ;
    RECT 67.89 31.39 68.1 31.46 ;
    RECT 67.89 31.75 68.1 31.82 ;
    RECT 68.35 31.03 68.56 31.1 ;
    RECT 68.35 31.39 68.56 31.46 ;
    RECT 68.35 31.75 68.56 31.82 ;
    RECT 28.05 31.03 28.26 31.1 ;
    RECT 28.05 31.39 28.26 31.46 ;
    RECT 28.05 31.75 28.26 31.82 ;
    RECT 28.51 31.03 28.72 31.1 ;
    RECT 28.51 31.39 28.72 31.46 ;
    RECT 28.51 31.75 28.72 31.82 ;
    RECT 24.73 31.03 24.94 31.1 ;
    RECT 24.73 31.39 24.94 31.46 ;
    RECT 24.73 31.75 24.94 31.82 ;
    RECT 25.19 31.03 25.4 31.1 ;
    RECT 25.19 31.39 25.4 31.46 ;
    RECT 25.19 31.75 25.4 31.82 ;
    RECT 21.41 31.03 21.62 31.1 ;
    RECT 21.41 31.39 21.62 31.46 ;
    RECT 21.41 31.75 21.62 31.82 ;
    RECT 21.87 31.03 22.08 31.1 ;
    RECT 21.87 31.39 22.08 31.46 ;
    RECT 21.87 31.75 22.08 31.82 ;
    RECT 18.09 31.03 18.3 31.1 ;
    RECT 18.09 31.39 18.3 31.46 ;
    RECT 18.09 31.75 18.3 31.82 ;
    RECT 18.55 31.03 18.76 31.1 ;
    RECT 18.55 31.39 18.76 31.46 ;
    RECT 18.55 31.75 18.76 31.82 ;
    RECT 120.825 31.39 120.895 31.46 ;
    RECT 14.77 31.03 14.98 31.1 ;
    RECT 14.77 31.39 14.98 31.46 ;
    RECT 14.77 31.75 14.98 31.82 ;
    RECT 15.23 31.03 15.44 31.1 ;
    RECT 15.23 31.39 15.44 31.46 ;
    RECT 15.23 31.75 15.44 31.82 ;
    RECT 11.45 31.03 11.66 31.1 ;
    RECT 11.45 31.39 11.66 31.46 ;
    RECT 11.45 31.75 11.66 31.82 ;
    RECT 11.91 31.03 12.12 31.1 ;
    RECT 11.91 31.39 12.12 31.46 ;
    RECT 11.91 31.75 12.12 31.82 ;
    RECT 8.13 31.03 8.34 31.1 ;
    RECT 8.13 31.39 8.34 31.46 ;
    RECT 8.13 31.75 8.34 31.82 ;
    RECT 8.59 31.03 8.8 31.1 ;
    RECT 8.59 31.39 8.8 31.46 ;
    RECT 8.59 31.75 8.8 31.82 ;
    RECT 4.81 31.03 5.02 31.1 ;
    RECT 4.81 31.39 5.02 31.46 ;
    RECT 4.81 31.75 5.02 31.82 ;
    RECT 5.27 31.03 5.48 31.1 ;
    RECT 5.27 31.39 5.48 31.46 ;
    RECT 5.27 31.75 5.48 31.82 ;
    RECT 1.49 31.03 1.7 31.1 ;
    RECT 1.49 31.39 1.7 31.46 ;
    RECT 1.49 31.75 1.7 31.82 ;
    RECT 1.95 31.03 2.16 31.1 ;
    RECT 1.95 31.39 2.16 31.46 ;
    RECT 1.95 31.75 2.16 31.82 ;
    RECT 64.57 31.03 64.78 31.1 ;
    RECT 64.57 31.39 64.78 31.46 ;
    RECT 64.57 31.75 64.78 31.82 ;
    RECT 65.03 31.03 65.24 31.1 ;
    RECT 65.03 31.39 65.24 31.46 ;
    RECT 65.03 31.75 65.24 31.82 ;
    RECT 61.25 70.65 61.46 70.72 ;
    RECT 61.25 71.01 61.46 71.08 ;
    RECT 61.25 71.37 61.46 71.44 ;
    RECT 61.71 70.65 61.92 70.72 ;
    RECT 61.71 71.01 61.92 71.08 ;
    RECT 61.71 71.37 61.92 71.44 ;
    RECT 57.93 70.65 58.14 70.72 ;
    RECT 57.93 71.01 58.14 71.08 ;
    RECT 57.93 71.37 58.14 71.44 ;
    RECT 58.39 70.65 58.6 70.72 ;
    RECT 58.39 71.01 58.6 71.08 ;
    RECT 58.39 71.37 58.6 71.44 ;
    RECT 54.61 70.65 54.82 70.72 ;
    RECT 54.61 71.01 54.82 71.08 ;
    RECT 54.61 71.37 54.82 71.44 ;
    RECT 55.07 70.65 55.28 70.72 ;
    RECT 55.07 71.01 55.28 71.08 ;
    RECT 55.07 71.37 55.28 71.44 ;
    RECT 51.29 70.65 51.5 70.72 ;
    RECT 51.29 71.01 51.5 71.08 ;
    RECT 51.29 71.37 51.5 71.44 ;
    RECT 51.75 70.65 51.96 70.72 ;
    RECT 51.75 71.01 51.96 71.08 ;
    RECT 51.75 71.37 51.96 71.44 ;
    RECT 47.97 70.65 48.18 70.72 ;
    RECT 47.97 71.01 48.18 71.08 ;
    RECT 47.97 71.37 48.18 71.44 ;
    RECT 48.43 70.65 48.64 70.72 ;
    RECT 48.43 71.01 48.64 71.08 ;
    RECT 48.43 71.37 48.64 71.44 ;
    RECT 44.65 70.65 44.86 70.72 ;
    RECT 44.65 71.01 44.86 71.08 ;
    RECT 44.65 71.37 44.86 71.44 ;
    RECT 45.11 70.65 45.32 70.72 ;
    RECT 45.11 71.01 45.32 71.08 ;
    RECT 45.11 71.37 45.32 71.44 ;
    RECT 41.33 70.65 41.54 70.72 ;
    RECT 41.33 71.01 41.54 71.08 ;
    RECT 41.33 71.37 41.54 71.44 ;
    RECT 41.79 70.65 42.0 70.72 ;
    RECT 41.79 71.01 42.0 71.08 ;
    RECT 41.79 71.37 42.0 71.44 ;
    RECT 38.01 70.65 38.22 70.72 ;
    RECT 38.01 71.01 38.22 71.08 ;
    RECT 38.01 71.37 38.22 71.44 ;
    RECT 38.47 70.65 38.68 70.72 ;
    RECT 38.47 71.01 38.68 71.08 ;
    RECT 38.47 71.37 38.68 71.44 ;
    RECT 0.4 71.01 0.47 71.08 ;
    RECT 34.69 70.65 34.9 70.72 ;
    RECT 34.69 71.01 34.9 71.08 ;
    RECT 34.69 71.37 34.9 71.44 ;
    RECT 35.15 70.65 35.36 70.72 ;
    RECT 35.15 71.01 35.36 71.08 ;
    RECT 35.15 71.37 35.36 71.44 ;
    RECT 117.69 70.65 117.9 70.72 ;
    RECT 117.69 71.01 117.9 71.08 ;
    RECT 117.69 71.37 117.9 71.44 ;
    RECT 118.15 70.65 118.36 70.72 ;
    RECT 118.15 71.01 118.36 71.08 ;
    RECT 118.15 71.37 118.36 71.44 ;
    RECT 114.37 70.65 114.58 70.72 ;
    RECT 114.37 71.01 114.58 71.08 ;
    RECT 114.37 71.37 114.58 71.44 ;
    RECT 114.83 70.65 115.04 70.72 ;
    RECT 114.83 71.01 115.04 71.08 ;
    RECT 114.83 71.37 115.04 71.44 ;
    RECT 111.05 70.65 111.26 70.72 ;
    RECT 111.05 71.01 111.26 71.08 ;
    RECT 111.05 71.37 111.26 71.44 ;
    RECT 111.51 70.65 111.72 70.72 ;
    RECT 111.51 71.01 111.72 71.08 ;
    RECT 111.51 71.37 111.72 71.44 ;
    RECT 107.73 70.65 107.94 70.72 ;
    RECT 107.73 71.01 107.94 71.08 ;
    RECT 107.73 71.37 107.94 71.44 ;
    RECT 108.19 70.65 108.4 70.72 ;
    RECT 108.19 71.01 108.4 71.08 ;
    RECT 108.19 71.37 108.4 71.44 ;
    RECT 104.41 70.65 104.62 70.72 ;
    RECT 104.41 71.01 104.62 71.08 ;
    RECT 104.41 71.37 104.62 71.44 ;
    RECT 104.87 70.65 105.08 70.72 ;
    RECT 104.87 71.01 105.08 71.08 ;
    RECT 104.87 71.37 105.08 71.44 ;
    RECT 101.09 70.65 101.3 70.72 ;
    RECT 101.09 71.01 101.3 71.08 ;
    RECT 101.09 71.37 101.3 71.44 ;
    RECT 101.55 70.65 101.76 70.72 ;
    RECT 101.55 71.01 101.76 71.08 ;
    RECT 101.55 71.37 101.76 71.44 ;
    RECT 97.77 70.65 97.98 70.72 ;
    RECT 97.77 71.01 97.98 71.08 ;
    RECT 97.77 71.37 97.98 71.44 ;
    RECT 98.23 70.65 98.44 70.72 ;
    RECT 98.23 71.01 98.44 71.08 ;
    RECT 98.23 71.37 98.44 71.44 ;
    RECT 94.45 70.65 94.66 70.72 ;
    RECT 94.45 71.01 94.66 71.08 ;
    RECT 94.45 71.37 94.66 71.44 ;
    RECT 94.91 70.65 95.12 70.72 ;
    RECT 94.91 71.01 95.12 71.08 ;
    RECT 94.91 71.37 95.12 71.44 ;
    RECT 91.13 70.65 91.34 70.72 ;
    RECT 91.13 71.01 91.34 71.08 ;
    RECT 91.13 71.37 91.34 71.44 ;
    RECT 91.59 70.65 91.8 70.72 ;
    RECT 91.59 71.01 91.8 71.08 ;
    RECT 91.59 71.37 91.8 71.44 ;
    RECT 87.81 70.65 88.02 70.72 ;
    RECT 87.81 71.01 88.02 71.08 ;
    RECT 87.81 71.37 88.02 71.44 ;
    RECT 88.27 70.65 88.48 70.72 ;
    RECT 88.27 71.01 88.48 71.08 ;
    RECT 88.27 71.37 88.48 71.44 ;
    RECT 84.49 70.65 84.7 70.72 ;
    RECT 84.49 71.01 84.7 71.08 ;
    RECT 84.49 71.37 84.7 71.44 ;
    RECT 84.95 70.65 85.16 70.72 ;
    RECT 84.95 71.01 85.16 71.08 ;
    RECT 84.95 71.37 85.16 71.44 ;
    RECT 81.17 70.65 81.38 70.72 ;
    RECT 81.17 71.01 81.38 71.08 ;
    RECT 81.17 71.37 81.38 71.44 ;
    RECT 81.63 70.65 81.84 70.72 ;
    RECT 81.63 71.01 81.84 71.08 ;
    RECT 81.63 71.37 81.84 71.44 ;
    RECT 77.85 70.65 78.06 70.72 ;
    RECT 77.85 71.01 78.06 71.08 ;
    RECT 77.85 71.37 78.06 71.44 ;
    RECT 78.31 70.65 78.52 70.72 ;
    RECT 78.31 71.01 78.52 71.08 ;
    RECT 78.31 71.37 78.52 71.44 ;
    RECT 74.53 70.65 74.74 70.72 ;
    RECT 74.53 71.01 74.74 71.08 ;
    RECT 74.53 71.37 74.74 71.44 ;
    RECT 74.99 70.65 75.2 70.72 ;
    RECT 74.99 71.01 75.2 71.08 ;
    RECT 74.99 71.37 75.2 71.44 ;
    RECT 71.21 70.65 71.42 70.72 ;
    RECT 71.21 71.01 71.42 71.08 ;
    RECT 71.21 71.37 71.42 71.44 ;
    RECT 71.67 70.65 71.88 70.72 ;
    RECT 71.67 71.01 71.88 71.08 ;
    RECT 71.67 71.37 71.88 71.44 ;
    RECT 31.37 70.65 31.58 70.72 ;
    RECT 31.37 71.01 31.58 71.08 ;
    RECT 31.37 71.37 31.58 71.44 ;
    RECT 31.83 70.65 32.04 70.72 ;
    RECT 31.83 71.01 32.04 71.08 ;
    RECT 31.83 71.37 32.04 71.44 ;
    RECT 67.89 70.65 68.1 70.72 ;
    RECT 67.89 71.01 68.1 71.08 ;
    RECT 67.89 71.37 68.1 71.44 ;
    RECT 68.35 70.65 68.56 70.72 ;
    RECT 68.35 71.01 68.56 71.08 ;
    RECT 68.35 71.37 68.56 71.44 ;
    RECT 28.05 70.65 28.26 70.72 ;
    RECT 28.05 71.01 28.26 71.08 ;
    RECT 28.05 71.37 28.26 71.44 ;
    RECT 28.51 70.65 28.72 70.72 ;
    RECT 28.51 71.01 28.72 71.08 ;
    RECT 28.51 71.37 28.72 71.44 ;
    RECT 24.73 70.65 24.94 70.72 ;
    RECT 24.73 71.01 24.94 71.08 ;
    RECT 24.73 71.37 24.94 71.44 ;
    RECT 25.19 70.65 25.4 70.72 ;
    RECT 25.19 71.01 25.4 71.08 ;
    RECT 25.19 71.37 25.4 71.44 ;
    RECT 21.41 70.65 21.62 70.72 ;
    RECT 21.41 71.01 21.62 71.08 ;
    RECT 21.41 71.37 21.62 71.44 ;
    RECT 21.87 70.65 22.08 70.72 ;
    RECT 21.87 71.01 22.08 71.08 ;
    RECT 21.87 71.37 22.08 71.44 ;
    RECT 18.09 70.65 18.3 70.72 ;
    RECT 18.09 71.01 18.3 71.08 ;
    RECT 18.09 71.37 18.3 71.44 ;
    RECT 18.55 70.65 18.76 70.72 ;
    RECT 18.55 71.01 18.76 71.08 ;
    RECT 18.55 71.37 18.76 71.44 ;
    RECT 120.825 71.01 120.895 71.08 ;
    RECT 14.77 70.65 14.98 70.72 ;
    RECT 14.77 71.01 14.98 71.08 ;
    RECT 14.77 71.37 14.98 71.44 ;
    RECT 15.23 70.65 15.44 70.72 ;
    RECT 15.23 71.01 15.44 71.08 ;
    RECT 15.23 71.37 15.44 71.44 ;
    RECT 11.45 70.65 11.66 70.72 ;
    RECT 11.45 71.01 11.66 71.08 ;
    RECT 11.45 71.37 11.66 71.44 ;
    RECT 11.91 70.65 12.12 70.72 ;
    RECT 11.91 71.01 12.12 71.08 ;
    RECT 11.91 71.37 12.12 71.44 ;
    RECT 8.13 70.65 8.34 70.72 ;
    RECT 8.13 71.01 8.34 71.08 ;
    RECT 8.13 71.37 8.34 71.44 ;
    RECT 8.59 70.65 8.8 70.72 ;
    RECT 8.59 71.01 8.8 71.08 ;
    RECT 8.59 71.37 8.8 71.44 ;
    RECT 4.81 70.65 5.02 70.72 ;
    RECT 4.81 71.01 5.02 71.08 ;
    RECT 4.81 71.37 5.02 71.44 ;
    RECT 5.27 70.65 5.48 70.72 ;
    RECT 5.27 71.01 5.48 71.08 ;
    RECT 5.27 71.37 5.48 71.44 ;
    RECT 1.49 70.65 1.7 70.72 ;
    RECT 1.49 71.01 1.7 71.08 ;
    RECT 1.49 71.37 1.7 71.44 ;
    RECT 1.95 70.65 2.16 70.72 ;
    RECT 1.95 71.01 2.16 71.08 ;
    RECT 1.95 71.37 2.16 71.44 ;
    RECT 64.57 70.65 64.78 70.72 ;
    RECT 64.57 71.01 64.78 71.08 ;
    RECT 64.57 71.37 64.78 71.44 ;
    RECT 65.03 70.65 65.24 70.72 ;
    RECT 65.03 71.01 65.24 71.08 ;
    RECT 65.03 71.37 65.24 71.44 ;
    RECT 61.25 30.31 61.46 30.38 ;
    RECT 61.25 30.67 61.46 30.74 ;
    RECT 61.25 31.03 61.46 31.1 ;
    RECT 61.71 30.31 61.92 30.38 ;
    RECT 61.71 30.67 61.92 30.74 ;
    RECT 61.71 31.03 61.92 31.1 ;
    RECT 57.93 30.31 58.14 30.38 ;
    RECT 57.93 30.67 58.14 30.74 ;
    RECT 57.93 31.03 58.14 31.1 ;
    RECT 58.39 30.31 58.6 30.38 ;
    RECT 58.39 30.67 58.6 30.74 ;
    RECT 58.39 31.03 58.6 31.1 ;
    RECT 54.61 30.31 54.82 30.38 ;
    RECT 54.61 30.67 54.82 30.74 ;
    RECT 54.61 31.03 54.82 31.1 ;
    RECT 55.07 30.31 55.28 30.38 ;
    RECT 55.07 30.67 55.28 30.74 ;
    RECT 55.07 31.03 55.28 31.1 ;
    RECT 51.29 30.31 51.5 30.38 ;
    RECT 51.29 30.67 51.5 30.74 ;
    RECT 51.29 31.03 51.5 31.1 ;
    RECT 51.75 30.31 51.96 30.38 ;
    RECT 51.75 30.67 51.96 30.74 ;
    RECT 51.75 31.03 51.96 31.1 ;
    RECT 47.97 30.31 48.18 30.38 ;
    RECT 47.97 30.67 48.18 30.74 ;
    RECT 47.97 31.03 48.18 31.1 ;
    RECT 48.43 30.31 48.64 30.38 ;
    RECT 48.43 30.67 48.64 30.74 ;
    RECT 48.43 31.03 48.64 31.1 ;
    RECT 44.65 30.31 44.86 30.38 ;
    RECT 44.65 30.67 44.86 30.74 ;
    RECT 44.65 31.03 44.86 31.1 ;
    RECT 45.11 30.31 45.32 30.38 ;
    RECT 45.11 30.67 45.32 30.74 ;
    RECT 45.11 31.03 45.32 31.1 ;
    RECT 41.33 30.31 41.54 30.38 ;
    RECT 41.33 30.67 41.54 30.74 ;
    RECT 41.33 31.03 41.54 31.1 ;
    RECT 41.79 30.31 42.0 30.38 ;
    RECT 41.79 30.67 42.0 30.74 ;
    RECT 41.79 31.03 42.0 31.1 ;
    RECT 38.01 30.31 38.22 30.38 ;
    RECT 38.01 30.67 38.22 30.74 ;
    RECT 38.01 31.03 38.22 31.1 ;
    RECT 38.47 30.31 38.68 30.38 ;
    RECT 38.47 30.67 38.68 30.74 ;
    RECT 38.47 31.03 38.68 31.1 ;
    RECT 0.4 30.67 0.47 30.74 ;
    RECT 34.69 30.31 34.9 30.38 ;
    RECT 34.69 30.67 34.9 30.74 ;
    RECT 34.69 31.03 34.9 31.1 ;
    RECT 35.15 30.31 35.36 30.38 ;
    RECT 35.15 30.67 35.36 30.74 ;
    RECT 35.15 31.03 35.36 31.1 ;
    RECT 117.69 30.31 117.9 30.38 ;
    RECT 117.69 30.67 117.9 30.74 ;
    RECT 117.69 31.03 117.9 31.1 ;
    RECT 118.15 30.31 118.36 30.38 ;
    RECT 118.15 30.67 118.36 30.74 ;
    RECT 118.15 31.03 118.36 31.1 ;
    RECT 114.37 30.31 114.58 30.38 ;
    RECT 114.37 30.67 114.58 30.74 ;
    RECT 114.37 31.03 114.58 31.1 ;
    RECT 114.83 30.31 115.04 30.38 ;
    RECT 114.83 30.67 115.04 30.74 ;
    RECT 114.83 31.03 115.04 31.1 ;
    RECT 111.05 30.31 111.26 30.38 ;
    RECT 111.05 30.67 111.26 30.74 ;
    RECT 111.05 31.03 111.26 31.1 ;
    RECT 111.51 30.31 111.72 30.38 ;
    RECT 111.51 30.67 111.72 30.74 ;
    RECT 111.51 31.03 111.72 31.1 ;
    RECT 107.73 30.31 107.94 30.38 ;
    RECT 107.73 30.67 107.94 30.74 ;
    RECT 107.73 31.03 107.94 31.1 ;
    RECT 108.19 30.31 108.4 30.38 ;
    RECT 108.19 30.67 108.4 30.74 ;
    RECT 108.19 31.03 108.4 31.1 ;
    RECT 104.41 30.31 104.62 30.38 ;
    RECT 104.41 30.67 104.62 30.74 ;
    RECT 104.41 31.03 104.62 31.1 ;
    RECT 104.87 30.31 105.08 30.38 ;
    RECT 104.87 30.67 105.08 30.74 ;
    RECT 104.87 31.03 105.08 31.1 ;
    RECT 101.09 30.31 101.3 30.38 ;
    RECT 101.09 30.67 101.3 30.74 ;
    RECT 101.09 31.03 101.3 31.1 ;
    RECT 101.55 30.31 101.76 30.38 ;
    RECT 101.55 30.67 101.76 30.74 ;
    RECT 101.55 31.03 101.76 31.1 ;
    RECT 97.77 30.31 97.98 30.38 ;
    RECT 97.77 30.67 97.98 30.74 ;
    RECT 97.77 31.03 97.98 31.1 ;
    RECT 98.23 30.31 98.44 30.38 ;
    RECT 98.23 30.67 98.44 30.74 ;
    RECT 98.23 31.03 98.44 31.1 ;
    RECT 94.45 30.31 94.66 30.38 ;
    RECT 94.45 30.67 94.66 30.74 ;
    RECT 94.45 31.03 94.66 31.1 ;
    RECT 94.91 30.31 95.12 30.38 ;
    RECT 94.91 30.67 95.12 30.74 ;
    RECT 94.91 31.03 95.12 31.1 ;
    RECT 91.13 30.31 91.34 30.38 ;
    RECT 91.13 30.67 91.34 30.74 ;
    RECT 91.13 31.03 91.34 31.1 ;
    RECT 91.59 30.31 91.8 30.38 ;
    RECT 91.59 30.67 91.8 30.74 ;
    RECT 91.59 31.03 91.8 31.1 ;
    RECT 87.81 30.31 88.02 30.38 ;
    RECT 87.81 30.67 88.02 30.74 ;
    RECT 87.81 31.03 88.02 31.1 ;
    RECT 88.27 30.31 88.48 30.38 ;
    RECT 88.27 30.67 88.48 30.74 ;
    RECT 88.27 31.03 88.48 31.1 ;
    RECT 84.49 30.31 84.7 30.38 ;
    RECT 84.49 30.67 84.7 30.74 ;
    RECT 84.49 31.03 84.7 31.1 ;
    RECT 84.95 30.31 85.16 30.38 ;
    RECT 84.95 30.67 85.16 30.74 ;
    RECT 84.95 31.03 85.16 31.1 ;
    RECT 81.17 30.31 81.38 30.38 ;
    RECT 81.17 30.67 81.38 30.74 ;
    RECT 81.17 31.03 81.38 31.1 ;
    RECT 81.63 30.31 81.84 30.38 ;
    RECT 81.63 30.67 81.84 30.74 ;
    RECT 81.63 31.03 81.84 31.1 ;
    RECT 77.85 30.31 78.06 30.38 ;
    RECT 77.85 30.67 78.06 30.74 ;
    RECT 77.85 31.03 78.06 31.1 ;
    RECT 78.31 30.31 78.52 30.38 ;
    RECT 78.31 30.67 78.52 30.74 ;
    RECT 78.31 31.03 78.52 31.1 ;
    RECT 74.53 30.31 74.74 30.38 ;
    RECT 74.53 30.67 74.74 30.74 ;
    RECT 74.53 31.03 74.74 31.1 ;
    RECT 74.99 30.31 75.2 30.38 ;
    RECT 74.99 30.67 75.2 30.74 ;
    RECT 74.99 31.03 75.2 31.1 ;
    RECT 71.21 30.31 71.42 30.38 ;
    RECT 71.21 30.67 71.42 30.74 ;
    RECT 71.21 31.03 71.42 31.1 ;
    RECT 71.67 30.31 71.88 30.38 ;
    RECT 71.67 30.67 71.88 30.74 ;
    RECT 71.67 31.03 71.88 31.1 ;
    RECT 31.37 30.31 31.58 30.38 ;
    RECT 31.37 30.67 31.58 30.74 ;
    RECT 31.37 31.03 31.58 31.1 ;
    RECT 31.83 30.31 32.04 30.38 ;
    RECT 31.83 30.67 32.04 30.74 ;
    RECT 31.83 31.03 32.04 31.1 ;
    RECT 67.89 30.31 68.1 30.38 ;
    RECT 67.89 30.67 68.1 30.74 ;
    RECT 67.89 31.03 68.1 31.1 ;
    RECT 68.35 30.31 68.56 30.38 ;
    RECT 68.35 30.67 68.56 30.74 ;
    RECT 68.35 31.03 68.56 31.1 ;
    RECT 28.05 30.31 28.26 30.38 ;
    RECT 28.05 30.67 28.26 30.74 ;
    RECT 28.05 31.03 28.26 31.1 ;
    RECT 28.51 30.31 28.72 30.38 ;
    RECT 28.51 30.67 28.72 30.74 ;
    RECT 28.51 31.03 28.72 31.1 ;
    RECT 24.73 30.31 24.94 30.38 ;
    RECT 24.73 30.67 24.94 30.74 ;
    RECT 24.73 31.03 24.94 31.1 ;
    RECT 25.19 30.31 25.4 30.38 ;
    RECT 25.19 30.67 25.4 30.74 ;
    RECT 25.19 31.03 25.4 31.1 ;
    RECT 21.41 30.31 21.62 30.38 ;
    RECT 21.41 30.67 21.62 30.74 ;
    RECT 21.41 31.03 21.62 31.1 ;
    RECT 21.87 30.31 22.08 30.38 ;
    RECT 21.87 30.67 22.08 30.74 ;
    RECT 21.87 31.03 22.08 31.1 ;
    RECT 18.09 30.31 18.3 30.38 ;
    RECT 18.09 30.67 18.3 30.74 ;
    RECT 18.09 31.03 18.3 31.1 ;
    RECT 18.55 30.31 18.76 30.38 ;
    RECT 18.55 30.67 18.76 30.74 ;
    RECT 18.55 31.03 18.76 31.1 ;
    RECT 120.825 30.67 120.895 30.74 ;
    RECT 14.77 30.31 14.98 30.38 ;
    RECT 14.77 30.67 14.98 30.74 ;
    RECT 14.77 31.03 14.98 31.1 ;
    RECT 15.23 30.31 15.44 30.38 ;
    RECT 15.23 30.67 15.44 30.74 ;
    RECT 15.23 31.03 15.44 31.1 ;
    RECT 11.45 30.31 11.66 30.38 ;
    RECT 11.45 30.67 11.66 30.74 ;
    RECT 11.45 31.03 11.66 31.1 ;
    RECT 11.91 30.31 12.12 30.38 ;
    RECT 11.91 30.67 12.12 30.74 ;
    RECT 11.91 31.03 12.12 31.1 ;
    RECT 8.13 30.31 8.34 30.38 ;
    RECT 8.13 30.67 8.34 30.74 ;
    RECT 8.13 31.03 8.34 31.1 ;
    RECT 8.59 30.31 8.8 30.38 ;
    RECT 8.59 30.67 8.8 30.74 ;
    RECT 8.59 31.03 8.8 31.1 ;
    RECT 4.81 30.31 5.02 30.38 ;
    RECT 4.81 30.67 5.02 30.74 ;
    RECT 4.81 31.03 5.02 31.1 ;
    RECT 5.27 30.31 5.48 30.38 ;
    RECT 5.27 30.67 5.48 30.74 ;
    RECT 5.27 31.03 5.48 31.1 ;
    RECT 1.49 30.31 1.7 30.38 ;
    RECT 1.49 30.67 1.7 30.74 ;
    RECT 1.49 31.03 1.7 31.1 ;
    RECT 1.95 30.31 2.16 30.38 ;
    RECT 1.95 30.67 2.16 30.74 ;
    RECT 1.95 31.03 2.16 31.1 ;
    RECT 64.57 30.31 64.78 30.38 ;
    RECT 64.57 30.67 64.78 30.74 ;
    RECT 64.57 31.03 64.78 31.1 ;
    RECT 65.03 30.31 65.24 30.38 ;
    RECT 65.03 30.67 65.24 30.74 ;
    RECT 65.03 31.03 65.24 31.1 ;
    RECT 61.25 69.93 61.46 70.0 ;
    RECT 61.25 70.29 61.46 70.36 ;
    RECT 61.25 70.65 61.46 70.72 ;
    RECT 61.71 69.93 61.92 70.0 ;
    RECT 61.71 70.29 61.92 70.36 ;
    RECT 61.71 70.65 61.92 70.72 ;
    RECT 57.93 69.93 58.14 70.0 ;
    RECT 57.93 70.29 58.14 70.36 ;
    RECT 57.93 70.65 58.14 70.72 ;
    RECT 58.39 69.93 58.6 70.0 ;
    RECT 58.39 70.29 58.6 70.36 ;
    RECT 58.39 70.65 58.6 70.72 ;
    RECT 54.61 69.93 54.82 70.0 ;
    RECT 54.61 70.29 54.82 70.36 ;
    RECT 54.61 70.65 54.82 70.72 ;
    RECT 55.07 69.93 55.28 70.0 ;
    RECT 55.07 70.29 55.28 70.36 ;
    RECT 55.07 70.65 55.28 70.72 ;
    RECT 51.29 69.93 51.5 70.0 ;
    RECT 51.29 70.29 51.5 70.36 ;
    RECT 51.29 70.65 51.5 70.72 ;
    RECT 51.75 69.93 51.96 70.0 ;
    RECT 51.75 70.29 51.96 70.36 ;
    RECT 51.75 70.65 51.96 70.72 ;
    RECT 47.97 69.93 48.18 70.0 ;
    RECT 47.97 70.29 48.18 70.36 ;
    RECT 47.97 70.65 48.18 70.72 ;
    RECT 48.43 69.93 48.64 70.0 ;
    RECT 48.43 70.29 48.64 70.36 ;
    RECT 48.43 70.65 48.64 70.72 ;
    RECT 44.65 69.93 44.86 70.0 ;
    RECT 44.65 70.29 44.86 70.36 ;
    RECT 44.65 70.65 44.86 70.72 ;
    RECT 45.11 69.93 45.32 70.0 ;
    RECT 45.11 70.29 45.32 70.36 ;
    RECT 45.11 70.65 45.32 70.72 ;
    RECT 41.33 69.93 41.54 70.0 ;
    RECT 41.33 70.29 41.54 70.36 ;
    RECT 41.33 70.65 41.54 70.72 ;
    RECT 41.79 69.93 42.0 70.0 ;
    RECT 41.79 70.29 42.0 70.36 ;
    RECT 41.79 70.65 42.0 70.72 ;
    RECT 38.01 69.93 38.22 70.0 ;
    RECT 38.01 70.29 38.22 70.36 ;
    RECT 38.01 70.65 38.22 70.72 ;
    RECT 38.47 69.93 38.68 70.0 ;
    RECT 38.47 70.29 38.68 70.36 ;
    RECT 38.47 70.65 38.68 70.72 ;
    RECT 0.4 70.29 0.47 70.36 ;
    RECT 34.69 69.93 34.9 70.0 ;
    RECT 34.69 70.29 34.9 70.36 ;
    RECT 34.69 70.65 34.9 70.72 ;
    RECT 35.15 69.93 35.36 70.0 ;
    RECT 35.15 70.29 35.36 70.36 ;
    RECT 35.15 70.65 35.36 70.72 ;
    RECT 117.69 69.93 117.9 70.0 ;
    RECT 117.69 70.29 117.9 70.36 ;
    RECT 117.69 70.65 117.9 70.72 ;
    RECT 118.15 69.93 118.36 70.0 ;
    RECT 118.15 70.29 118.36 70.36 ;
    RECT 118.15 70.65 118.36 70.72 ;
    RECT 114.37 69.93 114.58 70.0 ;
    RECT 114.37 70.29 114.58 70.36 ;
    RECT 114.37 70.65 114.58 70.72 ;
    RECT 114.83 69.93 115.04 70.0 ;
    RECT 114.83 70.29 115.04 70.36 ;
    RECT 114.83 70.65 115.04 70.72 ;
    RECT 111.05 69.93 111.26 70.0 ;
    RECT 111.05 70.29 111.26 70.36 ;
    RECT 111.05 70.65 111.26 70.72 ;
    RECT 111.51 69.93 111.72 70.0 ;
    RECT 111.51 70.29 111.72 70.36 ;
    RECT 111.51 70.65 111.72 70.72 ;
    RECT 107.73 69.93 107.94 70.0 ;
    RECT 107.73 70.29 107.94 70.36 ;
    RECT 107.73 70.65 107.94 70.72 ;
    RECT 108.19 69.93 108.4 70.0 ;
    RECT 108.19 70.29 108.4 70.36 ;
    RECT 108.19 70.65 108.4 70.72 ;
    RECT 104.41 69.93 104.62 70.0 ;
    RECT 104.41 70.29 104.62 70.36 ;
    RECT 104.41 70.65 104.62 70.72 ;
    RECT 104.87 69.93 105.08 70.0 ;
    RECT 104.87 70.29 105.08 70.36 ;
    RECT 104.87 70.65 105.08 70.72 ;
    RECT 101.09 69.93 101.3 70.0 ;
    RECT 101.09 70.29 101.3 70.36 ;
    RECT 101.09 70.65 101.3 70.72 ;
    RECT 101.55 69.93 101.76 70.0 ;
    RECT 101.55 70.29 101.76 70.36 ;
    RECT 101.55 70.65 101.76 70.72 ;
    RECT 97.77 69.93 97.98 70.0 ;
    RECT 97.77 70.29 97.98 70.36 ;
    RECT 97.77 70.65 97.98 70.72 ;
    RECT 98.23 69.93 98.44 70.0 ;
    RECT 98.23 70.29 98.44 70.36 ;
    RECT 98.23 70.65 98.44 70.72 ;
    RECT 94.45 69.93 94.66 70.0 ;
    RECT 94.45 70.29 94.66 70.36 ;
    RECT 94.45 70.65 94.66 70.72 ;
    RECT 94.91 69.93 95.12 70.0 ;
    RECT 94.91 70.29 95.12 70.36 ;
    RECT 94.91 70.65 95.12 70.72 ;
    RECT 91.13 69.93 91.34 70.0 ;
    RECT 91.13 70.29 91.34 70.36 ;
    RECT 91.13 70.65 91.34 70.72 ;
    RECT 91.59 69.93 91.8 70.0 ;
    RECT 91.59 70.29 91.8 70.36 ;
    RECT 91.59 70.65 91.8 70.72 ;
    RECT 87.81 69.93 88.02 70.0 ;
    RECT 87.81 70.29 88.02 70.36 ;
    RECT 87.81 70.65 88.02 70.72 ;
    RECT 88.27 69.93 88.48 70.0 ;
    RECT 88.27 70.29 88.48 70.36 ;
    RECT 88.27 70.65 88.48 70.72 ;
    RECT 84.49 69.93 84.7 70.0 ;
    RECT 84.49 70.29 84.7 70.36 ;
    RECT 84.49 70.65 84.7 70.72 ;
    RECT 84.95 69.93 85.16 70.0 ;
    RECT 84.95 70.29 85.16 70.36 ;
    RECT 84.95 70.65 85.16 70.72 ;
    RECT 81.17 69.93 81.38 70.0 ;
    RECT 81.17 70.29 81.38 70.36 ;
    RECT 81.17 70.65 81.38 70.72 ;
    RECT 81.63 69.93 81.84 70.0 ;
    RECT 81.63 70.29 81.84 70.36 ;
    RECT 81.63 70.65 81.84 70.72 ;
    RECT 77.85 69.93 78.06 70.0 ;
    RECT 77.85 70.29 78.06 70.36 ;
    RECT 77.85 70.65 78.06 70.72 ;
    RECT 78.31 69.93 78.52 70.0 ;
    RECT 78.31 70.29 78.52 70.36 ;
    RECT 78.31 70.65 78.52 70.72 ;
    RECT 74.53 69.93 74.74 70.0 ;
    RECT 74.53 70.29 74.74 70.36 ;
    RECT 74.53 70.65 74.74 70.72 ;
    RECT 74.99 69.93 75.2 70.0 ;
    RECT 74.99 70.29 75.2 70.36 ;
    RECT 74.99 70.65 75.2 70.72 ;
    RECT 71.21 69.93 71.42 70.0 ;
    RECT 71.21 70.29 71.42 70.36 ;
    RECT 71.21 70.65 71.42 70.72 ;
    RECT 71.67 69.93 71.88 70.0 ;
    RECT 71.67 70.29 71.88 70.36 ;
    RECT 71.67 70.65 71.88 70.72 ;
    RECT 31.37 69.93 31.58 70.0 ;
    RECT 31.37 70.29 31.58 70.36 ;
    RECT 31.37 70.65 31.58 70.72 ;
    RECT 31.83 69.93 32.04 70.0 ;
    RECT 31.83 70.29 32.04 70.36 ;
    RECT 31.83 70.65 32.04 70.72 ;
    RECT 67.89 69.93 68.1 70.0 ;
    RECT 67.89 70.29 68.1 70.36 ;
    RECT 67.89 70.65 68.1 70.72 ;
    RECT 68.35 69.93 68.56 70.0 ;
    RECT 68.35 70.29 68.56 70.36 ;
    RECT 68.35 70.65 68.56 70.72 ;
    RECT 28.05 69.93 28.26 70.0 ;
    RECT 28.05 70.29 28.26 70.36 ;
    RECT 28.05 70.65 28.26 70.72 ;
    RECT 28.51 69.93 28.72 70.0 ;
    RECT 28.51 70.29 28.72 70.36 ;
    RECT 28.51 70.65 28.72 70.72 ;
    RECT 24.73 69.93 24.94 70.0 ;
    RECT 24.73 70.29 24.94 70.36 ;
    RECT 24.73 70.65 24.94 70.72 ;
    RECT 25.19 69.93 25.4 70.0 ;
    RECT 25.19 70.29 25.4 70.36 ;
    RECT 25.19 70.65 25.4 70.72 ;
    RECT 21.41 69.93 21.62 70.0 ;
    RECT 21.41 70.29 21.62 70.36 ;
    RECT 21.41 70.65 21.62 70.72 ;
    RECT 21.87 69.93 22.08 70.0 ;
    RECT 21.87 70.29 22.08 70.36 ;
    RECT 21.87 70.65 22.08 70.72 ;
    RECT 18.09 69.93 18.3 70.0 ;
    RECT 18.09 70.29 18.3 70.36 ;
    RECT 18.09 70.65 18.3 70.72 ;
    RECT 18.55 69.93 18.76 70.0 ;
    RECT 18.55 70.29 18.76 70.36 ;
    RECT 18.55 70.65 18.76 70.72 ;
    RECT 120.825 70.29 120.895 70.36 ;
    RECT 14.77 69.93 14.98 70.0 ;
    RECT 14.77 70.29 14.98 70.36 ;
    RECT 14.77 70.65 14.98 70.72 ;
    RECT 15.23 69.93 15.44 70.0 ;
    RECT 15.23 70.29 15.44 70.36 ;
    RECT 15.23 70.65 15.44 70.72 ;
    RECT 11.45 69.93 11.66 70.0 ;
    RECT 11.45 70.29 11.66 70.36 ;
    RECT 11.45 70.65 11.66 70.72 ;
    RECT 11.91 69.93 12.12 70.0 ;
    RECT 11.91 70.29 12.12 70.36 ;
    RECT 11.91 70.65 12.12 70.72 ;
    RECT 8.13 69.93 8.34 70.0 ;
    RECT 8.13 70.29 8.34 70.36 ;
    RECT 8.13 70.65 8.34 70.72 ;
    RECT 8.59 69.93 8.8 70.0 ;
    RECT 8.59 70.29 8.8 70.36 ;
    RECT 8.59 70.65 8.8 70.72 ;
    RECT 4.81 69.93 5.02 70.0 ;
    RECT 4.81 70.29 5.02 70.36 ;
    RECT 4.81 70.65 5.02 70.72 ;
    RECT 5.27 69.93 5.48 70.0 ;
    RECT 5.27 70.29 5.48 70.36 ;
    RECT 5.27 70.65 5.48 70.72 ;
    RECT 1.49 69.93 1.7 70.0 ;
    RECT 1.49 70.29 1.7 70.36 ;
    RECT 1.49 70.65 1.7 70.72 ;
    RECT 1.95 69.93 2.16 70.0 ;
    RECT 1.95 70.29 2.16 70.36 ;
    RECT 1.95 70.65 2.16 70.72 ;
    RECT 64.57 69.93 64.78 70.0 ;
    RECT 64.57 70.29 64.78 70.36 ;
    RECT 64.57 70.65 64.78 70.72 ;
    RECT 65.03 69.93 65.24 70.0 ;
    RECT 65.03 70.29 65.24 70.36 ;
    RECT 65.03 70.65 65.24 70.72 ;
    RECT 61.25 29.59 61.46 29.66 ;
    RECT 61.25 29.95 61.46 30.02 ;
    RECT 61.25 30.31 61.46 30.38 ;
    RECT 61.71 29.59 61.92 29.66 ;
    RECT 61.71 29.95 61.92 30.02 ;
    RECT 61.71 30.31 61.92 30.38 ;
    RECT 57.93 29.59 58.14 29.66 ;
    RECT 57.93 29.95 58.14 30.02 ;
    RECT 57.93 30.31 58.14 30.38 ;
    RECT 58.39 29.59 58.6 29.66 ;
    RECT 58.39 29.95 58.6 30.02 ;
    RECT 58.39 30.31 58.6 30.38 ;
    RECT 54.61 29.59 54.82 29.66 ;
    RECT 54.61 29.95 54.82 30.02 ;
    RECT 54.61 30.31 54.82 30.38 ;
    RECT 55.07 29.59 55.28 29.66 ;
    RECT 55.07 29.95 55.28 30.02 ;
    RECT 55.07 30.31 55.28 30.38 ;
    RECT 51.29 29.59 51.5 29.66 ;
    RECT 51.29 29.95 51.5 30.02 ;
    RECT 51.29 30.31 51.5 30.38 ;
    RECT 51.75 29.59 51.96 29.66 ;
    RECT 51.75 29.95 51.96 30.02 ;
    RECT 51.75 30.31 51.96 30.38 ;
    RECT 47.97 29.59 48.18 29.66 ;
    RECT 47.97 29.95 48.18 30.02 ;
    RECT 47.97 30.31 48.18 30.38 ;
    RECT 48.43 29.59 48.64 29.66 ;
    RECT 48.43 29.95 48.64 30.02 ;
    RECT 48.43 30.31 48.64 30.38 ;
    RECT 44.65 29.59 44.86 29.66 ;
    RECT 44.65 29.95 44.86 30.02 ;
    RECT 44.65 30.31 44.86 30.38 ;
    RECT 45.11 29.59 45.32 29.66 ;
    RECT 45.11 29.95 45.32 30.02 ;
    RECT 45.11 30.31 45.32 30.38 ;
    RECT 41.33 29.59 41.54 29.66 ;
    RECT 41.33 29.95 41.54 30.02 ;
    RECT 41.33 30.31 41.54 30.38 ;
    RECT 41.79 29.59 42.0 29.66 ;
    RECT 41.79 29.95 42.0 30.02 ;
    RECT 41.79 30.31 42.0 30.38 ;
    RECT 38.01 29.59 38.22 29.66 ;
    RECT 38.01 29.95 38.22 30.02 ;
    RECT 38.01 30.31 38.22 30.38 ;
    RECT 38.47 29.59 38.68 29.66 ;
    RECT 38.47 29.95 38.68 30.02 ;
    RECT 38.47 30.31 38.68 30.38 ;
    RECT 0.4 29.95 0.47 30.02 ;
    RECT 34.69 29.59 34.9 29.66 ;
    RECT 34.69 29.95 34.9 30.02 ;
    RECT 34.69 30.31 34.9 30.38 ;
    RECT 35.15 29.59 35.36 29.66 ;
    RECT 35.15 29.95 35.36 30.02 ;
    RECT 35.15 30.31 35.36 30.38 ;
    RECT 117.69 29.59 117.9 29.66 ;
    RECT 117.69 29.95 117.9 30.02 ;
    RECT 117.69 30.31 117.9 30.38 ;
    RECT 118.15 29.59 118.36 29.66 ;
    RECT 118.15 29.95 118.36 30.02 ;
    RECT 118.15 30.31 118.36 30.38 ;
    RECT 114.37 29.59 114.58 29.66 ;
    RECT 114.37 29.95 114.58 30.02 ;
    RECT 114.37 30.31 114.58 30.38 ;
    RECT 114.83 29.59 115.04 29.66 ;
    RECT 114.83 29.95 115.04 30.02 ;
    RECT 114.83 30.31 115.04 30.38 ;
    RECT 111.05 29.59 111.26 29.66 ;
    RECT 111.05 29.95 111.26 30.02 ;
    RECT 111.05 30.31 111.26 30.38 ;
    RECT 111.51 29.59 111.72 29.66 ;
    RECT 111.51 29.95 111.72 30.02 ;
    RECT 111.51 30.31 111.72 30.38 ;
    RECT 107.73 29.59 107.94 29.66 ;
    RECT 107.73 29.95 107.94 30.02 ;
    RECT 107.73 30.31 107.94 30.38 ;
    RECT 108.19 29.59 108.4 29.66 ;
    RECT 108.19 29.95 108.4 30.02 ;
    RECT 108.19 30.31 108.4 30.38 ;
    RECT 104.41 29.59 104.62 29.66 ;
    RECT 104.41 29.95 104.62 30.02 ;
    RECT 104.41 30.31 104.62 30.38 ;
    RECT 104.87 29.59 105.08 29.66 ;
    RECT 104.87 29.95 105.08 30.02 ;
    RECT 104.87 30.31 105.08 30.38 ;
    RECT 101.09 29.59 101.3 29.66 ;
    RECT 101.09 29.95 101.3 30.02 ;
    RECT 101.09 30.31 101.3 30.38 ;
    RECT 101.55 29.59 101.76 29.66 ;
    RECT 101.55 29.95 101.76 30.02 ;
    RECT 101.55 30.31 101.76 30.38 ;
    RECT 97.77 29.59 97.98 29.66 ;
    RECT 97.77 29.95 97.98 30.02 ;
    RECT 97.77 30.31 97.98 30.38 ;
    RECT 98.23 29.59 98.44 29.66 ;
    RECT 98.23 29.95 98.44 30.02 ;
    RECT 98.23 30.31 98.44 30.38 ;
    RECT 94.45 29.59 94.66 29.66 ;
    RECT 94.45 29.95 94.66 30.02 ;
    RECT 94.45 30.31 94.66 30.38 ;
    RECT 94.91 29.59 95.12 29.66 ;
    RECT 94.91 29.95 95.12 30.02 ;
    RECT 94.91 30.31 95.12 30.38 ;
    RECT 91.13 29.59 91.34 29.66 ;
    RECT 91.13 29.95 91.34 30.02 ;
    RECT 91.13 30.31 91.34 30.38 ;
    RECT 91.59 29.59 91.8 29.66 ;
    RECT 91.59 29.95 91.8 30.02 ;
    RECT 91.59 30.31 91.8 30.38 ;
    RECT 87.81 29.59 88.02 29.66 ;
    RECT 87.81 29.95 88.02 30.02 ;
    RECT 87.81 30.31 88.02 30.38 ;
    RECT 88.27 29.59 88.48 29.66 ;
    RECT 88.27 29.95 88.48 30.02 ;
    RECT 88.27 30.31 88.48 30.38 ;
    RECT 84.49 29.59 84.7 29.66 ;
    RECT 84.49 29.95 84.7 30.02 ;
    RECT 84.49 30.31 84.7 30.38 ;
    RECT 84.95 29.59 85.16 29.66 ;
    RECT 84.95 29.95 85.16 30.02 ;
    RECT 84.95 30.31 85.16 30.38 ;
    RECT 81.17 29.59 81.38 29.66 ;
    RECT 81.17 29.95 81.38 30.02 ;
    RECT 81.17 30.31 81.38 30.38 ;
    RECT 81.63 29.59 81.84 29.66 ;
    RECT 81.63 29.95 81.84 30.02 ;
    RECT 81.63 30.31 81.84 30.38 ;
    RECT 77.85 29.59 78.06 29.66 ;
    RECT 77.85 29.95 78.06 30.02 ;
    RECT 77.85 30.31 78.06 30.38 ;
    RECT 78.31 29.59 78.52 29.66 ;
    RECT 78.31 29.95 78.52 30.02 ;
    RECT 78.31 30.31 78.52 30.38 ;
    RECT 74.53 29.59 74.74 29.66 ;
    RECT 74.53 29.95 74.74 30.02 ;
    RECT 74.53 30.31 74.74 30.38 ;
    RECT 74.99 29.59 75.2 29.66 ;
    RECT 74.99 29.95 75.2 30.02 ;
    RECT 74.99 30.31 75.2 30.38 ;
    RECT 71.21 29.59 71.42 29.66 ;
    RECT 71.21 29.95 71.42 30.02 ;
    RECT 71.21 30.31 71.42 30.38 ;
    RECT 71.67 29.59 71.88 29.66 ;
    RECT 71.67 29.95 71.88 30.02 ;
    RECT 71.67 30.31 71.88 30.38 ;
    RECT 31.37 29.59 31.58 29.66 ;
    RECT 31.37 29.95 31.58 30.02 ;
    RECT 31.37 30.31 31.58 30.38 ;
    RECT 31.83 29.59 32.04 29.66 ;
    RECT 31.83 29.95 32.04 30.02 ;
    RECT 31.83 30.31 32.04 30.38 ;
    RECT 67.89 29.59 68.1 29.66 ;
    RECT 67.89 29.95 68.1 30.02 ;
    RECT 67.89 30.31 68.1 30.38 ;
    RECT 68.35 29.59 68.56 29.66 ;
    RECT 68.35 29.95 68.56 30.02 ;
    RECT 68.35 30.31 68.56 30.38 ;
    RECT 28.05 29.59 28.26 29.66 ;
    RECT 28.05 29.95 28.26 30.02 ;
    RECT 28.05 30.31 28.26 30.38 ;
    RECT 28.51 29.59 28.72 29.66 ;
    RECT 28.51 29.95 28.72 30.02 ;
    RECT 28.51 30.31 28.72 30.38 ;
    RECT 24.73 29.59 24.94 29.66 ;
    RECT 24.73 29.95 24.94 30.02 ;
    RECT 24.73 30.31 24.94 30.38 ;
    RECT 25.19 29.59 25.4 29.66 ;
    RECT 25.19 29.95 25.4 30.02 ;
    RECT 25.19 30.31 25.4 30.38 ;
    RECT 21.41 29.59 21.62 29.66 ;
    RECT 21.41 29.95 21.62 30.02 ;
    RECT 21.41 30.31 21.62 30.38 ;
    RECT 21.87 29.59 22.08 29.66 ;
    RECT 21.87 29.95 22.08 30.02 ;
    RECT 21.87 30.31 22.08 30.38 ;
    RECT 18.09 29.59 18.3 29.66 ;
    RECT 18.09 29.95 18.3 30.02 ;
    RECT 18.09 30.31 18.3 30.38 ;
    RECT 18.55 29.59 18.76 29.66 ;
    RECT 18.55 29.95 18.76 30.02 ;
    RECT 18.55 30.31 18.76 30.38 ;
    RECT 120.825 29.95 120.895 30.02 ;
    RECT 14.77 29.59 14.98 29.66 ;
    RECT 14.77 29.95 14.98 30.02 ;
    RECT 14.77 30.31 14.98 30.38 ;
    RECT 15.23 29.59 15.44 29.66 ;
    RECT 15.23 29.95 15.44 30.02 ;
    RECT 15.23 30.31 15.44 30.38 ;
    RECT 11.45 29.59 11.66 29.66 ;
    RECT 11.45 29.95 11.66 30.02 ;
    RECT 11.45 30.31 11.66 30.38 ;
    RECT 11.91 29.59 12.12 29.66 ;
    RECT 11.91 29.95 12.12 30.02 ;
    RECT 11.91 30.31 12.12 30.38 ;
    RECT 8.13 29.59 8.34 29.66 ;
    RECT 8.13 29.95 8.34 30.02 ;
    RECT 8.13 30.31 8.34 30.38 ;
    RECT 8.59 29.59 8.8 29.66 ;
    RECT 8.59 29.95 8.8 30.02 ;
    RECT 8.59 30.31 8.8 30.38 ;
    RECT 4.81 29.59 5.02 29.66 ;
    RECT 4.81 29.95 5.02 30.02 ;
    RECT 4.81 30.31 5.02 30.38 ;
    RECT 5.27 29.59 5.48 29.66 ;
    RECT 5.27 29.95 5.48 30.02 ;
    RECT 5.27 30.31 5.48 30.38 ;
    RECT 1.49 29.59 1.7 29.66 ;
    RECT 1.49 29.95 1.7 30.02 ;
    RECT 1.49 30.31 1.7 30.38 ;
    RECT 1.95 29.59 2.16 29.66 ;
    RECT 1.95 29.95 2.16 30.02 ;
    RECT 1.95 30.31 2.16 30.38 ;
    RECT 64.57 29.59 64.78 29.66 ;
    RECT 64.57 29.95 64.78 30.02 ;
    RECT 64.57 30.31 64.78 30.38 ;
    RECT 65.03 29.59 65.24 29.66 ;
    RECT 65.03 29.95 65.24 30.02 ;
    RECT 65.03 30.31 65.24 30.38 ;
    RECT 61.25 69.21 61.46 69.28 ;
    RECT 61.25 69.57 61.46 69.64 ;
    RECT 61.25 69.93 61.46 70.0 ;
    RECT 61.71 69.21 61.92 69.28 ;
    RECT 61.71 69.57 61.92 69.64 ;
    RECT 61.71 69.93 61.92 70.0 ;
    RECT 57.93 69.21 58.14 69.28 ;
    RECT 57.93 69.57 58.14 69.64 ;
    RECT 57.93 69.93 58.14 70.0 ;
    RECT 58.39 69.21 58.6 69.28 ;
    RECT 58.39 69.57 58.6 69.64 ;
    RECT 58.39 69.93 58.6 70.0 ;
    RECT 54.61 69.21 54.82 69.28 ;
    RECT 54.61 69.57 54.82 69.64 ;
    RECT 54.61 69.93 54.82 70.0 ;
    RECT 55.07 69.21 55.28 69.28 ;
    RECT 55.07 69.57 55.28 69.64 ;
    RECT 55.07 69.93 55.28 70.0 ;
    RECT 51.29 69.21 51.5 69.28 ;
    RECT 51.29 69.57 51.5 69.64 ;
    RECT 51.29 69.93 51.5 70.0 ;
    RECT 51.75 69.21 51.96 69.28 ;
    RECT 51.75 69.57 51.96 69.64 ;
    RECT 51.75 69.93 51.96 70.0 ;
    RECT 47.97 69.21 48.18 69.28 ;
    RECT 47.97 69.57 48.18 69.64 ;
    RECT 47.97 69.93 48.18 70.0 ;
    RECT 48.43 69.21 48.64 69.28 ;
    RECT 48.43 69.57 48.64 69.64 ;
    RECT 48.43 69.93 48.64 70.0 ;
    RECT 44.65 69.21 44.86 69.28 ;
    RECT 44.65 69.57 44.86 69.64 ;
    RECT 44.65 69.93 44.86 70.0 ;
    RECT 45.11 69.21 45.32 69.28 ;
    RECT 45.11 69.57 45.32 69.64 ;
    RECT 45.11 69.93 45.32 70.0 ;
    RECT 41.33 69.21 41.54 69.28 ;
    RECT 41.33 69.57 41.54 69.64 ;
    RECT 41.33 69.93 41.54 70.0 ;
    RECT 41.79 69.21 42.0 69.28 ;
    RECT 41.79 69.57 42.0 69.64 ;
    RECT 41.79 69.93 42.0 70.0 ;
    RECT 38.01 69.21 38.22 69.28 ;
    RECT 38.01 69.57 38.22 69.64 ;
    RECT 38.01 69.93 38.22 70.0 ;
    RECT 38.47 69.21 38.68 69.28 ;
    RECT 38.47 69.57 38.68 69.64 ;
    RECT 38.47 69.93 38.68 70.0 ;
    RECT 0.4 69.57 0.47 69.64 ;
    RECT 34.69 69.21 34.9 69.28 ;
    RECT 34.69 69.57 34.9 69.64 ;
    RECT 34.69 69.93 34.9 70.0 ;
    RECT 35.15 69.21 35.36 69.28 ;
    RECT 35.15 69.57 35.36 69.64 ;
    RECT 35.15 69.93 35.36 70.0 ;
    RECT 117.69 69.21 117.9 69.28 ;
    RECT 117.69 69.57 117.9 69.64 ;
    RECT 117.69 69.93 117.9 70.0 ;
    RECT 118.15 69.21 118.36 69.28 ;
    RECT 118.15 69.57 118.36 69.64 ;
    RECT 118.15 69.93 118.36 70.0 ;
    RECT 114.37 69.21 114.58 69.28 ;
    RECT 114.37 69.57 114.58 69.64 ;
    RECT 114.37 69.93 114.58 70.0 ;
    RECT 114.83 69.21 115.04 69.28 ;
    RECT 114.83 69.57 115.04 69.64 ;
    RECT 114.83 69.93 115.04 70.0 ;
    RECT 111.05 69.21 111.26 69.28 ;
    RECT 111.05 69.57 111.26 69.64 ;
    RECT 111.05 69.93 111.26 70.0 ;
    RECT 111.51 69.21 111.72 69.28 ;
    RECT 111.51 69.57 111.72 69.64 ;
    RECT 111.51 69.93 111.72 70.0 ;
    RECT 107.73 69.21 107.94 69.28 ;
    RECT 107.73 69.57 107.94 69.64 ;
    RECT 107.73 69.93 107.94 70.0 ;
    RECT 108.19 69.21 108.4 69.28 ;
    RECT 108.19 69.57 108.4 69.64 ;
    RECT 108.19 69.93 108.4 70.0 ;
    RECT 104.41 69.21 104.62 69.28 ;
    RECT 104.41 69.57 104.62 69.64 ;
    RECT 104.41 69.93 104.62 70.0 ;
    RECT 104.87 69.21 105.08 69.28 ;
    RECT 104.87 69.57 105.08 69.64 ;
    RECT 104.87 69.93 105.08 70.0 ;
    RECT 101.09 69.21 101.3 69.28 ;
    RECT 101.09 69.57 101.3 69.64 ;
    RECT 101.09 69.93 101.3 70.0 ;
    RECT 101.55 69.21 101.76 69.28 ;
    RECT 101.55 69.57 101.76 69.64 ;
    RECT 101.55 69.93 101.76 70.0 ;
    RECT 97.77 69.21 97.98 69.28 ;
    RECT 97.77 69.57 97.98 69.64 ;
    RECT 97.77 69.93 97.98 70.0 ;
    RECT 98.23 69.21 98.44 69.28 ;
    RECT 98.23 69.57 98.44 69.64 ;
    RECT 98.23 69.93 98.44 70.0 ;
    RECT 94.45 69.21 94.66 69.28 ;
    RECT 94.45 69.57 94.66 69.64 ;
    RECT 94.45 69.93 94.66 70.0 ;
    RECT 94.91 69.21 95.12 69.28 ;
    RECT 94.91 69.57 95.12 69.64 ;
    RECT 94.91 69.93 95.12 70.0 ;
    RECT 91.13 69.21 91.34 69.28 ;
    RECT 91.13 69.57 91.34 69.64 ;
    RECT 91.13 69.93 91.34 70.0 ;
    RECT 91.59 69.21 91.8 69.28 ;
    RECT 91.59 69.57 91.8 69.64 ;
    RECT 91.59 69.93 91.8 70.0 ;
    RECT 87.81 69.21 88.02 69.28 ;
    RECT 87.81 69.57 88.02 69.64 ;
    RECT 87.81 69.93 88.02 70.0 ;
    RECT 88.27 69.21 88.48 69.28 ;
    RECT 88.27 69.57 88.48 69.64 ;
    RECT 88.27 69.93 88.48 70.0 ;
    RECT 84.49 69.21 84.7 69.28 ;
    RECT 84.49 69.57 84.7 69.64 ;
    RECT 84.49 69.93 84.7 70.0 ;
    RECT 84.95 69.21 85.16 69.28 ;
    RECT 84.95 69.57 85.16 69.64 ;
    RECT 84.95 69.93 85.16 70.0 ;
    RECT 81.17 69.21 81.38 69.28 ;
    RECT 81.17 69.57 81.38 69.64 ;
    RECT 81.17 69.93 81.38 70.0 ;
    RECT 81.63 69.21 81.84 69.28 ;
    RECT 81.63 69.57 81.84 69.64 ;
    RECT 81.63 69.93 81.84 70.0 ;
    RECT 77.85 69.21 78.06 69.28 ;
    RECT 77.85 69.57 78.06 69.64 ;
    RECT 77.85 69.93 78.06 70.0 ;
    RECT 78.31 69.21 78.52 69.28 ;
    RECT 78.31 69.57 78.52 69.64 ;
    RECT 78.31 69.93 78.52 70.0 ;
    RECT 74.53 69.21 74.74 69.28 ;
    RECT 74.53 69.57 74.74 69.64 ;
    RECT 74.53 69.93 74.74 70.0 ;
    RECT 74.99 69.21 75.2 69.28 ;
    RECT 74.99 69.57 75.2 69.64 ;
    RECT 74.99 69.93 75.2 70.0 ;
    RECT 71.21 69.21 71.42 69.28 ;
    RECT 71.21 69.57 71.42 69.64 ;
    RECT 71.21 69.93 71.42 70.0 ;
    RECT 71.67 69.21 71.88 69.28 ;
    RECT 71.67 69.57 71.88 69.64 ;
    RECT 71.67 69.93 71.88 70.0 ;
    RECT 31.37 69.21 31.58 69.28 ;
    RECT 31.37 69.57 31.58 69.64 ;
    RECT 31.37 69.93 31.58 70.0 ;
    RECT 31.83 69.21 32.04 69.28 ;
    RECT 31.83 69.57 32.04 69.64 ;
    RECT 31.83 69.93 32.04 70.0 ;
    RECT 67.89 69.21 68.1 69.28 ;
    RECT 67.89 69.57 68.1 69.64 ;
    RECT 67.89 69.93 68.1 70.0 ;
    RECT 68.35 69.21 68.56 69.28 ;
    RECT 68.35 69.57 68.56 69.64 ;
    RECT 68.35 69.93 68.56 70.0 ;
    RECT 28.05 69.21 28.26 69.28 ;
    RECT 28.05 69.57 28.26 69.64 ;
    RECT 28.05 69.93 28.26 70.0 ;
    RECT 28.51 69.21 28.72 69.28 ;
    RECT 28.51 69.57 28.72 69.64 ;
    RECT 28.51 69.93 28.72 70.0 ;
    RECT 24.73 69.21 24.94 69.28 ;
    RECT 24.73 69.57 24.94 69.64 ;
    RECT 24.73 69.93 24.94 70.0 ;
    RECT 25.19 69.21 25.4 69.28 ;
    RECT 25.19 69.57 25.4 69.64 ;
    RECT 25.19 69.93 25.4 70.0 ;
    RECT 21.41 69.21 21.62 69.28 ;
    RECT 21.41 69.57 21.62 69.64 ;
    RECT 21.41 69.93 21.62 70.0 ;
    RECT 21.87 69.21 22.08 69.28 ;
    RECT 21.87 69.57 22.08 69.64 ;
    RECT 21.87 69.93 22.08 70.0 ;
    RECT 18.09 69.21 18.3 69.28 ;
    RECT 18.09 69.57 18.3 69.64 ;
    RECT 18.09 69.93 18.3 70.0 ;
    RECT 18.55 69.21 18.76 69.28 ;
    RECT 18.55 69.57 18.76 69.64 ;
    RECT 18.55 69.93 18.76 70.0 ;
    RECT 120.825 69.57 120.895 69.64 ;
    RECT 14.77 69.21 14.98 69.28 ;
    RECT 14.77 69.57 14.98 69.64 ;
    RECT 14.77 69.93 14.98 70.0 ;
    RECT 15.23 69.21 15.44 69.28 ;
    RECT 15.23 69.57 15.44 69.64 ;
    RECT 15.23 69.93 15.44 70.0 ;
    RECT 11.45 69.21 11.66 69.28 ;
    RECT 11.45 69.57 11.66 69.64 ;
    RECT 11.45 69.93 11.66 70.0 ;
    RECT 11.91 69.21 12.12 69.28 ;
    RECT 11.91 69.57 12.12 69.64 ;
    RECT 11.91 69.93 12.12 70.0 ;
    RECT 8.13 69.21 8.34 69.28 ;
    RECT 8.13 69.57 8.34 69.64 ;
    RECT 8.13 69.93 8.34 70.0 ;
    RECT 8.59 69.21 8.8 69.28 ;
    RECT 8.59 69.57 8.8 69.64 ;
    RECT 8.59 69.93 8.8 70.0 ;
    RECT 4.81 69.21 5.02 69.28 ;
    RECT 4.81 69.57 5.02 69.64 ;
    RECT 4.81 69.93 5.02 70.0 ;
    RECT 5.27 69.21 5.48 69.28 ;
    RECT 5.27 69.57 5.48 69.64 ;
    RECT 5.27 69.93 5.48 70.0 ;
    RECT 1.49 69.21 1.7 69.28 ;
    RECT 1.49 69.57 1.7 69.64 ;
    RECT 1.49 69.93 1.7 70.0 ;
    RECT 1.95 69.21 2.16 69.28 ;
    RECT 1.95 69.57 2.16 69.64 ;
    RECT 1.95 69.93 2.16 70.0 ;
    RECT 64.57 69.21 64.78 69.28 ;
    RECT 64.57 69.57 64.78 69.64 ;
    RECT 64.57 69.93 64.78 70.0 ;
    RECT 65.03 69.21 65.24 69.28 ;
    RECT 65.03 69.57 65.24 69.64 ;
    RECT 65.03 69.93 65.24 70.0 ;
    RECT 61.25 28.87 61.46 28.94 ;
    RECT 61.25 29.23 61.46 29.3 ;
    RECT 61.25 29.59 61.46 29.66 ;
    RECT 61.71 28.87 61.92 28.94 ;
    RECT 61.71 29.23 61.92 29.3 ;
    RECT 61.71 29.59 61.92 29.66 ;
    RECT 57.93 28.87 58.14 28.94 ;
    RECT 57.93 29.23 58.14 29.3 ;
    RECT 57.93 29.59 58.14 29.66 ;
    RECT 58.39 28.87 58.6 28.94 ;
    RECT 58.39 29.23 58.6 29.3 ;
    RECT 58.39 29.59 58.6 29.66 ;
    RECT 54.61 28.87 54.82 28.94 ;
    RECT 54.61 29.23 54.82 29.3 ;
    RECT 54.61 29.59 54.82 29.66 ;
    RECT 55.07 28.87 55.28 28.94 ;
    RECT 55.07 29.23 55.28 29.3 ;
    RECT 55.07 29.59 55.28 29.66 ;
    RECT 51.29 28.87 51.5 28.94 ;
    RECT 51.29 29.23 51.5 29.3 ;
    RECT 51.29 29.59 51.5 29.66 ;
    RECT 51.75 28.87 51.96 28.94 ;
    RECT 51.75 29.23 51.96 29.3 ;
    RECT 51.75 29.59 51.96 29.66 ;
    RECT 47.97 28.87 48.18 28.94 ;
    RECT 47.97 29.23 48.18 29.3 ;
    RECT 47.97 29.59 48.18 29.66 ;
    RECT 48.43 28.87 48.64 28.94 ;
    RECT 48.43 29.23 48.64 29.3 ;
    RECT 48.43 29.59 48.64 29.66 ;
    RECT 44.65 28.87 44.86 28.94 ;
    RECT 44.65 29.23 44.86 29.3 ;
    RECT 44.65 29.59 44.86 29.66 ;
    RECT 45.11 28.87 45.32 28.94 ;
    RECT 45.11 29.23 45.32 29.3 ;
    RECT 45.11 29.59 45.32 29.66 ;
    RECT 41.33 28.87 41.54 28.94 ;
    RECT 41.33 29.23 41.54 29.3 ;
    RECT 41.33 29.59 41.54 29.66 ;
    RECT 41.79 28.87 42.0 28.94 ;
    RECT 41.79 29.23 42.0 29.3 ;
    RECT 41.79 29.59 42.0 29.66 ;
    RECT 38.01 28.87 38.22 28.94 ;
    RECT 38.01 29.23 38.22 29.3 ;
    RECT 38.01 29.59 38.22 29.66 ;
    RECT 38.47 28.87 38.68 28.94 ;
    RECT 38.47 29.23 38.68 29.3 ;
    RECT 38.47 29.59 38.68 29.66 ;
    RECT 0.4 29.23 0.47 29.3 ;
    RECT 34.69 28.87 34.9 28.94 ;
    RECT 34.69 29.23 34.9 29.3 ;
    RECT 34.69 29.59 34.9 29.66 ;
    RECT 35.15 28.87 35.36 28.94 ;
    RECT 35.15 29.23 35.36 29.3 ;
    RECT 35.15 29.59 35.36 29.66 ;
    RECT 117.69 28.87 117.9 28.94 ;
    RECT 117.69 29.23 117.9 29.3 ;
    RECT 117.69 29.59 117.9 29.66 ;
    RECT 118.15 28.87 118.36 28.94 ;
    RECT 118.15 29.23 118.36 29.3 ;
    RECT 118.15 29.59 118.36 29.66 ;
    RECT 114.37 28.87 114.58 28.94 ;
    RECT 114.37 29.23 114.58 29.3 ;
    RECT 114.37 29.59 114.58 29.66 ;
    RECT 114.83 28.87 115.04 28.94 ;
    RECT 114.83 29.23 115.04 29.3 ;
    RECT 114.83 29.59 115.04 29.66 ;
    RECT 111.05 28.87 111.26 28.94 ;
    RECT 111.05 29.23 111.26 29.3 ;
    RECT 111.05 29.59 111.26 29.66 ;
    RECT 111.51 28.87 111.72 28.94 ;
    RECT 111.51 29.23 111.72 29.3 ;
    RECT 111.51 29.59 111.72 29.66 ;
    RECT 107.73 28.87 107.94 28.94 ;
    RECT 107.73 29.23 107.94 29.3 ;
    RECT 107.73 29.59 107.94 29.66 ;
    RECT 108.19 28.87 108.4 28.94 ;
    RECT 108.19 29.23 108.4 29.3 ;
    RECT 108.19 29.59 108.4 29.66 ;
    RECT 104.41 28.87 104.62 28.94 ;
    RECT 104.41 29.23 104.62 29.3 ;
    RECT 104.41 29.59 104.62 29.66 ;
    RECT 104.87 28.87 105.08 28.94 ;
    RECT 104.87 29.23 105.08 29.3 ;
    RECT 104.87 29.59 105.08 29.66 ;
    RECT 101.09 28.87 101.3 28.94 ;
    RECT 101.09 29.23 101.3 29.3 ;
    RECT 101.09 29.59 101.3 29.66 ;
    RECT 101.55 28.87 101.76 28.94 ;
    RECT 101.55 29.23 101.76 29.3 ;
    RECT 101.55 29.59 101.76 29.66 ;
    RECT 97.77 28.87 97.98 28.94 ;
    RECT 97.77 29.23 97.98 29.3 ;
    RECT 97.77 29.59 97.98 29.66 ;
    RECT 98.23 28.87 98.44 28.94 ;
    RECT 98.23 29.23 98.44 29.3 ;
    RECT 98.23 29.59 98.44 29.66 ;
    RECT 94.45 28.87 94.66 28.94 ;
    RECT 94.45 29.23 94.66 29.3 ;
    RECT 94.45 29.59 94.66 29.66 ;
    RECT 94.91 28.87 95.12 28.94 ;
    RECT 94.91 29.23 95.12 29.3 ;
    RECT 94.91 29.59 95.12 29.66 ;
    RECT 91.13 28.87 91.34 28.94 ;
    RECT 91.13 29.23 91.34 29.3 ;
    RECT 91.13 29.59 91.34 29.66 ;
    RECT 91.59 28.87 91.8 28.94 ;
    RECT 91.59 29.23 91.8 29.3 ;
    RECT 91.59 29.59 91.8 29.66 ;
    RECT 87.81 28.87 88.02 28.94 ;
    RECT 87.81 29.23 88.02 29.3 ;
    RECT 87.81 29.59 88.02 29.66 ;
    RECT 88.27 28.87 88.48 28.94 ;
    RECT 88.27 29.23 88.48 29.3 ;
    RECT 88.27 29.59 88.48 29.66 ;
    RECT 84.49 28.87 84.7 28.94 ;
    RECT 84.49 29.23 84.7 29.3 ;
    RECT 84.49 29.59 84.7 29.66 ;
    RECT 84.95 28.87 85.16 28.94 ;
    RECT 84.95 29.23 85.16 29.3 ;
    RECT 84.95 29.59 85.16 29.66 ;
    RECT 81.17 28.87 81.38 28.94 ;
    RECT 81.17 29.23 81.38 29.3 ;
    RECT 81.17 29.59 81.38 29.66 ;
    RECT 81.63 28.87 81.84 28.94 ;
    RECT 81.63 29.23 81.84 29.3 ;
    RECT 81.63 29.59 81.84 29.66 ;
    RECT 77.85 28.87 78.06 28.94 ;
    RECT 77.85 29.23 78.06 29.3 ;
    RECT 77.85 29.59 78.06 29.66 ;
    RECT 78.31 28.87 78.52 28.94 ;
    RECT 78.31 29.23 78.52 29.3 ;
    RECT 78.31 29.59 78.52 29.66 ;
    RECT 74.53 28.87 74.74 28.94 ;
    RECT 74.53 29.23 74.74 29.3 ;
    RECT 74.53 29.59 74.74 29.66 ;
    RECT 74.99 28.87 75.2 28.94 ;
    RECT 74.99 29.23 75.2 29.3 ;
    RECT 74.99 29.59 75.2 29.66 ;
    RECT 71.21 28.87 71.42 28.94 ;
    RECT 71.21 29.23 71.42 29.3 ;
    RECT 71.21 29.59 71.42 29.66 ;
    RECT 71.67 28.87 71.88 28.94 ;
    RECT 71.67 29.23 71.88 29.3 ;
    RECT 71.67 29.59 71.88 29.66 ;
    RECT 31.37 28.87 31.58 28.94 ;
    RECT 31.37 29.23 31.58 29.3 ;
    RECT 31.37 29.59 31.58 29.66 ;
    RECT 31.83 28.87 32.04 28.94 ;
    RECT 31.83 29.23 32.04 29.3 ;
    RECT 31.83 29.59 32.04 29.66 ;
    RECT 67.89 28.87 68.1 28.94 ;
    RECT 67.89 29.23 68.1 29.3 ;
    RECT 67.89 29.59 68.1 29.66 ;
    RECT 68.35 28.87 68.56 28.94 ;
    RECT 68.35 29.23 68.56 29.3 ;
    RECT 68.35 29.59 68.56 29.66 ;
    RECT 28.05 28.87 28.26 28.94 ;
    RECT 28.05 29.23 28.26 29.3 ;
    RECT 28.05 29.59 28.26 29.66 ;
    RECT 28.51 28.87 28.72 28.94 ;
    RECT 28.51 29.23 28.72 29.3 ;
    RECT 28.51 29.59 28.72 29.66 ;
    RECT 24.73 28.87 24.94 28.94 ;
    RECT 24.73 29.23 24.94 29.3 ;
    RECT 24.73 29.59 24.94 29.66 ;
    RECT 25.19 28.87 25.4 28.94 ;
    RECT 25.19 29.23 25.4 29.3 ;
    RECT 25.19 29.59 25.4 29.66 ;
    RECT 21.41 28.87 21.62 28.94 ;
    RECT 21.41 29.23 21.62 29.3 ;
    RECT 21.41 29.59 21.62 29.66 ;
    RECT 21.87 28.87 22.08 28.94 ;
    RECT 21.87 29.23 22.08 29.3 ;
    RECT 21.87 29.59 22.08 29.66 ;
    RECT 18.09 28.87 18.3 28.94 ;
    RECT 18.09 29.23 18.3 29.3 ;
    RECT 18.09 29.59 18.3 29.66 ;
    RECT 18.55 28.87 18.76 28.94 ;
    RECT 18.55 29.23 18.76 29.3 ;
    RECT 18.55 29.59 18.76 29.66 ;
    RECT 120.825 29.23 120.895 29.3 ;
    RECT 14.77 28.87 14.98 28.94 ;
    RECT 14.77 29.23 14.98 29.3 ;
    RECT 14.77 29.59 14.98 29.66 ;
    RECT 15.23 28.87 15.44 28.94 ;
    RECT 15.23 29.23 15.44 29.3 ;
    RECT 15.23 29.59 15.44 29.66 ;
    RECT 11.45 28.87 11.66 28.94 ;
    RECT 11.45 29.23 11.66 29.3 ;
    RECT 11.45 29.59 11.66 29.66 ;
    RECT 11.91 28.87 12.12 28.94 ;
    RECT 11.91 29.23 12.12 29.3 ;
    RECT 11.91 29.59 12.12 29.66 ;
    RECT 8.13 28.87 8.34 28.94 ;
    RECT 8.13 29.23 8.34 29.3 ;
    RECT 8.13 29.59 8.34 29.66 ;
    RECT 8.59 28.87 8.8 28.94 ;
    RECT 8.59 29.23 8.8 29.3 ;
    RECT 8.59 29.59 8.8 29.66 ;
    RECT 4.81 28.87 5.02 28.94 ;
    RECT 4.81 29.23 5.02 29.3 ;
    RECT 4.81 29.59 5.02 29.66 ;
    RECT 5.27 28.87 5.48 28.94 ;
    RECT 5.27 29.23 5.48 29.3 ;
    RECT 5.27 29.59 5.48 29.66 ;
    RECT 1.49 28.87 1.7 28.94 ;
    RECT 1.49 29.23 1.7 29.3 ;
    RECT 1.49 29.59 1.7 29.66 ;
    RECT 1.95 28.87 2.16 28.94 ;
    RECT 1.95 29.23 2.16 29.3 ;
    RECT 1.95 29.59 2.16 29.66 ;
    RECT 64.57 28.87 64.78 28.94 ;
    RECT 64.57 29.23 64.78 29.3 ;
    RECT 64.57 29.59 64.78 29.66 ;
    RECT 65.03 28.87 65.24 28.94 ;
    RECT 65.03 29.23 65.24 29.3 ;
    RECT 65.03 29.59 65.24 29.66 ;
    RECT 61.25 68.49 61.46 68.56 ;
    RECT 61.25 68.85 61.46 68.92 ;
    RECT 61.25 69.21 61.46 69.28 ;
    RECT 61.71 68.49 61.92 68.56 ;
    RECT 61.71 68.85 61.92 68.92 ;
    RECT 61.71 69.21 61.92 69.28 ;
    RECT 57.93 68.49 58.14 68.56 ;
    RECT 57.93 68.85 58.14 68.92 ;
    RECT 57.93 69.21 58.14 69.28 ;
    RECT 58.39 68.49 58.6 68.56 ;
    RECT 58.39 68.85 58.6 68.92 ;
    RECT 58.39 69.21 58.6 69.28 ;
    RECT 54.61 68.49 54.82 68.56 ;
    RECT 54.61 68.85 54.82 68.92 ;
    RECT 54.61 69.21 54.82 69.28 ;
    RECT 55.07 68.49 55.28 68.56 ;
    RECT 55.07 68.85 55.28 68.92 ;
    RECT 55.07 69.21 55.28 69.28 ;
    RECT 51.29 68.49 51.5 68.56 ;
    RECT 51.29 68.85 51.5 68.92 ;
    RECT 51.29 69.21 51.5 69.28 ;
    RECT 51.75 68.49 51.96 68.56 ;
    RECT 51.75 68.85 51.96 68.92 ;
    RECT 51.75 69.21 51.96 69.28 ;
    RECT 47.97 68.49 48.18 68.56 ;
    RECT 47.97 68.85 48.18 68.92 ;
    RECT 47.97 69.21 48.18 69.28 ;
    RECT 48.43 68.49 48.64 68.56 ;
    RECT 48.43 68.85 48.64 68.92 ;
    RECT 48.43 69.21 48.64 69.28 ;
    RECT 44.65 68.49 44.86 68.56 ;
    RECT 44.65 68.85 44.86 68.92 ;
    RECT 44.65 69.21 44.86 69.28 ;
    RECT 45.11 68.49 45.32 68.56 ;
    RECT 45.11 68.85 45.32 68.92 ;
    RECT 45.11 69.21 45.32 69.28 ;
    RECT 41.33 68.49 41.54 68.56 ;
    RECT 41.33 68.85 41.54 68.92 ;
    RECT 41.33 69.21 41.54 69.28 ;
    RECT 41.79 68.49 42.0 68.56 ;
    RECT 41.79 68.85 42.0 68.92 ;
    RECT 41.79 69.21 42.0 69.28 ;
    RECT 38.01 68.49 38.22 68.56 ;
    RECT 38.01 68.85 38.22 68.92 ;
    RECT 38.01 69.21 38.22 69.28 ;
    RECT 38.47 68.49 38.68 68.56 ;
    RECT 38.47 68.85 38.68 68.92 ;
    RECT 38.47 69.21 38.68 69.28 ;
    RECT 0.4 68.85 0.47 68.92 ;
    RECT 34.69 68.49 34.9 68.56 ;
    RECT 34.69 68.85 34.9 68.92 ;
    RECT 34.69 69.21 34.9 69.28 ;
    RECT 35.15 68.49 35.36 68.56 ;
    RECT 35.15 68.85 35.36 68.92 ;
    RECT 35.15 69.21 35.36 69.28 ;
    RECT 117.69 68.49 117.9 68.56 ;
    RECT 117.69 68.85 117.9 68.92 ;
    RECT 117.69 69.21 117.9 69.28 ;
    RECT 118.15 68.49 118.36 68.56 ;
    RECT 118.15 68.85 118.36 68.92 ;
    RECT 118.15 69.21 118.36 69.28 ;
    RECT 114.37 68.49 114.58 68.56 ;
    RECT 114.37 68.85 114.58 68.92 ;
    RECT 114.37 69.21 114.58 69.28 ;
    RECT 114.83 68.49 115.04 68.56 ;
    RECT 114.83 68.85 115.04 68.92 ;
    RECT 114.83 69.21 115.04 69.28 ;
    RECT 111.05 68.49 111.26 68.56 ;
    RECT 111.05 68.85 111.26 68.92 ;
    RECT 111.05 69.21 111.26 69.28 ;
    RECT 111.51 68.49 111.72 68.56 ;
    RECT 111.51 68.85 111.72 68.92 ;
    RECT 111.51 69.21 111.72 69.28 ;
    RECT 107.73 68.49 107.94 68.56 ;
    RECT 107.73 68.85 107.94 68.92 ;
    RECT 107.73 69.21 107.94 69.28 ;
    RECT 108.19 68.49 108.4 68.56 ;
    RECT 108.19 68.85 108.4 68.92 ;
    RECT 108.19 69.21 108.4 69.28 ;
    RECT 104.41 68.49 104.62 68.56 ;
    RECT 104.41 68.85 104.62 68.92 ;
    RECT 104.41 69.21 104.62 69.28 ;
    RECT 104.87 68.49 105.08 68.56 ;
    RECT 104.87 68.85 105.08 68.92 ;
    RECT 104.87 69.21 105.08 69.28 ;
    RECT 101.09 68.49 101.3 68.56 ;
    RECT 101.09 68.85 101.3 68.92 ;
    RECT 101.09 69.21 101.3 69.28 ;
    RECT 101.55 68.49 101.76 68.56 ;
    RECT 101.55 68.85 101.76 68.92 ;
    RECT 101.55 69.21 101.76 69.28 ;
    RECT 97.77 68.49 97.98 68.56 ;
    RECT 97.77 68.85 97.98 68.92 ;
    RECT 97.77 69.21 97.98 69.28 ;
    RECT 98.23 68.49 98.44 68.56 ;
    RECT 98.23 68.85 98.44 68.92 ;
    RECT 98.23 69.21 98.44 69.28 ;
    RECT 94.45 68.49 94.66 68.56 ;
    RECT 94.45 68.85 94.66 68.92 ;
    RECT 94.45 69.21 94.66 69.28 ;
    RECT 94.91 68.49 95.12 68.56 ;
    RECT 94.91 68.85 95.12 68.92 ;
    RECT 94.91 69.21 95.12 69.28 ;
    RECT 91.13 68.49 91.34 68.56 ;
    RECT 91.13 68.85 91.34 68.92 ;
    RECT 91.13 69.21 91.34 69.28 ;
    RECT 91.59 68.49 91.8 68.56 ;
    RECT 91.59 68.85 91.8 68.92 ;
    RECT 91.59 69.21 91.8 69.28 ;
    RECT 87.81 68.49 88.02 68.56 ;
    RECT 87.81 68.85 88.02 68.92 ;
    RECT 87.81 69.21 88.02 69.28 ;
    RECT 88.27 68.49 88.48 68.56 ;
    RECT 88.27 68.85 88.48 68.92 ;
    RECT 88.27 69.21 88.48 69.28 ;
    RECT 84.49 68.49 84.7 68.56 ;
    RECT 84.49 68.85 84.7 68.92 ;
    RECT 84.49 69.21 84.7 69.28 ;
    RECT 84.95 68.49 85.16 68.56 ;
    RECT 84.95 68.85 85.16 68.92 ;
    RECT 84.95 69.21 85.16 69.28 ;
    RECT 81.17 68.49 81.38 68.56 ;
    RECT 81.17 68.85 81.38 68.92 ;
    RECT 81.17 69.21 81.38 69.28 ;
    RECT 81.63 68.49 81.84 68.56 ;
    RECT 81.63 68.85 81.84 68.92 ;
    RECT 81.63 69.21 81.84 69.28 ;
    RECT 77.85 68.49 78.06 68.56 ;
    RECT 77.85 68.85 78.06 68.92 ;
    RECT 77.85 69.21 78.06 69.28 ;
    RECT 78.31 68.49 78.52 68.56 ;
    RECT 78.31 68.85 78.52 68.92 ;
    RECT 78.31 69.21 78.52 69.28 ;
    RECT 74.53 68.49 74.74 68.56 ;
    RECT 74.53 68.85 74.74 68.92 ;
    RECT 74.53 69.21 74.74 69.28 ;
    RECT 74.99 68.49 75.2 68.56 ;
    RECT 74.99 68.85 75.2 68.92 ;
    RECT 74.99 69.21 75.2 69.28 ;
    RECT 71.21 68.49 71.42 68.56 ;
    RECT 71.21 68.85 71.42 68.92 ;
    RECT 71.21 69.21 71.42 69.28 ;
    RECT 71.67 68.49 71.88 68.56 ;
    RECT 71.67 68.85 71.88 68.92 ;
    RECT 71.67 69.21 71.88 69.28 ;
    RECT 31.37 68.49 31.58 68.56 ;
    RECT 31.37 68.85 31.58 68.92 ;
    RECT 31.37 69.21 31.58 69.28 ;
    RECT 31.83 68.49 32.04 68.56 ;
    RECT 31.83 68.85 32.04 68.92 ;
    RECT 31.83 69.21 32.04 69.28 ;
    RECT 67.89 68.49 68.1 68.56 ;
    RECT 67.89 68.85 68.1 68.92 ;
    RECT 67.89 69.21 68.1 69.28 ;
    RECT 68.35 68.49 68.56 68.56 ;
    RECT 68.35 68.85 68.56 68.92 ;
    RECT 68.35 69.21 68.56 69.28 ;
    RECT 28.05 68.49 28.26 68.56 ;
    RECT 28.05 68.85 28.26 68.92 ;
    RECT 28.05 69.21 28.26 69.28 ;
    RECT 28.51 68.49 28.72 68.56 ;
    RECT 28.51 68.85 28.72 68.92 ;
    RECT 28.51 69.21 28.72 69.28 ;
    RECT 24.73 68.49 24.94 68.56 ;
    RECT 24.73 68.85 24.94 68.92 ;
    RECT 24.73 69.21 24.94 69.28 ;
    RECT 25.19 68.49 25.4 68.56 ;
    RECT 25.19 68.85 25.4 68.92 ;
    RECT 25.19 69.21 25.4 69.28 ;
    RECT 21.41 68.49 21.62 68.56 ;
    RECT 21.41 68.85 21.62 68.92 ;
    RECT 21.41 69.21 21.62 69.28 ;
    RECT 21.87 68.49 22.08 68.56 ;
    RECT 21.87 68.85 22.08 68.92 ;
    RECT 21.87 69.21 22.08 69.28 ;
    RECT 18.09 68.49 18.3 68.56 ;
    RECT 18.09 68.85 18.3 68.92 ;
    RECT 18.09 69.21 18.3 69.28 ;
    RECT 18.55 68.49 18.76 68.56 ;
    RECT 18.55 68.85 18.76 68.92 ;
    RECT 18.55 69.21 18.76 69.28 ;
    RECT 120.825 68.85 120.895 68.92 ;
    RECT 14.77 68.49 14.98 68.56 ;
    RECT 14.77 68.85 14.98 68.92 ;
    RECT 14.77 69.21 14.98 69.28 ;
    RECT 15.23 68.49 15.44 68.56 ;
    RECT 15.23 68.85 15.44 68.92 ;
    RECT 15.23 69.21 15.44 69.28 ;
    RECT 11.45 68.49 11.66 68.56 ;
    RECT 11.45 68.85 11.66 68.92 ;
    RECT 11.45 69.21 11.66 69.28 ;
    RECT 11.91 68.49 12.12 68.56 ;
    RECT 11.91 68.85 12.12 68.92 ;
    RECT 11.91 69.21 12.12 69.28 ;
    RECT 8.13 68.49 8.34 68.56 ;
    RECT 8.13 68.85 8.34 68.92 ;
    RECT 8.13 69.21 8.34 69.28 ;
    RECT 8.59 68.49 8.8 68.56 ;
    RECT 8.59 68.85 8.8 68.92 ;
    RECT 8.59 69.21 8.8 69.28 ;
    RECT 4.81 68.49 5.02 68.56 ;
    RECT 4.81 68.85 5.02 68.92 ;
    RECT 4.81 69.21 5.02 69.28 ;
    RECT 5.27 68.49 5.48 68.56 ;
    RECT 5.27 68.85 5.48 68.92 ;
    RECT 5.27 69.21 5.48 69.28 ;
    RECT 1.49 68.49 1.7 68.56 ;
    RECT 1.49 68.85 1.7 68.92 ;
    RECT 1.49 69.21 1.7 69.28 ;
    RECT 1.95 68.49 2.16 68.56 ;
    RECT 1.95 68.85 2.16 68.92 ;
    RECT 1.95 69.21 2.16 69.28 ;
    RECT 64.57 68.49 64.78 68.56 ;
    RECT 64.57 68.85 64.78 68.92 ;
    RECT 64.57 69.21 64.78 69.28 ;
    RECT 65.03 68.49 65.24 68.56 ;
    RECT 65.03 68.85 65.24 68.92 ;
    RECT 65.03 69.21 65.24 69.28 ;
    RECT 61.25 67.77 61.46 67.84 ;
    RECT 61.25 68.13 61.46 68.2 ;
    RECT 61.25 68.49 61.46 68.56 ;
    RECT 61.71 67.77 61.92 67.84 ;
    RECT 61.71 68.13 61.92 68.2 ;
    RECT 61.71 68.49 61.92 68.56 ;
    RECT 57.93 67.77 58.14 67.84 ;
    RECT 57.93 68.13 58.14 68.2 ;
    RECT 57.93 68.49 58.14 68.56 ;
    RECT 58.39 67.77 58.6 67.84 ;
    RECT 58.39 68.13 58.6 68.2 ;
    RECT 58.39 68.49 58.6 68.56 ;
    RECT 54.61 67.77 54.82 67.84 ;
    RECT 54.61 68.13 54.82 68.2 ;
    RECT 54.61 68.49 54.82 68.56 ;
    RECT 55.07 67.77 55.28 67.84 ;
    RECT 55.07 68.13 55.28 68.2 ;
    RECT 55.07 68.49 55.28 68.56 ;
    RECT 51.29 67.77 51.5 67.84 ;
    RECT 51.29 68.13 51.5 68.2 ;
    RECT 51.29 68.49 51.5 68.56 ;
    RECT 51.75 67.77 51.96 67.84 ;
    RECT 51.75 68.13 51.96 68.2 ;
    RECT 51.75 68.49 51.96 68.56 ;
    RECT 47.97 67.77 48.18 67.84 ;
    RECT 47.97 68.13 48.18 68.2 ;
    RECT 47.97 68.49 48.18 68.56 ;
    RECT 48.43 67.77 48.64 67.84 ;
    RECT 48.43 68.13 48.64 68.2 ;
    RECT 48.43 68.49 48.64 68.56 ;
    RECT 44.65 67.77 44.86 67.84 ;
    RECT 44.65 68.13 44.86 68.2 ;
    RECT 44.65 68.49 44.86 68.56 ;
    RECT 45.11 67.77 45.32 67.84 ;
    RECT 45.11 68.13 45.32 68.2 ;
    RECT 45.11 68.49 45.32 68.56 ;
    RECT 41.33 67.77 41.54 67.84 ;
    RECT 41.33 68.13 41.54 68.2 ;
    RECT 41.33 68.49 41.54 68.56 ;
    RECT 41.79 67.77 42.0 67.84 ;
    RECT 41.79 68.13 42.0 68.2 ;
    RECT 41.79 68.49 42.0 68.56 ;
    RECT 38.01 67.77 38.22 67.84 ;
    RECT 38.01 68.13 38.22 68.2 ;
    RECT 38.01 68.49 38.22 68.56 ;
    RECT 38.47 67.77 38.68 67.84 ;
    RECT 38.47 68.13 38.68 68.2 ;
    RECT 38.47 68.49 38.68 68.56 ;
    RECT 0.4 68.13 0.47 68.2 ;
    RECT 34.69 67.77 34.9 67.84 ;
    RECT 34.69 68.13 34.9 68.2 ;
    RECT 34.69 68.49 34.9 68.56 ;
    RECT 35.15 67.77 35.36 67.84 ;
    RECT 35.15 68.13 35.36 68.2 ;
    RECT 35.15 68.49 35.36 68.56 ;
    RECT 117.69 67.77 117.9 67.84 ;
    RECT 117.69 68.13 117.9 68.2 ;
    RECT 117.69 68.49 117.9 68.56 ;
    RECT 118.15 67.77 118.36 67.84 ;
    RECT 118.15 68.13 118.36 68.2 ;
    RECT 118.15 68.49 118.36 68.56 ;
    RECT 114.37 67.77 114.58 67.84 ;
    RECT 114.37 68.13 114.58 68.2 ;
    RECT 114.37 68.49 114.58 68.56 ;
    RECT 114.83 67.77 115.04 67.84 ;
    RECT 114.83 68.13 115.04 68.2 ;
    RECT 114.83 68.49 115.04 68.56 ;
    RECT 111.05 67.77 111.26 67.84 ;
    RECT 111.05 68.13 111.26 68.2 ;
    RECT 111.05 68.49 111.26 68.56 ;
    RECT 111.51 67.77 111.72 67.84 ;
    RECT 111.51 68.13 111.72 68.2 ;
    RECT 111.51 68.49 111.72 68.56 ;
    RECT 107.73 67.77 107.94 67.84 ;
    RECT 107.73 68.13 107.94 68.2 ;
    RECT 107.73 68.49 107.94 68.56 ;
    RECT 108.19 67.77 108.4 67.84 ;
    RECT 108.19 68.13 108.4 68.2 ;
    RECT 108.19 68.49 108.4 68.56 ;
    RECT 104.41 67.77 104.62 67.84 ;
    RECT 104.41 68.13 104.62 68.2 ;
    RECT 104.41 68.49 104.62 68.56 ;
    RECT 104.87 67.77 105.08 67.84 ;
    RECT 104.87 68.13 105.08 68.2 ;
    RECT 104.87 68.49 105.08 68.56 ;
    RECT 101.09 67.77 101.3 67.84 ;
    RECT 101.09 68.13 101.3 68.2 ;
    RECT 101.09 68.49 101.3 68.56 ;
    RECT 101.55 67.77 101.76 67.84 ;
    RECT 101.55 68.13 101.76 68.2 ;
    RECT 101.55 68.49 101.76 68.56 ;
    RECT 97.77 67.77 97.98 67.84 ;
    RECT 97.77 68.13 97.98 68.2 ;
    RECT 97.77 68.49 97.98 68.56 ;
    RECT 98.23 67.77 98.44 67.84 ;
    RECT 98.23 68.13 98.44 68.2 ;
    RECT 98.23 68.49 98.44 68.56 ;
    RECT 94.45 67.77 94.66 67.84 ;
    RECT 94.45 68.13 94.66 68.2 ;
    RECT 94.45 68.49 94.66 68.56 ;
    RECT 94.91 67.77 95.12 67.84 ;
    RECT 94.91 68.13 95.12 68.2 ;
    RECT 94.91 68.49 95.12 68.56 ;
    RECT 91.13 67.77 91.34 67.84 ;
    RECT 91.13 68.13 91.34 68.2 ;
    RECT 91.13 68.49 91.34 68.56 ;
    RECT 91.59 67.77 91.8 67.84 ;
    RECT 91.59 68.13 91.8 68.2 ;
    RECT 91.59 68.49 91.8 68.56 ;
    RECT 87.81 67.77 88.02 67.84 ;
    RECT 87.81 68.13 88.02 68.2 ;
    RECT 87.81 68.49 88.02 68.56 ;
    RECT 88.27 67.77 88.48 67.84 ;
    RECT 88.27 68.13 88.48 68.2 ;
    RECT 88.27 68.49 88.48 68.56 ;
    RECT 84.49 67.77 84.7 67.84 ;
    RECT 84.49 68.13 84.7 68.2 ;
    RECT 84.49 68.49 84.7 68.56 ;
    RECT 84.95 67.77 85.16 67.84 ;
    RECT 84.95 68.13 85.16 68.2 ;
    RECT 84.95 68.49 85.16 68.56 ;
    RECT 81.17 67.77 81.38 67.84 ;
    RECT 81.17 68.13 81.38 68.2 ;
    RECT 81.17 68.49 81.38 68.56 ;
    RECT 81.63 67.77 81.84 67.84 ;
    RECT 81.63 68.13 81.84 68.2 ;
    RECT 81.63 68.49 81.84 68.56 ;
    RECT 77.85 67.77 78.06 67.84 ;
    RECT 77.85 68.13 78.06 68.2 ;
    RECT 77.85 68.49 78.06 68.56 ;
    RECT 78.31 67.77 78.52 67.84 ;
    RECT 78.31 68.13 78.52 68.2 ;
    RECT 78.31 68.49 78.52 68.56 ;
    RECT 74.53 67.77 74.74 67.84 ;
    RECT 74.53 68.13 74.74 68.2 ;
    RECT 74.53 68.49 74.74 68.56 ;
    RECT 74.99 67.77 75.2 67.84 ;
    RECT 74.99 68.13 75.2 68.2 ;
    RECT 74.99 68.49 75.2 68.56 ;
    RECT 71.21 67.77 71.42 67.84 ;
    RECT 71.21 68.13 71.42 68.2 ;
    RECT 71.21 68.49 71.42 68.56 ;
    RECT 71.67 67.77 71.88 67.84 ;
    RECT 71.67 68.13 71.88 68.2 ;
    RECT 71.67 68.49 71.88 68.56 ;
    RECT 31.37 67.77 31.58 67.84 ;
    RECT 31.37 68.13 31.58 68.2 ;
    RECT 31.37 68.49 31.58 68.56 ;
    RECT 31.83 67.77 32.04 67.84 ;
    RECT 31.83 68.13 32.04 68.2 ;
    RECT 31.83 68.49 32.04 68.56 ;
    RECT 67.89 67.77 68.1 67.84 ;
    RECT 67.89 68.13 68.1 68.2 ;
    RECT 67.89 68.49 68.1 68.56 ;
    RECT 68.35 67.77 68.56 67.84 ;
    RECT 68.35 68.13 68.56 68.2 ;
    RECT 68.35 68.49 68.56 68.56 ;
    RECT 28.05 67.77 28.26 67.84 ;
    RECT 28.05 68.13 28.26 68.2 ;
    RECT 28.05 68.49 28.26 68.56 ;
    RECT 28.51 67.77 28.72 67.84 ;
    RECT 28.51 68.13 28.72 68.2 ;
    RECT 28.51 68.49 28.72 68.56 ;
    RECT 24.73 67.77 24.94 67.84 ;
    RECT 24.73 68.13 24.94 68.2 ;
    RECT 24.73 68.49 24.94 68.56 ;
    RECT 25.19 67.77 25.4 67.84 ;
    RECT 25.19 68.13 25.4 68.2 ;
    RECT 25.19 68.49 25.4 68.56 ;
    RECT 21.41 67.77 21.62 67.84 ;
    RECT 21.41 68.13 21.62 68.2 ;
    RECT 21.41 68.49 21.62 68.56 ;
    RECT 21.87 67.77 22.08 67.84 ;
    RECT 21.87 68.13 22.08 68.2 ;
    RECT 21.87 68.49 22.08 68.56 ;
    RECT 18.09 67.77 18.3 67.84 ;
    RECT 18.09 68.13 18.3 68.2 ;
    RECT 18.09 68.49 18.3 68.56 ;
    RECT 18.55 67.77 18.76 67.84 ;
    RECT 18.55 68.13 18.76 68.2 ;
    RECT 18.55 68.49 18.76 68.56 ;
    RECT 120.825 68.13 120.895 68.2 ;
    RECT 14.77 67.77 14.98 67.84 ;
    RECT 14.77 68.13 14.98 68.2 ;
    RECT 14.77 68.49 14.98 68.56 ;
    RECT 15.23 67.77 15.44 67.84 ;
    RECT 15.23 68.13 15.44 68.2 ;
    RECT 15.23 68.49 15.44 68.56 ;
    RECT 11.45 67.77 11.66 67.84 ;
    RECT 11.45 68.13 11.66 68.2 ;
    RECT 11.45 68.49 11.66 68.56 ;
    RECT 11.91 67.77 12.12 67.84 ;
    RECT 11.91 68.13 12.12 68.2 ;
    RECT 11.91 68.49 12.12 68.56 ;
    RECT 8.13 67.77 8.34 67.84 ;
    RECT 8.13 68.13 8.34 68.2 ;
    RECT 8.13 68.49 8.34 68.56 ;
    RECT 8.59 67.77 8.8 67.84 ;
    RECT 8.59 68.13 8.8 68.2 ;
    RECT 8.59 68.49 8.8 68.56 ;
    RECT 4.81 67.77 5.02 67.84 ;
    RECT 4.81 68.13 5.02 68.2 ;
    RECT 4.81 68.49 5.02 68.56 ;
    RECT 5.27 67.77 5.48 67.84 ;
    RECT 5.27 68.13 5.48 68.2 ;
    RECT 5.27 68.49 5.48 68.56 ;
    RECT 1.49 67.77 1.7 67.84 ;
    RECT 1.49 68.13 1.7 68.2 ;
    RECT 1.49 68.49 1.7 68.56 ;
    RECT 1.95 67.77 2.16 67.84 ;
    RECT 1.95 68.13 2.16 68.2 ;
    RECT 1.95 68.49 2.16 68.56 ;
    RECT 64.57 67.77 64.78 67.84 ;
    RECT 64.57 68.13 64.78 68.2 ;
    RECT 64.57 68.49 64.78 68.56 ;
    RECT 65.03 67.77 65.24 67.84 ;
    RECT 65.03 68.13 65.24 68.2 ;
    RECT 65.03 68.49 65.24 68.56 ;
    RECT 61.25 67.05 61.46 67.12 ;
    RECT 61.25 67.41 61.46 67.48 ;
    RECT 61.25 67.77 61.46 67.84 ;
    RECT 61.71 67.05 61.92 67.12 ;
    RECT 61.71 67.41 61.92 67.48 ;
    RECT 61.71 67.77 61.92 67.84 ;
    RECT 57.93 67.05 58.14 67.12 ;
    RECT 57.93 67.41 58.14 67.48 ;
    RECT 57.93 67.77 58.14 67.84 ;
    RECT 58.39 67.05 58.6 67.12 ;
    RECT 58.39 67.41 58.6 67.48 ;
    RECT 58.39 67.77 58.6 67.84 ;
    RECT 54.61 67.05 54.82 67.12 ;
    RECT 54.61 67.41 54.82 67.48 ;
    RECT 54.61 67.77 54.82 67.84 ;
    RECT 55.07 67.05 55.28 67.12 ;
    RECT 55.07 67.41 55.28 67.48 ;
    RECT 55.07 67.77 55.28 67.84 ;
    RECT 51.29 67.05 51.5 67.12 ;
    RECT 51.29 67.41 51.5 67.48 ;
    RECT 51.29 67.77 51.5 67.84 ;
    RECT 51.75 67.05 51.96 67.12 ;
    RECT 51.75 67.41 51.96 67.48 ;
    RECT 51.75 67.77 51.96 67.84 ;
    RECT 47.97 67.05 48.18 67.12 ;
    RECT 47.97 67.41 48.18 67.48 ;
    RECT 47.97 67.77 48.18 67.84 ;
    RECT 48.43 67.05 48.64 67.12 ;
    RECT 48.43 67.41 48.64 67.48 ;
    RECT 48.43 67.77 48.64 67.84 ;
    RECT 44.65 67.05 44.86 67.12 ;
    RECT 44.65 67.41 44.86 67.48 ;
    RECT 44.65 67.77 44.86 67.84 ;
    RECT 45.11 67.05 45.32 67.12 ;
    RECT 45.11 67.41 45.32 67.48 ;
    RECT 45.11 67.77 45.32 67.84 ;
    RECT 41.33 67.05 41.54 67.12 ;
    RECT 41.33 67.41 41.54 67.48 ;
    RECT 41.33 67.77 41.54 67.84 ;
    RECT 41.79 67.05 42.0 67.12 ;
    RECT 41.79 67.41 42.0 67.48 ;
    RECT 41.79 67.77 42.0 67.84 ;
    RECT 38.01 67.05 38.22 67.12 ;
    RECT 38.01 67.41 38.22 67.48 ;
    RECT 38.01 67.77 38.22 67.84 ;
    RECT 38.47 67.05 38.68 67.12 ;
    RECT 38.47 67.41 38.68 67.48 ;
    RECT 38.47 67.77 38.68 67.84 ;
    RECT 0.4 67.41 0.47 67.48 ;
    RECT 34.69 67.05 34.9 67.12 ;
    RECT 34.69 67.41 34.9 67.48 ;
    RECT 34.69 67.77 34.9 67.84 ;
    RECT 35.15 67.05 35.36 67.12 ;
    RECT 35.15 67.41 35.36 67.48 ;
    RECT 35.15 67.77 35.36 67.84 ;
    RECT 117.69 67.05 117.9 67.12 ;
    RECT 117.69 67.41 117.9 67.48 ;
    RECT 117.69 67.77 117.9 67.84 ;
    RECT 118.15 67.05 118.36 67.12 ;
    RECT 118.15 67.41 118.36 67.48 ;
    RECT 118.15 67.77 118.36 67.84 ;
    RECT 114.37 67.05 114.58 67.12 ;
    RECT 114.37 67.41 114.58 67.48 ;
    RECT 114.37 67.77 114.58 67.84 ;
    RECT 114.83 67.05 115.04 67.12 ;
    RECT 114.83 67.41 115.04 67.48 ;
    RECT 114.83 67.77 115.04 67.84 ;
    RECT 111.05 67.05 111.26 67.12 ;
    RECT 111.05 67.41 111.26 67.48 ;
    RECT 111.05 67.77 111.26 67.84 ;
    RECT 111.51 67.05 111.72 67.12 ;
    RECT 111.51 67.41 111.72 67.48 ;
    RECT 111.51 67.77 111.72 67.84 ;
    RECT 107.73 67.05 107.94 67.12 ;
    RECT 107.73 67.41 107.94 67.48 ;
    RECT 107.73 67.77 107.94 67.84 ;
    RECT 108.19 67.05 108.4 67.12 ;
    RECT 108.19 67.41 108.4 67.48 ;
    RECT 108.19 67.77 108.4 67.84 ;
    RECT 104.41 67.05 104.62 67.12 ;
    RECT 104.41 67.41 104.62 67.48 ;
    RECT 104.41 67.77 104.62 67.84 ;
    RECT 104.87 67.05 105.08 67.12 ;
    RECT 104.87 67.41 105.08 67.48 ;
    RECT 104.87 67.77 105.08 67.84 ;
    RECT 101.09 67.05 101.3 67.12 ;
    RECT 101.09 67.41 101.3 67.48 ;
    RECT 101.09 67.77 101.3 67.84 ;
    RECT 101.55 67.05 101.76 67.12 ;
    RECT 101.55 67.41 101.76 67.48 ;
    RECT 101.55 67.77 101.76 67.84 ;
    RECT 97.77 67.05 97.98 67.12 ;
    RECT 97.77 67.41 97.98 67.48 ;
    RECT 97.77 67.77 97.98 67.84 ;
    RECT 98.23 67.05 98.44 67.12 ;
    RECT 98.23 67.41 98.44 67.48 ;
    RECT 98.23 67.77 98.44 67.84 ;
    RECT 94.45 67.05 94.66 67.12 ;
    RECT 94.45 67.41 94.66 67.48 ;
    RECT 94.45 67.77 94.66 67.84 ;
    RECT 94.91 67.05 95.12 67.12 ;
    RECT 94.91 67.41 95.12 67.48 ;
    RECT 94.91 67.77 95.12 67.84 ;
    RECT 91.13 67.05 91.34 67.12 ;
    RECT 91.13 67.41 91.34 67.48 ;
    RECT 91.13 67.77 91.34 67.84 ;
    RECT 91.59 67.05 91.8 67.12 ;
    RECT 91.59 67.41 91.8 67.48 ;
    RECT 91.59 67.77 91.8 67.84 ;
    RECT 87.81 67.05 88.02 67.12 ;
    RECT 87.81 67.41 88.02 67.48 ;
    RECT 87.81 67.77 88.02 67.84 ;
    RECT 88.27 67.05 88.48 67.12 ;
    RECT 88.27 67.41 88.48 67.48 ;
    RECT 88.27 67.77 88.48 67.84 ;
    RECT 84.49 67.05 84.7 67.12 ;
    RECT 84.49 67.41 84.7 67.48 ;
    RECT 84.49 67.77 84.7 67.84 ;
    RECT 84.95 67.05 85.16 67.12 ;
    RECT 84.95 67.41 85.16 67.48 ;
    RECT 84.95 67.77 85.16 67.84 ;
    RECT 81.17 67.05 81.38 67.12 ;
    RECT 81.17 67.41 81.38 67.48 ;
    RECT 81.17 67.77 81.38 67.84 ;
    RECT 81.63 67.05 81.84 67.12 ;
    RECT 81.63 67.41 81.84 67.48 ;
    RECT 81.63 67.77 81.84 67.84 ;
    RECT 77.85 67.05 78.06 67.12 ;
    RECT 77.85 67.41 78.06 67.48 ;
    RECT 77.85 67.77 78.06 67.84 ;
    RECT 78.31 67.05 78.52 67.12 ;
    RECT 78.31 67.41 78.52 67.48 ;
    RECT 78.31 67.77 78.52 67.84 ;
    RECT 74.53 67.05 74.74 67.12 ;
    RECT 74.53 67.41 74.74 67.48 ;
    RECT 74.53 67.77 74.74 67.84 ;
    RECT 74.99 67.05 75.2 67.12 ;
    RECT 74.99 67.41 75.2 67.48 ;
    RECT 74.99 67.77 75.2 67.84 ;
    RECT 71.21 67.05 71.42 67.12 ;
    RECT 71.21 67.41 71.42 67.48 ;
    RECT 71.21 67.77 71.42 67.84 ;
    RECT 71.67 67.05 71.88 67.12 ;
    RECT 71.67 67.41 71.88 67.48 ;
    RECT 71.67 67.77 71.88 67.84 ;
    RECT 31.37 67.05 31.58 67.12 ;
    RECT 31.37 67.41 31.58 67.48 ;
    RECT 31.37 67.77 31.58 67.84 ;
    RECT 31.83 67.05 32.04 67.12 ;
    RECT 31.83 67.41 32.04 67.48 ;
    RECT 31.83 67.77 32.04 67.84 ;
    RECT 67.89 67.05 68.1 67.12 ;
    RECT 67.89 67.41 68.1 67.48 ;
    RECT 67.89 67.77 68.1 67.84 ;
    RECT 68.35 67.05 68.56 67.12 ;
    RECT 68.35 67.41 68.56 67.48 ;
    RECT 68.35 67.77 68.56 67.84 ;
    RECT 28.05 67.05 28.26 67.12 ;
    RECT 28.05 67.41 28.26 67.48 ;
    RECT 28.05 67.77 28.26 67.84 ;
    RECT 28.51 67.05 28.72 67.12 ;
    RECT 28.51 67.41 28.72 67.48 ;
    RECT 28.51 67.77 28.72 67.84 ;
    RECT 24.73 67.05 24.94 67.12 ;
    RECT 24.73 67.41 24.94 67.48 ;
    RECT 24.73 67.77 24.94 67.84 ;
    RECT 25.19 67.05 25.4 67.12 ;
    RECT 25.19 67.41 25.4 67.48 ;
    RECT 25.19 67.77 25.4 67.84 ;
    RECT 21.41 67.05 21.62 67.12 ;
    RECT 21.41 67.41 21.62 67.48 ;
    RECT 21.41 67.77 21.62 67.84 ;
    RECT 21.87 67.05 22.08 67.12 ;
    RECT 21.87 67.41 22.08 67.48 ;
    RECT 21.87 67.77 22.08 67.84 ;
    RECT 18.09 67.05 18.3 67.12 ;
    RECT 18.09 67.41 18.3 67.48 ;
    RECT 18.09 67.77 18.3 67.84 ;
    RECT 18.55 67.05 18.76 67.12 ;
    RECT 18.55 67.41 18.76 67.48 ;
    RECT 18.55 67.77 18.76 67.84 ;
    RECT 120.825 67.41 120.895 67.48 ;
    RECT 14.77 67.05 14.98 67.12 ;
    RECT 14.77 67.41 14.98 67.48 ;
    RECT 14.77 67.77 14.98 67.84 ;
    RECT 15.23 67.05 15.44 67.12 ;
    RECT 15.23 67.41 15.44 67.48 ;
    RECT 15.23 67.77 15.44 67.84 ;
    RECT 11.45 67.05 11.66 67.12 ;
    RECT 11.45 67.41 11.66 67.48 ;
    RECT 11.45 67.77 11.66 67.84 ;
    RECT 11.91 67.05 12.12 67.12 ;
    RECT 11.91 67.41 12.12 67.48 ;
    RECT 11.91 67.77 12.12 67.84 ;
    RECT 8.13 67.05 8.34 67.12 ;
    RECT 8.13 67.41 8.34 67.48 ;
    RECT 8.13 67.77 8.34 67.84 ;
    RECT 8.59 67.05 8.8 67.12 ;
    RECT 8.59 67.41 8.8 67.48 ;
    RECT 8.59 67.77 8.8 67.84 ;
    RECT 4.81 67.05 5.02 67.12 ;
    RECT 4.81 67.41 5.02 67.48 ;
    RECT 4.81 67.77 5.02 67.84 ;
    RECT 5.27 67.05 5.48 67.12 ;
    RECT 5.27 67.41 5.48 67.48 ;
    RECT 5.27 67.77 5.48 67.84 ;
    RECT 1.49 67.05 1.7 67.12 ;
    RECT 1.49 67.41 1.7 67.48 ;
    RECT 1.49 67.77 1.7 67.84 ;
    RECT 1.95 67.05 2.16 67.12 ;
    RECT 1.95 67.41 2.16 67.48 ;
    RECT 1.95 67.77 2.16 67.84 ;
    RECT 64.57 67.05 64.78 67.12 ;
    RECT 64.57 67.41 64.78 67.48 ;
    RECT 64.57 67.77 64.78 67.84 ;
    RECT 65.03 67.05 65.24 67.12 ;
    RECT 65.03 67.41 65.24 67.48 ;
    RECT 65.03 67.77 65.24 67.84 ;
    RECT 61.25 66.33 61.46 66.4 ;
    RECT 61.25 66.69 61.46 66.76 ;
    RECT 61.25 67.05 61.46 67.12 ;
    RECT 61.71 66.33 61.92 66.4 ;
    RECT 61.71 66.69 61.92 66.76 ;
    RECT 61.71 67.05 61.92 67.12 ;
    RECT 57.93 66.33 58.14 66.4 ;
    RECT 57.93 66.69 58.14 66.76 ;
    RECT 57.93 67.05 58.14 67.12 ;
    RECT 58.39 66.33 58.6 66.4 ;
    RECT 58.39 66.69 58.6 66.76 ;
    RECT 58.39 67.05 58.6 67.12 ;
    RECT 54.61 66.33 54.82 66.4 ;
    RECT 54.61 66.69 54.82 66.76 ;
    RECT 54.61 67.05 54.82 67.12 ;
    RECT 55.07 66.33 55.28 66.4 ;
    RECT 55.07 66.69 55.28 66.76 ;
    RECT 55.07 67.05 55.28 67.12 ;
    RECT 51.29 66.33 51.5 66.4 ;
    RECT 51.29 66.69 51.5 66.76 ;
    RECT 51.29 67.05 51.5 67.12 ;
    RECT 51.75 66.33 51.96 66.4 ;
    RECT 51.75 66.69 51.96 66.76 ;
    RECT 51.75 67.05 51.96 67.12 ;
    RECT 47.97 66.33 48.18 66.4 ;
    RECT 47.97 66.69 48.18 66.76 ;
    RECT 47.97 67.05 48.18 67.12 ;
    RECT 48.43 66.33 48.64 66.4 ;
    RECT 48.43 66.69 48.64 66.76 ;
    RECT 48.43 67.05 48.64 67.12 ;
    RECT 44.65 66.33 44.86 66.4 ;
    RECT 44.65 66.69 44.86 66.76 ;
    RECT 44.65 67.05 44.86 67.12 ;
    RECT 45.11 66.33 45.32 66.4 ;
    RECT 45.11 66.69 45.32 66.76 ;
    RECT 45.11 67.05 45.32 67.12 ;
    RECT 41.33 66.33 41.54 66.4 ;
    RECT 41.33 66.69 41.54 66.76 ;
    RECT 41.33 67.05 41.54 67.12 ;
    RECT 41.79 66.33 42.0 66.4 ;
    RECT 41.79 66.69 42.0 66.76 ;
    RECT 41.79 67.05 42.0 67.12 ;
    RECT 38.01 66.33 38.22 66.4 ;
    RECT 38.01 66.69 38.22 66.76 ;
    RECT 38.01 67.05 38.22 67.12 ;
    RECT 38.47 66.33 38.68 66.4 ;
    RECT 38.47 66.69 38.68 66.76 ;
    RECT 38.47 67.05 38.68 67.12 ;
    RECT 0.4 66.69 0.47 66.76 ;
    RECT 34.69 66.33 34.9 66.4 ;
    RECT 34.69 66.69 34.9 66.76 ;
    RECT 34.69 67.05 34.9 67.12 ;
    RECT 35.15 66.33 35.36 66.4 ;
    RECT 35.15 66.69 35.36 66.76 ;
    RECT 35.15 67.05 35.36 67.12 ;
    RECT 117.69 66.33 117.9 66.4 ;
    RECT 117.69 66.69 117.9 66.76 ;
    RECT 117.69 67.05 117.9 67.12 ;
    RECT 118.15 66.33 118.36 66.4 ;
    RECT 118.15 66.69 118.36 66.76 ;
    RECT 118.15 67.05 118.36 67.12 ;
    RECT 114.37 66.33 114.58 66.4 ;
    RECT 114.37 66.69 114.58 66.76 ;
    RECT 114.37 67.05 114.58 67.12 ;
    RECT 114.83 66.33 115.04 66.4 ;
    RECT 114.83 66.69 115.04 66.76 ;
    RECT 114.83 67.05 115.04 67.12 ;
    RECT 111.05 66.33 111.26 66.4 ;
    RECT 111.05 66.69 111.26 66.76 ;
    RECT 111.05 67.05 111.26 67.12 ;
    RECT 111.51 66.33 111.72 66.4 ;
    RECT 111.51 66.69 111.72 66.76 ;
    RECT 111.51 67.05 111.72 67.12 ;
    RECT 107.73 66.33 107.94 66.4 ;
    RECT 107.73 66.69 107.94 66.76 ;
    RECT 107.73 67.05 107.94 67.12 ;
    RECT 108.19 66.33 108.4 66.4 ;
    RECT 108.19 66.69 108.4 66.76 ;
    RECT 108.19 67.05 108.4 67.12 ;
    RECT 104.41 66.33 104.62 66.4 ;
    RECT 104.41 66.69 104.62 66.76 ;
    RECT 104.41 67.05 104.62 67.12 ;
    RECT 104.87 66.33 105.08 66.4 ;
    RECT 104.87 66.69 105.08 66.76 ;
    RECT 104.87 67.05 105.08 67.12 ;
    RECT 101.09 66.33 101.3 66.4 ;
    RECT 101.09 66.69 101.3 66.76 ;
    RECT 101.09 67.05 101.3 67.12 ;
    RECT 101.55 66.33 101.76 66.4 ;
    RECT 101.55 66.69 101.76 66.76 ;
    RECT 101.55 67.05 101.76 67.12 ;
    RECT 97.77 66.33 97.98 66.4 ;
    RECT 97.77 66.69 97.98 66.76 ;
    RECT 97.77 67.05 97.98 67.12 ;
    RECT 98.23 66.33 98.44 66.4 ;
    RECT 98.23 66.69 98.44 66.76 ;
    RECT 98.23 67.05 98.44 67.12 ;
    RECT 94.45 66.33 94.66 66.4 ;
    RECT 94.45 66.69 94.66 66.76 ;
    RECT 94.45 67.05 94.66 67.12 ;
    RECT 94.91 66.33 95.12 66.4 ;
    RECT 94.91 66.69 95.12 66.76 ;
    RECT 94.91 67.05 95.12 67.12 ;
    RECT 91.13 66.33 91.34 66.4 ;
    RECT 91.13 66.69 91.34 66.76 ;
    RECT 91.13 67.05 91.34 67.12 ;
    RECT 91.59 66.33 91.8 66.4 ;
    RECT 91.59 66.69 91.8 66.76 ;
    RECT 91.59 67.05 91.8 67.12 ;
    RECT 87.81 66.33 88.02 66.4 ;
    RECT 87.81 66.69 88.02 66.76 ;
    RECT 87.81 67.05 88.02 67.12 ;
    RECT 88.27 66.33 88.48 66.4 ;
    RECT 88.27 66.69 88.48 66.76 ;
    RECT 88.27 67.05 88.48 67.12 ;
    RECT 84.49 66.33 84.7 66.4 ;
    RECT 84.49 66.69 84.7 66.76 ;
    RECT 84.49 67.05 84.7 67.12 ;
    RECT 84.95 66.33 85.16 66.4 ;
    RECT 84.95 66.69 85.16 66.76 ;
    RECT 84.95 67.05 85.16 67.12 ;
    RECT 81.17 66.33 81.38 66.4 ;
    RECT 81.17 66.69 81.38 66.76 ;
    RECT 81.17 67.05 81.38 67.12 ;
    RECT 81.63 66.33 81.84 66.4 ;
    RECT 81.63 66.69 81.84 66.76 ;
    RECT 81.63 67.05 81.84 67.12 ;
    RECT 77.85 66.33 78.06 66.4 ;
    RECT 77.85 66.69 78.06 66.76 ;
    RECT 77.85 67.05 78.06 67.12 ;
    RECT 78.31 66.33 78.52 66.4 ;
    RECT 78.31 66.69 78.52 66.76 ;
    RECT 78.31 67.05 78.52 67.12 ;
    RECT 74.53 66.33 74.74 66.4 ;
    RECT 74.53 66.69 74.74 66.76 ;
    RECT 74.53 67.05 74.74 67.12 ;
    RECT 74.99 66.33 75.2 66.4 ;
    RECT 74.99 66.69 75.2 66.76 ;
    RECT 74.99 67.05 75.2 67.12 ;
    RECT 71.21 66.33 71.42 66.4 ;
    RECT 71.21 66.69 71.42 66.76 ;
    RECT 71.21 67.05 71.42 67.12 ;
    RECT 71.67 66.33 71.88 66.4 ;
    RECT 71.67 66.69 71.88 66.76 ;
    RECT 71.67 67.05 71.88 67.12 ;
    RECT 31.37 66.33 31.58 66.4 ;
    RECT 31.37 66.69 31.58 66.76 ;
    RECT 31.37 67.05 31.58 67.12 ;
    RECT 31.83 66.33 32.04 66.4 ;
    RECT 31.83 66.69 32.04 66.76 ;
    RECT 31.83 67.05 32.04 67.12 ;
    RECT 67.89 66.33 68.1 66.4 ;
    RECT 67.89 66.69 68.1 66.76 ;
    RECT 67.89 67.05 68.1 67.12 ;
    RECT 68.35 66.33 68.56 66.4 ;
    RECT 68.35 66.69 68.56 66.76 ;
    RECT 68.35 67.05 68.56 67.12 ;
    RECT 28.05 66.33 28.26 66.4 ;
    RECT 28.05 66.69 28.26 66.76 ;
    RECT 28.05 67.05 28.26 67.12 ;
    RECT 28.51 66.33 28.72 66.4 ;
    RECT 28.51 66.69 28.72 66.76 ;
    RECT 28.51 67.05 28.72 67.12 ;
    RECT 24.73 66.33 24.94 66.4 ;
    RECT 24.73 66.69 24.94 66.76 ;
    RECT 24.73 67.05 24.94 67.12 ;
    RECT 25.19 66.33 25.4 66.4 ;
    RECT 25.19 66.69 25.4 66.76 ;
    RECT 25.19 67.05 25.4 67.12 ;
    RECT 21.41 66.33 21.62 66.4 ;
    RECT 21.41 66.69 21.62 66.76 ;
    RECT 21.41 67.05 21.62 67.12 ;
    RECT 21.87 66.33 22.08 66.4 ;
    RECT 21.87 66.69 22.08 66.76 ;
    RECT 21.87 67.05 22.08 67.12 ;
    RECT 18.09 66.33 18.3 66.4 ;
    RECT 18.09 66.69 18.3 66.76 ;
    RECT 18.09 67.05 18.3 67.12 ;
    RECT 18.55 66.33 18.76 66.4 ;
    RECT 18.55 66.69 18.76 66.76 ;
    RECT 18.55 67.05 18.76 67.12 ;
    RECT 120.825 66.69 120.895 66.76 ;
    RECT 14.77 66.33 14.98 66.4 ;
    RECT 14.77 66.69 14.98 66.76 ;
    RECT 14.77 67.05 14.98 67.12 ;
    RECT 15.23 66.33 15.44 66.4 ;
    RECT 15.23 66.69 15.44 66.76 ;
    RECT 15.23 67.05 15.44 67.12 ;
    RECT 11.45 66.33 11.66 66.4 ;
    RECT 11.45 66.69 11.66 66.76 ;
    RECT 11.45 67.05 11.66 67.12 ;
    RECT 11.91 66.33 12.12 66.4 ;
    RECT 11.91 66.69 12.12 66.76 ;
    RECT 11.91 67.05 12.12 67.12 ;
    RECT 8.13 66.33 8.34 66.4 ;
    RECT 8.13 66.69 8.34 66.76 ;
    RECT 8.13 67.05 8.34 67.12 ;
    RECT 8.59 66.33 8.8 66.4 ;
    RECT 8.59 66.69 8.8 66.76 ;
    RECT 8.59 67.05 8.8 67.12 ;
    RECT 4.81 66.33 5.02 66.4 ;
    RECT 4.81 66.69 5.02 66.76 ;
    RECT 4.81 67.05 5.02 67.12 ;
    RECT 5.27 66.33 5.48 66.4 ;
    RECT 5.27 66.69 5.48 66.76 ;
    RECT 5.27 67.05 5.48 67.12 ;
    RECT 1.49 66.33 1.7 66.4 ;
    RECT 1.49 66.69 1.7 66.76 ;
    RECT 1.49 67.05 1.7 67.12 ;
    RECT 1.95 66.33 2.16 66.4 ;
    RECT 1.95 66.69 2.16 66.76 ;
    RECT 1.95 67.05 2.16 67.12 ;
    RECT 64.57 66.33 64.78 66.4 ;
    RECT 64.57 66.69 64.78 66.76 ;
    RECT 64.57 67.05 64.78 67.12 ;
    RECT 65.03 66.33 65.24 66.4 ;
    RECT 65.03 66.69 65.24 66.76 ;
    RECT 65.03 67.05 65.24 67.12 ;
    RECT 61.25 65.61 61.46 65.68 ;
    RECT 61.25 65.97 61.46 66.04 ;
    RECT 61.25 66.33 61.46 66.4 ;
    RECT 61.71 65.61 61.92 65.68 ;
    RECT 61.71 65.97 61.92 66.04 ;
    RECT 61.71 66.33 61.92 66.4 ;
    RECT 57.93 65.61 58.14 65.68 ;
    RECT 57.93 65.97 58.14 66.04 ;
    RECT 57.93 66.33 58.14 66.4 ;
    RECT 58.39 65.61 58.6 65.68 ;
    RECT 58.39 65.97 58.6 66.04 ;
    RECT 58.39 66.33 58.6 66.4 ;
    RECT 54.61 65.61 54.82 65.68 ;
    RECT 54.61 65.97 54.82 66.04 ;
    RECT 54.61 66.33 54.82 66.4 ;
    RECT 55.07 65.61 55.28 65.68 ;
    RECT 55.07 65.97 55.28 66.04 ;
    RECT 55.07 66.33 55.28 66.4 ;
    RECT 51.29 65.61 51.5 65.68 ;
    RECT 51.29 65.97 51.5 66.04 ;
    RECT 51.29 66.33 51.5 66.4 ;
    RECT 51.75 65.61 51.96 65.68 ;
    RECT 51.75 65.97 51.96 66.04 ;
    RECT 51.75 66.33 51.96 66.4 ;
    RECT 47.97 65.61 48.18 65.68 ;
    RECT 47.97 65.97 48.18 66.04 ;
    RECT 47.97 66.33 48.18 66.4 ;
    RECT 48.43 65.61 48.64 65.68 ;
    RECT 48.43 65.97 48.64 66.04 ;
    RECT 48.43 66.33 48.64 66.4 ;
    RECT 44.65 65.61 44.86 65.68 ;
    RECT 44.65 65.97 44.86 66.04 ;
    RECT 44.65 66.33 44.86 66.4 ;
    RECT 45.11 65.61 45.32 65.68 ;
    RECT 45.11 65.97 45.32 66.04 ;
    RECT 45.11 66.33 45.32 66.4 ;
    RECT 41.33 65.61 41.54 65.68 ;
    RECT 41.33 65.97 41.54 66.04 ;
    RECT 41.33 66.33 41.54 66.4 ;
    RECT 41.79 65.61 42.0 65.68 ;
    RECT 41.79 65.97 42.0 66.04 ;
    RECT 41.79 66.33 42.0 66.4 ;
    RECT 38.01 65.61 38.22 65.68 ;
    RECT 38.01 65.97 38.22 66.04 ;
    RECT 38.01 66.33 38.22 66.4 ;
    RECT 38.47 65.61 38.68 65.68 ;
    RECT 38.47 65.97 38.68 66.04 ;
    RECT 38.47 66.33 38.68 66.4 ;
    RECT 0.4 65.97 0.47 66.04 ;
    RECT 34.69 65.61 34.9 65.68 ;
    RECT 34.69 65.97 34.9 66.04 ;
    RECT 34.69 66.33 34.9 66.4 ;
    RECT 35.15 65.61 35.36 65.68 ;
    RECT 35.15 65.97 35.36 66.04 ;
    RECT 35.15 66.33 35.36 66.4 ;
    RECT 117.69 65.61 117.9 65.68 ;
    RECT 117.69 65.97 117.9 66.04 ;
    RECT 117.69 66.33 117.9 66.4 ;
    RECT 118.15 65.61 118.36 65.68 ;
    RECT 118.15 65.97 118.36 66.04 ;
    RECT 118.15 66.33 118.36 66.4 ;
    RECT 114.37 65.61 114.58 65.68 ;
    RECT 114.37 65.97 114.58 66.04 ;
    RECT 114.37 66.33 114.58 66.4 ;
    RECT 114.83 65.61 115.04 65.68 ;
    RECT 114.83 65.97 115.04 66.04 ;
    RECT 114.83 66.33 115.04 66.4 ;
    RECT 111.05 65.61 111.26 65.68 ;
    RECT 111.05 65.97 111.26 66.04 ;
    RECT 111.05 66.33 111.26 66.4 ;
    RECT 111.51 65.61 111.72 65.68 ;
    RECT 111.51 65.97 111.72 66.04 ;
    RECT 111.51 66.33 111.72 66.4 ;
    RECT 107.73 65.61 107.94 65.68 ;
    RECT 107.73 65.97 107.94 66.04 ;
    RECT 107.73 66.33 107.94 66.4 ;
    RECT 108.19 65.61 108.4 65.68 ;
    RECT 108.19 65.97 108.4 66.04 ;
    RECT 108.19 66.33 108.4 66.4 ;
    RECT 104.41 65.61 104.62 65.68 ;
    RECT 104.41 65.97 104.62 66.04 ;
    RECT 104.41 66.33 104.62 66.4 ;
    RECT 104.87 65.61 105.08 65.68 ;
    RECT 104.87 65.97 105.08 66.04 ;
    RECT 104.87 66.33 105.08 66.4 ;
    RECT 101.09 65.61 101.3 65.68 ;
    RECT 101.09 65.97 101.3 66.04 ;
    RECT 101.09 66.33 101.3 66.4 ;
    RECT 101.55 65.61 101.76 65.68 ;
    RECT 101.55 65.97 101.76 66.04 ;
    RECT 101.55 66.33 101.76 66.4 ;
    RECT 97.77 65.61 97.98 65.68 ;
    RECT 97.77 65.97 97.98 66.04 ;
    RECT 97.77 66.33 97.98 66.4 ;
    RECT 98.23 65.61 98.44 65.68 ;
    RECT 98.23 65.97 98.44 66.04 ;
    RECT 98.23 66.33 98.44 66.4 ;
    RECT 94.45 65.61 94.66 65.68 ;
    RECT 94.45 65.97 94.66 66.04 ;
    RECT 94.45 66.33 94.66 66.4 ;
    RECT 94.91 65.61 95.12 65.68 ;
    RECT 94.91 65.97 95.12 66.04 ;
    RECT 94.91 66.33 95.12 66.4 ;
    RECT 91.13 65.61 91.34 65.68 ;
    RECT 91.13 65.97 91.34 66.04 ;
    RECT 91.13 66.33 91.34 66.4 ;
    RECT 91.59 65.61 91.8 65.68 ;
    RECT 91.59 65.97 91.8 66.04 ;
    RECT 91.59 66.33 91.8 66.4 ;
    RECT 87.81 65.61 88.02 65.68 ;
    RECT 87.81 65.97 88.02 66.04 ;
    RECT 87.81 66.33 88.02 66.4 ;
    RECT 88.27 65.61 88.48 65.68 ;
    RECT 88.27 65.97 88.48 66.04 ;
    RECT 88.27 66.33 88.48 66.4 ;
    RECT 84.49 65.61 84.7 65.68 ;
    RECT 84.49 65.97 84.7 66.04 ;
    RECT 84.49 66.33 84.7 66.4 ;
    RECT 84.95 65.61 85.16 65.68 ;
    RECT 84.95 65.97 85.16 66.04 ;
    RECT 84.95 66.33 85.16 66.4 ;
    RECT 81.17 65.61 81.38 65.68 ;
    RECT 81.17 65.97 81.38 66.04 ;
    RECT 81.17 66.33 81.38 66.4 ;
    RECT 81.63 65.61 81.84 65.68 ;
    RECT 81.63 65.97 81.84 66.04 ;
    RECT 81.63 66.33 81.84 66.4 ;
    RECT 77.85 65.61 78.06 65.68 ;
    RECT 77.85 65.97 78.06 66.04 ;
    RECT 77.85 66.33 78.06 66.4 ;
    RECT 78.31 65.61 78.52 65.68 ;
    RECT 78.31 65.97 78.52 66.04 ;
    RECT 78.31 66.33 78.52 66.4 ;
    RECT 74.53 65.61 74.74 65.68 ;
    RECT 74.53 65.97 74.74 66.04 ;
    RECT 74.53 66.33 74.74 66.4 ;
    RECT 74.99 65.61 75.2 65.68 ;
    RECT 74.99 65.97 75.2 66.04 ;
    RECT 74.99 66.33 75.2 66.4 ;
    RECT 71.21 65.61 71.42 65.68 ;
    RECT 71.21 65.97 71.42 66.04 ;
    RECT 71.21 66.33 71.42 66.4 ;
    RECT 71.67 65.61 71.88 65.68 ;
    RECT 71.67 65.97 71.88 66.04 ;
    RECT 71.67 66.33 71.88 66.4 ;
    RECT 31.37 65.61 31.58 65.68 ;
    RECT 31.37 65.97 31.58 66.04 ;
    RECT 31.37 66.33 31.58 66.4 ;
    RECT 31.83 65.61 32.04 65.68 ;
    RECT 31.83 65.97 32.04 66.04 ;
    RECT 31.83 66.33 32.04 66.4 ;
    RECT 67.89 65.61 68.1 65.68 ;
    RECT 67.89 65.97 68.1 66.04 ;
    RECT 67.89 66.33 68.1 66.4 ;
    RECT 68.35 65.61 68.56 65.68 ;
    RECT 68.35 65.97 68.56 66.04 ;
    RECT 68.35 66.33 68.56 66.4 ;
    RECT 28.05 65.61 28.26 65.68 ;
    RECT 28.05 65.97 28.26 66.04 ;
    RECT 28.05 66.33 28.26 66.4 ;
    RECT 28.51 65.61 28.72 65.68 ;
    RECT 28.51 65.97 28.72 66.04 ;
    RECT 28.51 66.33 28.72 66.4 ;
    RECT 24.73 65.61 24.94 65.68 ;
    RECT 24.73 65.97 24.94 66.04 ;
    RECT 24.73 66.33 24.94 66.4 ;
    RECT 25.19 65.61 25.4 65.68 ;
    RECT 25.19 65.97 25.4 66.04 ;
    RECT 25.19 66.33 25.4 66.4 ;
    RECT 21.41 65.61 21.62 65.68 ;
    RECT 21.41 65.97 21.62 66.04 ;
    RECT 21.41 66.33 21.62 66.4 ;
    RECT 21.87 65.61 22.08 65.68 ;
    RECT 21.87 65.97 22.08 66.04 ;
    RECT 21.87 66.33 22.08 66.4 ;
    RECT 18.09 65.61 18.3 65.68 ;
    RECT 18.09 65.97 18.3 66.04 ;
    RECT 18.09 66.33 18.3 66.4 ;
    RECT 18.55 65.61 18.76 65.68 ;
    RECT 18.55 65.97 18.76 66.04 ;
    RECT 18.55 66.33 18.76 66.4 ;
    RECT 120.825 65.97 120.895 66.04 ;
    RECT 14.77 65.61 14.98 65.68 ;
    RECT 14.77 65.97 14.98 66.04 ;
    RECT 14.77 66.33 14.98 66.4 ;
    RECT 15.23 65.61 15.44 65.68 ;
    RECT 15.23 65.97 15.44 66.04 ;
    RECT 15.23 66.33 15.44 66.4 ;
    RECT 11.45 65.61 11.66 65.68 ;
    RECT 11.45 65.97 11.66 66.04 ;
    RECT 11.45 66.33 11.66 66.4 ;
    RECT 11.91 65.61 12.12 65.68 ;
    RECT 11.91 65.97 12.12 66.04 ;
    RECT 11.91 66.33 12.12 66.4 ;
    RECT 8.13 65.61 8.34 65.68 ;
    RECT 8.13 65.97 8.34 66.04 ;
    RECT 8.13 66.33 8.34 66.4 ;
    RECT 8.59 65.61 8.8 65.68 ;
    RECT 8.59 65.97 8.8 66.04 ;
    RECT 8.59 66.33 8.8 66.4 ;
    RECT 4.81 65.61 5.02 65.68 ;
    RECT 4.81 65.97 5.02 66.04 ;
    RECT 4.81 66.33 5.02 66.4 ;
    RECT 5.27 65.61 5.48 65.68 ;
    RECT 5.27 65.97 5.48 66.04 ;
    RECT 5.27 66.33 5.48 66.4 ;
    RECT 1.49 65.61 1.7 65.68 ;
    RECT 1.49 65.97 1.7 66.04 ;
    RECT 1.49 66.33 1.7 66.4 ;
    RECT 1.95 65.61 2.16 65.68 ;
    RECT 1.95 65.97 2.16 66.04 ;
    RECT 1.95 66.33 2.16 66.4 ;
    RECT 64.57 65.61 64.78 65.68 ;
    RECT 64.57 65.97 64.78 66.04 ;
    RECT 64.57 66.33 64.78 66.4 ;
    RECT 65.03 65.61 65.24 65.68 ;
    RECT 65.03 65.97 65.24 66.04 ;
    RECT 65.03 66.33 65.24 66.4 ;
    RECT 61.25 28.15 61.46 28.22 ;
    RECT 61.25 28.51 61.46 28.58 ;
    RECT 61.25 28.87 61.46 28.94 ;
    RECT 61.71 28.15 61.92 28.22 ;
    RECT 61.71 28.51 61.92 28.58 ;
    RECT 61.71 28.87 61.92 28.94 ;
    RECT 57.93 28.15 58.14 28.22 ;
    RECT 57.93 28.51 58.14 28.58 ;
    RECT 57.93 28.87 58.14 28.94 ;
    RECT 58.39 28.15 58.6 28.22 ;
    RECT 58.39 28.51 58.6 28.58 ;
    RECT 58.39 28.87 58.6 28.94 ;
    RECT 54.61 28.15 54.82 28.22 ;
    RECT 54.61 28.51 54.82 28.58 ;
    RECT 54.61 28.87 54.82 28.94 ;
    RECT 55.07 28.15 55.28 28.22 ;
    RECT 55.07 28.51 55.28 28.58 ;
    RECT 55.07 28.87 55.28 28.94 ;
    RECT 51.29 28.15 51.5 28.22 ;
    RECT 51.29 28.51 51.5 28.58 ;
    RECT 51.29 28.87 51.5 28.94 ;
    RECT 51.75 28.15 51.96 28.22 ;
    RECT 51.75 28.51 51.96 28.58 ;
    RECT 51.75 28.87 51.96 28.94 ;
    RECT 47.97 28.15 48.18 28.22 ;
    RECT 47.97 28.51 48.18 28.58 ;
    RECT 47.97 28.87 48.18 28.94 ;
    RECT 48.43 28.15 48.64 28.22 ;
    RECT 48.43 28.51 48.64 28.58 ;
    RECT 48.43 28.87 48.64 28.94 ;
    RECT 44.65 28.15 44.86 28.22 ;
    RECT 44.65 28.51 44.86 28.58 ;
    RECT 44.65 28.87 44.86 28.94 ;
    RECT 45.11 28.15 45.32 28.22 ;
    RECT 45.11 28.51 45.32 28.58 ;
    RECT 45.11 28.87 45.32 28.94 ;
    RECT 41.33 28.15 41.54 28.22 ;
    RECT 41.33 28.51 41.54 28.58 ;
    RECT 41.33 28.87 41.54 28.94 ;
    RECT 41.79 28.15 42.0 28.22 ;
    RECT 41.79 28.51 42.0 28.58 ;
    RECT 41.79 28.87 42.0 28.94 ;
    RECT 38.01 28.15 38.22 28.22 ;
    RECT 38.01 28.51 38.22 28.58 ;
    RECT 38.01 28.87 38.22 28.94 ;
    RECT 38.47 28.15 38.68 28.22 ;
    RECT 38.47 28.51 38.68 28.58 ;
    RECT 38.47 28.87 38.68 28.94 ;
    RECT 0.4 28.51 0.47 28.58 ;
    RECT 34.69 28.15 34.9 28.22 ;
    RECT 34.69 28.51 34.9 28.58 ;
    RECT 34.69 28.87 34.9 28.94 ;
    RECT 35.15 28.15 35.36 28.22 ;
    RECT 35.15 28.51 35.36 28.58 ;
    RECT 35.15 28.87 35.36 28.94 ;
    RECT 117.69 28.15 117.9 28.22 ;
    RECT 117.69 28.51 117.9 28.58 ;
    RECT 117.69 28.87 117.9 28.94 ;
    RECT 118.15 28.15 118.36 28.22 ;
    RECT 118.15 28.51 118.36 28.58 ;
    RECT 118.15 28.87 118.36 28.94 ;
    RECT 114.37 28.15 114.58 28.22 ;
    RECT 114.37 28.51 114.58 28.58 ;
    RECT 114.37 28.87 114.58 28.94 ;
    RECT 114.83 28.15 115.04 28.22 ;
    RECT 114.83 28.51 115.04 28.58 ;
    RECT 114.83 28.87 115.04 28.94 ;
    RECT 111.05 28.15 111.26 28.22 ;
    RECT 111.05 28.51 111.26 28.58 ;
    RECT 111.05 28.87 111.26 28.94 ;
    RECT 111.51 28.15 111.72 28.22 ;
    RECT 111.51 28.51 111.72 28.58 ;
    RECT 111.51 28.87 111.72 28.94 ;
    RECT 107.73 28.15 107.94 28.22 ;
    RECT 107.73 28.51 107.94 28.58 ;
    RECT 107.73 28.87 107.94 28.94 ;
    RECT 108.19 28.15 108.4 28.22 ;
    RECT 108.19 28.51 108.4 28.58 ;
    RECT 108.19 28.87 108.4 28.94 ;
    RECT 104.41 28.15 104.62 28.22 ;
    RECT 104.41 28.51 104.62 28.58 ;
    RECT 104.41 28.87 104.62 28.94 ;
    RECT 104.87 28.15 105.08 28.22 ;
    RECT 104.87 28.51 105.08 28.58 ;
    RECT 104.87 28.87 105.08 28.94 ;
    RECT 101.09 28.15 101.3 28.22 ;
    RECT 101.09 28.51 101.3 28.58 ;
    RECT 101.09 28.87 101.3 28.94 ;
    RECT 101.55 28.15 101.76 28.22 ;
    RECT 101.55 28.51 101.76 28.58 ;
    RECT 101.55 28.87 101.76 28.94 ;
    RECT 97.77 28.15 97.98 28.22 ;
    RECT 97.77 28.51 97.98 28.58 ;
    RECT 97.77 28.87 97.98 28.94 ;
    RECT 98.23 28.15 98.44 28.22 ;
    RECT 98.23 28.51 98.44 28.58 ;
    RECT 98.23 28.87 98.44 28.94 ;
    RECT 94.45 28.15 94.66 28.22 ;
    RECT 94.45 28.51 94.66 28.58 ;
    RECT 94.45 28.87 94.66 28.94 ;
    RECT 94.91 28.15 95.12 28.22 ;
    RECT 94.91 28.51 95.12 28.58 ;
    RECT 94.91 28.87 95.12 28.94 ;
    RECT 91.13 28.15 91.34 28.22 ;
    RECT 91.13 28.51 91.34 28.58 ;
    RECT 91.13 28.87 91.34 28.94 ;
    RECT 91.59 28.15 91.8 28.22 ;
    RECT 91.59 28.51 91.8 28.58 ;
    RECT 91.59 28.87 91.8 28.94 ;
    RECT 87.81 28.15 88.02 28.22 ;
    RECT 87.81 28.51 88.02 28.58 ;
    RECT 87.81 28.87 88.02 28.94 ;
    RECT 88.27 28.15 88.48 28.22 ;
    RECT 88.27 28.51 88.48 28.58 ;
    RECT 88.27 28.87 88.48 28.94 ;
    RECT 84.49 28.15 84.7 28.22 ;
    RECT 84.49 28.51 84.7 28.58 ;
    RECT 84.49 28.87 84.7 28.94 ;
    RECT 84.95 28.15 85.16 28.22 ;
    RECT 84.95 28.51 85.16 28.58 ;
    RECT 84.95 28.87 85.16 28.94 ;
    RECT 81.17 28.15 81.38 28.22 ;
    RECT 81.17 28.51 81.38 28.58 ;
    RECT 81.17 28.87 81.38 28.94 ;
    RECT 81.63 28.15 81.84 28.22 ;
    RECT 81.63 28.51 81.84 28.58 ;
    RECT 81.63 28.87 81.84 28.94 ;
    RECT 77.85 28.15 78.06 28.22 ;
    RECT 77.85 28.51 78.06 28.58 ;
    RECT 77.85 28.87 78.06 28.94 ;
    RECT 78.31 28.15 78.52 28.22 ;
    RECT 78.31 28.51 78.52 28.58 ;
    RECT 78.31 28.87 78.52 28.94 ;
    RECT 74.53 28.15 74.74 28.22 ;
    RECT 74.53 28.51 74.74 28.58 ;
    RECT 74.53 28.87 74.74 28.94 ;
    RECT 74.99 28.15 75.2 28.22 ;
    RECT 74.99 28.51 75.2 28.58 ;
    RECT 74.99 28.87 75.2 28.94 ;
    RECT 71.21 28.15 71.42 28.22 ;
    RECT 71.21 28.51 71.42 28.58 ;
    RECT 71.21 28.87 71.42 28.94 ;
    RECT 71.67 28.15 71.88 28.22 ;
    RECT 71.67 28.51 71.88 28.58 ;
    RECT 71.67 28.87 71.88 28.94 ;
    RECT 31.37 28.15 31.58 28.22 ;
    RECT 31.37 28.51 31.58 28.58 ;
    RECT 31.37 28.87 31.58 28.94 ;
    RECT 31.83 28.15 32.04 28.22 ;
    RECT 31.83 28.51 32.04 28.58 ;
    RECT 31.83 28.87 32.04 28.94 ;
    RECT 67.89 28.15 68.1 28.22 ;
    RECT 67.89 28.51 68.1 28.58 ;
    RECT 67.89 28.87 68.1 28.94 ;
    RECT 68.35 28.15 68.56 28.22 ;
    RECT 68.35 28.51 68.56 28.58 ;
    RECT 68.35 28.87 68.56 28.94 ;
    RECT 28.05 28.15 28.26 28.22 ;
    RECT 28.05 28.51 28.26 28.58 ;
    RECT 28.05 28.87 28.26 28.94 ;
    RECT 28.51 28.15 28.72 28.22 ;
    RECT 28.51 28.51 28.72 28.58 ;
    RECT 28.51 28.87 28.72 28.94 ;
    RECT 24.73 28.15 24.94 28.22 ;
    RECT 24.73 28.51 24.94 28.58 ;
    RECT 24.73 28.87 24.94 28.94 ;
    RECT 25.19 28.15 25.4 28.22 ;
    RECT 25.19 28.51 25.4 28.58 ;
    RECT 25.19 28.87 25.4 28.94 ;
    RECT 21.41 28.15 21.62 28.22 ;
    RECT 21.41 28.51 21.62 28.58 ;
    RECT 21.41 28.87 21.62 28.94 ;
    RECT 21.87 28.15 22.08 28.22 ;
    RECT 21.87 28.51 22.08 28.58 ;
    RECT 21.87 28.87 22.08 28.94 ;
    RECT 18.09 28.15 18.3 28.22 ;
    RECT 18.09 28.51 18.3 28.58 ;
    RECT 18.09 28.87 18.3 28.94 ;
    RECT 18.55 28.15 18.76 28.22 ;
    RECT 18.55 28.51 18.76 28.58 ;
    RECT 18.55 28.87 18.76 28.94 ;
    RECT 120.825 28.51 120.895 28.58 ;
    RECT 14.77 28.15 14.98 28.22 ;
    RECT 14.77 28.51 14.98 28.58 ;
    RECT 14.77 28.87 14.98 28.94 ;
    RECT 15.23 28.15 15.44 28.22 ;
    RECT 15.23 28.51 15.44 28.58 ;
    RECT 15.23 28.87 15.44 28.94 ;
    RECT 11.45 28.15 11.66 28.22 ;
    RECT 11.45 28.51 11.66 28.58 ;
    RECT 11.45 28.87 11.66 28.94 ;
    RECT 11.91 28.15 12.12 28.22 ;
    RECT 11.91 28.51 12.12 28.58 ;
    RECT 11.91 28.87 12.12 28.94 ;
    RECT 8.13 28.15 8.34 28.22 ;
    RECT 8.13 28.51 8.34 28.58 ;
    RECT 8.13 28.87 8.34 28.94 ;
    RECT 8.59 28.15 8.8 28.22 ;
    RECT 8.59 28.51 8.8 28.58 ;
    RECT 8.59 28.87 8.8 28.94 ;
    RECT 4.81 28.15 5.02 28.22 ;
    RECT 4.81 28.51 5.02 28.58 ;
    RECT 4.81 28.87 5.02 28.94 ;
    RECT 5.27 28.15 5.48 28.22 ;
    RECT 5.27 28.51 5.48 28.58 ;
    RECT 5.27 28.87 5.48 28.94 ;
    RECT 1.49 28.15 1.7 28.22 ;
    RECT 1.49 28.51 1.7 28.58 ;
    RECT 1.49 28.87 1.7 28.94 ;
    RECT 1.95 28.15 2.16 28.22 ;
    RECT 1.95 28.51 2.16 28.58 ;
    RECT 1.95 28.87 2.16 28.94 ;
    RECT 64.57 28.15 64.78 28.22 ;
    RECT 64.57 28.51 64.78 28.58 ;
    RECT 64.57 28.87 64.78 28.94 ;
    RECT 65.03 28.15 65.24 28.22 ;
    RECT 65.03 28.51 65.24 28.58 ;
    RECT 65.03 28.87 65.24 28.94 ;
    RECT 61.25 27.43 61.46 27.5 ;
    RECT 61.25 27.79 61.46 27.86 ;
    RECT 61.25 28.15 61.46 28.22 ;
    RECT 61.71 27.43 61.92 27.5 ;
    RECT 61.71 27.79 61.92 27.86 ;
    RECT 61.71 28.15 61.92 28.22 ;
    RECT 57.93 27.43 58.14 27.5 ;
    RECT 57.93 27.79 58.14 27.86 ;
    RECT 57.93 28.15 58.14 28.22 ;
    RECT 58.39 27.43 58.6 27.5 ;
    RECT 58.39 27.79 58.6 27.86 ;
    RECT 58.39 28.15 58.6 28.22 ;
    RECT 54.61 27.43 54.82 27.5 ;
    RECT 54.61 27.79 54.82 27.86 ;
    RECT 54.61 28.15 54.82 28.22 ;
    RECT 55.07 27.43 55.28 27.5 ;
    RECT 55.07 27.79 55.28 27.86 ;
    RECT 55.07 28.15 55.28 28.22 ;
    RECT 51.29 27.43 51.5 27.5 ;
    RECT 51.29 27.79 51.5 27.86 ;
    RECT 51.29 28.15 51.5 28.22 ;
    RECT 51.75 27.43 51.96 27.5 ;
    RECT 51.75 27.79 51.96 27.86 ;
    RECT 51.75 28.15 51.96 28.22 ;
    RECT 47.97 27.43 48.18 27.5 ;
    RECT 47.97 27.79 48.18 27.86 ;
    RECT 47.97 28.15 48.18 28.22 ;
    RECT 48.43 27.43 48.64 27.5 ;
    RECT 48.43 27.79 48.64 27.86 ;
    RECT 48.43 28.15 48.64 28.22 ;
    RECT 44.65 27.43 44.86 27.5 ;
    RECT 44.65 27.79 44.86 27.86 ;
    RECT 44.65 28.15 44.86 28.22 ;
    RECT 45.11 27.43 45.32 27.5 ;
    RECT 45.11 27.79 45.32 27.86 ;
    RECT 45.11 28.15 45.32 28.22 ;
    RECT 41.33 27.43 41.54 27.5 ;
    RECT 41.33 27.79 41.54 27.86 ;
    RECT 41.33 28.15 41.54 28.22 ;
    RECT 41.79 27.43 42.0 27.5 ;
    RECT 41.79 27.79 42.0 27.86 ;
    RECT 41.79 28.15 42.0 28.22 ;
    RECT 38.01 27.43 38.22 27.5 ;
    RECT 38.01 27.79 38.22 27.86 ;
    RECT 38.01 28.15 38.22 28.22 ;
    RECT 38.47 27.43 38.68 27.5 ;
    RECT 38.47 27.79 38.68 27.86 ;
    RECT 38.47 28.15 38.68 28.22 ;
    RECT 0.4 27.79 0.47 27.86 ;
    RECT 34.69 27.43 34.9 27.5 ;
    RECT 34.69 27.79 34.9 27.86 ;
    RECT 34.69 28.15 34.9 28.22 ;
    RECT 35.15 27.43 35.36 27.5 ;
    RECT 35.15 27.79 35.36 27.86 ;
    RECT 35.15 28.15 35.36 28.22 ;
    RECT 117.69 27.43 117.9 27.5 ;
    RECT 117.69 27.79 117.9 27.86 ;
    RECT 117.69 28.15 117.9 28.22 ;
    RECT 118.15 27.43 118.36 27.5 ;
    RECT 118.15 27.79 118.36 27.86 ;
    RECT 118.15 28.15 118.36 28.22 ;
    RECT 114.37 27.43 114.58 27.5 ;
    RECT 114.37 27.79 114.58 27.86 ;
    RECT 114.37 28.15 114.58 28.22 ;
    RECT 114.83 27.43 115.04 27.5 ;
    RECT 114.83 27.79 115.04 27.86 ;
    RECT 114.83 28.15 115.04 28.22 ;
    RECT 111.05 27.43 111.26 27.5 ;
    RECT 111.05 27.79 111.26 27.86 ;
    RECT 111.05 28.15 111.26 28.22 ;
    RECT 111.51 27.43 111.72 27.5 ;
    RECT 111.51 27.79 111.72 27.86 ;
    RECT 111.51 28.15 111.72 28.22 ;
    RECT 107.73 27.43 107.94 27.5 ;
    RECT 107.73 27.79 107.94 27.86 ;
    RECT 107.73 28.15 107.94 28.22 ;
    RECT 108.19 27.43 108.4 27.5 ;
    RECT 108.19 27.79 108.4 27.86 ;
    RECT 108.19 28.15 108.4 28.22 ;
    RECT 104.41 27.43 104.62 27.5 ;
    RECT 104.41 27.79 104.62 27.86 ;
    RECT 104.41 28.15 104.62 28.22 ;
    RECT 104.87 27.43 105.08 27.5 ;
    RECT 104.87 27.79 105.08 27.86 ;
    RECT 104.87 28.15 105.08 28.22 ;
    RECT 101.09 27.43 101.3 27.5 ;
    RECT 101.09 27.79 101.3 27.86 ;
    RECT 101.09 28.15 101.3 28.22 ;
    RECT 101.55 27.43 101.76 27.5 ;
    RECT 101.55 27.79 101.76 27.86 ;
    RECT 101.55 28.15 101.76 28.22 ;
    RECT 97.77 27.43 97.98 27.5 ;
    RECT 97.77 27.79 97.98 27.86 ;
    RECT 97.77 28.15 97.98 28.22 ;
    RECT 98.23 27.43 98.44 27.5 ;
    RECT 98.23 27.79 98.44 27.86 ;
    RECT 98.23 28.15 98.44 28.22 ;
    RECT 94.45 27.43 94.66 27.5 ;
    RECT 94.45 27.79 94.66 27.86 ;
    RECT 94.45 28.15 94.66 28.22 ;
    RECT 94.91 27.43 95.12 27.5 ;
    RECT 94.91 27.79 95.12 27.86 ;
    RECT 94.91 28.15 95.12 28.22 ;
    RECT 91.13 27.43 91.34 27.5 ;
    RECT 91.13 27.79 91.34 27.86 ;
    RECT 91.13 28.15 91.34 28.22 ;
    RECT 91.59 27.43 91.8 27.5 ;
    RECT 91.59 27.79 91.8 27.86 ;
    RECT 91.59 28.15 91.8 28.22 ;
    RECT 87.81 27.43 88.02 27.5 ;
    RECT 87.81 27.79 88.02 27.86 ;
    RECT 87.81 28.15 88.02 28.22 ;
    RECT 88.27 27.43 88.48 27.5 ;
    RECT 88.27 27.79 88.48 27.86 ;
    RECT 88.27 28.15 88.48 28.22 ;
    RECT 84.49 27.43 84.7 27.5 ;
    RECT 84.49 27.79 84.7 27.86 ;
    RECT 84.49 28.15 84.7 28.22 ;
    RECT 84.95 27.43 85.16 27.5 ;
    RECT 84.95 27.79 85.16 27.86 ;
    RECT 84.95 28.15 85.16 28.22 ;
    RECT 81.17 27.43 81.38 27.5 ;
    RECT 81.17 27.79 81.38 27.86 ;
    RECT 81.17 28.15 81.38 28.22 ;
    RECT 81.63 27.43 81.84 27.5 ;
    RECT 81.63 27.79 81.84 27.86 ;
    RECT 81.63 28.15 81.84 28.22 ;
    RECT 77.85 27.43 78.06 27.5 ;
    RECT 77.85 27.79 78.06 27.86 ;
    RECT 77.85 28.15 78.06 28.22 ;
    RECT 78.31 27.43 78.52 27.5 ;
    RECT 78.31 27.79 78.52 27.86 ;
    RECT 78.31 28.15 78.52 28.22 ;
    RECT 74.53 27.43 74.74 27.5 ;
    RECT 74.53 27.79 74.74 27.86 ;
    RECT 74.53 28.15 74.74 28.22 ;
    RECT 74.99 27.43 75.2 27.5 ;
    RECT 74.99 27.79 75.2 27.86 ;
    RECT 74.99 28.15 75.2 28.22 ;
    RECT 71.21 27.43 71.42 27.5 ;
    RECT 71.21 27.79 71.42 27.86 ;
    RECT 71.21 28.15 71.42 28.22 ;
    RECT 71.67 27.43 71.88 27.5 ;
    RECT 71.67 27.79 71.88 27.86 ;
    RECT 71.67 28.15 71.88 28.22 ;
    RECT 31.37 27.43 31.58 27.5 ;
    RECT 31.37 27.79 31.58 27.86 ;
    RECT 31.37 28.15 31.58 28.22 ;
    RECT 31.83 27.43 32.04 27.5 ;
    RECT 31.83 27.79 32.04 27.86 ;
    RECT 31.83 28.15 32.04 28.22 ;
    RECT 67.89 27.43 68.1 27.5 ;
    RECT 67.89 27.79 68.1 27.86 ;
    RECT 67.89 28.15 68.1 28.22 ;
    RECT 68.35 27.43 68.56 27.5 ;
    RECT 68.35 27.79 68.56 27.86 ;
    RECT 68.35 28.15 68.56 28.22 ;
    RECT 28.05 27.43 28.26 27.5 ;
    RECT 28.05 27.79 28.26 27.86 ;
    RECT 28.05 28.15 28.26 28.22 ;
    RECT 28.51 27.43 28.72 27.5 ;
    RECT 28.51 27.79 28.72 27.86 ;
    RECT 28.51 28.15 28.72 28.22 ;
    RECT 24.73 27.43 24.94 27.5 ;
    RECT 24.73 27.79 24.94 27.86 ;
    RECT 24.73 28.15 24.94 28.22 ;
    RECT 25.19 27.43 25.4 27.5 ;
    RECT 25.19 27.79 25.4 27.86 ;
    RECT 25.19 28.15 25.4 28.22 ;
    RECT 21.41 27.43 21.62 27.5 ;
    RECT 21.41 27.79 21.62 27.86 ;
    RECT 21.41 28.15 21.62 28.22 ;
    RECT 21.87 27.43 22.08 27.5 ;
    RECT 21.87 27.79 22.08 27.86 ;
    RECT 21.87 28.15 22.08 28.22 ;
    RECT 18.09 27.43 18.3 27.5 ;
    RECT 18.09 27.79 18.3 27.86 ;
    RECT 18.09 28.15 18.3 28.22 ;
    RECT 18.55 27.43 18.76 27.5 ;
    RECT 18.55 27.79 18.76 27.86 ;
    RECT 18.55 28.15 18.76 28.22 ;
    RECT 120.825 27.79 120.895 27.86 ;
    RECT 14.77 27.43 14.98 27.5 ;
    RECT 14.77 27.79 14.98 27.86 ;
    RECT 14.77 28.15 14.98 28.22 ;
    RECT 15.23 27.43 15.44 27.5 ;
    RECT 15.23 27.79 15.44 27.86 ;
    RECT 15.23 28.15 15.44 28.22 ;
    RECT 11.45 27.43 11.66 27.5 ;
    RECT 11.45 27.79 11.66 27.86 ;
    RECT 11.45 28.15 11.66 28.22 ;
    RECT 11.91 27.43 12.12 27.5 ;
    RECT 11.91 27.79 12.12 27.86 ;
    RECT 11.91 28.15 12.12 28.22 ;
    RECT 8.13 27.43 8.34 27.5 ;
    RECT 8.13 27.79 8.34 27.86 ;
    RECT 8.13 28.15 8.34 28.22 ;
    RECT 8.59 27.43 8.8 27.5 ;
    RECT 8.59 27.79 8.8 27.86 ;
    RECT 8.59 28.15 8.8 28.22 ;
    RECT 4.81 27.43 5.02 27.5 ;
    RECT 4.81 27.79 5.02 27.86 ;
    RECT 4.81 28.15 5.02 28.22 ;
    RECT 5.27 27.43 5.48 27.5 ;
    RECT 5.27 27.79 5.48 27.86 ;
    RECT 5.27 28.15 5.48 28.22 ;
    RECT 1.49 27.43 1.7 27.5 ;
    RECT 1.49 27.79 1.7 27.86 ;
    RECT 1.49 28.15 1.7 28.22 ;
    RECT 1.95 27.43 2.16 27.5 ;
    RECT 1.95 27.79 2.16 27.86 ;
    RECT 1.95 28.15 2.16 28.22 ;
    RECT 64.57 27.43 64.78 27.5 ;
    RECT 64.57 27.79 64.78 27.86 ;
    RECT 64.57 28.15 64.78 28.22 ;
    RECT 65.03 27.43 65.24 27.5 ;
    RECT 65.03 27.79 65.24 27.86 ;
    RECT 65.03 28.15 65.24 28.22 ;
    RECT 61.25 26.71 61.46 26.78 ;
    RECT 61.25 27.07 61.46 27.14 ;
    RECT 61.25 27.43 61.46 27.5 ;
    RECT 61.71 26.71 61.92 26.78 ;
    RECT 61.71 27.07 61.92 27.14 ;
    RECT 61.71 27.43 61.92 27.5 ;
    RECT 57.93 26.71 58.14 26.78 ;
    RECT 57.93 27.07 58.14 27.14 ;
    RECT 57.93 27.43 58.14 27.5 ;
    RECT 58.39 26.71 58.6 26.78 ;
    RECT 58.39 27.07 58.6 27.14 ;
    RECT 58.39 27.43 58.6 27.5 ;
    RECT 54.61 26.71 54.82 26.78 ;
    RECT 54.61 27.07 54.82 27.14 ;
    RECT 54.61 27.43 54.82 27.5 ;
    RECT 55.07 26.71 55.28 26.78 ;
    RECT 55.07 27.07 55.28 27.14 ;
    RECT 55.07 27.43 55.28 27.5 ;
    RECT 51.29 26.71 51.5 26.78 ;
    RECT 51.29 27.07 51.5 27.14 ;
    RECT 51.29 27.43 51.5 27.5 ;
    RECT 51.75 26.71 51.96 26.78 ;
    RECT 51.75 27.07 51.96 27.14 ;
    RECT 51.75 27.43 51.96 27.5 ;
    RECT 47.97 26.71 48.18 26.78 ;
    RECT 47.97 27.07 48.18 27.14 ;
    RECT 47.97 27.43 48.18 27.5 ;
    RECT 48.43 26.71 48.64 26.78 ;
    RECT 48.43 27.07 48.64 27.14 ;
    RECT 48.43 27.43 48.64 27.5 ;
    RECT 44.65 26.71 44.86 26.78 ;
    RECT 44.65 27.07 44.86 27.14 ;
    RECT 44.65 27.43 44.86 27.5 ;
    RECT 45.11 26.71 45.32 26.78 ;
    RECT 45.11 27.07 45.32 27.14 ;
    RECT 45.11 27.43 45.32 27.5 ;
    RECT 41.33 26.71 41.54 26.78 ;
    RECT 41.33 27.07 41.54 27.14 ;
    RECT 41.33 27.43 41.54 27.5 ;
    RECT 41.79 26.71 42.0 26.78 ;
    RECT 41.79 27.07 42.0 27.14 ;
    RECT 41.79 27.43 42.0 27.5 ;
    RECT 38.01 26.71 38.22 26.78 ;
    RECT 38.01 27.07 38.22 27.14 ;
    RECT 38.01 27.43 38.22 27.5 ;
    RECT 38.47 26.71 38.68 26.78 ;
    RECT 38.47 27.07 38.68 27.14 ;
    RECT 38.47 27.43 38.68 27.5 ;
    RECT 0.4 27.07 0.47 27.14 ;
    RECT 34.69 26.71 34.9 26.78 ;
    RECT 34.69 27.07 34.9 27.14 ;
    RECT 34.69 27.43 34.9 27.5 ;
    RECT 35.15 26.71 35.36 26.78 ;
    RECT 35.15 27.07 35.36 27.14 ;
    RECT 35.15 27.43 35.36 27.5 ;
    RECT 117.69 26.71 117.9 26.78 ;
    RECT 117.69 27.07 117.9 27.14 ;
    RECT 117.69 27.43 117.9 27.5 ;
    RECT 118.15 26.71 118.36 26.78 ;
    RECT 118.15 27.07 118.36 27.14 ;
    RECT 118.15 27.43 118.36 27.5 ;
    RECT 114.37 26.71 114.58 26.78 ;
    RECT 114.37 27.07 114.58 27.14 ;
    RECT 114.37 27.43 114.58 27.5 ;
    RECT 114.83 26.71 115.04 26.78 ;
    RECT 114.83 27.07 115.04 27.14 ;
    RECT 114.83 27.43 115.04 27.5 ;
    RECT 111.05 26.71 111.26 26.78 ;
    RECT 111.05 27.07 111.26 27.14 ;
    RECT 111.05 27.43 111.26 27.5 ;
    RECT 111.51 26.71 111.72 26.78 ;
    RECT 111.51 27.07 111.72 27.14 ;
    RECT 111.51 27.43 111.72 27.5 ;
    RECT 107.73 26.71 107.94 26.78 ;
    RECT 107.73 27.07 107.94 27.14 ;
    RECT 107.73 27.43 107.94 27.5 ;
    RECT 108.19 26.71 108.4 26.78 ;
    RECT 108.19 27.07 108.4 27.14 ;
    RECT 108.19 27.43 108.4 27.5 ;
    RECT 104.41 26.71 104.62 26.78 ;
    RECT 104.41 27.07 104.62 27.14 ;
    RECT 104.41 27.43 104.62 27.5 ;
    RECT 104.87 26.71 105.08 26.78 ;
    RECT 104.87 27.07 105.08 27.14 ;
    RECT 104.87 27.43 105.08 27.5 ;
    RECT 101.09 26.71 101.3 26.78 ;
    RECT 101.09 27.07 101.3 27.14 ;
    RECT 101.09 27.43 101.3 27.5 ;
    RECT 101.55 26.71 101.76 26.78 ;
    RECT 101.55 27.07 101.76 27.14 ;
    RECT 101.55 27.43 101.76 27.5 ;
    RECT 97.77 26.71 97.98 26.78 ;
    RECT 97.77 27.07 97.98 27.14 ;
    RECT 97.77 27.43 97.98 27.5 ;
    RECT 98.23 26.71 98.44 26.78 ;
    RECT 98.23 27.07 98.44 27.14 ;
    RECT 98.23 27.43 98.44 27.5 ;
    RECT 94.45 26.71 94.66 26.78 ;
    RECT 94.45 27.07 94.66 27.14 ;
    RECT 94.45 27.43 94.66 27.5 ;
    RECT 94.91 26.71 95.12 26.78 ;
    RECT 94.91 27.07 95.12 27.14 ;
    RECT 94.91 27.43 95.12 27.5 ;
    RECT 91.13 26.71 91.34 26.78 ;
    RECT 91.13 27.07 91.34 27.14 ;
    RECT 91.13 27.43 91.34 27.5 ;
    RECT 91.59 26.71 91.8 26.78 ;
    RECT 91.59 27.07 91.8 27.14 ;
    RECT 91.59 27.43 91.8 27.5 ;
    RECT 87.81 26.71 88.02 26.78 ;
    RECT 87.81 27.07 88.02 27.14 ;
    RECT 87.81 27.43 88.02 27.5 ;
    RECT 88.27 26.71 88.48 26.78 ;
    RECT 88.27 27.07 88.48 27.14 ;
    RECT 88.27 27.43 88.48 27.5 ;
    RECT 84.49 26.71 84.7 26.78 ;
    RECT 84.49 27.07 84.7 27.14 ;
    RECT 84.49 27.43 84.7 27.5 ;
    RECT 84.95 26.71 85.16 26.78 ;
    RECT 84.95 27.07 85.16 27.14 ;
    RECT 84.95 27.43 85.16 27.5 ;
    RECT 81.17 26.71 81.38 26.78 ;
    RECT 81.17 27.07 81.38 27.14 ;
    RECT 81.17 27.43 81.38 27.5 ;
    RECT 81.63 26.71 81.84 26.78 ;
    RECT 81.63 27.07 81.84 27.14 ;
    RECT 81.63 27.43 81.84 27.5 ;
    RECT 77.85 26.71 78.06 26.78 ;
    RECT 77.85 27.07 78.06 27.14 ;
    RECT 77.85 27.43 78.06 27.5 ;
    RECT 78.31 26.71 78.52 26.78 ;
    RECT 78.31 27.07 78.52 27.14 ;
    RECT 78.31 27.43 78.52 27.5 ;
    RECT 74.53 26.71 74.74 26.78 ;
    RECT 74.53 27.07 74.74 27.14 ;
    RECT 74.53 27.43 74.74 27.5 ;
    RECT 74.99 26.71 75.2 26.78 ;
    RECT 74.99 27.07 75.2 27.14 ;
    RECT 74.99 27.43 75.2 27.5 ;
    RECT 71.21 26.71 71.42 26.78 ;
    RECT 71.21 27.07 71.42 27.14 ;
    RECT 71.21 27.43 71.42 27.5 ;
    RECT 71.67 26.71 71.88 26.78 ;
    RECT 71.67 27.07 71.88 27.14 ;
    RECT 71.67 27.43 71.88 27.5 ;
    RECT 31.37 26.71 31.58 26.78 ;
    RECT 31.37 27.07 31.58 27.14 ;
    RECT 31.37 27.43 31.58 27.5 ;
    RECT 31.83 26.71 32.04 26.78 ;
    RECT 31.83 27.07 32.04 27.14 ;
    RECT 31.83 27.43 32.04 27.5 ;
    RECT 67.89 26.71 68.1 26.78 ;
    RECT 67.89 27.07 68.1 27.14 ;
    RECT 67.89 27.43 68.1 27.5 ;
    RECT 68.35 26.71 68.56 26.78 ;
    RECT 68.35 27.07 68.56 27.14 ;
    RECT 68.35 27.43 68.56 27.5 ;
    RECT 28.05 26.71 28.26 26.78 ;
    RECT 28.05 27.07 28.26 27.14 ;
    RECT 28.05 27.43 28.26 27.5 ;
    RECT 28.51 26.71 28.72 26.78 ;
    RECT 28.51 27.07 28.72 27.14 ;
    RECT 28.51 27.43 28.72 27.5 ;
    RECT 24.73 26.71 24.94 26.78 ;
    RECT 24.73 27.07 24.94 27.14 ;
    RECT 24.73 27.43 24.94 27.5 ;
    RECT 25.19 26.71 25.4 26.78 ;
    RECT 25.19 27.07 25.4 27.14 ;
    RECT 25.19 27.43 25.4 27.5 ;
    RECT 21.41 26.71 21.62 26.78 ;
    RECT 21.41 27.07 21.62 27.14 ;
    RECT 21.41 27.43 21.62 27.5 ;
    RECT 21.87 26.71 22.08 26.78 ;
    RECT 21.87 27.07 22.08 27.14 ;
    RECT 21.87 27.43 22.08 27.5 ;
    RECT 18.09 26.71 18.3 26.78 ;
    RECT 18.09 27.07 18.3 27.14 ;
    RECT 18.09 27.43 18.3 27.5 ;
    RECT 18.55 26.71 18.76 26.78 ;
    RECT 18.55 27.07 18.76 27.14 ;
    RECT 18.55 27.43 18.76 27.5 ;
    RECT 120.825 27.07 120.895 27.14 ;
    RECT 14.77 26.71 14.98 26.78 ;
    RECT 14.77 27.07 14.98 27.14 ;
    RECT 14.77 27.43 14.98 27.5 ;
    RECT 15.23 26.71 15.44 26.78 ;
    RECT 15.23 27.07 15.44 27.14 ;
    RECT 15.23 27.43 15.44 27.5 ;
    RECT 11.45 26.71 11.66 26.78 ;
    RECT 11.45 27.07 11.66 27.14 ;
    RECT 11.45 27.43 11.66 27.5 ;
    RECT 11.91 26.71 12.12 26.78 ;
    RECT 11.91 27.07 12.12 27.14 ;
    RECT 11.91 27.43 12.12 27.5 ;
    RECT 8.13 26.71 8.34 26.78 ;
    RECT 8.13 27.07 8.34 27.14 ;
    RECT 8.13 27.43 8.34 27.5 ;
    RECT 8.59 26.71 8.8 26.78 ;
    RECT 8.59 27.07 8.8 27.14 ;
    RECT 8.59 27.43 8.8 27.5 ;
    RECT 4.81 26.71 5.02 26.78 ;
    RECT 4.81 27.07 5.02 27.14 ;
    RECT 4.81 27.43 5.02 27.5 ;
    RECT 5.27 26.71 5.48 26.78 ;
    RECT 5.27 27.07 5.48 27.14 ;
    RECT 5.27 27.43 5.48 27.5 ;
    RECT 1.49 26.71 1.7 26.78 ;
    RECT 1.49 27.07 1.7 27.14 ;
    RECT 1.49 27.43 1.7 27.5 ;
    RECT 1.95 26.71 2.16 26.78 ;
    RECT 1.95 27.07 2.16 27.14 ;
    RECT 1.95 27.43 2.16 27.5 ;
    RECT 64.57 26.71 64.78 26.78 ;
    RECT 64.57 27.07 64.78 27.14 ;
    RECT 64.57 27.43 64.78 27.5 ;
    RECT 65.03 26.71 65.24 26.78 ;
    RECT 65.03 27.07 65.24 27.14 ;
    RECT 65.03 27.43 65.24 27.5 ;
    RECT 61.25 25.99 61.46 26.06 ;
    RECT 61.25 26.35 61.46 26.42 ;
    RECT 61.25 26.71 61.46 26.78 ;
    RECT 61.71 25.99 61.92 26.06 ;
    RECT 61.71 26.35 61.92 26.42 ;
    RECT 61.71 26.71 61.92 26.78 ;
    RECT 57.93 25.99 58.14 26.06 ;
    RECT 57.93 26.35 58.14 26.42 ;
    RECT 57.93 26.71 58.14 26.78 ;
    RECT 58.39 25.99 58.6 26.06 ;
    RECT 58.39 26.35 58.6 26.42 ;
    RECT 58.39 26.71 58.6 26.78 ;
    RECT 54.61 25.99 54.82 26.06 ;
    RECT 54.61 26.35 54.82 26.42 ;
    RECT 54.61 26.71 54.82 26.78 ;
    RECT 55.07 25.99 55.28 26.06 ;
    RECT 55.07 26.35 55.28 26.42 ;
    RECT 55.07 26.71 55.28 26.78 ;
    RECT 51.29 25.99 51.5 26.06 ;
    RECT 51.29 26.35 51.5 26.42 ;
    RECT 51.29 26.71 51.5 26.78 ;
    RECT 51.75 25.99 51.96 26.06 ;
    RECT 51.75 26.35 51.96 26.42 ;
    RECT 51.75 26.71 51.96 26.78 ;
    RECT 47.97 25.99 48.18 26.06 ;
    RECT 47.97 26.35 48.18 26.42 ;
    RECT 47.97 26.71 48.18 26.78 ;
    RECT 48.43 25.99 48.64 26.06 ;
    RECT 48.43 26.35 48.64 26.42 ;
    RECT 48.43 26.71 48.64 26.78 ;
    RECT 44.65 25.99 44.86 26.06 ;
    RECT 44.65 26.35 44.86 26.42 ;
    RECT 44.65 26.71 44.86 26.78 ;
    RECT 45.11 25.99 45.32 26.06 ;
    RECT 45.11 26.35 45.32 26.42 ;
    RECT 45.11 26.71 45.32 26.78 ;
    RECT 41.33 25.99 41.54 26.06 ;
    RECT 41.33 26.35 41.54 26.42 ;
    RECT 41.33 26.71 41.54 26.78 ;
    RECT 41.79 25.99 42.0 26.06 ;
    RECT 41.79 26.35 42.0 26.42 ;
    RECT 41.79 26.71 42.0 26.78 ;
    RECT 38.01 25.99 38.22 26.06 ;
    RECT 38.01 26.35 38.22 26.42 ;
    RECT 38.01 26.71 38.22 26.78 ;
    RECT 38.47 25.99 38.68 26.06 ;
    RECT 38.47 26.35 38.68 26.42 ;
    RECT 38.47 26.71 38.68 26.78 ;
    RECT 0.4 26.35 0.47 26.42 ;
    RECT 34.69 25.99 34.9 26.06 ;
    RECT 34.69 26.35 34.9 26.42 ;
    RECT 34.69 26.71 34.9 26.78 ;
    RECT 35.15 25.99 35.36 26.06 ;
    RECT 35.15 26.35 35.36 26.42 ;
    RECT 35.15 26.71 35.36 26.78 ;
    RECT 117.69 25.99 117.9 26.06 ;
    RECT 117.69 26.35 117.9 26.42 ;
    RECT 117.69 26.71 117.9 26.78 ;
    RECT 118.15 25.99 118.36 26.06 ;
    RECT 118.15 26.35 118.36 26.42 ;
    RECT 118.15 26.71 118.36 26.78 ;
    RECT 114.37 25.99 114.58 26.06 ;
    RECT 114.37 26.35 114.58 26.42 ;
    RECT 114.37 26.71 114.58 26.78 ;
    RECT 114.83 25.99 115.04 26.06 ;
    RECT 114.83 26.35 115.04 26.42 ;
    RECT 114.83 26.71 115.04 26.78 ;
    RECT 111.05 25.99 111.26 26.06 ;
    RECT 111.05 26.35 111.26 26.42 ;
    RECT 111.05 26.71 111.26 26.78 ;
    RECT 111.51 25.99 111.72 26.06 ;
    RECT 111.51 26.35 111.72 26.42 ;
    RECT 111.51 26.71 111.72 26.78 ;
    RECT 107.73 25.99 107.94 26.06 ;
    RECT 107.73 26.35 107.94 26.42 ;
    RECT 107.73 26.71 107.94 26.78 ;
    RECT 108.19 25.99 108.4 26.06 ;
    RECT 108.19 26.35 108.4 26.42 ;
    RECT 108.19 26.71 108.4 26.78 ;
    RECT 104.41 25.99 104.62 26.06 ;
    RECT 104.41 26.35 104.62 26.42 ;
    RECT 104.41 26.71 104.62 26.78 ;
    RECT 104.87 25.99 105.08 26.06 ;
    RECT 104.87 26.35 105.08 26.42 ;
    RECT 104.87 26.71 105.08 26.78 ;
    RECT 101.09 25.99 101.3 26.06 ;
    RECT 101.09 26.35 101.3 26.42 ;
    RECT 101.09 26.71 101.3 26.78 ;
    RECT 101.55 25.99 101.76 26.06 ;
    RECT 101.55 26.35 101.76 26.42 ;
    RECT 101.55 26.71 101.76 26.78 ;
    RECT 97.77 25.99 97.98 26.06 ;
    RECT 97.77 26.35 97.98 26.42 ;
    RECT 97.77 26.71 97.98 26.78 ;
    RECT 98.23 25.99 98.44 26.06 ;
    RECT 98.23 26.35 98.44 26.42 ;
    RECT 98.23 26.71 98.44 26.78 ;
    RECT 94.45 25.99 94.66 26.06 ;
    RECT 94.45 26.35 94.66 26.42 ;
    RECT 94.45 26.71 94.66 26.78 ;
    RECT 94.91 25.99 95.12 26.06 ;
    RECT 94.91 26.35 95.12 26.42 ;
    RECT 94.91 26.71 95.12 26.78 ;
    RECT 91.13 25.99 91.34 26.06 ;
    RECT 91.13 26.35 91.34 26.42 ;
    RECT 91.13 26.71 91.34 26.78 ;
    RECT 91.59 25.99 91.8 26.06 ;
    RECT 91.59 26.35 91.8 26.42 ;
    RECT 91.59 26.71 91.8 26.78 ;
    RECT 87.81 25.99 88.02 26.06 ;
    RECT 87.81 26.35 88.02 26.42 ;
    RECT 87.81 26.71 88.02 26.78 ;
    RECT 88.27 25.99 88.48 26.06 ;
    RECT 88.27 26.35 88.48 26.42 ;
    RECT 88.27 26.71 88.48 26.78 ;
    RECT 84.49 25.99 84.7 26.06 ;
    RECT 84.49 26.35 84.7 26.42 ;
    RECT 84.49 26.71 84.7 26.78 ;
    RECT 84.95 25.99 85.16 26.06 ;
    RECT 84.95 26.35 85.16 26.42 ;
    RECT 84.95 26.71 85.16 26.78 ;
    RECT 81.17 25.99 81.38 26.06 ;
    RECT 81.17 26.35 81.38 26.42 ;
    RECT 81.17 26.71 81.38 26.78 ;
    RECT 81.63 25.99 81.84 26.06 ;
    RECT 81.63 26.35 81.84 26.42 ;
    RECT 81.63 26.71 81.84 26.78 ;
    RECT 77.85 25.99 78.06 26.06 ;
    RECT 77.85 26.35 78.06 26.42 ;
    RECT 77.85 26.71 78.06 26.78 ;
    RECT 78.31 25.99 78.52 26.06 ;
    RECT 78.31 26.35 78.52 26.42 ;
    RECT 78.31 26.71 78.52 26.78 ;
    RECT 74.53 25.99 74.74 26.06 ;
    RECT 74.53 26.35 74.74 26.42 ;
    RECT 74.53 26.71 74.74 26.78 ;
    RECT 74.99 25.99 75.2 26.06 ;
    RECT 74.99 26.35 75.2 26.42 ;
    RECT 74.99 26.71 75.2 26.78 ;
    RECT 71.21 25.99 71.42 26.06 ;
    RECT 71.21 26.35 71.42 26.42 ;
    RECT 71.21 26.71 71.42 26.78 ;
    RECT 71.67 25.99 71.88 26.06 ;
    RECT 71.67 26.35 71.88 26.42 ;
    RECT 71.67 26.71 71.88 26.78 ;
    RECT 31.37 25.99 31.58 26.06 ;
    RECT 31.37 26.35 31.58 26.42 ;
    RECT 31.37 26.71 31.58 26.78 ;
    RECT 31.83 25.99 32.04 26.06 ;
    RECT 31.83 26.35 32.04 26.42 ;
    RECT 31.83 26.71 32.04 26.78 ;
    RECT 67.89 25.99 68.1 26.06 ;
    RECT 67.89 26.35 68.1 26.42 ;
    RECT 67.89 26.71 68.1 26.78 ;
    RECT 68.35 25.99 68.56 26.06 ;
    RECT 68.35 26.35 68.56 26.42 ;
    RECT 68.35 26.71 68.56 26.78 ;
    RECT 28.05 25.99 28.26 26.06 ;
    RECT 28.05 26.35 28.26 26.42 ;
    RECT 28.05 26.71 28.26 26.78 ;
    RECT 28.51 25.99 28.72 26.06 ;
    RECT 28.51 26.35 28.72 26.42 ;
    RECT 28.51 26.71 28.72 26.78 ;
    RECT 24.73 25.99 24.94 26.06 ;
    RECT 24.73 26.35 24.94 26.42 ;
    RECT 24.73 26.71 24.94 26.78 ;
    RECT 25.19 25.99 25.4 26.06 ;
    RECT 25.19 26.35 25.4 26.42 ;
    RECT 25.19 26.71 25.4 26.78 ;
    RECT 21.41 25.99 21.62 26.06 ;
    RECT 21.41 26.35 21.62 26.42 ;
    RECT 21.41 26.71 21.62 26.78 ;
    RECT 21.87 25.99 22.08 26.06 ;
    RECT 21.87 26.35 22.08 26.42 ;
    RECT 21.87 26.71 22.08 26.78 ;
    RECT 18.09 25.99 18.3 26.06 ;
    RECT 18.09 26.35 18.3 26.42 ;
    RECT 18.09 26.71 18.3 26.78 ;
    RECT 18.55 25.99 18.76 26.06 ;
    RECT 18.55 26.35 18.76 26.42 ;
    RECT 18.55 26.71 18.76 26.78 ;
    RECT 120.825 26.35 120.895 26.42 ;
    RECT 14.77 25.99 14.98 26.06 ;
    RECT 14.77 26.35 14.98 26.42 ;
    RECT 14.77 26.71 14.98 26.78 ;
    RECT 15.23 25.99 15.44 26.06 ;
    RECT 15.23 26.35 15.44 26.42 ;
    RECT 15.23 26.71 15.44 26.78 ;
    RECT 11.45 25.99 11.66 26.06 ;
    RECT 11.45 26.35 11.66 26.42 ;
    RECT 11.45 26.71 11.66 26.78 ;
    RECT 11.91 25.99 12.12 26.06 ;
    RECT 11.91 26.35 12.12 26.42 ;
    RECT 11.91 26.71 12.12 26.78 ;
    RECT 8.13 25.99 8.34 26.06 ;
    RECT 8.13 26.35 8.34 26.42 ;
    RECT 8.13 26.71 8.34 26.78 ;
    RECT 8.59 25.99 8.8 26.06 ;
    RECT 8.59 26.35 8.8 26.42 ;
    RECT 8.59 26.71 8.8 26.78 ;
    RECT 4.81 25.99 5.02 26.06 ;
    RECT 4.81 26.35 5.02 26.42 ;
    RECT 4.81 26.71 5.02 26.78 ;
    RECT 5.27 25.99 5.48 26.06 ;
    RECT 5.27 26.35 5.48 26.42 ;
    RECT 5.27 26.71 5.48 26.78 ;
    RECT 1.49 25.99 1.7 26.06 ;
    RECT 1.49 26.35 1.7 26.42 ;
    RECT 1.49 26.71 1.7 26.78 ;
    RECT 1.95 25.99 2.16 26.06 ;
    RECT 1.95 26.35 2.16 26.42 ;
    RECT 1.95 26.71 2.16 26.78 ;
    RECT 64.57 25.99 64.78 26.06 ;
    RECT 64.57 26.35 64.78 26.42 ;
    RECT 64.57 26.71 64.78 26.78 ;
    RECT 65.03 25.99 65.24 26.06 ;
    RECT 65.03 26.35 65.24 26.42 ;
    RECT 65.03 26.71 65.24 26.78 ;
    RECT 61.25 25.27 61.46 25.34 ;
    RECT 61.25 25.63 61.46 25.7 ;
    RECT 61.25 25.99 61.46 26.06 ;
    RECT 61.71 25.27 61.92 25.34 ;
    RECT 61.71 25.63 61.92 25.7 ;
    RECT 61.71 25.99 61.92 26.06 ;
    RECT 57.93 25.27 58.14 25.34 ;
    RECT 57.93 25.63 58.14 25.7 ;
    RECT 57.93 25.99 58.14 26.06 ;
    RECT 58.39 25.27 58.6 25.34 ;
    RECT 58.39 25.63 58.6 25.7 ;
    RECT 58.39 25.99 58.6 26.06 ;
    RECT 54.61 25.27 54.82 25.34 ;
    RECT 54.61 25.63 54.82 25.7 ;
    RECT 54.61 25.99 54.82 26.06 ;
    RECT 55.07 25.27 55.28 25.34 ;
    RECT 55.07 25.63 55.28 25.7 ;
    RECT 55.07 25.99 55.28 26.06 ;
    RECT 51.29 25.27 51.5 25.34 ;
    RECT 51.29 25.63 51.5 25.7 ;
    RECT 51.29 25.99 51.5 26.06 ;
    RECT 51.75 25.27 51.96 25.34 ;
    RECT 51.75 25.63 51.96 25.7 ;
    RECT 51.75 25.99 51.96 26.06 ;
    RECT 47.97 25.27 48.18 25.34 ;
    RECT 47.97 25.63 48.18 25.7 ;
    RECT 47.97 25.99 48.18 26.06 ;
    RECT 48.43 25.27 48.64 25.34 ;
    RECT 48.43 25.63 48.64 25.7 ;
    RECT 48.43 25.99 48.64 26.06 ;
    RECT 44.65 25.27 44.86 25.34 ;
    RECT 44.65 25.63 44.86 25.7 ;
    RECT 44.65 25.99 44.86 26.06 ;
    RECT 45.11 25.27 45.32 25.34 ;
    RECT 45.11 25.63 45.32 25.7 ;
    RECT 45.11 25.99 45.32 26.06 ;
    RECT 41.33 25.27 41.54 25.34 ;
    RECT 41.33 25.63 41.54 25.7 ;
    RECT 41.33 25.99 41.54 26.06 ;
    RECT 41.79 25.27 42.0 25.34 ;
    RECT 41.79 25.63 42.0 25.7 ;
    RECT 41.79 25.99 42.0 26.06 ;
    RECT 38.01 25.27 38.22 25.34 ;
    RECT 38.01 25.63 38.22 25.7 ;
    RECT 38.01 25.99 38.22 26.06 ;
    RECT 38.47 25.27 38.68 25.34 ;
    RECT 38.47 25.63 38.68 25.7 ;
    RECT 38.47 25.99 38.68 26.06 ;
    RECT 0.4 25.63 0.47 25.7 ;
    RECT 34.69 25.27 34.9 25.34 ;
    RECT 34.69 25.63 34.9 25.7 ;
    RECT 34.69 25.99 34.9 26.06 ;
    RECT 35.15 25.27 35.36 25.34 ;
    RECT 35.15 25.63 35.36 25.7 ;
    RECT 35.15 25.99 35.36 26.06 ;
    RECT 117.69 25.27 117.9 25.34 ;
    RECT 117.69 25.63 117.9 25.7 ;
    RECT 117.69 25.99 117.9 26.06 ;
    RECT 118.15 25.27 118.36 25.34 ;
    RECT 118.15 25.63 118.36 25.7 ;
    RECT 118.15 25.99 118.36 26.06 ;
    RECT 114.37 25.27 114.58 25.34 ;
    RECT 114.37 25.63 114.58 25.7 ;
    RECT 114.37 25.99 114.58 26.06 ;
    RECT 114.83 25.27 115.04 25.34 ;
    RECT 114.83 25.63 115.04 25.7 ;
    RECT 114.83 25.99 115.04 26.06 ;
    RECT 111.05 25.27 111.26 25.34 ;
    RECT 111.05 25.63 111.26 25.7 ;
    RECT 111.05 25.99 111.26 26.06 ;
    RECT 111.51 25.27 111.72 25.34 ;
    RECT 111.51 25.63 111.72 25.7 ;
    RECT 111.51 25.99 111.72 26.06 ;
    RECT 107.73 25.27 107.94 25.34 ;
    RECT 107.73 25.63 107.94 25.7 ;
    RECT 107.73 25.99 107.94 26.06 ;
    RECT 108.19 25.27 108.4 25.34 ;
    RECT 108.19 25.63 108.4 25.7 ;
    RECT 108.19 25.99 108.4 26.06 ;
    RECT 104.41 25.27 104.62 25.34 ;
    RECT 104.41 25.63 104.62 25.7 ;
    RECT 104.41 25.99 104.62 26.06 ;
    RECT 104.87 25.27 105.08 25.34 ;
    RECT 104.87 25.63 105.08 25.7 ;
    RECT 104.87 25.99 105.08 26.06 ;
    RECT 101.09 25.27 101.3 25.34 ;
    RECT 101.09 25.63 101.3 25.7 ;
    RECT 101.09 25.99 101.3 26.06 ;
    RECT 101.55 25.27 101.76 25.34 ;
    RECT 101.55 25.63 101.76 25.7 ;
    RECT 101.55 25.99 101.76 26.06 ;
    RECT 97.77 25.27 97.98 25.34 ;
    RECT 97.77 25.63 97.98 25.7 ;
    RECT 97.77 25.99 97.98 26.06 ;
    RECT 98.23 25.27 98.44 25.34 ;
    RECT 98.23 25.63 98.44 25.7 ;
    RECT 98.23 25.99 98.44 26.06 ;
    RECT 94.45 25.27 94.66 25.34 ;
    RECT 94.45 25.63 94.66 25.7 ;
    RECT 94.45 25.99 94.66 26.06 ;
    RECT 94.91 25.27 95.12 25.34 ;
    RECT 94.91 25.63 95.12 25.7 ;
    RECT 94.91 25.99 95.12 26.06 ;
    RECT 91.13 25.27 91.34 25.34 ;
    RECT 91.13 25.63 91.34 25.7 ;
    RECT 91.13 25.99 91.34 26.06 ;
    RECT 91.59 25.27 91.8 25.34 ;
    RECT 91.59 25.63 91.8 25.7 ;
    RECT 91.59 25.99 91.8 26.06 ;
    RECT 87.81 25.27 88.02 25.34 ;
    RECT 87.81 25.63 88.02 25.7 ;
    RECT 87.81 25.99 88.02 26.06 ;
    RECT 88.27 25.27 88.48 25.34 ;
    RECT 88.27 25.63 88.48 25.7 ;
    RECT 88.27 25.99 88.48 26.06 ;
    RECT 84.49 25.27 84.7 25.34 ;
    RECT 84.49 25.63 84.7 25.7 ;
    RECT 84.49 25.99 84.7 26.06 ;
    RECT 84.95 25.27 85.16 25.34 ;
    RECT 84.95 25.63 85.16 25.7 ;
    RECT 84.95 25.99 85.16 26.06 ;
    RECT 81.17 25.27 81.38 25.34 ;
    RECT 81.17 25.63 81.38 25.7 ;
    RECT 81.17 25.99 81.38 26.06 ;
    RECT 81.63 25.27 81.84 25.34 ;
    RECT 81.63 25.63 81.84 25.7 ;
    RECT 81.63 25.99 81.84 26.06 ;
    RECT 77.85 25.27 78.06 25.34 ;
    RECT 77.85 25.63 78.06 25.7 ;
    RECT 77.85 25.99 78.06 26.06 ;
    RECT 78.31 25.27 78.52 25.34 ;
    RECT 78.31 25.63 78.52 25.7 ;
    RECT 78.31 25.99 78.52 26.06 ;
    RECT 74.53 25.27 74.74 25.34 ;
    RECT 74.53 25.63 74.74 25.7 ;
    RECT 74.53 25.99 74.74 26.06 ;
    RECT 74.99 25.27 75.2 25.34 ;
    RECT 74.99 25.63 75.2 25.7 ;
    RECT 74.99 25.99 75.2 26.06 ;
    RECT 71.21 25.27 71.42 25.34 ;
    RECT 71.21 25.63 71.42 25.7 ;
    RECT 71.21 25.99 71.42 26.06 ;
    RECT 71.67 25.27 71.88 25.34 ;
    RECT 71.67 25.63 71.88 25.7 ;
    RECT 71.67 25.99 71.88 26.06 ;
    RECT 31.37 25.27 31.58 25.34 ;
    RECT 31.37 25.63 31.58 25.7 ;
    RECT 31.37 25.99 31.58 26.06 ;
    RECT 31.83 25.27 32.04 25.34 ;
    RECT 31.83 25.63 32.04 25.7 ;
    RECT 31.83 25.99 32.04 26.06 ;
    RECT 67.89 25.27 68.1 25.34 ;
    RECT 67.89 25.63 68.1 25.7 ;
    RECT 67.89 25.99 68.1 26.06 ;
    RECT 68.35 25.27 68.56 25.34 ;
    RECT 68.35 25.63 68.56 25.7 ;
    RECT 68.35 25.99 68.56 26.06 ;
    RECT 28.05 25.27 28.26 25.34 ;
    RECT 28.05 25.63 28.26 25.7 ;
    RECT 28.05 25.99 28.26 26.06 ;
    RECT 28.51 25.27 28.72 25.34 ;
    RECT 28.51 25.63 28.72 25.7 ;
    RECT 28.51 25.99 28.72 26.06 ;
    RECT 24.73 25.27 24.94 25.34 ;
    RECT 24.73 25.63 24.94 25.7 ;
    RECT 24.73 25.99 24.94 26.06 ;
    RECT 25.19 25.27 25.4 25.34 ;
    RECT 25.19 25.63 25.4 25.7 ;
    RECT 25.19 25.99 25.4 26.06 ;
    RECT 21.41 25.27 21.62 25.34 ;
    RECT 21.41 25.63 21.62 25.7 ;
    RECT 21.41 25.99 21.62 26.06 ;
    RECT 21.87 25.27 22.08 25.34 ;
    RECT 21.87 25.63 22.08 25.7 ;
    RECT 21.87 25.99 22.08 26.06 ;
    RECT 18.09 25.27 18.3 25.34 ;
    RECT 18.09 25.63 18.3 25.7 ;
    RECT 18.09 25.99 18.3 26.06 ;
    RECT 18.55 25.27 18.76 25.34 ;
    RECT 18.55 25.63 18.76 25.7 ;
    RECT 18.55 25.99 18.76 26.06 ;
    RECT 120.825 25.63 120.895 25.7 ;
    RECT 14.77 25.27 14.98 25.34 ;
    RECT 14.77 25.63 14.98 25.7 ;
    RECT 14.77 25.99 14.98 26.06 ;
    RECT 15.23 25.27 15.44 25.34 ;
    RECT 15.23 25.63 15.44 25.7 ;
    RECT 15.23 25.99 15.44 26.06 ;
    RECT 11.45 25.27 11.66 25.34 ;
    RECT 11.45 25.63 11.66 25.7 ;
    RECT 11.45 25.99 11.66 26.06 ;
    RECT 11.91 25.27 12.12 25.34 ;
    RECT 11.91 25.63 12.12 25.7 ;
    RECT 11.91 25.99 12.12 26.06 ;
    RECT 8.13 25.27 8.34 25.34 ;
    RECT 8.13 25.63 8.34 25.7 ;
    RECT 8.13 25.99 8.34 26.06 ;
    RECT 8.59 25.27 8.8 25.34 ;
    RECT 8.59 25.63 8.8 25.7 ;
    RECT 8.59 25.99 8.8 26.06 ;
    RECT 4.81 25.27 5.02 25.34 ;
    RECT 4.81 25.63 5.02 25.7 ;
    RECT 4.81 25.99 5.02 26.06 ;
    RECT 5.27 25.27 5.48 25.34 ;
    RECT 5.27 25.63 5.48 25.7 ;
    RECT 5.27 25.99 5.48 26.06 ;
    RECT 1.49 25.27 1.7 25.34 ;
    RECT 1.49 25.63 1.7 25.7 ;
    RECT 1.49 25.99 1.7 26.06 ;
    RECT 1.95 25.27 2.16 25.34 ;
    RECT 1.95 25.63 2.16 25.7 ;
    RECT 1.95 25.99 2.16 26.06 ;
    RECT 64.57 25.27 64.78 25.34 ;
    RECT 64.57 25.63 64.78 25.7 ;
    RECT 64.57 25.99 64.78 26.06 ;
    RECT 65.03 25.27 65.24 25.34 ;
    RECT 65.03 25.63 65.24 25.7 ;
    RECT 65.03 25.99 65.24 26.06 ;
    RECT 61.25 64.89 61.46 64.96 ;
    RECT 61.25 65.25 61.46 65.32 ;
    RECT 61.25 65.61 61.46 65.68 ;
    RECT 61.71 64.89 61.92 64.96 ;
    RECT 61.71 65.25 61.92 65.32 ;
    RECT 61.71 65.61 61.92 65.68 ;
    RECT 57.93 64.89 58.14 64.96 ;
    RECT 57.93 65.25 58.14 65.32 ;
    RECT 57.93 65.61 58.14 65.68 ;
    RECT 58.39 64.89 58.6 64.96 ;
    RECT 58.39 65.25 58.6 65.32 ;
    RECT 58.39 65.61 58.6 65.68 ;
    RECT 54.61 64.89 54.82 64.96 ;
    RECT 54.61 65.25 54.82 65.32 ;
    RECT 54.61 65.61 54.82 65.68 ;
    RECT 55.07 64.89 55.28 64.96 ;
    RECT 55.07 65.25 55.28 65.32 ;
    RECT 55.07 65.61 55.28 65.68 ;
    RECT 51.29 64.89 51.5 64.96 ;
    RECT 51.29 65.25 51.5 65.32 ;
    RECT 51.29 65.61 51.5 65.68 ;
    RECT 51.75 64.89 51.96 64.96 ;
    RECT 51.75 65.25 51.96 65.32 ;
    RECT 51.75 65.61 51.96 65.68 ;
    RECT 47.97 64.89 48.18 64.96 ;
    RECT 47.97 65.25 48.18 65.32 ;
    RECT 47.97 65.61 48.18 65.68 ;
    RECT 48.43 64.89 48.64 64.96 ;
    RECT 48.43 65.25 48.64 65.32 ;
    RECT 48.43 65.61 48.64 65.68 ;
    RECT 44.65 64.89 44.86 64.96 ;
    RECT 44.65 65.25 44.86 65.32 ;
    RECT 44.65 65.61 44.86 65.68 ;
    RECT 45.11 64.89 45.32 64.96 ;
    RECT 45.11 65.25 45.32 65.32 ;
    RECT 45.11 65.61 45.32 65.68 ;
    RECT 41.33 64.89 41.54 64.96 ;
    RECT 41.33 65.25 41.54 65.32 ;
    RECT 41.33 65.61 41.54 65.68 ;
    RECT 41.79 64.89 42.0 64.96 ;
    RECT 41.79 65.25 42.0 65.32 ;
    RECT 41.79 65.61 42.0 65.68 ;
    RECT 38.01 64.89 38.22 64.96 ;
    RECT 38.01 65.25 38.22 65.32 ;
    RECT 38.01 65.61 38.22 65.68 ;
    RECT 38.47 64.89 38.68 64.96 ;
    RECT 38.47 65.25 38.68 65.32 ;
    RECT 38.47 65.61 38.68 65.68 ;
    RECT 0.4 65.25 0.47 65.32 ;
    RECT 34.69 64.89 34.9 64.96 ;
    RECT 34.69 65.25 34.9 65.32 ;
    RECT 34.69 65.61 34.9 65.68 ;
    RECT 35.15 64.89 35.36 64.96 ;
    RECT 35.15 65.25 35.36 65.32 ;
    RECT 35.15 65.61 35.36 65.68 ;
    RECT 117.69 64.89 117.9 64.96 ;
    RECT 117.69 65.25 117.9 65.32 ;
    RECT 117.69 65.61 117.9 65.68 ;
    RECT 118.15 64.89 118.36 64.96 ;
    RECT 118.15 65.25 118.36 65.32 ;
    RECT 118.15 65.61 118.36 65.68 ;
    RECT 114.37 64.89 114.58 64.96 ;
    RECT 114.37 65.25 114.58 65.32 ;
    RECT 114.37 65.61 114.58 65.68 ;
    RECT 114.83 64.89 115.04 64.96 ;
    RECT 114.83 65.25 115.04 65.32 ;
    RECT 114.83 65.61 115.04 65.68 ;
    RECT 111.05 64.89 111.26 64.96 ;
    RECT 111.05 65.25 111.26 65.32 ;
    RECT 111.05 65.61 111.26 65.68 ;
    RECT 111.51 64.89 111.72 64.96 ;
    RECT 111.51 65.25 111.72 65.32 ;
    RECT 111.51 65.61 111.72 65.68 ;
    RECT 107.73 64.89 107.94 64.96 ;
    RECT 107.73 65.25 107.94 65.32 ;
    RECT 107.73 65.61 107.94 65.68 ;
    RECT 108.19 64.89 108.4 64.96 ;
    RECT 108.19 65.25 108.4 65.32 ;
    RECT 108.19 65.61 108.4 65.68 ;
    RECT 104.41 64.89 104.62 64.96 ;
    RECT 104.41 65.25 104.62 65.32 ;
    RECT 104.41 65.61 104.62 65.68 ;
    RECT 104.87 64.89 105.08 64.96 ;
    RECT 104.87 65.25 105.08 65.32 ;
    RECT 104.87 65.61 105.08 65.68 ;
    RECT 101.09 64.89 101.3 64.96 ;
    RECT 101.09 65.25 101.3 65.32 ;
    RECT 101.09 65.61 101.3 65.68 ;
    RECT 101.55 64.89 101.76 64.96 ;
    RECT 101.55 65.25 101.76 65.32 ;
    RECT 101.55 65.61 101.76 65.68 ;
    RECT 97.77 64.89 97.98 64.96 ;
    RECT 97.77 65.25 97.98 65.32 ;
    RECT 97.77 65.61 97.98 65.68 ;
    RECT 98.23 64.89 98.44 64.96 ;
    RECT 98.23 65.25 98.44 65.32 ;
    RECT 98.23 65.61 98.44 65.68 ;
    RECT 94.45 64.89 94.66 64.96 ;
    RECT 94.45 65.25 94.66 65.32 ;
    RECT 94.45 65.61 94.66 65.68 ;
    RECT 94.91 64.89 95.12 64.96 ;
    RECT 94.91 65.25 95.12 65.32 ;
    RECT 94.91 65.61 95.12 65.68 ;
    RECT 91.13 64.89 91.34 64.96 ;
    RECT 91.13 65.25 91.34 65.32 ;
    RECT 91.13 65.61 91.34 65.68 ;
    RECT 91.59 64.89 91.8 64.96 ;
    RECT 91.59 65.25 91.8 65.32 ;
    RECT 91.59 65.61 91.8 65.68 ;
    RECT 87.81 64.89 88.02 64.96 ;
    RECT 87.81 65.25 88.02 65.32 ;
    RECT 87.81 65.61 88.02 65.68 ;
    RECT 88.27 64.89 88.48 64.96 ;
    RECT 88.27 65.25 88.48 65.32 ;
    RECT 88.27 65.61 88.48 65.68 ;
    RECT 84.49 64.89 84.7 64.96 ;
    RECT 84.49 65.25 84.7 65.32 ;
    RECT 84.49 65.61 84.7 65.68 ;
    RECT 84.95 64.89 85.16 64.96 ;
    RECT 84.95 65.25 85.16 65.32 ;
    RECT 84.95 65.61 85.16 65.68 ;
    RECT 81.17 64.89 81.38 64.96 ;
    RECT 81.17 65.25 81.38 65.32 ;
    RECT 81.17 65.61 81.38 65.68 ;
    RECT 81.63 64.89 81.84 64.96 ;
    RECT 81.63 65.25 81.84 65.32 ;
    RECT 81.63 65.61 81.84 65.68 ;
    RECT 77.85 64.89 78.06 64.96 ;
    RECT 77.85 65.25 78.06 65.32 ;
    RECT 77.85 65.61 78.06 65.68 ;
    RECT 78.31 64.89 78.52 64.96 ;
    RECT 78.31 65.25 78.52 65.32 ;
    RECT 78.31 65.61 78.52 65.68 ;
    RECT 74.53 64.89 74.74 64.96 ;
    RECT 74.53 65.25 74.74 65.32 ;
    RECT 74.53 65.61 74.74 65.68 ;
    RECT 74.99 64.89 75.2 64.96 ;
    RECT 74.99 65.25 75.2 65.32 ;
    RECT 74.99 65.61 75.2 65.68 ;
    RECT 71.21 64.89 71.42 64.96 ;
    RECT 71.21 65.25 71.42 65.32 ;
    RECT 71.21 65.61 71.42 65.68 ;
    RECT 71.67 64.89 71.88 64.96 ;
    RECT 71.67 65.25 71.88 65.32 ;
    RECT 71.67 65.61 71.88 65.68 ;
    RECT 31.37 64.89 31.58 64.96 ;
    RECT 31.37 65.25 31.58 65.32 ;
    RECT 31.37 65.61 31.58 65.68 ;
    RECT 31.83 64.89 32.04 64.96 ;
    RECT 31.83 65.25 32.04 65.32 ;
    RECT 31.83 65.61 32.04 65.68 ;
    RECT 67.89 64.89 68.1 64.96 ;
    RECT 67.89 65.25 68.1 65.32 ;
    RECT 67.89 65.61 68.1 65.68 ;
    RECT 68.35 64.89 68.56 64.96 ;
    RECT 68.35 65.25 68.56 65.32 ;
    RECT 68.35 65.61 68.56 65.68 ;
    RECT 28.05 64.89 28.26 64.96 ;
    RECT 28.05 65.25 28.26 65.32 ;
    RECT 28.05 65.61 28.26 65.68 ;
    RECT 28.51 64.89 28.72 64.96 ;
    RECT 28.51 65.25 28.72 65.32 ;
    RECT 28.51 65.61 28.72 65.68 ;
    RECT 24.73 64.89 24.94 64.96 ;
    RECT 24.73 65.25 24.94 65.32 ;
    RECT 24.73 65.61 24.94 65.68 ;
    RECT 25.19 64.89 25.4 64.96 ;
    RECT 25.19 65.25 25.4 65.32 ;
    RECT 25.19 65.61 25.4 65.68 ;
    RECT 21.41 64.89 21.62 64.96 ;
    RECT 21.41 65.25 21.62 65.32 ;
    RECT 21.41 65.61 21.62 65.68 ;
    RECT 21.87 64.89 22.08 64.96 ;
    RECT 21.87 65.25 22.08 65.32 ;
    RECT 21.87 65.61 22.08 65.68 ;
    RECT 18.09 64.89 18.3 64.96 ;
    RECT 18.09 65.25 18.3 65.32 ;
    RECT 18.09 65.61 18.3 65.68 ;
    RECT 18.55 64.89 18.76 64.96 ;
    RECT 18.55 65.25 18.76 65.32 ;
    RECT 18.55 65.61 18.76 65.68 ;
    RECT 120.825 65.25 120.895 65.32 ;
    RECT 14.77 64.89 14.98 64.96 ;
    RECT 14.77 65.25 14.98 65.32 ;
    RECT 14.77 65.61 14.98 65.68 ;
    RECT 15.23 64.89 15.44 64.96 ;
    RECT 15.23 65.25 15.44 65.32 ;
    RECT 15.23 65.61 15.44 65.68 ;
    RECT 11.45 64.89 11.66 64.96 ;
    RECT 11.45 65.25 11.66 65.32 ;
    RECT 11.45 65.61 11.66 65.68 ;
    RECT 11.91 64.89 12.12 64.96 ;
    RECT 11.91 65.25 12.12 65.32 ;
    RECT 11.91 65.61 12.12 65.68 ;
    RECT 8.13 64.89 8.34 64.96 ;
    RECT 8.13 65.25 8.34 65.32 ;
    RECT 8.13 65.61 8.34 65.68 ;
    RECT 8.59 64.89 8.8 64.96 ;
    RECT 8.59 65.25 8.8 65.32 ;
    RECT 8.59 65.61 8.8 65.68 ;
    RECT 4.81 64.89 5.02 64.96 ;
    RECT 4.81 65.25 5.02 65.32 ;
    RECT 4.81 65.61 5.02 65.68 ;
    RECT 5.27 64.89 5.48 64.96 ;
    RECT 5.27 65.25 5.48 65.32 ;
    RECT 5.27 65.61 5.48 65.68 ;
    RECT 1.49 64.89 1.7 64.96 ;
    RECT 1.49 65.25 1.7 65.32 ;
    RECT 1.49 65.61 1.7 65.68 ;
    RECT 1.95 64.89 2.16 64.96 ;
    RECT 1.95 65.25 2.16 65.32 ;
    RECT 1.95 65.61 2.16 65.68 ;
    RECT 64.57 64.89 64.78 64.96 ;
    RECT 64.57 65.25 64.78 65.32 ;
    RECT 64.57 65.61 64.78 65.68 ;
    RECT 65.03 64.89 65.24 64.96 ;
    RECT 65.03 65.25 65.24 65.32 ;
    RECT 65.03 65.61 65.24 65.68 ;
    RECT 61.25 56.23 61.46 56.3 ;
    RECT 61.25 56.59 61.46 56.66 ;
    RECT 61.25 56.95 61.46 57.02 ;
    RECT 61.71 56.23 61.92 56.3 ;
    RECT 61.71 56.59 61.92 56.66 ;
    RECT 61.71 56.95 61.92 57.02 ;
    RECT 57.93 56.23 58.14 56.3 ;
    RECT 57.93 56.59 58.14 56.66 ;
    RECT 57.93 56.95 58.14 57.02 ;
    RECT 58.39 56.23 58.6 56.3 ;
    RECT 58.39 56.59 58.6 56.66 ;
    RECT 58.39 56.95 58.6 57.02 ;
    RECT 54.61 56.23 54.82 56.3 ;
    RECT 54.61 56.59 54.82 56.66 ;
    RECT 54.61 56.95 54.82 57.02 ;
    RECT 55.07 56.23 55.28 56.3 ;
    RECT 55.07 56.59 55.28 56.66 ;
    RECT 55.07 56.95 55.28 57.02 ;
    RECT 51.29 56.23 51.5 56.3 ;
    RECT 51.29 56.59 51.5 56.66 ;
    RECT 51.29 56.95 51.5 57.02 ;
    RECT 51.75 56.23 51.96 56.3 ;
    RECT 51.75 56.59 51.96 56.66 ;
    RECT 51.75 56.95 51.96 57.02 ;
    RECT 47.97 56.23 48.18 56.3 ;
    RECT 47.97 56.59 48.18 56.66 ;
    RECT 47.97 56.95 48.18 57.02 ;
    RECT 48.43 56.23 48.64 56.3 ;
    RECT 48.43 56.59 48.64 56.66 ;
    RECT 48.43 56.95 48.64 57.02 ;
    RECT 44.65 56.23 44.86 56.3 ;
    RECT 44.65 56.59 44.86 56.66 ;
    RECT 44.65 56.95 44.86 57.02 ;
    RECT 45.11 56.23 45.32 56.3 ;
    RECT 45.11 56.59 45.32 56.66 ;
    RECT 45.11 56.95 45.32 57.02 ;
    RECT 41.33 56.23 41.54 56.3 ;
    RECT 41.33 56.59 41.54 56.66 ;
    RECT 41.33 56.95 41.54 57.02 ;
    RECT 41.79 56.23 42.0 56.3 ;
    RECT 41.79 56.59 42.0 56.66 ;
    RECT 41.79 56.95 42.0 57.02 ;
    RECT 38.01 56.23 38.22 56.3 ;
    RECT 38.01 56.59 38.22 56.66 ;
    RECT 38.01 56.95 38.22 57.02 ;
    RECT 38.47 56.23 38.68 56.3 ;
    RECT 38.47 56.59 38.68 56.66 ;
    RECT 38.47 56.95 38.68 57.02 ;
    RECT 34.69 56.23 34.9 56.3 ;
    RECT 34.69 56.59 34.9 56.66 ;
    RECT 34.69 56.95 34.9 57.02 ;
    RECT 35.15 56.23 35.36 56.3 ;
    RECT 35.15 56.59 35.36 56.66 ;
    RECT 35.15 56.95 35.36 57.02 ;
    RECT 117.69 56.23 117.9 56.3 ;
    RECT 117.69 56.59 117.9 56.66 ;
    RECT 117.69 56.95 117.9 57.02 ;
    RECT 118.15 56.23 118.36 56.3 ;
    RECT 118.15 56.59 118.36 56.66 ;
    RECT 118.15 56.95 118.36 57.02 ;
    RECT 114.37 56.23 114.58 56.3 ;
    RECT 114.37 56.59 114.58 56.66 ;
    RECT 114.37 56.95 114.58 57.02 ;
    RECT 114.83 56.23 115.04 56.3 ;
    RECT 114.83 56.59 115.04 56.66 ;
    RECT 114.83 56.95 115.04 57.02 ;
    RECT 111.05 56.23 111.26 56.3 ;
    RECT 111.05 56.59 111.26 56.66 ;
    RECT 111.05 56.95 111.26 57.02 ;
    RECT 111.51 56.23 111.72 56.3 ;
    RECT 111.51 56.59 111.72 56.66 ;
    RECT 111.51 56.95 111.72 57.02 ;
    RECT 107.73 56.23 107.94 56.3 ;
    RECT 107.73 56.59 107.94 56.66 ;
    RECT 107.73 56.95 107.94 57.02 ;
    RECT 108.19 56.23 108.4 56.3 ;
    RECT 108.19 56.59 108.4 56.66 ;
    RECT 108.19 56.95 108.4 57.02 ;
    RECT 104.41 56.23 104.62 56.3 ;
    RECT 104.41 56.59 104.62 56.66 ;
    RECT 104.41 56.95 104.62 57.02 ;
    RECT 104.87 56.23 105.08 56.3 ;
    RECT 104.87 56.59 105.08 56.66 ;
    RECT 104.87 56.95 105.08 57.02 ;
    RECT 101.09 56.23 101.3 56.3 ;
    RECT 101.09 56.59 101.3 56.66 ;
    RECT 101.09 56.95 101.3 57.02 ;
    RECT 101.55 56.23 101.76 56.3 ;
    RECT 101.55 56.59 101.76 56.66 ;
    RECT 101.55 56.95 101.76 57.02 ;
    RECT 120.825 56.59 120.895 56.66 ;
    RECT 97.77 56.23 97.98 56.3 ;
    RECT 97.77 56.59 97.98 56.66 ;
    RECT 97.77 56.95 97.98 57.02 ;
    RECT 98.23 56.23 98.44 56.3 ;
    RECT 98.23 56.59 98.44 56.66 ;
    RECT 98.23 56.95 98.44 57.02 ;
    RECT 94.45 56.23 94.66 56.3 ;
    RECT 94.45 56.59 94.66 56.66 ;
    RECT 94.45 56.95 94.66 57.02 ;
    RECT 94.91 56.23 95.12 56.3 ;
    RECT 94.91 56.59 95.12 56.66 ;
    RECT 94.91 56.95 95.12 57.02 ;
    RECT 91.13 56.23 91.34 56.3 ;
    RECT 91.13 56.59 91.34 56.66 ;
    RECT 91.13 56.95 91.34 57.02 ;
    RECT 91.59 56.23 91.8 56.3 ;
    RECT 91.59 56.59 91.8 56.66 ;
    RECT 91.59 56.95 91.8 57.02 ;
    RECT 87.81 56.23 88.02 56.3 ;
    RECT 87.81 56.59 88.02 56.66 ;
    RECT 87.81 56.95 88.02 57.02 ;
    RECT 88.27 56.23 88.48 56.3 ;
    RECT 88.27 56.59 88.48 56.66 ;
    RECT 88.27 56.95 88.48 57.02 ;
    RECT 84.49 56.23 84.7 56.3 ;
    RECT 84.49 56.59 84.7 56.66 ;
    RECT 84.49 56.95 84.7 57.02 ;
    RECT 84.95 56.23 85.16 56.3 ;
    RECT 84.95 56.59 85.16 56.66 ;
    RECT 84.95 56.95 85.16 57.02 ;
    RECT 81.17 56.23 81.38 56.3 ;
    RECT 81.17 56.59 81.38 56.66 ;
    RECT 81.17 56.95 81.38 57.02 ;
    RECT 81.63 56.23 81.84 56.3 ;
    RECT 81.63 56.59 81.84 56.66 ;
    RECT 81.63 56.95 81.84 57.02 ;
    RECT 77.85 56.23 78.06 56.3 ;
    RECT 77.85 56.59 78.06 56.66 ;
    RECT 77.85 56.95 78.06 57.02 ;
    RECT 78.31 56.23 78.52 56.3 ;
    RECT 78.31 56.59 78.52 56.66 ;
    RECT 78.31 56.95 78.52 57.02 ;
    RECT 74.53 56.23 74.74 56.3 ;
    RECT 74.53 56.59 74.74 56.66 ;
    RECT 74.53 56.95 74.74 57.02 ;
    RECT 74.99 56.23 75.2 56.3 ;
    RECT 74.99 56.59 75.2 56.66 ;
    RECT 74.99 56.95 75.2 57.02 ;
    RECT 71.21 56.23 71.42 56.3 ;
    RECT 71.21 56.59 71.42 56.66 ;
    RECT 71.21 56.95 71.42 57.02 ;
    RECT 71.67 56.23 71.88 56.3 ;
    RECT 71.67 56.59 71.88 56.66 ;
    RECT 71.67 56.95 71.88 57.02 ;
    RECT 0.4 56.59 0.47 56.66 ;
    RECT 31.37 56.23 31.58 56.3 ;
    RECT 31.37 56.59 31.58 56.66 ;
    RECT 31.37 56.95 31.58 57.02 ;
    RECT 31.83 56.23 32.04 56.3 ;
    RECT 31.83 56.59 32.04 56.66 ;
    RECT 31.83 56.95 32.04 57.02 ;
    RECT 67.89 56.23 68.1 56.3 ;
    RECT 67.89 56.59 68.1 56.66 ;
    RECT 67.89 56.95 68.1 57.02 ;
    RECT 68.35 56.23 68.56 56.3 ;
    RECT 68.35 56.59 68.56 56.66 ;
    RECT 68.35 56.95 68.56 57.02 ;
    RECT 28.05 56.23 28.26 56.3 ;
    RECT 28.05 56.59 28.26 56.66 ;
    RECT 28.05 56.95 28.26 57.02 ;
    RECT 28.51 56.23 28.72 56.3 ;
    RECT 28.51 56.59 28.72 56.66 ;
    RECT 28.51 56.95 28.72 57.02 ;
    RECT 24.73 56.23 24.94 56.3 ;
    RECT 24.73 56.59 24.94 56.66 ;
    RECT 24.73 56.95 24.94 57.02 ;
    RECT 25.19 56.23 25.4 56.3 ;
    RECT 25.19 56.59 25.4 56.66 ;
    RECT 25.19 56.95 25.4 57.02 ;
    RECT 21.41 56.23 21.62 56.3 ;
    RECT 21.41 56.59 21.62 56.66 ;
    RECT 21.41 56.95 21.62 57.02 ;
    RECT 21.87 56.23 22.08 56.3 ;
    RECT 21.87 56.59 22.08 56.66 ;
    RECT 21.87 56.95 22.08 57.02 ;
    RECT 18.09 56.23 18.3 56.3 ;
    RECT 18.09 56.59 18.3 56.66 ;
    RECT 18.09 56.95 18.3 57.02 ;
    RECT 18.55 56.23 18.76 56.3 ;
    RECT 18.55 56.59 18.76 56.66 ;
    RECT 18.55 56.95 18.76 57.02 ;
    RECT 14.77 56.23 14.98 56.3 ;
    RECT 14.77 56.59 14.98 56.66 ;
    RECT 14.77 56.95 14.98 57.02 ;
    RECT 15.23 56.23 15.44 56.3 ;
    RECT 15.23 56.59 15.44 56.66 ;
    RECT 15.23 56.95 15.44 57.02 ;
    RECT 11.45 56.23 11.66 56.3 ;
    RECT 11.45 56.59 11.66 56.66 ;
    RECT 11.45 56.95 11.66 57.02 ;
    RECT 11.91 56.23 12.12 56.3 ;
    RECT 11.91 56.59 12.12 56.66 ;
    RECT 11.91 56.95 12.12 57.02 ;
    RECT 8.13 56.23 8.34 56.3 ;
    RECT 8.13 56.59 8.34 56.66 ;
    RECT 8.13 56.95 8.34 57.02 ;
    RECT 8.59 56.23 8.8 56.3 ;
    RECT 8.59 56.59 8.8 56.66 ;
    RECT 8.59 56.95 8.8 57.02 ;
    RECT 4.81 56.23 5.02 56.3 ;
    RECT 4.81 56.59 5.02 56.66 ;
    RECT 4.81 56.95 5.02 57.02 ;
    RECT 5.27 56.23 5.48 56.3 ;
    RECT 5.27 56.59 5.48 56.66 ;
    RECT 5.27 56.95 5.48 57.02 ;
    RECT 1.49 56.23 1.7 56.3 ;
    RECT 1.49 56.59 1.7 56.66 ;
    RECT 1.49 56.95 1.7 57.02 ;
    RECT 1.95 56.23 2.16 56.3 ;
    RECT 1.95 56.59 2.16 56.66 ;
    RECT 1.95 56.95 2.16 57.02 ;
    RECT 64.57 56.23 64.78 56.3 ;
    RECT 64.57 56.59 64.78 56.66 ;
    RECT 64.57 56.95 64.78 57.02 ;
    RECT 65.03 56.23 65.24 56.3 ;
    RECT 65.03 56.59 65.24 56.66 ;
    RECT 65.03 56.95 65.24 57.02 ;
    RECT 61.25 24.55 61.46 24.62 ;
    RECT 61.25 24.91 61.46 24.98 ;
    RECT 61.25 25.27 61.46 25.34 ;
    RECT 61.71 24.55 61.92 24.62 ;
    RECT 61.71 24.91 61.92 24.98 ;
    RECT 61.71 25.27 61.92 25.34 ;
    RECT 57.93 24.55 58.14 24.62 ;
    RECT 57.93 24.91 58.14 24.98 ;
    RECT 57.93 25.27 58.14 25.34 ;
    RECT 58.39 24.55 58.6 24.62 ;
    RECT 58.39 24.91 58.6 24.98 ;
    RECT 58.39 25.27 58.6 25.34 ;
    RECT 54.61 24.55 54.82 24.62 ;
    RECT 54.61 24.91 54.82 24.98 ;
    RECT 54.61 25.27 54.82 25.34 ;
    RECT 55.07 24.55 55.28 24.62 ;
    RECT 55.07 24.91 55.28 24.98 ;
    RECT 55.07 25.27 55.28 25.34 ;
    RECT 51.29 24.55 51.5 24.62 ;
    RECT 51.29 24.91 51.5 24.98 ;
    RECT 51.29 25.27 51.5 25.34 ;
    RECT 51.75 24.55 51.96 24.62 ;
    RECT 51.75 24.91 51.96 24.98 ;
    RECT 51.75 25.27 51.96 25.34 ;
    RECT 47.97 24.55 48.18 24.62 ;
    RECT 47.97 24.91 48.18 24.98 ;
    RECT 47.97 25.27 48.18 25.34 ;
    RECT 48.43 24.55 48.64 24.62 ;
    RECT 48.43 24.91 48.64 24.98 ;
    RECT 48.43 25.27 48.64 25.34 ;
    RECT 44.65 24.55 44.86 24.62 ;
    RECT 44.65 24.91 44.86 24.98 ;
    RECT 44.65 25.27 44.86 25.34 ;
    RECT 45.11 24.55 45.32 24.62 ;
    RECT 45.11 24.91 45.32 24.98 ;
    RECT 45.11 25.27 45.32 25.34 ;
    RECT 41.33 24.55 41.54 24.62 ;
    RECT 41.33 24.91 41.54 24.98 ;
    RECT 41.33 25.27 41.54 25.34 ;
    RECT 41.79 24.55 42.0 24.62 ;
    RECT 41.79 24.91 42.0 24.98 ;
    RECT 41.79 25.27 42.0 25.34 ;
    RECT 38.01 24.55 38.22 24.62 ;
    RECT 38.01 24.91 38.22 24.98 ;
    RECT 38.01 25.27 38.22 25.34 ;
    RECT 38.47 24.55 38.68 24.62 ;
    RECT 38.47 24.91 38.68 24.98 ;
    RECT 38.47 25.27 38.68 25.34 ;
    RECT 0.4 24.91 0.47 24.98 ;
    RECT 34.69 24.55 34.9 24.62 ;
    RECT 34.69 24.91 34.9 24.98 ;
    RECT 34.69 25.27 34.9 25.34 ;
    RECT 35.15 24.55 35.36 24.62 ;
    RECT 35.15 24.91 35.36 24.98 ;
    RECT 35.15 25.27 35.36 25.34 ;
    RECT 117.69 24.55 117.9 24.62 ;
    RECT 117.69 24.91 117.9 24.98 ;
    RECT 117.69 25.27 117.9 25.34 ;
    RECT 118.15 24.55 118.36 24.62 ;
    RECT 118.15 24.91 118.36 24.98 ;
    RECT 118.15 25.27 118.36 25.34 ;
    RECT 114.37 24.55 114.58 24.62 ;
    RECT 114.37 24.91 114.58 24.98 ;
    RECT 114.37 25.27 114.58 25.34 ;
    RECT 114.83 24.55 115.04 24.62 ;
    RECT 114.83 24.91 115.04 24.98 ;
    RECT 114.83 25.27 115.04 25.34 ;
    RECT 111.05 24.55 111.26 24.62 ;
    RECT 111.05 24.91 111.26 24.98 ;
    RECT 111.05 25.27 111.26 25.34 ;
    RECT 111.51 24.55 111.72 24.62 ;
    RECT 111.51 24.91 111.72 24.98 ;
    RECT 111.51 25.27 111.72 25.34 ;
    RECT 107.73 24.55 107.94 24.62 ;
    RECT 107.73 24.91 107.94 24.98 ;
    RECT 107.73 25.27 107.94 25.34 ;
    RECT 108.19 24.55 108.4 24.62 ;
    RECT 108.19 24.91 108.4 24.98 ;
    RECT 108.19 25.27 108.4 25.34 ;
    RECT 104.41 24.55 104.62 24.62 ;
    RECT 104.41 24.91 104.62 24.98 ;
    RECT 104.41 25.27 104.62 25.34 ;
    RECT 104.87 24.55 105.08 24.62 ;
    RECT 104.87 24.91 105.08 24.98 ;
    RECT 104.87 25.27 105.08 25.34 ;
    RECT 101.09 24.55 101.3 24.62 ;
    RECT 101.09 24.91 101.3 24.98 ;
    RECT 101.09 25.27 101.3 25.34 ;
    RECT 101.55 24.55 101.76 24.62 ;
    RECT 101.55 24.91 101.76 24.98 ;
    RECT 101.55 25.27 101.76 25.34 ;
    RECT 97.77 24.55 97.98 24.62 ;
    RECT 97.77 24.91 97.98 24.98 ;
    RECT 97.77 25.27 97.98 25.34 ;
    RECT 98.23 24.55 98.44 24.62 ;
    RECT 98.23 24.91 98.44 24.98 ;
    RECT 98.23 25.27 98.44 25.34 ;
    RECT 94.45 24.55 94.66 24.62 ;
    RECT 94.45 24.91 94.66 24.98 ;
    RECT 94.45 25.27 94.66 25.34 ;
    RECT 94.91 24.55 95.12 24.62 ;
    RECT 94.91 24.91 95.12 24.98 ;
    RECT 94.91 25.27 95.12 25.34 ;
    RECT 91.13 24.55 91.34 24.62 ;
    RECT 91.13 24.91 91.34 24.98 ;
    RECT 91.13 25.27 91.34 25.34 ;
    RECT 91.59 24.55 91.8 24.62 ;
    RECT 91.59 24.91 91.8 24.98 ;
    RECT 91.59 25.27 91.8 25.34 ;
    RECT 87.81 24.55 88.02 24.62 ;
    RECT 87.81 24.91 88.02 24.98 ;
    RECT 87.81 25.27 88.02 25.34 ;
    RECT 88.27 24.55 88.48 24.62 ;
    RECT 88.27 24.91 88.48 24.98 ;
    RECT 88.27 25.27 88.48 25.34 ;
    RECT 84.49 24.55 84.7 24.62 ;
    RECT 84.49 24.91 84.7 24.98 ;
    RECT 84.49 25.27 84.7 25.34 ;
    RECT 84.95 24.55 85.16 24.62 ;
    RECT 84.95 24.91 85.16 24.98 ;
    RECT 84.95 25.27 85.16 25.34 ;
    RECT 81.17 24.55 81.38 24.62 ;
    RECT 81.17 24.91 81.38 24.98 ;
    RECT 81.17 25.27 81.38 25.34 ;
    RECT 81.63 24.55 81.84 24.62 ;
    RECT 81.63 24.91 81.84 24.98 ;
    RECT 81.63 25.27 81.84 25.34 ;
    RECT 77.85 24.55 78.06 24.62 ;
    RECT 77.85 24.91 78.06 24.98 ;
    RECT 77.85 25.27 78.06 25.34 ;
    RECT 78.31 24.55 78.52 24.62 ;
    RECT 78.31 24.91 78.52 24.98 ;
    RECT 78.31 25.27 78.52 25.34 ;
    RECT 74.53 24.55 74.74 24.62 ;
    RECT 74.53 24.91 74.74 24.98 ;
    RECT 74.53 25.27 74.74 25.34 ;
    RECT 74.99 24.55 75.2 24.62 ;
    RECT 74.99 24.91 75.2 24.98 ;
    RECT 74.99 25.27 75.2 25.34 ;
    RECT 71.21 24.55 71.42 24.62 ;
    RECT 71.21 24.91 71.42 24.98 ;
    RECT 71.21 25.27 71.42 25.34 ;
    RECT 71.67 24.55 71.88 24.62 ;
    RECT 71.67 24.91 71.88 24.98 ;
    RECT 71.67 25.27 71.88 25.34 ;
    RECT 31.37 24.55 31.58 24.62 ;
    RECT 31.37 24.91 31.58 24.98 ;
    RECT 31.37 25.27 31.58 25.34 ;
    RECT 31.83 24.55 32.04 24.62 ;
    RECT 31.83 24.91 32.04 24.98 ;
    RECT 31.83 25.27 32.04 25.34 ;
    RECT 67.89 24.55 68.1 24.62 ;
    RECT 67.89 24.91 68.1 24.98 ;
    RECT 67.89 25.27 68.1 25.34 ;
    RECT 68.35 24.55 68.56 24.62 ;
    RECT 68.35 24.91 68.56 24.98 ;
    RECT 68.35 25.27 68.56 25.34 ;
    RECT 28.05 24.55 28.26 24.62 ;
    RECT 28.05 24.91 28.26 24.98 ;
    RECT 28.05 25.27 28.26 25.34 ;
    RECT 28.51 24.55 28.72 24.62 ;
    RECT 28.51 24.91 28.72 24.98 ;
    RECT 28.51 25.27 28.72 25.34 ;
    RECT 24.73 24.55 24.94 24.62 ;
    RECT 24.73 24.91 24.94 24.98 ;
    RECT 24.73 25.27 24.94 25.34 ;
    RECT 25.19 24.55 25.4 24.62 ;
    RECT 25.19 24.91 25.4 24.98 ;
    RECT 25.19 25.27 25.4 25.34 ;
    RECT 21.41 24.55 21.62 24.62 ;
    RECT 21.41 24.91 21.62 24.98 ;
    RECT 21.41 25.27 21.62 25.34 ;
    RECT 21.87 24.55 22.08 24.62 ;
    RECT 21.87 24.91 22.08 24.98 ;
    RECT 21.87 25.27 22.08 25.34 ;
    RECT 18.09 24.55 18.3 24.62 ;
    RECT 18.09 24.91 18.3 24.98 ;
    RECT 18.09 25.27 18.3 25.34 ;
    RECT 18.55 24.55 18.76 24.62 ;
    RECT 18.55 24.91 18.76 24.98 ;
    RECT 18.55 25.27 18.76 25.34 ;
    RECT 120.825 24.91 120.895 24.98 ;
    RECT 14.77 24.55 14.98 24.62 ;
    RECT 14.77 24.91 14.98 24.98 ;
    RECT 14.77 25.27 14.98 25.34 ;
    RECT 15.23 24.55 15.44 24.62 ;
    RECT 15.23 24.91 15.44 24.98 ;
    RECT 15.23 25.27 15.44 25.34 ;
    RECT 11.45 24.55 11.66 24.62 ;
    RECT 11.45 24.91 11.66 24.98 ;
    RECT 11.45 25.27 11.66 25.34 ;
    RECT 11.91 24.55 12.12 24.62 ;
    RECT 11.91 24.91 12.12 24.98 ;
    RECT 11.91 25.27 12.12 25.34 ;
    RECT 8.13 24.55 8.34 24.62 ;
    RECT 8.13 24.91 8.34 24.98 ;
    RECT 8.13 25.27 8.34 25.34 ;
    RECT 8.59 24.55 8.8 24.62 ;
    RECT 8.59 24.91 8.8 24.98 ;
    RECT 8.59 25.27 8.8 25.34 ;
    RECT 4.81 24.55 5.02 24.62 ;
    RECT 4.81 24.91 5.02 24.98 ;
    RECT 4.81 25.27 5.02 25.34 ;
    RECT 5.27 24.55 5.48 24.62 ;
    RECT 5.27 24.91 5.48 24.98 ;
    RECT 5.27 25.27 5.48 25.34 ;
    RECT 1.49 24.55 1.7 24.62 ;
    RECT 1.49 24.91 1.7 24.98 ;
    RECT 1.49 25.27 1.7 25.34 ;
    RECT 1.95 24.55 2.16 24.62 ;
    RECT 1.95 24.91 2.16 24.98 ;
    RECT 1.95 25.27 2.16 25.34 ;
    RECT 64.57 24.55 64.78 24.62 ;
    RECT 64.57 24.91 64.78 24.98 ;
    RECT 64.57 25.27 64.78 25.34 ;
    RECT 65.03 24.55 65.24 24.62 ;
    RECT 65.03 24.91 65.24 24.98 ;
    RECT 65.03 25.27 65.24 25.34 ;
    RECT 61.25 64.17 61.46 64.24 ;
    RECT 61.25 64.53 61.46 64.6 ;
    RECT 61.25 64.89 61.46 64.96 ;
    RECT 61.71 64.17 61.92 64.24 ;
    RECT 61.71 64.53 61.92 64.6 ;
    RECT 61.71 64.89 61.92 64.96 ;
    RECT 57.93 64.17 58.14 64.24 ;
    RECT 57.93 64.53 58.14 64.6 ;
    RECT 57.93 64.89 58.14 64.96 ;
    RECT 58.39 64.17 58.6 64.24 ;
    RECT 58.39 64.53 58.6 64.6 ;
    RECT 58.39 64.89 58.6 64.96 ;
    RECT 54.61 64.17 54.82 64.24 ;
    RECT 54.61 64.53 54.82 64.6 ;
    RECT 54.61 64.89 54.82 64.96 ;
    RECT 55.07 64.17 55.28 64.24 ;
    RECT 55.07 64.53 55.28 64.6 ;
    RECT 55.07 64.89 55.28 64.96 ;
    RECT 51.29 64.17 51.5 64.24 ;
    RECT 51.29 64.53 51.5 64.6 ;
    RECT 51.29 64.89 51.5 64.96 ;
    RECT 51.75 64.17 51.96 64.24 ;
    RECT 51.75 64.53 51.96 64.6 ;
    RECT 51.75 64.89 51.96 64.96 ;
    RECT 47.97 64.17 48.18 64.24 ;
    RECT 47.97 64.53 48.18 64.6 ;
    RECT 47.97 64.89 48.18 64.96 ;
    RECT 48.43 64.17 48.64 64.24 ;
    RECT 48.43 64.53 48.64 64.6 ;
    RECT 48.43 64.89 48.64 64.96 ;
    RECT 44.65 64.17 44.86 64.24 ;
    RECT 44.65 64.53 44.86 64.6 ;
    RECT 44.65 64.89 44.86 64.96 ;
    RECT 45.11 64.17 45.32 64.24 ;
    RECT 45.11 64.53 45.32 64.6 ;
    RECT 45.11 64.89 45.32 64.96 ;
    RECT 41.33 64.17 41.54 64.24 ;
    RECT 41.33 64.53 41.54 64.6 ;
    RECT 41.33 64.89 41.54 64.96 ;
    RECT 41.79 64.17 42.0 64.24 ;
    RECT 41.79 64.53 42.0 64.6 ;
    RECT 41.79 64.89 42.0 64.96 ;
    RECT 38.01 64.17 38.22 64.24 ;
    RECT 38.01 64.53 38.22 64.6 ;
    RECT 38.01 64.89 38.22 64.96 ;
    RECT 38.47 64.17 38.68 64.24 ;
    RECT 38.47 64.53 38.68 64.6 ;
    RECT 38.47 64.89 38.68 64.96 ;
    RECT 0.4 64.53 0.47 64.6 ;
    RECT 34.69 64.17 34.9 64.24 ;
    RECT 34.69 64.53 34.9 64.6 ;
    RECT 34.69 64.89 34.9 64.96 ;
    RECT 35.15 64.17 35.36 64.24 ;
    RECT 35.15 64.53 35.36 64.6 ;
    RECT 35.15 64.89 35.36 64.96 ;
    RECT 117.69 64.17 117.9 64.24 ;
    RECT 117.69 64.53 117.9 64.6 ;
    RECT 117.69 64.89 117.9 64.96 ;
    RECT 118.15 64.17 118.36 64.24 ;
    RECT 118.15 64.53 118.36 64.6 ;
    RECT 118.15 64.89 118.36 64.96 ;
    RECT 114.37 64.17 114.58 64.24 ;
    RECT 114.37 64.53 114.58 64.6 ;
    RECT 114.37 64.89 114.58 64.96 ;
    RECT 114.83 64.17 115.04 64.24 ;
    RECT 114.83 64.53 115.04 64.6 ;
    RECT 114.83 64.89 115.04 64.96 ;
    RECT 111.05 64.17 111.26 64.24 ;
    RECT 111.05 64.53 111.26 64.6 ;
    RECT 111.05 64.89 111.26 64.96 ;
    RECT 111.51 64.17 111.72 64.24 ;
    RECT 111.51 64.53 111.72 64.6 ;
    RECT 111.51 64.89 111.72 64.96 ;
    RECT 107.73 64.17 107.94 64.24 ;
    RECT 107.73 64.53 107.94 64.6 ;
    RECT 107.73 64.89 107.94 64.96 ;
    RECT 108.19 64.17 108.4 64.24 ;
    RECT 108.19 64.53 108.4 64.6 ;
    RECT 108.19 64.89 108.4 64.96 ;
    RECT 104.41 64.17 104.62 64.24 ;
    RECT 104.41 64.53 104.62 64.6 ;
    RECT 104.41 64.89 104.62 64.96 ;
    RECT 104.87 64.17 105.08 64.24 ;
    RECT 104.87 64.53 105.08 64.6 ;
    RECT 104.87 64.89 105.08 64.96 ;
    RECT 101.09 64.17 101.3 64.24 ;
    RECT 101.09 64.53 101.3 64.6 ;
    RECT 101.09 64.89 101.3 64.96 ;
    RECT 101.55 64.17 101.76 64.24 ;
    RECT 101.55 64.53 101.76 64.6 ;
    RECT 101.55 64.89 101.76 64.96 ;
    RECT 97.77 64.17 97.98 64.24 ;
    RECT 97.77 64.53 97.98 64.6 ;
    RECT 97.77 64.89 97.98 64.96 ;
    RECT 98.23 64.17 98.44 64.24 ;
    RECT 98.23 64.53 98.44 64.6 ;
    RECT 98.23 64.89 98.44 64.96 ;
    RECT 94.45 64.17 94.66 64.24 ;
    RECT 94.45 64.53 94.66 64.6 ;
    RECT 94.45 64.89 94.66 64.96 ;
    RECT 94.91 64.17 95.12 64.24 ;
    RECT 94.91 64.53 95.12 64.6 ;
    RECT 94.91 64.89 95.12 64.96 ;
    RECT 91.13 64.17 91.34 64.24 ;
    RECT 91.13 64.53 91.34 64.6 ;
    RECT 91.13 64.89 91.34 64.96 ;
    RECT 91.59 64.17 91.8 64.24 ;
    RECT 91.59 64.53 91.8 64.6 ;
    RECT 91.59 64.89 91.8 64.96 ;
    RECT 87.81 64.17 88.02 64.24 ;
    RECT 87.81 64.53 88.02 64.6 ;
    RECT 87.81 64.89 88.02 64.96 ;
    RECT 88.27 64.17 88.48 64.24 ;
    RECT 88.27 64.53 88.48 64.6 ;
    RECT 88.27 64.89 88.48 64.96 ;
    RECT 84.49 64.17 84.7 64.24 ;
    RECT 84.49 64.53 84.7 64.6 ;
    RECT 84.49 64.89 84.7 64.96 ;
    RECT 84.95 64.17 85.16 64.24 ;
    RECT 84.95 64.53 85.16 64.6 ;
    RECT 84.95 64.89 85.16 64.96 ;
    RECT 81.17 64.17 81.38 64.24 ;
    RECT 81.17 64.53 81.38 64.6 ;
    RECT 81.17 64.89 81.38 64.96 ;
    RECT 81.63 64.17 81.84 64.24 ;
    RECT 81.63 64.53 81.84 64.6 ;
    RECT 81.63 64.89 81.84 64.96 ;
    RECT 77.85 64.17 78.06 64.24 ;
    RECT 77.85 64.53 78.06 64.6 ;
    RECT 77.85 64.89 78.06 64.96 ;
    RECT 78.31 64.17 78.52 64.24 ;
    RECT 78.31 64.53 78.52 64.6 ;
    RECT 78.31 64.89 78.52 64.96 ;
    RECT 74.53 64.17 74.74 64.24 ;
    RECT 74.53 64.53 74.74 64.6 ;
    RECT 74.53 64.89 74.74 64.96 ;
    RECT 74.99 64.17 75.2 64.24 ;
    RECT 74.99 64.53 75.2 64.6 ;
    RECT 74.99 64.89 75.2 64.96 ;
    RECT 71.21 64.17 71.42 64.24 ;
    RECT 71.21 64.53 71.42 64.6 ;
    RECT 71.21 64.89 71.42 64.96 ;
    RECT 71.67 64.17 71.88 64.24 ;
    RECT 71.67 64.53 71.88 64.6 ;
    RECT 71.67 64.89 71.88 64.96 ;
    RECT 31.37 64.17 31.58 64.24 ;
    RECT 31.37 64.53 31.58 64.6 ;
    RECT 31.37 64.89 31.58 64.96 ;
    RECT 31.83 64.17 32.04 64.24 ;
    RECT 31.83 64.53 32.04 64.6 ;
    RECT 31.83 64.89 32.04 64.96 ;
    RECT 67.89 64.17 68.1 64.24 ;
    RECT 67.89 64.53 68.1 64.6 ;
    RECT 67.89 64.89 68.1 64.96 ;
    RECT 68.35 64.17 68.56 64.24 ;
    RECT 68.35 64.53 68.56 64.6 ;
    RECT 68.35 64.89 68.56 64.96 ;
    RECT 28.05 64.17 28.26 64.24 ;
    RECT 28.05 64.53 28.26 64.6 ;
    RECT 28.05 64.89 28.26 64.96 ;
    RECT 28.51 64.17 28.72 64.24 ;
    RECT 28.51 64.53 28.72 64.6 ;
    RECT 28.51 64.89 28.72 64.96 ;
    RECT 24.73 64.17 24.94 64.24 ;
    RECT 24.73 64.53 24.94 64.6 ;
    RECT 24.73 64.89 24.94 64.96 ;
    RECT 25.19 64.17 25.4 64.24 ;
    RECT 25.19 64.53 25.4 64.6 ;
    RECT 25.19 64.89 25.4 64.96 ;
    RECT 21.41 64.17 21.62 64.24 ;
    RECT 21.41 64.53 21.62 64.6 ;
    RECT 21.41 64.89 21.62 64.96 ;
    RECT 21.87 64.17 22.08 64.24 ;
    RECT 21.87 64.53 22.08 64.6 ;
    RECT 21.87 64.89 22.08 64.96 ;
    RECT 18.09 64.17 18.3 64.24 ;
    RECT 18.09 64.53 18.3 64.6 ;
    RECT 18.09 64.89 18.3 64.96 ;
    RECT 18.55 64.17 18.76 64.24 ;
    RECT 18.55 64.53 18.76 64.6 ;
    RECT 18.55 64.89 18.76 64.96 ;
    RECT 120.825 64.53 120.895 64.6 ;
    RECT 14.77 64.17 14.98 64.24 ;
    RECT 14.77 64.53 14.98 64.6 ;
    RECT 14.77 64.89 14.98 64.96 ;
    RECT 15.23 64.17 15.44 64.24 ;
    RECT 15.23 64.53 15.44 64.6 ;
    RECT 15.23 64.89 15.44 64.96 ;
    RECT 11.45 64.17 11.66 64.24 ;
    RECT 11.45 64.53 11.66 64.6 ;
    RECT 11.45 64.89 11.66 64.96 ;
    RECT 11.91 64.17 12.12 64.24 ;
    RECT 11.91 64.53 12.12 64.6 ;
    RECT 11.91 64.89 12.12 64.96 ;
    RECT 8.13 64.17 8.34 64.24 ;
    RECT 8.13 64.53 8.34 64.6 ;
    RECT 8.13 64.89 8.34 64.96 ;
    RECT 8.59 64.17 8.8 64.24 ;
    RECT 8.59 64.53 8.8 64.6 ;
    RECT 8.59 64.89 8.8 64.96 ;
    RECT 4.81 64.17 5.02 64.24 ;
    RECT 4.81 64.53 5.02 64.6 ;
    RECT 4.81 64.89 5.02 64.96 ;
    RECT 5.27 64.17 5.48 64.24 ;
    RECT 5.27 64.53 5.48 64.6 ;
    RECT 5.27 64.89 5.48 64.96 ;
    RECT 1.49 64.17 1.7 64.24 ;
    RECT 1.49 64.53 1.7 64.6 ;
    RECT 1.49 64.89 1.7 64.96 ;
    RECT 1.95 64.17 2.16 64.24 ;
    RECT 1.95 64.53 2.16 64.6 ;
    RECT 1.95 64.89 2.16 64.96 ;
    RECT 64.57 64.17 64.78 64.24 ;
    RECT 64.57 64.53 64.78 64.6 ;
    RECT 64.57 64.89 64.78 64.96 ;
    RECT 65.03 64.17 65.24 64.24 ;
    RECT 65.03 64.53 65.24 64.6 ;
    RECT 65.03 64.89 65.24 64.96 ;
    RECT 61.25 23.83 61.46 23.9 ;
    RECT 61.25 24.19 61.46 24.26 ;
    RECT 61.25 24.55 61.46 24.62 ;
    RECT 61.71 23.83 61.92 23.9 ;
    RECT 61.71 24.19 61.92 24.26 ;
    RECT 61.71 24.55 61.92 24.62 ;
    RECT 57.93 23.83 58.14 23.9 ;
    RECT 57.93 24.19 58.14 24.26 ;
    RECT 57.93 24.55 58.14 24.62 ;
    RECT 58.39 23.83 58.6 23.9 ;
    RECT 58.39 24.19 58.6 24.26 ;
    RECT 58.39 24.55 58.6 24.62 ;
    RECT 54.61 23.83 54.82 23.9 ;
    RECT 54.61 24.19 54.82 24.26 ;
    RECT 54.61 24.55 54.82 24.62 ;
    RECT 55.07 23.83 55.28 23.9 ;
    RECT 55.07 24.19 55.28 24.26 ;
    RECT 55.07 24.55 55.28 24.62 ;
    RECT 51.29 23.83 51.5 23.9 ;
    RECT 51.29 24.19 51.5 24.26 ;
    RECT 51.29 24.55 51.5 24.62 ;
    RECT 51.75 23.83 51.96 23.9 ;
    RECT 51.75 24.19 51.96 24.26 ;
    RECT 51.75 24.55 51.96 24.62 ;
    RECT 47.97 23.83 48.18 23.9 ;
    RECT 47.97 24.19 48.18 24.26 ;
    RECT 47.97 24.55 48.18 24.62 ;
    RECT 48.43 23.83 48.64 23.9 ;
    RECT 48.43 24.19 48.64 24.26 ;
    RECT 48.43 24.55 48.64 24.62 ;
    RECT 44.65 23.83 44.86 23.9 ;
    RECT 44.65 24.19 44.86 24.26 ;
    RECT 44.65 24.55 44.86 24.62 ;
    RECT 45.11 23.83 45.32 23.9 ;
    RECT 45.11 24.19 45.32 24.26 ;
    RECT 45.11 24.55 45.32 24.62 ;
    RECT 41.33 23.83 41.54 23.9 ;
    RECT 41.33 24.19 41.54 24.26 ;
    RECT 41.33 24.55 41.54 24.62 ;
    RECT 41.79 23.83 42.0 23.9 ;
    RECT 41.79 24.19 42.0 24.26 ;
    RECT 41.79 24.55 42.0 24.62 ;
    RECT 38.01 23.83 38.22 23.9 ;
    RECT 38.01 24.19 38.22 24.26 ;
    RECT 38.01 24.55 38.22 24.62 ;
    RECT 38.47 23.83 38.68 23.9 ;
    RECT 38.47 24.19 38.68 24.26 ;
    RECT 38.47 24.55 38.68 24.62 ;
    RECT 0.4 24.19 0.47 24.26 ;
    RECT 34.69 23.83 34.9 23.9 ;
    RECT 34.69 24.19 34.9 24.26 ;
    RECT 34.69 24.55 34.9 24.62 ;
    RECT 35.15 23.83 35.36 23.9 ;
    RECT 35.15 24.19 35.36 24.26 ;
    RECT 35.15 24.55 35.36 24.62 ;
    RECT 117.69 23.83 117.9 23.9 ;
    RECT 117.69 24.19 117.9 24.26 ;
    RECT 117.69 24.55 117.9 24.62 ;
    RECT 118.15 23.83 118.36 23.9 ;
    RECT 118.15 24.19 118.36 24.26 ;
    RECT 118.15 24.55 118.36 24.62 ;
    RECT 114.37 23.83 114.58 23.9 ;
    RECT 114.37 24.19 114.58 24.26 ;
    RECT 114.37 24.55 114.58 24.62 ;
    RECT 114.83 23.83 115.04 23.9 ;
    RECT 114.83 24.19 115.04 24.26 ;
    RECT 114.83 24.55 115.04 24.62 ;
    RECT 111.05 23.83 111.26 23.9 ;
    RECT 111.05 24.19 111.26 24.26 ;
    RECT 111.05 24.55 111.26 24.62 ;
    RECT 111.51 23.83 111.72 23.9 ;
    RECT 111.51 24.19 111.72 24.26 ;
    RECT 111.51 24.55 111.72 24.62 ;
    RECT 107.73 23.83 107.94 23.9 ;
    RECT 107.73 24.19 107.94 24.26 ;
    RECT 107.73 24.55 107.94 24.62 ;
    RECT 108.19 23.83 108.4 23.9 ;
    RECT 108.19 24.19 108.4 24.26 ;
    RECT 108.19 24.55 108.4 24.62 ;
    RECT 104.41 23.83 104.62 23.9 ;
    RECT 104.41 24.19 104.62 24.26 ;
    RECT 104.41 24.55 104.62 24.62 ;
    RECT 104.87 23.83 105.08 23.9 ;
    RECT 104.87 24.19 105.08 24.26 ;
    RECT 104.87 24.55 105.08 24.62 ;
    RECT 101.09 23.83 101.3 23.9 ;
    RECT 101.09 24.19 101.3 24.26 ;
    RECT 101.09 24.55 101.3 24.62 ;
    RECT 101.55 23.83 101.76 23.9 ;
    RECT 101.55 24.19 101.76 24.26 ;
    RECT 101.55 24.55 101.76 24.62 ;
    RECT 97.77 23.83 97.98 23.9 ;
    RECT 97.77 24.19 97.98 24.26 ;
    RECT 97.77 24.55 97.98 24.62 ;
    RECT 98.23 23.83 98.44 23.9 ;
    RECT 98.23 24.19 98.44 24.26 ;
    RECT 98.23 24.55 98.44 24.62 ;
    RECT 94.45 23.83 94.66 23.9 ;
    RECT 94.45 24.19 94.66 24.26 ;
    RECT 94.45 24.55 94.66 24.62 ;
    RECT 94.91 23.83 95.12 23.9 ;
    RECT 94.91 24.19 95.12 24.26 ;
    RECT 94.91 24.55 95.12 24.62 ;
    RECT 91.13 23.83 91.34 23.9 ;
    RECT 91.13 24.19 91.34 24.26 ;
    RECT 91.13 24.55 91.34 24.62 ;
    RECT 91.59 23.83 91.8 23.9 ;
    RECT 91.59 24.19 91.8 24.26 ;
    RECT 91.59 24.55 91.8 24.62 ;
    RECT 87.81 23.83 88.02 23.9 ;
    RECT 87.81 24.19 88.02 24.26 ;
    RECT 87.81 24.55 88.02 24.62 ;
    RECT 88.27 23.83 88.48 23.9 ;
    RECT 88.27 24.19 88.48 24.26 ;
    RECT 88.27 24.55 88.48 24.62 ;
    RECT 84.49 23.83 84.7 23.9 ;
    RECT 84.49 24.19 84.7 24.26 ;
    RECT 84.49 24.55 84.7 24.62 ;
    RECT 84.95 23.83 85.16 23.9 ;
    RECT 84.95 24.19 85.16 24.26 ;
    RECT 84.95 24.55 85.16 24.62 ;
    RECT 81.17 23.83 81.38 23.9 ;
    RECT 81.17 24.19 81.38 24.26 ;
    RECT 81.17 24.55 81.38 24.62 ;
    RECT 81.63 23.83 81.84 23.9 ;
    RECT 81.63 24.19 81.84 24.26 ;
    RECT 81.63 24.55 81.84 24.62 ;
    RECT 77.85 23.83 78.06 23.9 ;
    RECT 77.85 24.19 78.06 24.26 ;
    RECT 77.85 24.55 78.06 24.62 ;
    RECT 78.31 23.83 78.52 23.9 ;
    RECT 78.31 24.19 78.52 24.26 ;
    RECT 78.31 24.55 78.52 24.62 ;
    RECT 74.53 23.83 74.74 23.9 ;
    RECT 74.53 24.19 74.74 24.26 ;
    RECT 74.53 24.55 74.74 24.62 ;
    RECT 74.99 23.83 75.2 23.9 ;
    RECT 74.99 24.19 75.2 24.26 ;
    RECT 74.99 24.55 75.2 24.62 ;
    RECT 71.21 23.83 71.42 23.9 ;
    RECT 71.21 24.19 71.42 24.26 ;
    RECT 71.21 24.55 71.42 24.62 ;
    RECT 71.67 23.83 71.88 23.9 ;
    RECT 71.67 24.19 71.88 24.26 ;
    RECT 71.67 24.55 71.88 24.62 ;
    RECT 31.37 23.83 31.58 23.9 ;
    RECT 31.37 24.19 31.58 24.26 ;
    RECT 31.37 24.55 31.58 24.62 ;
    RECT 31.83 23.83 32.04 23.9 ;
    RECT 31.83 24.19 32.04 24.26 ;
    RECT 31.83 24.55 32.04 24.62 ;
    RECT 67.89 23.83 68.1 23.9 ;
    RECT 67.89 24.19 68.1 24.26 ;
    RECT 67.89 24.55 68.1 24.62 ;
    RECT 68.35 23.83 68.56 23.9 ;
    RECT 68.35 24.19 68.56 24.26 ;
    RECT 68.35 24.55 68.56 24.62 ;
    RECT 28.05 23.83 28.26 23.9 ;
    RECT 28.05 24.19 28.26 24.26 ;
    RECT 28.05 24.55 28.26 24.62 ;
    RECT 28.51 23.83 28.72 23.9 ;
    RECT 28.51 24.19 28.72 24.26 ;
    RECT 28.51 24.55 28.72 24.62 ;
    RECT 24.73 23.83 24.94 23.9 ;
    RECT 24.73 24.19 24.94 24.26 ;
    RECT 24.73 24.55 24.94 24.62 ;
    RECT 25.19 23.83 25.4 23.9 ;
    RECT 25.19 24.19 25.4 24.26 ;
    RECT 25.19 24.55 25.4 24.62 ;
    RECT 21.41 23.83 21.62 23.9 ;
    RECT 21.41 24.19 21.62 24.26 ;
    RECT 21.41 24.55 21.62 24.62 ;
    RECT 21.87 23.83 22.08 23.9 ;
    RECT 21.87 24.19 22.08 24.26 ;
    RECT 21.87 24.55 22.08 24.62 ;
    RECT 18.09 23.83 18.3 23.9 ;
    RECT 18.09 24.19 18.3 24.26 ;
    RECT 18.09 24.55 18.3 24.62 ;
    RECT 18.55 23.83 18.76 23.9 ;
    RECT 18.55 24.19 18.76 24.26 ;
    RECT 18.55 24.55 18.76 24.62 ;
    RECT 120.825 24.19 120.895 24.26 ;
    RECT 14.77 23.83 14.98 23.9 ;
    RECT 14.77 24.19 14.98 24.26 ;
    RECT 14.77 24.55 14.98 24.62 ;
    RECT 15.23 23.83 15.44 23.9 ;
    RECT 15.23 24.19 15.44 24.26 ;
    RECT 15.23 24.55 15.44 24.62 ;
    RECT 11.45 23.83 11.66 23.9 ;
    RECT 11.45 24.19 11.66 24.26 ;
    RECT 11.45 24.55 11.66 24.62 ;
    RECT 11.91 23.83 12.12 23.9 ;
    RECT 11.91 24.19 12.12 24.26 ;
    RECT 11.91 24.55 12.12 24.62 ;
    RECT 8.13 23.83 8.34 23.9 ;
    RECT 8.13 24.19 8.34 24.26 ;
    RECT 8.13 24.55 8.34 24.62 ;
    RECT 8.59 23.83 8.8 23.9 ;
    RECT 8.59 24.19 8.8 24.26 ;
    RECT 8.59 24.55 8.8 24.62 ;
    RECT 4.81 23.83 5.02 23.9 ;
    RECT 4.81 24.19 5.02 24.26 ;
    RECT 4.81 24.55 5.02 24.62 ;
    RECT 5.27 23.83 5.48 23.9 ;
    RECT 5.27 24.19 5.48 24.26 ;
    RECT 5.27 24.55 5.48 24.62 ;
    RECT 1.49 23.83 1.7 23.9 ;
    RECT 1.49 24.19 1.7 24.26 ;
    RECT 1.49 24.55 1.7 24.62 ;
    RECT 1.95 23.83 2.16 23.9 ;
    RECT 1.95 24.19 2.16 24.26 ;
    RECT 1.95 24.55 2.16 24.62 ;
    RECT 64.57 23.83 64.78 23.9 ;
    RECT 64.57 24.19 64.78 24.26 ;
    RECT 64.57 24.55 64.78 24.62 ;
    RECT 65.03 23.83 65.24 23.9 ;
    RECT 65.03 24.19 65.24 24.26 ;
    RECT 65.03 24.55 65.24 24.62 ;
    RECT 61.25 63.45 61.46 63.52 ;
    RECT 61.25 63.81 61.46 63.88 ;
    RECT 61.25 64.17 61.46 64.24 ;
    RECT 61.71 63.45 61.92 63.52 ;
    RECT 61.71 63.81 61.92 63.88 ;
    RECT 61.71 64.17 61.92 64.24 ;
    RECT 57.93 63.45 58.14 63.52 ;
    RECT 57.93 63.81 58.14 63.88 ;
    RECT 57.93 64.17 58.14 64.24 ;
    RECT 58.39 63.45 58.6 63.52 ;
    RECT 58.39 63.81 58.6 63.88 ;
    RECT 58.39 64.17 58.6 64.24 ;
    RECT 54.61 63.45 54.82 63.52 ;
    RECT 54.61 63.81 54.82 63.88 ;
    RECT 54.61 64.17 54.82 64.24 ;
    RECT 55.07 63.45 55.28 63.52 ;
    RECT 55.07 63.81 55.28 63.88 ;
    RECT 55.07 64.17 55.28 64.24 ;
    RECT 51.29 63.45 51.5 63.52 ;
    RECT 51.29 63.81 51.5 63.88 ;
    RECT 51.29 64.17 51.5 64.24 ;
    RECT 51.75 63.45 51.96 63.52 ;
    RECT 51.75 63.81 51.96 63.88 ;
    RECT 51.75 64.17 51.96 64.24 ;
    RECT 47.97 63.45 48.18 63.52 ;
    RECT 47.97 63.81 48.18 63.88 ;
    RECT 47.97 64.17 48.18 64.24 ;
    RECT 48.43 63.45 48.64 63.52 ;
    RECT 48.43 63.81 48.64 63.88 ;
    RECT 48.43 64.17 48.64 64.24 ;
    RECT 44.65 63.45 44.86 63.52 ;
    RECT 44.65 63.81 44.86 63.88 ;
    RECT 44.65 64.17 44.86 64.24 ;
    RECT 45.11 63.45 45.32 63.52 ;
    RECT 45.11 63.81 45.32 63.88 ;
    RECT 45.11 64.17 45.32 64.24 ;
    RECT 41.33 63.45 41.54 63.52 ;
    RECT 41.33 63.81 41.54 63.88 ;
    RECT 41.33 64.17 41.54 64.24 ;
    RECT 41.79 63.45 42.0 63.52 ;
    RECT 41.79 63.81 42.0 63.88 ;
    RECT 41.79 64.17 42.0 64.24 ;
    RECT 38.01 63.45 38.22 63.52 ;
    RECT 38.01 63.81 38.22 63.88 ;
    RECT 38.01 64.17 38.22 64.24 ;
    RECT 38.47 63.45 38.68 63.52 ;
    RECT 38.47 63.81 38.68 63.88 ;
    RECT 38.47 64.17 38.68 64.24 ;
    RECT 0.4 63.81 0.47 63.88 ;
    RECT 34.69 63.45 34.9 63.52 ;
    RECT 34.69 63.81 34.9 63.88 ;
    RECT 34.69 64.17 34.9 64.24 ;
    RECT 35.15 63.45 35.36 63.52 ;
    RECT 35.15 63.81 35.36 63.88 ;
    RECT 35.15 64.17 35.36 64.24 ;
    RECT 117.69 63.45 117.9 63.52 ;
    RECT 117.69 63.81 117.9 63.88 ;
    RECT 117.69 64.17 117.9 64.24 ;
    RECT 118.15 63.45 118.36 63.52 ;
    RECT 118.15 63.81 118.36 63.88 ;
    RECT 118.15 64.17 118.36 64.24 ;
    RECT 114.37 63.45 114.58 63.52 ;
    RECT 114.37 63.81 114.58 63.88 ;
    RECT 114.37 64.17 114.58 64.24 ;
    RECT 114.83 63.45 115.04 63.52 ;
    RECT 114.83 63.81 115.04 63.88 ;
    RECT 114.83 64.17 115.04 64.24 ;
    RECT 111.05 63.45 111.26 63.52 ;
    RECT 111.05 63.81 111.26 63.88 ;
    RECT 111.05 64.17 111.26 64.24 ;
    RECT 111.51 63.45 111.72 63.52 ;
    RECT 111.51 63.81 111.72 63.88 ;
    RECT 111.51 64.17 111.72 64.24 ;
    RECT 107.73 63.45 107.94 63.52 ;
    RECT 107.73 63.81 107.94 63.88 ;
    RECT 107.73 64.17 107.94 64.24 ;
    RECT 108.19 63.45 108.4 63.52 ;
    RECT 108.19 63.81 108.4 63.88 ;
    RECT 108.19 64.17 108.4 64.24 ;
    RECT 104.41 63.45 104.62 63.52 ;
    RECT 104.41 63.81 104.62 63.88 ;
    RECT 104.41 64.17 104.62 64.24 ;
    RECT 104.87 63.45 105.08 63.52 ;
    RECT 104.87 63.81 105.08 63.88 ;
    RECT 104.87 64.17 105.08 64.24 ;
    RECT 101.09 63.45 101.3 63.52 ;
    RECT 101.09 63.81 101.3 63.88 ;
    RECT 101.09 64.17 101.3 64.24 ;
    RECT 101.55 63.45 101.76 63.52 ;
    RECT 101.55 63.81 101.76 63.88 ;
    RECT 101.55 64.17 101.76 64.24 ;
    RECT 97.77 63.45 97.98 63.52 ;
    RECT 97.77 63.81 97.98 63.88 ;
    RECT 97.77 64.17 97.98 64.24 ;
    RECT 98.23 63.45 98.44 63.52 ;
    RECT 98.23 63.81 98.44 63.88 ;
    RECT 98.23 64.17 98.44 64.24 ;
    RECT 94.45 63.45 94.66 63.52 ;
    RECT 94.45 63.81 94.66 63.88 ;
    RECT 94.45 64.17 94.66 64.24 ;
    RECT 94.91 63.45 95.12 63.52 ;
    RECT 94.91 63.81 95.12 63.88 ;
    RECT 94.91 64.17 95.12 64.24 ;
    RECT 91.13 63.45 91.34 63.52 ;
    RECT 91.13 63.81 91.34 63.88 ;
    RECT 91.13 64.17 91.34 64.24 ;
    RECT 91.59 63.45 91.8 63.52 ;
    RECT 91.59 63.81 91.8 63.88 ;
    RECT 91.59 64.17 91.8 64.24 ;
    RECT 87.81 63.45 88.02 63.52 ;
    RECT 87.81 63.81 88.02 63.88 ;
    RECT 87.81 64.17 88.02 64.24 ;
    RECT 88.27 63.45 88.48 63.52 ;
    RECT 88.27 63.81 88.48 63.88 ;
    RECT 88.27 64.17 88.48 64.24 ;
    RECT 84.49 63.45 84.7 63.52 ;
    RECT 84.49 63.81 84.7 63.88 ;
    RECT 84.49 64.17 84.7 64.24 ;
    RECT 84.95 63.45 85.16 63.52 ;
    RECT 84.95 63.81 85.16 63.88 ;
    RECT 84.95 64.17 85.16 64.24 ;
    RECT 81.17 63.45 81.38 63.52 ;
    RECT 81.17 63.81 81.38 63.88 ;
    RECT 81.17 64.17 81.38 64.24 ;
    RECT 81.63 63.45 81.84 63.52 ;
    RECT 81.63 63.81 81.84 63.88 ;
    RECT 81.63 64.17 81.84 64.24 ;
    RECT 77.85 63.45 78.06 63.52 ;
    RECT 77.85 63.81 78.06 63.88 ;
    RECT 77.85 64.17 78.06 64.24 ;
    RECT 78.31 63.45 78.52 63.52 ;
    RECT 78.31 63.81 78.52 63.88 ;
    RECT 78.31 64.17 78.52 64.24 ;
    RECT 74.53 63.45 74.74 63.52 ;
    RECT 74.53 63.81 74.74 63.88 ;
    RECT 74.53 64.17 74.74 64.24 ;
    RECT 74.99 63.45 75.2 63.52 ;
    RECT 74.99 63.81 75.2 63.88 ;
    RECT 74.99 64.17 75.2 64.24 ;
    RECT 71.21 63.45 71.42 63.52 ;
    RECT 71.21 63.81 71.42 63.88 ;
    RECT 71.21 64.17 71.42 64.24 ;
    RECT 71.67 63.45 71.88 63.52 ;
    RECT 71.67 63.81 71.88 63.88 ;
    RECT 71.67 64.17 71.88 64.24 ;
    RECT 31.37 63.45 31.58 63.52 ;
    RECT 31.37 63.81 31.58 63.88 ;
    RECT 31.37 64.17 31.58 64.24 ;
    RECT 31.83 63.45 32.04 63.52 ;
    RECT 31.83 63.81 32.04 63.88 ;
    RECT 31.83 64.17 32.04 64.24 ;
    RECT 67.89 63.45 68.1 63.52 ;
    RECT 67.89 63.81 68.1 63.88 ;
    RECT 67.89 64.17 68.1 64.24 ;
    RECT 68.35 63.45 68.56 63.52 ;
    RECT 68.35 63.81 68.56 63.88 ;
    RECT 68.35 64.17 68.56 64.24 ;
    RECT 28.05 63.45 28.26 63.52 ;
    RECT 28.05 63.81 28.26 63.88 ;
    RECT 28.05 64.17 28.26 64.24 ;
    RECT 28.51 63.45 28.72 63.52 ;
    RECT 28.51 63.81 28.72 63.88 ;
    RECT 28.51 64.17 28.72 64.24 ;
    RECT 24.73 63.45 24.94 63.52 ;
    RECT 24.73 63.81 24.94 63.88 ;
    RECT 24.73 64.17 24.94 64.24 ;
    RECT 25.19 63.45 25.4 63.52 ;
    RECT 25.19 63.81 25.4 63.88 ;
    RECT 25.19 64.17 25.4 64.24 ;
    RECT 21.41 63.45 21.62 63.52 ;
    RECT 21.41 63.81 21.62 63.88 ;
    RECT 21.41 64.17 21.62 64.24 ;
    RECT 21.87 63.45 22.08 63.52 ;
    RECT 21.87 63.81 22.08 63.88 ;
    RECT 21.87 64.17 22.08 64.24 ;
    RECT 18.09 63.45 18.3 63.52 ;
    RECT 18.09 63.81 18.3 63.88 ;
    RECT 18.09 64.17 18.3 64.24 ;
    RECT 18.55 63.45 18.76 63.52 ;
    RECT 18.55 63.81 18.76 63.88 ;
    RECT 18.55 64.17 18.76 64.24 ;
    RECT 120.825 63.81 120.895 63.88 ;
    RECT 14.77 63.45 14.98 63.52 ;
    RECT 14.77 63.81 14.98 63.88 ;
    RECT 14.77 64.17 14.98 64.24 ;
    RECT 15.23 63.45 15.44 63.52 ;
    RECT 15.23 63.81 15.44 63.88 ;
    RECT 15.23 64.17 15.44 64.24 ;
    RECT 11.45 63.45 11.66 63.52 ;
    RECT 11.45 63.81 11.66 63.88 ;
    RECT 11.45 64.17 11.66 64.24 ;
    RECT 11.91 63.45 12.12 63.52 ;
    RECT 11.91 63.81 12.12 63.88 ;
    RECT 11.91 64.17 12.12 64.24 ;
    RECT 8.13 63.45 8.34 63.52 ;
    RECT 8.13 63.81 8.34 63.88 ;
    RECT 8.13 64.17 8.34 64.24 ;
    RECT 8.59 63.45 8.8 63.52 ;
    RECT 8.59 63.81 8.8 63.88 ;
    RECT 8.59 64.17 8.8 64.24 ;
    RECT 4.81 63.45 5.02 63.52 ;
    RECT 4.81 63.81 5.02 63.88 ;
    RECT 4.81 64.17 5.02 64.24 ;
    RECT 5.27 63.45 5.48 63.52 ;
    RECT 5.27 63.81 5.48 63.88 ;
    RECT 5.27 64.17 5.48 64.24 ;
    RECT 1.49 63.45 1.7 63.52 ;
    RECT 1.49 63.81 1.7 63.88 ;
    RECT 1.49 64.17 1.7 64.24 ;
    RECT 1.95 63.45 2.16 63.52 ;
    RECT 1.95 63.81 2.16 63.88 ;
    RECT 1.95 64.17 2.16 64.24 ;
    RECT 64.57 63.45 64.78 63.52 ;
    RECT 64.57 63.81 64.78 63.88 ;
    RECT 64.57 64.17 64.78 64.24 ;
    RECT 65.03 63.45 65.24 63.52 ;
    RECT 65.03 63.81 65.24 63.88 ;
    RECT 65.03 64.17 65.24 64.24 ;
    RECT 61.25 23.11 61.46 23.18 ;
    RECT 61.25 23.47 61.46 23.54 ;
    RECT 61.25 23.83 61.46 23.9 ;
    RECT 61.71 23.11 61.92 23.18 ;
    RECT 61.71 23.47 61.92 23.54 ;
    RECT 61.71 23.83 61.92 23.9 ;
    RECT 57.93 23.11 58.14 23.18 ;
    RECT 57.93 23.47 58.14 23.54 ;
    RECT 57.93 23.83 58.14 23.9 ;
    RECT 58.39 23.11 58.6 23.18 ;
    RECT 58.39 23.47 58.6 23.54 ;
    RECT 58.39 23.83 58.6 23.9 ;
    RECT 54.61 23.11 54.82 23.18 ;
    RECT 54.61 23.47 54.82 23.54 ;
    RECT 54.61 23.83 54.82 23.9 ;
    RECT 55.07 23.11 55.28 23.18 ;
    RECT 55.07 23.47 55.28 23.54 ;
    RECT 55.07 23.83 55.28 23.9 ;
    RECT 51.29 23.11 51.5 23.18 ;
    RECT 51.29 23.47 51.5 23.54 ;
    RECT 51.29 23.83 51.5 23.9 ;
    RECT 51.75 23.11 51.96 23.18 ;
    RECT 51.75 23.47 51.96 23.54 ;
    RECT 51.75 23.83 51.96 23.9 ;
    RECT 47.97 23.11 48.18 23.18 ;
    RECT 47.97 23.47 48.18 23.54 ;
    RECT 47.97 23.83 48.18 23.9 ;
    RECT 48.43 23.11 48.64 23.18 ;
    RECT 48.43 23.47 48.64 23.54 ;
    RECT 48.43 23.83 48.64 23.9 ;
    RECT 44.65 23.11 44.86 23.18 ;
    RECT 44.65 23.47 44.86 23.54 ;
    RECT 44.65 23.83 44.86 23.9 ;
    RECT 45.11 23.11 45.32 23.18 ;
    RECT 45.11 23.47 45.32 23.54 ;
    RECT 45.11 23.83 45.32 23.9 ;
    RECT 41.33 23.11 41.54 23.18 ;
    RECT 41.33 23.47 41.54 23.54 ;
    RECT 41.33 23.83 41.54 23.9 ;
    RECT 41.79 23.11 42.0 23.18 ;
    RECT 41.79 23.47 42.0 23.54 ;
    RECT 41.79 23.83 42.0 23.9 ;
    RECT 38.01 23.11 38.22 23.18 ;
    RECT 38.01 23.47 38.22 23.54 ;
    RECT 38.01 23.83 38.22 23.9 ;
    RECT 38.47 23.11 38.68 23.18 ;
    RECT 38.47 23.47 38.68 23.54 ;
    RECT 38.47 23.83 38.68 23.9 ;
    RECT 0.4 23.47 0.47 23.54 ;
    RECT 34.69 23.11 34.9 23.18 ;
    RECT 34.69 23.47 34.9 23.54 ;
    RECT 34.69 23.83 34.9 23.9 ;
    RECT 35.15 23.11 35.36 23.18 ;
    RECT 35.15 23.47 35.36 23.54 ;
    RECT 35.15 23.83 35.36 23.9 ;
    RECT 117.69 23.11 117.9 23.18 ;
    RECT 117.69 23.47 117.9 23.54 ;
    RECT 117.69 23.83 117.9 23.9 ;
    RECT 118.15 23.11 118.36 23.18 ;
    RECT 118.15 23.47 118.36 23.54 ;
    RECT 118.15 23.83 118.36 23.9 ;
    RECT 114.37 23.11 114.58 23.18 ;
    RECT 114.37 23.47 114.58 23.54 ;
    RECT 114.37 23.83 114.58 23.9 ;
    RECT 114.83 23.11 115.04 23.18 ;
    RECT 114.83 23.47 115.04 23.54 ;
    RECT 114.83 23.83 115.04 23.9 ;
    RECT 111.05 23.11 111.26 23.18 ;
    RECT 111.05 23.47 111.26 23.54 ;
    RECT 111.05 23.83 111.26 23.9 ;
    RECT 111.51 23.11 111.72 23.18 ;
    RECT 111.51 23.47 111.72 23.54 ;
    RECT 111.51 23.83 111.72 23.9 ;
    RECT 107.73 23.11 107.94 23.18 ;
    RECT 107.73 23.47 107.94 23.54 ;
    RECT 107.73 23.83 107.94 23.9 ;
    RECT 108.19 23.11 108.4 23.18 ;
    RECT 108.19 23.47 108.4 23.54 ;
    RECT 108.19 23.83 108.4 23.9 ;
    RECT 104.41 23.11 104.62 23.18 ;
    RECT 104.41 23.47 104.62 23.54 ;
    RECT 104.41 23.83 104.62 23.9 ;
    RECT 104.87 23.11 105.08 23.18 ;
    RECT 104.87 23.47 105.08 23.54 ;
    RECT 104.87 23.83 105.08 23.9 ;
    RECT 101.09 23.11 101.3 23.18 ;
    RECT 101.09 23.47 101.3 23.54 ;
    RECT 101.09 23.83 101.3 23.9 ;
    RECT 101.55 23.11 101.76 23.18 ;
    RECT 101.55 23.47 101.76 23.54 ;
    RECT 101.55 23.83 101.76 23.9 ;
    RECT 97.77 23.11 97.98 23.18 ;
    RECT 97.77 23.47 97.98 23.54 ;
    RECT 97.77 23.83 97.98 23.9 ;
    RECT 98.23 23.11 98.44 23.18 ;
    RECT 98.23 23.47 98.44 23.54 ;
    RECT 98.23 23.83 98.44 23.9 ;
    RECT 94.45 23.11 94.66 23.18 ;
    RECT 94.45 23.47 94.66 23.54 ;
    RECT 94.45 23.83 94.66 23.9 ;
    RECT 94.91 23.11 95.12 23.18 ;
    RECT 94.91 23.47 95.12 23.54 ;
    RECT 94.91 23.83 95.12 23.9 ;
    RECT 91.13 23.11 91.34 23.18 ;
    RECT 91.13 23.47 91.34 23.54 ;
    RECT 91.13 23.83 91.34 23.9 ;
    RECT 91.59 23.11 91.8 23.18 ;
    RECT 91.59 23.47 91.8 23.54 ;
    RECT 91.59 23.83 91.8 23.9 ;
    RECT 87.81 23.11 88.02 23.18 ;
    RECT 87.81 23.47 88.02 23.54 ;
    RECT 87.81 23.83 88.02 23.9 ;
    RECT 88.27 23.11 88.48 23.18 ;
    RECT 88.27 23.47 88.48 23.54 ;
    RECT 88.27 23.83 88.48 23.9 ;
    RECT 84.49 23.11 84.7 23.18 ;
    RECT 84.49 23.47 84.7 23.54 ;
    RECT 84.49 23.83 84.7 23.9 ;
    RECT 84.95 23.11 85.16 23.18 ;
    RECT 84.95 23.47 85.16 23.54 ;
    RECT 84.95 23.83 85.16 23.9 ;
    RECT 81.17 23.11 81.38 23.18 ;
    RECT 81.17 23.47 81.38 23.54 ;
    RECT 81.17 23.83 81.38 23.9 ;
    RECT 81.63 23.11 81.84 23.18 ;
    RECT 81.63 23.47 81.84 23.54 ;
    RECT 81.63 23.83 81.84 23.9 ;
    RECT 77.85 23.11 78.06 23.18 ;
    RECT 77.85 23.47 78.06 23.54 ;
    RECT 77.85 23.83 78.06 23.9 ;
    RECT 78.31 23.11 78.52 23.18 ;
    RECT 78.31 23.47 78.52 23.54 ;
    RECT 78.31 23.83 78.52 23.9 ;
    RECT 74.53 23.11 74.74 23.18 ;
    RECT 74.53 23.47 74.74 23.54 ;
    RECT 74.53 23.83 74.74 23.9 ;
    RECT 74.99 23.11 75.2 23.18 ;
    RECT 74.99 23.47 75.2 23.54 ;
    RECT 74.99 23.83 75.2 23.9 ;
    RECT 71.21 23.11 71.42 23.18 ;
    RECT 71.21 23.47 71.42 23.54 ;
    RECT 71.21 23.83 71.42 23.9 ;
    RECT 71.67 23.11 71.88 23.18 ;
    RECT 71.67 23.47 71.88 23.54 ;
    RECT 71.67 23.83 71.88 23.9 ;
    RECT 31.37 23.11 31.58 23.18 ;
    RECT 31.37 23.47 31.58 23.54 ;
    RECT 31.37 23.83 31.58 23.9 ;
    RECT 31.83 23.11 32.04 23.18 ;
    RECT 31.83 23.47 32.04 23.54 ;
    RECT 31.83 23.83 32.04 23.9 ;
    RECT 67.89 23.11 68.1 23.18 ;
    RECT 67.89 23.47 68.1 23.54 ;
    RECT 67.89 23.83 68.1 23.9 ;
    RECT 68.35 23.11 68.56 23.18 ;
    RECT 68.35 23.47 68.56 23.54 ;
    RECT 68.35 23.83 68.56 23.9 ;
    RECT 28.05 23.11 28.26 23.18 ;
    RECT 28.05 23.47 28.26 23.54 ;
    RECT 28.05 23.83 28.26 23.9 ;
    RECT 28.51 23.11 28.72 23.18 ;
    RECT 28.51 23.47 28.72 23.54 ;
    RECT 28.51 23.83 28.72 23.9 ;
    RECT 24.73 23.11 24.94 23.18 ;
    RECT 24.73 23.47 24.94 23.54 ;
    RECT 24.73 23.83 24.94 23.9 ;
    RECT 25.19 23.11 25.4 23.18 ;
    RECT 25.19 23.47 25.4 23.54 ;
    RECT 25.19 23.83 25.4 23.9 ;
    RECT 21.41 23.11 21.62 23.18 ;
    RECT 21.41 23.47 21.62 23.54 ;
    RECT 21.41 23.83 21.62 23.9 ;
    RECT 21.87 23.11 22.08 23.18 ;
    RECT 21.87 23.47 22.08 23.54 ;
    RECT 21.87 23.83 22.08 23.9 ;
    RECT 18.09 23.11 18.3 23.18 ;
    RECT 18.09 23.47 18.3 23.54 ;
    RECT 18.09 23.83 18.3 23.9 ;
    RECT 18.55 23.11 18.76 23.18 ;
    RECT 18.55 23.47 18.76 23.54 ;
    RECT 18.55 23.83 18.76 23.9 ;
    RECT 120.825 23.47 120.895 23.54 ;
    RECT 14.77 23.11 14.98 23.18 ;
    RECT 14.77 23.47 14.98 23.54 ;
    RECT 14.77 23.83 14.98 23.9 ;
    RECT 15.23 23.11 15.44 23.18 ;
    RECT 15.23 23.47 15.44 23.54 ;
    RECT 15.23 23.83 15.44 23.9 ;
    RECT 11.45 23.11 11.66 23.18 ;
    RECT 11.45 23.47 11.66 23.54 ;
    RECT 11.45 23.83 11.66 23.9 ;
    RECT 11.91 23.11 12.12 23.18 ;
    RECT 11.91 23.47 12.12 23.54 ;
    RECT 11.91 23.83 12.12 23.9 ;
    RECT 8.13 23.11 8.34 23.18 ;
    RECT 8.13 23.47 8.34 23.54 ;
    RECT 8.13 23.83 8.34 23.9 ;
    RECT 8.59 23.11 8.8 23.18 ;
    RECT 8.59 23.47 8.8 23.54 ;
    RECT 8.59 23.83 8.8 23.9 ;
    RECT 4.81 23.11 5.02 23.18 ;
    RECT 4.81 23.47 5.02 23.54 ;
    RECT 4.81 23.83 5.02 23.9 ;
    RECT 5.27 23.11 5.48 23.18 ;
    RECT 5.27 23.47 5.48 23.54 ;
    RECT 5.27 23.83 5.48 23.9 ;
    RECT 1.49 23.11 1.7 23.18 ;
    RECT 1.49 23.47 1.7 23.54 ;
    RECT 1.49 23.83 1.7 23.9 ;
    RECT 1.95 23.11 2.16 23.18 ;
    RECT 1.95 23.47 2.16 23.54 ;
    RECT 1.95 23.83 2.16 23.9 ;
    RECT 64.57 23.11 64.78 23.18 ;
    RECT 64.57 23.47 64.78 23.54 ;
    RECT 64.57 23.83 64.78 23.9 ;
    RECT 65.03 23.11 65.24 23.18 ;
    RECT 65.03 23.47 65.24 23.54 ;
    RECT 65.03 23.83 65.24 23.9 ;
    RECT 61.25 62.73 61.46 62.8 ;
    RECT 61.25 63.09 61.46 63.16 ;
    RECT 61.25 63.45 61.46 63.52 ;
    RECT 61.71 62.73 61.92 62.8 ;
    RECT 61.71 63.09 61.92 63.16 ;
    RECT 61.71 63.45 61.92 63.52 ;
    RECT 57.93 62.73 58.14 62.8 ;
    RECT 57.93 63.09 58.14 63.16 ;
    RECT 57.93 63.45 58.14 63.52 ;
    RECT 58.39 62.73 58.6 62.8 ;
    RECT 58.39 63.09 58.6 63.16 ;
    RECT 58.39 63.45 58.6 63.52 ;
    RECT 54.61 62.73 54.82 62.8 ;
    RECT 54.61 63.09 54.82 63.16 ;
    RECT 54.61 63.45 54.82 63.52 ;
    RECT 55.07 62.73 55.28 62.8 ;
    RECT 55.07 63.09 55.28 63.16 ;
    RECT 55.07 63.45 55.28 63.52 ;
    RECT 51.29 62.73 51.5 62.8 ;
    RECT 51.29 63.09 51.5 63.16 ;
    RECT 51.29 63.45 51.5 63.52 ;
    RECT 51.75 62.73 51.96 62.8 ;
    RECT 51.75 63.09 51.96 63.16 ;
    RECT 51.75 63.45 51.96 63.52 ;
    RECT 47.97 62.73 48.18 62.8 ;
    RECT 47.97 63.09 48.18 63.16 ;
    RECT 47.97 63.45 48.18 63.52 ;
    RECT 48.43 62.73 48.64 62.8 ;
    RECT 48.43 63.09 48.64 63.16 ;
    RECT 48.43 63.45 48.64 63.52 ;
    RECT 44.65 62.73 44.86 62.8 ;
    RECT 44.65 63.09 44.86 63.16 ;
    RECT 44.65 63.45 44.86 63.52 ;
    RECT 45.11 62.73 45.32 62.8 ;
    RECT 45.11 63.09 45.32 63.16 ;
    RECT 45.11 63.45 45.32 63.52 ;
    RECT 41.33 62.73 41.54 62.8 ;
    RECT 41.33 63.09 41.54 63.16 ;
    RECT 41.33 63.45 41.54 63.52 ;
    RECT 41.79 62.73 42.0 62.8 ;
    RECT 41.79 63.09 42.0 63.16 ;
    RECT 41.79 63.45 42.0 63.52 ;
    RECT 38.01 62.73 38.22 62.8 ;
    RECT 38.01 63.09 38.22 63.16 ;
    RECT 38.01 63.45 38.22 63.52 ;
    RECT 38.47 62.73 38.68 62.8 ;
    RECT 38.47 63.09 38.68 63.16 ;
    RECT 38.47 63.45 38.68 63.52 ;
    RECT 0.4 63.09 0.47 63.16 ;
    RECT 34.69 62.73 34.9 62.8 ;
    RECT 34.69 63.09 34.9 63.16 ;
    RECT 34.69 63.45 34.9 63.52 ;
    RECT 35.15 62.73 35.36 62.8 ;
    RECT 35.15 63.09 35.36 63.16 ;
    RECT 35.15 63.45 35.36 63.52 ;
    RECT 117.69 62.73 117.9 62.8 ;
    RECT 117.69 63.09 117.9 63.16 ;
    RECT 117.69 63.45 117.9 63.52 ;
    RECT 118.15 62.73 118.36 62.8 ;
    RECT 118.15 63.09 118.36 63.16 ;
    RECT 118.15 63.45 118.36 63.52 ;
    RECT 114.37 62.73 114.58 62.8 ;
    RECT 114.37 63.09 114.58 63.16 ;
    RECT 114.37 63.45 114.58 63.52 ;
    RECT 114.83 62.73 115.04 62.8 ;
    RECT 114.83 63.09 115.04 63.16 ;
    RECT 114.83 63.45 115.04 63.52 ;
    RECT 111.05 62.73 111.26 62.8 ;
    RECT 111.05 63.09 111.26 63.16 ;
    RECT 111.05 63.45 111.26 63.52 ;
    RECT 111.51 62.73 111.72 62.8 ;
    RECT 111.51 63.09 111.72 63.16 ;
    RECT 111.51 63.45 111.72 63.52 ;
    RECT 107.73 62.73 107.94 62.8 ;
    RECT 107.73 63.09 107.94 63.16 ;
    RECT 107.73 63.45 107.94 63.52 ;
    RECT 108.19 62.73 108.4 62.8 ;
    RECT 108.19 63.09 108.4 63.16 ;
    RECT 108.19 63.45 108.4 63.52 ;
    RECT 104.41 62.73 104.62 62.8 ;
    RECT 104.41 63.09 104.62 63.16 ;
    RECT 104.41 63.45 104.62 63.52 ;
    RECT 104.87 62.73 105.08 62.8 ;
    RECT 104.87 63.09 105.08 63.16 ;
    RECT 104.87 63.45 105.08 63.52 ;
    RECT 101.09 62.73 101.3 62.8 ;
    RECT 101.09 63.09 101.3 63.16 ;
    RECT 101.09 63.45 101.3 63.52 ;
    RECT 101.55 62.73 101.76 62.8 ;
    RECT 101.55 63.09 101.76 63.16 ;
    RECT 101.55 63.45 101.76 63.52 ;
    RECT 97.77 62.73 97.98 62.8 ;
    RECT 97.77 63.09 97.98 63.16 ;
    RECT 97.77 63.45 97.98 63.52 ;
    RECT 98.23 62.73 98.44 62.8 ;
    RECT 98.23 63.09 98.44 63.16 ;
    RECT 98.23 63.45 98.44 63.52 ;
    RECT 94.45 62.73 94.66 62.8 ;
    RECT 94.45 63.09 94.66 63.16 ;
    RECT 94.45 63.45 94.66 63.52 ;
    RECT 94.91 62.73 95.12 62.8 ;
    RECT 94.91 63.09 95.12 63.16 ;
    RECT 94.91 63.45 95.12 63.52 ;
    RECT 91.13 62.73 91.34 62.8 ;
    RECT 91.13 63.09 91.34 63.16 ;
    RECT 91.13 63.45 91.34 63.52 ;
    RECT 91.59 62.73 91.8 62.8 ;
    RECT 91.59 63.09 91.8 63.16 ;
    RECT 91.59 63.45 91.8 63.52 ;
    RECT 87.81 62.73 88.02 62.8 ;
    RECT 87.81 63.09 88.02 63.16 ;
    RECT 87.81 63.45 88.02 63.52 ;
    RECT 88.27 62.73 88.48 62.8 ;
    RECT 88.27 63.09 88.48 63.16 ;
    RECT 88.27 63.45 88.48 63.52 ;
    RECT 84.49 62.73 84.7 62.8 ;
    RECT 84.49 63.09 84.7 63.16 ;
    RECT 84.49 63.45 84.7 63.52 ;
    RECT 84.95 62.73 85.16 62.8 ;
    RECT 84.95 63.09 85.16 63.16 ;
    RECT 84.95 63.45 85.16 63.52 ;
    RECT 81.17 62.73 81.38 62.8 ;
    RECT 81.17 63.09 81.38 63.16 ;
    RECT 81.17 63.45 81.38 63.52 ;
    RECT 81.63 62.73 81.84 62.8 ;
    RECT 81.63 63.09 81.84 63.16 ;
    RECT 81.63 63.45 81.84 63.52 ;
    RECT 77.85 62.73 78.06 62.8 ;
    RECT 77.85 63.09 78.06 63.16 ;
    RECT 77.85 63.45 78.06 63.52 ;
    RECT 78.31 62.73 78.52 62.8 ;
    RECT 78.31 63.09 78.52 63.16 ;
    RECT 78.31 63.45 78.52 63.52 ;
    RECT 74.53 62.73 74.74 62.8 ;
    RECT 74.53 63.09 74.74 63.16 ;
    RECT 74.53 63.45 74.74 63.52 ;
    RECT 74.99 62.73 75.2 62.8 ;
    RECT 74.99 63.09 75.2 63.16 ;
    RECT 74.99 63.45 75.2 63.52 ;
    RECT 71.21 62.73 71.42 62.8 ;
    RECT 71.21 63.09 71.42 63.16 ;
    RECT 71.21 63.45 71.42 63.52 ;
    RECT 71.67 62.73 71.88 62.8 ;
    RECT 71.67 63.09 71.88 63.16 ;
    RECT 71.67 63.45 71.88 63.52 ;
    RECT 31.37 62.73 31.58 62.8 ;
    RECT 31.37 63.09 31.58 63.16 ;
    RECT 31.37 63.45 31.58 63.52 ;
    RECT 31.83 62.73 32.04 62.8 ;
    RECT 31.83 63.09 32.04 63.16 ;
    RECT 31.83 63.45 32.04 63.52 ;
    RECT 67.89 62.73 68.1 62.8 ;
    RECT 67.89 63.09 68.1 63.16 ;
    RECT 67.89 63.45 68.1 63.52 ;
    RECT 68.35 62.73 68.56 62.8 ;
    RECT 68.35 63.09 68.56 63.16 ;
    RECT 68.35 63.45 68.56 63.52 ;
    RECT 28.05 62.73 28.26 62.8 ;
    RECT 28.05 63.09 28.26 63.16 ;
    RECT 28.05 63.45 28.26 63.52 ;
    RECT 28.51 62.73 28.72 62.8 ;
    RECT 28.51 63.09 28.72 63.16 ;
    RECT 28.51 63.45 28.72 63.52 ;
    RECT 24.73 62.73 24.94 62.8 ;
    RECT 24.73 63.09 24.94 63.16 ;
    RECT 24.73 63.45 24.94 63.52 ;
    RECT 25.19 62.73 25.4 62.8 ;
    RECT 25.19 63.09 25.4 63.16 ;
    RECT 25.19 63.45 25.4 63.52 ;
    RECT 21.41 62.73 21.62 62.8 ;
    RECT 21.41 63.09 21.62 63.16 ;
    RECT 21.41 63.45 21.62 63.52 ;
    RECT 21.87 62.73 22.08 62.8 ;
    RECT 21.87 63.09 22.08 63.16 ;
    RECT 21.87 63.45 22.08 63.52 ;
    RECT 18.09 62.73 18.3 62.8 ;
    RECT 18.09 63.09 18.3 63.16 ;
    RECT 18.09 63.45 18.3 63.52 ;
    RECT 18.55 62.73 18.76 62.8 ;
    RECT 18.55 63.09 18.76 63.16 ;
    RECT 18.55 63.45 18.76 63.52 ;
    RECT 120.825 63.09 120.895 63.16 ;
    RECT 14.77 62.73 14.98 62.8 ;
    RECT 14.77 63.09 14.98 63.16 ;
    RECT 14.77 63.45 14.98 63.52 ;
    RECT 15.23 62.73 15.44 62.8 ;
    RECT 15.23 63.09 15.44 63.16 ;
    RECT 15.23 63.45 15.44 63.52 ;
    RECT 11.45 62.73 11.66 62.8 ;
    RECT 11.45 63.09 11.66 63.16 ;
    RECT 11.45 63.45 11.66 63.52 ;
    RECT 11.91 62.73 12.12 62.8 ;
    RECT 11.91 63.09 12.12 63.16 ;
    RECT 11.91 63.45 12.12 63.52 ;
    RECT 8.13 62.73 8.34 62.8 ;
    RECT 8.13 63.09 8.34 63.16 ;
    RECT 8.13 63.45 8.34 63.52 ;
    RECT 8.59 62.73 8.8 62.8 ;
    RECT 8.59 63.09 8.8 63.16 ;
    RECT 8.59 63.45 8.8 63.52 ;
    RECT 4.81 62.73 5.02 62.8 ;
    RECT 4.81 63.09 5.02 63.16 ;
    RECT 4.81 63.45 5.02 63.52 ;
    RECT 5.27 62.73 5.48 62.8 ;
    RECT 5.27 63.09 5.48 63.16 ;
    RECT 5.27 63.45 5.48 63.52 ;
    RECT 1.49 62.73 1.7 62.8 ;
    RECT 1.49 63.09 1.7 63.16 ;
    RECT 1.49 63.45 1.7 63.52 ;
    RECT 1.95 62.73 2.16 62.8 ;
    RECT 1.95 63.09 2.16 63.16 ;
    RECT 1.95 63.45 2.16 63.52 ;
    RECT 64.57 62.73 64.78 62.8 ;
    RECT 64.57 63.09 64.78 63.16 ;
    RECT 64.57 63.45 64.78 63.52 ;
    RECT 65.03 62.73 65.24 62.8 ;
    RECT 65.03 63.09 65.24 63.16 ;
    RECT 65.03 63.45 65.24 63.52 ;
    RECT 61.25 22.39 61.46 22.46 ;
    RECT 61.25 22.75 61.46 22.82 ;
    RECT 61.25 23.11 61.46 23.18 ;
    RECT 61.71 22.39 61.92 22.46 ;
    RECT 61.71 22.75 61.92 22.82 ;
    RECT 61.71 23.11 61.92 23.18 ;
    RECT 57.93 22.39 58.14 22.46 ;
    RECT 57.93 22.75 58.14 22.82 ;
    RECT 57.93 23.11 58.14 23.18 ;
    RECT 58.39 22.39 58.6 22.46 ;
    RECT 58.39 22.75 58.6 22.82 ;
    RECT 58.39 23.11 58.6 23.18 ;
    RECT 54.61 22.39 54.82 22.46 ;
    RECT 54.61 22.75 54.82 22.82 ;
    RECT 54.61 23.11 54.82 23.18 ;
    RECT 55.07 22.39 55.28 22.46 ;
    RECT 55.07 22.75 55.28 22.82 ;
    RECT 55.07 23.11 55.28 23.18 ;
    RECT 51.29 22.39 51.5 22.46 ;
    RECT 51.29 22.75 51.5 22.82 ;
    RECT 51.29 23.11 51.5 23.18 ;
    RECT 51.75 22.39 51.96 22.46 ;
    RECT 51.75 22.75 51.96 22.82 ;
    RECT 51.75 23.11 51.96 23.18 ;
    RECT 47.97 22.39 48.18 22.46 ;
    RECT 47.97 22.75 48.18 22.82 ;
    RECT 47.97 23.11 48.18 23.18 ;
    RECT 48.43 22.39 48.64 22.46 ;
    RECT 48.43 22.75 48.64 22.82 ;
    RECT 48.43 23.11 48.64 23.18 ;
    RECT 44.65 22.39 44.86 22.46 ;
    RECT 44.65 22.75 44.86 22.82 ;
    RECT 44.65 23.11 44.86 23.18 ;
    RECT 45.11 22.39 45.32 22.46 ;
    RECT 45.11 22.75 45.32 22.82 ;
    RECT 45.11 23.11 45.32 23.18 ;
    RECT 41.33 22.39 41.54 22.46 ;
    RECT 41.33 22.75 41.54 22.82 ;
    RECT 41.33 23.11 41.54 23.18 ;
    RECT 41.79 22.39 42.0 22.46 ;
    RECT 41.79 22.75 42.0 22.82 ;
    RECT 41.79 23.11 42.0 23.18 ;
    RECT 38.01 22.39 38.22 22.46 ;
    RECT 38.01 22.75 38.22 22.82 ;
    RECT 38.01 23.11 38.22 23.18 ;
    RECT 38.47 22.39 38.68 22.46 ;
    RECT 38.47 22.75 38.68 22.82 ;
    RECT 38.47 23.11 38.68 23.18 ;
    RECT 0.4 22.75 0.47 22.82 ;
    RECT 34.69 22.39 34.9 22.46 ;
    RECT 34.69 22.75 34.9 22.82 ;
    RECT 34.69 23.11 34.9 23.18 ;
    RECT 35.15 22.39 35.36 22.46 ;
    RECT 35.15 22.75 35.36 22.82 ;
    RECT 35.15 23.11 35.36 23.18 ;
    RECT 117.69 22.39 117.9 22.46 ;
    RECT 117.69 22.75 117.9 22.82 ;
    RECT 117.69 23.11 117.9 23.18 ;
    RECT 118.15 22.39 118.36 22.46 ;
    RECT 118.15 22.75 118.36 22.82 ;
    RECT 118.15 23.11 118.36 23.18 ;
    RECT 114.37 22.39 114.58 22.46 ;
    RECT 114.37 22.75 114.58 22.82 ;
    RECT 114.37 23.11 114.58 23.18 ;
    RECT 114.83 22.39 115.04 22.46 ;
    RECT 114.83 22.75 115.04 22.82 ;
    RECT 114.83 23.11 115.04 23.18 ;
    RECT 111.05 22.39 111.26 22.46 ;
    RECT 111.05 22.75 111.26 22.82 ;
    RECT 111.05 23.11 111.26 23.18 ;
    RECT 111.51 22.39 111.72 22.46 ;
    RECT 111.51 22.75 111.72 22.82 ;
    RECT 111.51 23.11 111.72 23.18 ;
    RECT 107.73 22.39 107.94 22.46 ;
    RECT 107.73 22.75 107.94 22.82 ;
    RECT 107.73 23.11 107.94 23.18 ;
    RECT 108.19 22.39 108.4 22.46 ;
    RECT 108.19 22.75 108.4 22.82 ;
    RECT 108.19 23.11 108.4 23.18 ;
    RECT 104.41 22.39 104.62 22.46 ;
    RECT 104.41 22.75 104.62 22.82 ;
    RECT 104.41 23.11 104.62 23.18 ;
    RECT 104.87 22.39 105.08 22.46 ;
    RECT 104.87 22.75 105.08 22.82 ;
    RECT 104.87 23.11 105.08 23.18 ;
    RECT 101.09 22.39 101.3 22.46 ;
    RECT 101.09 22.75 101.3 22.82 ;
    RECT 101.09 23.11 101.3 23.18 ;
    RECT 101.55 22.39 101.76 22.46 ;
    RECT 101.55 22.75 101.76 22.82 ;
    RECT 101.55 23.11 101.76 23.18 ;
    RECT 97.77 22.39 97.98 22.46 ;
    RECT 97.77 22.75 97.98 22.82 ;
    RECT 97.77 23.11 97.98 23.18 ;
    RECT 98.23 22.39 98.44 22.46 ;
    RECT 98.23 22.75 98.44 22.82 ;
    RECT 98.23 23.11 98.44 23.18 ;
    RECT 94.45 22.39 94.66 22.46 ;
    RECT 94.45 22.75 94.66 22.82 ;
    RECT 94.45 23.11 94.66 23.18 ;
    RECT 94.91 22.39 95.12 22.46 ;
    RECT 94.91 22.75 95.12 22.82 ;
    RECT 94.91 23.11 95.12 23.18 ;
    RECT 91.13 22.39 91.34 22.46 ;
    RECT 91.13 22.75 91.34 22.82 ;
    RECT 91.13 23.11 91.34 23.18 ;
    RECT 91.59 22.39 91.8 22.46 ;
    RECT 91.59 22.75 91.8 22.82 ;
    RECT 91.59 23.11 91.8 23.18 ;
    RECT 87.81 22.39 88.02 22.46 ;
    RECT 87.81 22.75 88.02 22.82 ;
    RECT 87.81 23.11 88.02 23.18 ;
    RECT 88.27 22.39 88.48 22.46 ;
    RECT 88.27 22.75 88.48 22.82 ;
    RECT 88.27 23.11 88.48 23.18 ;
    RECT 84.49 22.39 84.7 22.46 ;
    RECT 84.49 22.75 84.7 22.82 ;
    RECT 84.49 23.11 84.7 23.18 ;
    RECT 84.95 22.39 85.16 22.46 ;
    RECT 84.95 22.75 85.16 22.82 ;
    RECT 84.95 23.11 85.16 23.18 ;
    RECT 81.17 22.39 81.38 22.46 ;
    RECT 81.17 22.75 81.38 22.82 ;
    RECT 81.17 23.11 81.38 23.18 ;
    RECT 81.63 22.39 81.84 22.46 ;
    RECT 81.63 22.75 81.84 22.82 ;
    RECT 81.63 23.11 81.84 23.18 ;
    RECT 77.85 22.39 78.06 22.46 ;
    RECT 77.85 22.75 78.06 22.82 ;
    RECT 77.85 23.11 78.06 23.18 ;
    RECT 78.31 22.39 78.52 22.46 ;
    RECT 78.31 22.75 78.52 22.82 ;
    RECT 78.31 23.11 78.52 23.18 ;
    RECT 74.53 22.39 74.74 22.46 ;
    RECT 74.53 22.75 74.74 22.82 ;
    RECT 74.53 23.11 74.74 23.18 ;
    RECT 74.99 22.39 75.2 22.46 ;
    RECT 74.99 22.75 75.2 22.82 ;
    RECT 74.99 23.11 75.2 23.18 ;
    RECT 71.21 22.39 71.42 22.46 ;
    RECT 71.21 22.75 71.42 22.82 ;
    RECT 71.21 23.11 71.42 23.18 ;
    RECT 71.67 22.39 71.88 22.46 ;
    RECT 71.67 22.75 71.88 22.82 ;
    RECT 71.67 23.11 71.88 23.18 ;
    RECT 31.37 22.39 31.58 22.46 ;
    RECT 31.37 22.75 31.58 22.82 ;
    RECT 31.37 23.11 31.58 23.18 ;
    RECT 31.83 22.39 32.04 22.46 ;
    RECT 31.83 22.75 32.04 22.82 ;
    RECT 31.83 23.11 32.04 23.18 ;
    RECT 67.89 22.39 68.1 22.46 ;
    RECT 67.89 22.75 68.1 22.82 ;
    RECT 67.89 23.11 68.1 23.18 ;
    RECT 68.35 22.39 68.56 22.46 ;
    RECT 68.35 22.75 68.56 22.82 ;
    RECT 68.35 23.11 68.56 23.18 ;
    RECT 28.05 22.39 28.26 22.46 ;
    RECT 28.05 22.75 28.26 22.82 ;
    RECT 28.05 23.11 28.26 23.18 ;
    RECT 28.51 22.39 28.72 22.46 ;
    RECT 28.51 22.75 28.72 22.82 ;
    RECT 28.51 23.11 28.72 23.18 ;
    RECT 24.73 22.39 24.94 22.46 ;
    RECT 24.73 22.75 24.94 22.82 ;
    RECT 24.73 23.11 24.94 23.18 ;
    RECT 25.19 22.39 25.4 22.46 ;
    RECT 25.19 22.75 25.4 22.82 ;
    RECT 25.19 23.11 25.4 23.18 ;
    RECT 21.41 22.39 21.62 22.46 ;
    RECT 21.41 22.75 21.62 22.82 ;
    RECT 21.41 23.11 21.62 23.18 ;
    RECT 21.87 22.39 22.08 22.46 ;
    RECT 21.87 22.75 22.08 22.82 ;
    RECT 21.87 23.11 22.08 23.18 ;
    RECT 18.09 22.39 18.3 22.46 ;
    RECT 18.09 22.75 18.3 22.82 ;
    RECT 18.09 23.11 18.3 23.18 ;
    RECT 18.55 22.39 18.76 22.46 ;
    RECT 18.55 22.75 18.76 22.82 ;
    RECT 18.55 23.11 18.76 23.18 ;
    RECT 120.825 22.75 120.895 22.82 ;
    RECT 14.77 22.39 14.98 22.46 ;
    RECT 14.77 22.75 14.98 22.82 ;
    RECT 14.77 23.11 14.98 23.18 ;
    RECT 15.23 22.39 15.44 22.46 ;
    RECT 15.23 22.75 15.44 22.82 ;
    RECT 15.23 23.11 15.44 23.18 ;
    RECT 11.45 22.39 11.66 22.46 ;
    RECT 11.45 22.75 11.66 22.82 ;
    RECT 11.45 23.11 11.66 23.18 ;
    RECT 11.91 22.39 12.12 22.46 ;
    RECT 11.91 22.75 12.12 22.82 ;
    RECT 11.91 23.11 12.12 23.18 ;
    RECT 8.13 22.39 8.34 22.46 ;
    RECT 8.13 22.75 8.34 22.82 ;
    RECT 8.13 23.11 8.34 23.18 ;
    RECT 8.59 22.39 8.8 22.46 ;
    RECT 8.59 22.75 8.8 22.82 ;
    RECT 8.59 23.11 8.8 23.18 ;
    RECT 4.81 22.39 5.02 22.46 ;
    RECT 4.81 22.75 5.02 22.82 ;
    RECT 4.81 23.11 5.02 23.18 ;
    RECT 5.27 22.39 5.48 22.46 ;
    RECT 5.27 22.75 5.48 22.82 ;
    RECT 5.27 23.11 5.48 23.18 ;
    RECT 1.49 22.39 1.7 22.46 ;
    RECT 1.49 22.75 1.7 22.82 ;
    RECT 1.49 23.11 1.7 23.18 ;
    RECT 1.95 22.39 2.16 22.46 ;
    RECT 1.95 22.75 2.16 22.82 ;
    RECT 1.95 23.11 2.16 23.18 ;
    RECT 64.57 22.39 64.78 22.46 ;
    RECT 64.57 22.75 64.78 22.82 ;
    RECT 64.57 23.11 64.78 23.18 ;
    RECT 65.03 22.39 65.24 22.46 ;
    RECT 65.03 22.75 65.24 22.82 ;
    RECT 65.03 23.11 65.24 23.18 ;
    RECT 61.25 62.01 61.46 62.08 ;
    RECT 61.25 62.37 61.46 62.44 ;
    RECT 61.25 62.73 61.46 62.8 ;
    RECT 61.71 62.01 61.92 62.08 ;
    RECT 61.71 62.37 61.92 62.44 ;
    RECT 61.71 62.73 61.92 62.8 ;
    RECT 57.93 62.01 58.14 62.08 ;
    RECT 57.93 62.37 58.14 62.44 ;
    RECT 57.93 62.73 58.14 62.8 ;
    RECT 58.39 62.01 58.6 62.08 ;
    RECT 58.39 62.37 58.6 62.44 ;
    RECT 58.39 62.73 58.6 62.8 ;
    RECT 54.61 62.01 54.82 62.08 ;
    RECT 54.61 62.37 54.82 62.44 ;
    RECT 54.61 62.73 54.82 62.8 ;
    RECT 55.07 62.01 55.28 62.08 ;
    RECT 55.07 62.37 55.28 62.44 ;
    RECT 55.07 62.73 55.28 62.8 ;
    RECT 51.29 62.01 51.5 62.08 ;
    RECT 51.29 62.37 51.5 62.44 ;
    RECT 51.29 62.73 51.5 62.8 ;
    RECT 51.75 62.01 51.96 62.08 ;
    RECT 51.75 62.37 51.96 62.44 ;
    RECT 51.75 62.73 51.96 62.8 ;
    RECT 47.97 62.01 48.18 62.08 ;
    RECT 47.97 62.37 48.18 62.44 ;
    RECT 47.97 62.73 48.18 62.8 ;
    RECT 48.43 62.01 48.64 62.08 ;
    RECT 48.43 62.37 48.64 62.44 ;
    RECT 48.43 62.73 48.64 62.8 ;
    RECT 44.65 62.01 44.86 62.08 ;
    RECT 44.65 62.37 44.86 62.44 ;
    RECT 44.65 62.73 44.86 62.8 ;
    RECT 45.11 62.01 45.32 62.08 ;
    RECT 45.11 62.37 45.32 62.44 ;
    RECT 45.11 62.73 45.32 62.8 ;
    RECT 41.33 62.01 41.54 62.08 ;
    RECT 41.33 62.37 41.54 62.44 ;
    RECT 41.33 62.73 41.54 62.8 ;
    RECT 41.79 62.01 42.0 62.08 ;
    RECT 41.79 62.37 42.0 62.44 ;
    RECT 41.79 62.73 42.0 62.8 ;
    RECT 38.01 62.01 38.22 62.08 ;
    RECT 38.01 62.37 38.22 62.44 ;
    RECT 38.01 62.73 38.22 62.8 ;
    RECT 38.47 62.01 38.68 62.08 ;
    RECT 38.47 62.37 38.68 62.44 ;
    RECT 38.47 62.73 38.68 62.8 ;
    RECT 0.4 62.37 0.47 62.44 ;
    RECT 34.69 62.01 34.9 62.08 ;
    RECT 34.69 62.37 34.9 62.44 ;
    RECT 34.69 62.73 34.9 62.8 ;
    RECT 35.15 62.01 35.36 62.08 ;
    RECT 35.15 62.37 35.36 62.44 ;
    RECT 35.15 62.73 35.36 62.8 ;
    RECT 117.69 62.01 117.9 62.08 ;
    RECT 117.69 62.37 117.9 62.44 ;
    RECT 117.69 62.73 117.9 62.8 ;
    RECT 118.15 62.01 118.36 62.08 ;
    RECT 118.15 62.37 118.36 62.44 ;
    RECT 118.15 62.73 118.36 62.8 ;
    RECT 114.37 62.01 114.58 62.08 ;
    RECT 114.37 62.37 114.58 62.44 ;
    RECT 114.37 62.73 114.58 62.8 ;
    RECT 114.83 62.01 115.04 62.08 ;
    RECT 114.83 62.37 115.04 62.44 ;
    RECT 114.83 62.73 115.04 62.8 ;
    RECT 111.05 62.01 111.26 62.08 ;
    RECT 111.05 62.37 111.26 62.44 ;
    RECT 111.05 62.73 111.26 62.8 ;
    RECT 111.51 62.01 111.72 62.08 ;
    RECT 111.51 62.37 111.72 62.44 ;
    RECT 111.51 62.73 111.72 62.8 ;
    RECT 107.73 62.01 107.94 62.08 ;
    RECT 107.73 62.37 107.94 62.44 ;
    RECT 107.73 62.73 107.94 62.8 ;
    RECT 108.19 62.01 108.4 62.08 ;
    RECT 108.19 62.37 108.4 62.44 ;
    RECT 108.19 62.73 108.4 62.8 ;
    RECT 104.41 62.01 104.62 62.08 ;
    RECT 104.41 62.37 104.62 62.44 ;
    RECT 104.41 62.73 104.62 62.8 ;
    RECT 104.87 62.01 105.08 62.08 ;
    RECT 104.87 62.37 105.08 62.44 ;
    RECT 104.87 62.73 105.08 62.8 ;
    RECT 101.09 62.01 101.3 62.08 ;
    RECT 101.09 62.37 101.3 62.44 ;
    RECT 101.09 62.73 101.3 62.8 ;
    RECT 101.55 62.01 101.76 62.08 ;
    RECT 101.55 62.37 101.76 62.44 ;
    RECT 101.55 62.73 101.76 62.8 ;
    RECT 97.77 62.01 97.98 62.08 ;
    RECT 97.77 62.37 97.98 62.44 ;
    RECT 97.77 62.73 97.98 62.8 ;
    RECT 98.23 62.01 98.44 62.08 ;
    RECT 98.23 62.37 98.44 62.44 ;
    RECT 98.23 62.73 98.44 62.8 ;
    RECT 94.45 62.01 94.66 62.08 ;
    RECT 94.45 62.37 94.66 62.44 ;
    RECT 94.45 62.73 94.66 62.8 ;
    RECT 94.91 62.01 95.12 62.08 ;
    RECT 94.91 62.37 95.12 62.44 ;
    RECT 94.91 62.73 95.12 62.8 ;
    RECT 91.13 62.01 91.34 62.08 ;
    RECT 91.13 62.37 91.34 62.44 ;
    RECT 91.13 62.73 91.34 62.8 ;
    RECT 91.59 62.01 91.8 62.08 ;
    RECT 91.59 62.37 91.8 62.44 ;
    RECT 91.59 62.73 91.8 62.8 ;
    RECT 87.81 62.01 88.02 62.08 ;
    RECT 87.81 62.37 88.02 62.44 ;
    RECT 87.81 62.73 88.02 62.8 ;
    RECT 88.27 62.01 88.48 62.08 ;
    RECT 88.27 62.37 88.48 62.44 ;
    RECT 88.27 62.73 88.48 62.8 ;
    RECT 84.49 62.01 84.7 62.08 ;
    RECT 84.49 62.37 84.7 62.44 ;
    RECT 84.49 62.73 84.7 62.8 ;
    RECT 84.95 62.01 85.16 62.08 ;
    RECT 84.95 62.37 85.16 62.44 ;
    RECT 84.95 62.73 85.16 62.8 ;
    RECT 81.17 62.01 81.38 62.08 ;
    RECT 81.17 62.37 81.38 62.44 ;
    RECT 81.17 62.73 81.38 62.8 ;
    RECT 81.63 62.01 81.84 62.08 ;
    RECT 81.63 62.37 81.84 62.44 ;
    RECT 81.63 62.73 81.84 62.8 ;
    RECT 77.85 62.01 78.06 62.08 ;
    RECT 77.85 62.37 78.06 62.44 ;
    RECT 77.85 62.73 78.06 62.8 ;
    RECT 78.31 62.01 78.52 62.08 ;
    RECT 78.31 62.37 78.52 62.44 ;
    RECT 78.31 62.73 78.52 62.8 ;
    RECT 74.53 62.01 74.74 62.08 ;
    RECT 74.53 62.37 74.74 62.44 ;
    RECT 74.53 62.73 74.74 62.8 ;
    RECT 74.99 62.01 75.2 62.08 ;
    RECT 74.99 62.37 75.2 62.44 ;
    RECT 74.99 62.73 75.2 62.8 ;
    RECT 71.21 62.01 71.42 62.08 ;
    RECT 71.21 62.37 71.42 62.44 ;
    RECT 71.21 62.73 71.42 62.8 ;
    RECT 71.67 62.01 71.88 62.08 ;
    RECT 71.67 62.37 71.88 62.44 ;
    RECT 71.67 62.73 71.88 62.8 ;
    RECT 31.37 62.01 31.58 62.08 ;
    RECT 31.37 62.37 31.58 62.44 ;
    RECT 31.37 62.73 31.58 62.8 ;
    RECT 31.83 62.01 32.04 62.08 ;
    RECT 31.83 62.37 32.04 62.44 ;
    RECT 31.83 62.73 32.04 62.8 ;
    RECT 67.89 62.01 68.1 62.08 ;
    RECT 67.89 62.37 68.1 62.44 ;
    RECT 67.89 62.73 68.1 62.8 ;
    RECT 68.35 62.01 68.56 62.08 ;
    RECT 68.35 62.37 68.56 62.44 ;
    RECT 68.35 62.73 68.56 62.8 ;
    RECT 28.05 62.01 28.26 62.08 ;
    RECT 28.05 62.37 28.26 62.44 ;
    RECT 28.05 62.73 28.26 62.8 ;
    RECT 28.51 62.01 28.72 62.08 ;
    RECT 28.51 62.37 28.72 62.44 ;
    RECT 28.51 62.73 28.72 62.8 ;
    RECT 24.73 62.01 24.94 62.08 ;
    RECT 24.73 62.37 24.94 62.44 ;
    RECT 24.73 62.73 24.94 62.8 ;
    RECT 25.19 62.01 25.4 62.08 ;
    RECT 25.19 62.37 25.4 62.44 ;
    RECT 25.19 62.73 25.4 62.8 ;
    RECT 21.41 62.01 21.62 62.08 ;
    RECT 21.41 62.37 21.62 62.44 ;
    RECT 21.41 62.73 21.62 62.8 ;
    RECT 21.87 62.01 22.08 62.08 ;
    RECT 21.87 62.37 22.08 62.44 ;
    RECT 21.87 62.73 22.08 62.8 ;
    RECT 18.09 62.01 18.3 62.08 ;
    RECT 18.09 62.37 18.3 62.44 ;
    RECT 18.09 62.73 18.3 62.8 ;
    RECT 18.55 62.01 18.76 62.08 ;
    RECT 18.55 62.37 18.76 62.44 ;
    RECT 18.55 62.73 18.76 62.8 ;
    RECT 120.825 62.37 120.895 62.44 ;
    RECT 14.77 62.01 14.98 62.08 ;
    RECT 14.77 62.37 14.98 62.44 ;
    RECT 14.77 62.73 14.98 62.8 ;
    RECT 15.23 62.01 15.44 62.08 ;
    RECT 15.23 62.37 15.44 62.44 ;
    RECT 15.23 62.73 15.44 62.8 ;
    RECT 11.45 62.01 11.66 62.08 ;
    RECT 11.45 62.37 11.66 62.44 ;
    RECT 11.45 62.73 11.66 62.8 ;
    RECT 11.91 62.01 12.12 62.08 ;
    RECT 11.91 62.37 12.12 62.44 ;
    RECT 11.91 62.73 12.12 62.8 ;
    RECT 8.13 62.01 8.34 62.08 ;
    RECT 8.13 62.37 8.34 62.44 ;
    RECT 8.13 62.73 8.34 62.8 ;
    RECT 8.59 62.01 8.8 62.08 ;
    RECT 8.59 62.37 8.8 62.44 ;
    RECT 8.59 62.73 8.8 62.8 ;
    RECT 4.81 62.01 5.02 62.08 ;
    RECT 4.81 62.37 5.02 62.44 ;
    RECT 4.81 62.73 5.02 62.8 ;
    RECT 5.27 62.01 5.48 62.08 ;
    RECT 5.27 62.37 5.48 62.44 ;
    RECT 5.27 62.73 5.48 62.8 ;
    RECT 1.49 62.01 1.7 62.08 ;
    RECT 1.49 62.37 1.7 62.44 ;
    RECT 1.49 62.73 1.7 62.8 ;
    RECT 1.95 62.01 2.16 62.08 ;
    RECT 1.95 62.37 2.16 62.44 ;
    RECT 1.95 62.73 2.16 62.8 ;
    RECT 64.57 62.01 64.78 62.08 ;
    RECT 64.57 62.37 64.78 62.44 ;
    RECT 64.57 62.73 64.78 62.8 ;
    RECT 65.03 62.01 65.24 62.08 ;
    RECT 65.03 62.37 65.24 62.44 ;
    RECT 65.03 62.73 65.24 62.8 ;
    RECT 61.25 21.67 61.46 21.74 ;
    RECT 61.25 22.03 61.46 22.1 ;
    RECT 61.25 22.39 61.46 22.46 ;
    RECT 61.71 21.67 61.92 21.74 ;
    RECT 61.71 22.03 61.92 22.1 ;
    RECT 61.71 22.39 61.92 22.46 ;
    RECT 57.93 21.67 58.14 21.74 ;
    RECT 57.93 22.03 58.14 22.1 ;
    RECT 57.93 22.39 58.14 22.46 ;
    RECT 58.39 21.67 58.6 21.74 ;
    RECT 58.39 22.03 58.6 22.1 ;
    RECT 58.39 22.39 58.6 22.46 ;
    RECT 54.61 21.67 54.82 21.74 ;
    RECT 54.61 22.03 54.82 22.1 ;
    RECT 54.61 22.39 54.82 22.46 ;
    RECT 55.07 21.67 55.28 21.74 ;
    RECT 55.07 22.03 55.28 22.1 ;
    RECT 55.07 22.39 55.28 22.46 ;
    RECT 51.29 21.67 51.5 21.74 ;
    RECT 51.29 22.03 51.5 22.1 ;
    RECT 51.29 22.39 51.5 22.46 ;
    RECT 51.75 21.67 51.96 21.74 ;
    RECT 51.75 22.03 51.96 22.1 ;
    RECT 51.75 22.39 51.96 22.46 ;
    RECT 47.97 21.67 48.18 21.74 ;
    RECT 47.97 22.03 48.18 22.1 ;
    RECT 47.97 22.39 48.18 22.46 ;
    RECT 48.43 21.67 48.64 21.74 ;
    RECT 48.43 22.03 48.64 22.1 ;
    RECT 48.43 22.39 48.64 22.46 ;
    RECT 44.65 21.67 44.86 21.74 ;
    RECT 44.65 22.03 44.86 22.1 ;
    RECT 44.65 22.39 44.86 22.46 ;
    RECT 45.11 21.67 45.32 21.74 ;
    RECT 45.11 22.03 45.32 22.1 ;
    RECT 45.11 22.39 45.32 22.46 ;
    RECT 41.33 21.67 41.54 21.74 ;
    RECT 41.33 22.03 41.54 22.1 ;
    RECT 41.33 22.39 41.54 22.46 ;
    RECT 41.79 21.67 42.0 21.74 ;
    RECT 41.79 22.03 42.0 22.1 ;
    RECT 41.79 22.39 42.0 22.46 ;
    RECT 38.01 21.67 38.22 21.74 ;
    RECT 38.01 22.03 38.22 22.1 ;
    RECT 38.01 22.39 38.22 22.46 ;
    RECT 38.47 21.67 38.68 21.74 ;
    RECT 38.47 22.03 38.68 22.1 ;
    RECT 38.47 22.39 38.68 22.46 ;
    RECT 0.4 22.03 0.47 22.1 ;
    RECT 34.69 21.67 34.9 21.74 ;
    RECT 34.69 22.03 34.9 22.1 ;
    RECT 34.69 22.39 34.9 22.46 ;
    RECT 35.15 21.67 35.36 21.74 ;
    RECT 35.15 22.03 35.36 22.1 ;
    RECT 35.15 22.39 35.36 22.46 ;
    RECT 117.69 21.67 117.9 21.74 ;
    RECT 117.69 22.03 117.9 22.1 ;
    RECT 117.69 22.39 117.9 22.46 ;
    RECT 118.15 21.67 118.36 21.74 ;
    RECT 118.15 22.03 118.36 22.1 ;
    RECT 118.15 22.39 118.36 22.46 ;
    RECT 114.37 21.67 114.58 21.74 ;
    RECT 114.37 22.03 114.58 22.1 ;
    RECT 114.37 22.39 114.58 22.46 ;
    RECT 114.83 21.67 115.04 21.74 ;
    RECT 114.83 22.03 115.04 22.1 ;
    RECT 114.83 22.39 115.04 22.46 ;
    RECT 111.05 21.67 111.26 21.74 ;
    RECT 111.05 22.03 111.26 22.1 ;
    RECT 111.05 22.39 111.26 22.46 ;
    RECT 111.51 21.67 111.72 21.74 ;
    RECT 111.51 22.03 111.72 22.1 ;
    RECT 111.51 22.39 111.72 22.46 ;
    RECT 107.73 21.67 107.94 21.74 ;
    RECT 107.73 22.03 107.94 22.1 ;
    RECT 107.73 22.39 107.94 22.46 ;
    RECT 108.19 21.67 108.4 21.74 ;
    RECT 108.19 22.03 108.4 22.1 ;
    RECT 108.19 22.39 108.4 22.46 ;
    RECT 104.41 21.67 104.62 21.74 ;
    RECT 104.41 22.03 104.62 22.1 ;
    RECT 104.41 22.39 104.62 22.46 ;
    RECT 104.87 21.67 105.08 21.74 ;
    RECT 104.87 22.03 105.08 22.1 ;
    RECT 104.87 22.39 105.08 22.46 ;
    RECT 101.09 21.67 101.3 21.74 ;
    RECT 101.09 22.03 101.3 22.1 ;
    RECT 101.09 22.39 101.3 22.46 ;
    RECT 101.55 21.67 101.76 21.74 ;
    RECT 101.55 22.03 101.76 22.1 ;
    RECT 101.55 22.39 101.76 22.46 ;
    RECT 97.77 21.67 97.98 21.74 ;
    RECT 97.77 22.03 97.98 22.1 ;
    RECT 97.77 22.39 97.98 22.46 ;
    RECT 98.23 21.67 98.44 21.74 ;
    RECT 98.23 22.03 98.44 22.1 ;
    RECT 98.23 22.39 98.44 22.46 ;
    RECT 94.45 21.67 94.66 21.74 ;
    RECT 94.45 22.03 94.66 22.1 ;
    RECT 94.45 22.39 94.66 22.46 ;
    RECT 94.91 21.67 95.12 21.74 ;
    RECT 94.91 22.03 95.12 22.1 ;
    RECT 94.91 22.39 95.12 22.46 ;
    RECT 91.13 21.67 91.34 21.74 ;
    RECT 91.13 22.03 91.34 22.1 ;
    RECT 91.13 22.39 91.34 22.46 ;
    RECT 91.59 21.67 91.8 21.74 ;
    RECT 91.59 22.03 91.8 22.1 ;
    RECT 91.59 22.39 91.8 22.46 ;
    RECT 87.81 21.67 88.02 21.74 ;
    RECT 87.81 22.03 88.02 22.1 ;
    RECT 87.81 22.39 88.02 22.46 ;
    RECT 88.27 21.67 88.48 21.74 ;
    RECT 88.27 22.03 88.48 22.1 ;
    RECT 88.27 22.39 88.48 22.46 ;
    RECT 84.49 21.67 84.7 21.74 ;
    RECT 84.49 22.03 84.7 22.1 ;
    RECT 84.49 22.39 84.7 22.46 ;
    RECT 84.95 21.67 85.16 21.74 ;
    RECT 84.95 22.03 85.16 22.1 ;
    RECT 84.95 22.39 85.16 22.46 ;
    RECT 81.17 21.67 81.38 21.74 ;
    RECT 81.17 22.03 81.38 22.1 ;
    RECT 81.17 22.39 81.38 22.46 ;
    RECT 81.63 21.67 81.84 21.74 ;
    RECT 81.63 22.03 81.84 22.1 ;
    RECT 81.63 22.39 81.84 22.46 ;
    RECT 77.85 21.67 78.06 21.74 ;
    RECT 77.85 22.03 78.06 22.1 ;
    RECT 77.85 22.39 78.06 22.46 ;
    RECT 78.31 21.67 78.52 21.74 ;
    RECT 78.31 22.03 78.52 22.1 ;
    RECT 78.31 22.39 78.52 22.46 ;
    RECT 74.53 21.67 74.74 21.74 ;
    RECT 74.53 22.03 74.74 22.1 ;
    RECT 74.53 22.39 74.74 22.46 ;
    RECT 74.99 21.67 75.2 21.74 ;
    RECT 74.99 22.03 75.2 22.1 ;
    RECT 74.99 22.39 75.2 22.46 ;
    RECT 71.21 21.67 71.42 21.74 ;
    RECT 71.21 22.03 71.42 22.1 ;
    RECT 71.21 22.39 71.42 22.46 ;
    RECT 71.67 21.67 71.88 21.74 ;
    RECT 71.67 22.03 71.88 22.1 ;
    RECT 71.67 22.39 71.88 22.46 ;
    RECT 31.37 21.67 31.58 21.74 ;
    RECT 31.37 22.03 31.58 22.1 ;
    RECT 31.37 22.39 31.58 22.46 ;
    RECT 31.83 21.67 32.04 21.74 ;
    RECT 31.83 22.03 32.04 22.1 ;
    RECT 31.83 22.39 32.04 22.46 ;
    RECT 67.89 21.67 68.1 21.74 ;
    RECT 67.89 22.03 68.1 22.1 ;
    RECT 67.89 22.39 68.1 22.46 ;
    RECT 68.35 21.67 68.56 21.74 ;
    RECT 68.35 22.03 68.56 22.1 ;
    RECT 68.35 22.39 68.56 22.46 ;
    RECT 28.05 21.67 28.26 21.74 ;
    RECT 28.05 22.03 28.26 22.1 ;
    RECT 28.05 22.39 28.26 22.46 ;
    RECT 28.51 21.67 28.72 21.74 ;
    RECT 28.51 22.03 28.72 22.1 ;
    RECT 28.51 22.39 28.72 22.46 ;
    RECT 24.73 21.67 24.94 21.74 ;
    RECT 24.73 22.03 24.94 22.1 ;
    RECT 24.73 22.39 24.94 22.46 ;
    RECT 25.19 21.67 25.4 21.74 ;
    RECT 25.19 22.03 25.4 22.1 ;
    RECT 25.19 22.39 25.4 22.46 ;
    RECT 21.41 21.67 21.62 21.74 ;
    RECT 21.41 22.03 21.62 22.1 ;
    RECT 21.41 22.39 21.62 22.46 ;
    RECT 21.87 21.67 22.08 21.74 ;
    RECT 21.87 22.03 22.08 22.1 ;
    RECT 21.87 22.39 22.08 22.46 ;
    RECT 18.09 21.67 18.3 21.74 ;
    RECT 18.09 22.03 18.3 22.1 ;
    RECT 18.09 22.39 18.3 22.46 ;
    RECT 18.55 21.67 18.76 21.74 ;
    RECT 18.55 22.03 18.76 22.1 ;
    RECT 18.55 22.39 18.76 22.46 ;
    RECT 120.825 22.03 120.895 22.1 ;
    RECT 14.77 21.67 14.98 21.74 ;
    RECT 14.77 22.03 14.98 22.1 ;
    RECT 14.77 22.39 14.98 22.46 ;
    RECT 15.23 21.67 15.44 21.74 ;
    RECT 15.23 22.03 15.44 22.1 ;
    RECT 15.23 22.39 15.44 22.46 ;
    RECT 11.45 21.67 11.66 21.74 ;
    RECT 11.45 22.03 11.66 22.1 ;
    RECT 11.45 22.39 11.66 22.46 ;
    RECT 11.91 21.67 12.12 21.74 ;
    RECT 11.91 22.03 12.12 22.1 ;
    RECT 11.91 22.39 12.12 22.46 ;
    RECT 8.13 21.67 8.34 21.74 ;
    RECT 8.13 22.03 8.34 22.1 ;
    RECT 8.13 22.39 8.34 22.46 ;
    RECT 8.59 21.67 8.8 21.74 ;
    RECT 8.59 22.03 8.8 22.1 ;
    RECT 8.59 22.39 8.8 22.46 ;
    RECT 4.81 21.67 5.02 21.74 ;
    RECT 4.81 22.03 5.02 22.1 ;
    RECT 4.81 22.39 5.02 22.46 ;
    RECT 5.27 21.67 5.48 21.74 ;
    RECT 5.27 22.03 5.48 22.1 ;
    RECT 5.27 22.39 5.48 22.46 ;
    RECT 1.49 21.67 1.7 21.74 ;
    RECT 1.49 22.03 1.7 22.1 ;
    RECT 1.49 22.39 1.7 22.46 ;
    RECT 1.95 21.67 2.16 21.74 ;
    RECT 1.95 22.03 2.16 22.1 ;
    RECT 1.95 22.39 2.16 22.46 ;
    RECT 64.57 21.67 64.78 21.74 ;
    RECT 64.57 22.03 64.78 22.1 ;
    RECT 64.57 22.39 64.78 22.46 ;
    RECT 65.03 21.67 65.24 21.74 ;
    RECT 65.03 22.03 65.24 22.1 ;
    RECT 65.03 22.39 65.24 22.46 ;
    RECT 61.25 61.29 61.46 61.36 ;
    RECT 61.25 61.65 61.46 61.72 ;
    RECT 61.25 62.01 61.46 62.08 ;
    RECT 61.71 61.29 61.92 61.36 ;
    RECT 61.71 61.65 61.92 61.72 ;
    RECT 61.71 62.01 61.92 62.08 ;
    RECT 57.93 61.29 58.14 61.36 ;
    RECT 57.93 61.65 58.14 61.72 ;
    RECT 57.93 62.01 58.14 62.08 ;
    RECT 58.39 61.29 58.6 61.36 ;
    RECT 58.39 61.65 58.6 61.72 ;
    RECT 58.39 62.01 58.6 62.08 ;
    RECT 54.61 61.29 54.82 61.36 ;
    RECT 54.61 61.65 54.82 61.72 ;
    RECT 54.61 62.01 54.82 62.08 ;
    RECT 55.07 61.29 55.28 61.36 ;
    RECT 55.07 61.65 55.28 61.72 ;
    RECT 55.07 62.01 55.28 62.08 ;
    RECT 51.29 61.29 51.5 61.36 ;
    RECT 51.29 61.65 51.5 61.72 ;
    RECT 51.29 62.01 51.5 62.08 ;
    RECT 51.75 61.29 51.96 61.36 ;
    RECT 51.75 61.65 51.96 61.72 ;
    RECT 51.75 62.01 51.96 62.08 ;
    RECT 47.97 61.29 48.18 61.36 ;
    RECT 47.97 61.65 48.18 61.72 ;
    RECT 47.97 62.01 48.18 62.08 ;
    RECT 48.43 61.29 48.64 61.36 ;
    RECT 48.43 61.65 48.64 61.72 ;
    RECT 48.43 62.01 48.64 62.08 ;
    RECT 44.65 61.29 44.86 61.36 ;
    RECT 44.65 61.65 44.86 61.72 ;
    RECT 44.65 62.01 44.86 62.08 ;
    RECT 45.11 61.29 45.32 61.36 ;
    RECT 45.11 61.65 45.32 61.72 ;
    RECT 45.11 62.01 45.32 62.08 ;
    RECT 41.33 61.29 41.54 61.36 ;
    RECT 41.33 61.65 41.54 61.72 ;
    RECT 41.33 62.01 41.54 62.08 ;
    RECT 41.79 61.29 42.0 61.36 ;
    RECT 41.79 61.65 42.0 61.72 ;
    RECT 41.79 62.01 42.0 62.08 ;
    RECT 38.01 61.29 38.22 61.36 ;
    RECT 38.01 61.65 38.22 61.72 ;
    RECT 38.01 62.01 38.22 62.08 ;
    RECT 38.47 61.29 38.68 61.36 ;
    RECT 38.47 61.65 38.68 61.72 ;
    RECT 38.47 62.01 38.68 62.08 ;
    RECT 0.4 61.65 0.47 61.72 ;
    RECT 34.69 61.29 34.9 61.36 ;
    RECT 34.69 61.65 34.9 61.72 ;
    RECT 34.69 62.01 34.9 62.08 ;
    RECT 35.15 61.29 35.36 61.36 ;
    RECT 35.15 61.65 35.36 61.72 ;
    RECT 35.15 62.01 35.36 62.08 ;
    RECT 117.69 61.29 117.9 61.36 ;
    RECT 117.69 61.65 117.9 61.72 ;
    RECT 117.69 62.01 117.9 62.08 ;
    RECT 118.15 61.29 118.36 61.36 ;
    RECT 118.15 61.65 118.36 61.72 ;
    RECT 118.15 62.01 118.36 62.08 ;
    RECT 114.37 61.29 114.58 61.36 ;
    RECT 114.37 61.65 114.58 61.72 ;
    RECT 114.37 62.01 114.58 62.08 ;
    RECT 114.83 61.29 115.04 61.36 ;
    RECT 114.83 61.65 115.04 61.72 ;
    RECT 114.83 62.01 115.04 62.08 ;
    RECT 111.05 61.29 111.26 61.36 ;
    RECT 111.05 61.65 111.26 61.72 ;
    RECT 111.05 62.01 111.26 62.08 ;
    RECT 111.51 61.29 111.72 61.36 ;
    RECT 111.51 61.65 111.72 61.72 ;
    RECT 111.51 62.01 111.72 62.08 ;
    RECT 107.73 61.29 107.94 61.36 ;
    RECT 107.73 61.65 107.94 61.72 ;
    RECT 107.73 62.01 107.94 62.08 ;
    RECT 108.19 61.29 108.4 61.36 ;
    RECT 108.19 61.65 108.4 61.72 ;
    RECT 108.19 62.01 108.4 62.08 ;
    RECT 104.41 61.29 104.62 61.36 ;
    RECT 104.41 61.65 104.62 61.72 ;
    RECT 104.41 62.01 104.62 62.08 ;
    RECT 104.87 61.29 105.08 61.36 ;
    RECT 104.87 61.65 105.08 61.72 ;
    RECT 104.87 62.01 105.08 62.08 ;
    RECT 101.09 61.29 101.3 61.36 ;
    RECT 101.09 61.65 101.3 61.72 ;
    RECT 101.09 62.01 101.3 62.08 ;
    RECT 101.55 61.29 101.76 61.36 ;
    RECT 101.55 61.65 101.76 61.72 ;
    RECT 101.55 62.01 101.76 62.08 ;
    RECT 97.77 61.29 97.98 61.36 ;
    RECT 97.77 61.65 97.98 61.72 ;
    RECT 97.77 62.01 97.98 62.08 ;
    RECT 98.23 61.29 98.44 61.36 ;
    RECT 98.23 61.65 98.44 61.72 ;
    RECT 98.23 62.01 98.44 62.08 ;
    RECT 94.45 61.29 94.66 61.36 ;
    RECT 94.45 61.65 94.66 61.72 ;
    RECT 94.45 62.01 94.66 62.08 ;
    RECT 94.91 61.29 95.12 61.36 ;
    RECT 94.91 61.65 95.12 61.72 ;
    RECT 94.91 62.01 95.12 62.08 ;
    RECT 91.13 61.29 91.34 61.36 ;
    RECT 91.13 61.65 91.34 61.72 ;
    RECT 91.13 62.01 91.34 62.08 ;
    RECT 91.59 61.29 91.8 61.36 ;
    RECT 91.59 61.65 91.8 61.72 ;
    RECT 91.59 62.01 91.8 62.08 ;
    RECT 87.81 61.29 88.02 61.36 ;
    RECT 87.81 61.65 88.02 61.72 ;
    RECT 87.81 62.01 88.02 62.08 ;
    RECT 88.27 61.29 88.48 61.36 ;
    RECT 88.27 61.65 88.48 61.72 ;
    RECT 88.27 62.01 88.48 62.08 ;
    RECT 84.49 61.29 84.7 61.36 ;
    RECT 84.49 61.65 84.7 61.72 ;
    RECT 84.49 62.01 84.7 62.08 ;
    RECT 84.95 61.29 85.16 61.36 ;
    RECT 84.95 61.65 85.16 61.72 ;
    RECT 84.95 62.01 85.16 62.08 ;
    RECT 81.17 61.29 81.38 61.36 ;
    RECT 81.17 61.65 81.38 61.72 ;
    RECT 81.17 62.01 81.38 62.08 ;
    RECT 81.63 61.29 81.84 61.36 ;
    RECT 81.63 61.65 81.84 61.72 ;
    RECT 81.63 62.01 81.84 62.08 ;
    RECT 77.85 61.29 78.06 61.36 ;
    RECT 77.85 61.65 78.06 61.72 ;
    RECT 77.85 62.01 78.06 62.08 ;
    RECT 78.31 61.29 78.52 61.36 ;
    RECT 78.31 61.65 78.52 61.72 ;
    RECT 78.31 62.01 78.52 62.08 ;
    RECT 74.53 61.29 74.74 61.36 ;
    RECT 74.53 61.65 74.74 61.72 ;
    RECT 74.53 62.01 74.74 62.08 ;
    RECT 74.99 61.29 75.2 61.36 ;
    RECT 74.99 61.65 75.2 61.72 ;
    RECT 74.99 62.01 75.2 62.08 ;
    RECT 71.21 61.29 71.42 61.36 ;
    RECT 71.21 61.65 71.42 61.72 ;
    RECT 71.21 62.01 71.42 62.08 ;
    RECT 71.67 61.29 71.88 61.36 ;
    RECT 71.67 61.65 71.88 61.72 ;
    RECT 71.67 62.01 71.88 62.08 ;
    RECT 31.37 61.29 31.58 61.36 ;
    RECT 31.37 61.65 31.58 61.72 ;
    RECT 31.37 62.01 31.58 62.08 ;
    RECT 31.83 61.29 32.04 61.36 ;
    RECT 31.83 61.65 32.04 61.72 ;
    RECT 31.83 62.01 32.04 62.08 ;
    RECT 67.89 61.29 68.1 61.36 ;
    RECT 67.89 61.65 68.1 61.72 ;
    RECT 67.89 62.01 68.1 62.08 ;
    RECT 68.35 61.29 68.56 61.36 ;
    RECT 68.35 61.65 68.56 61.72 ;
    RECT 68.35 62.01 68.56 62.08 ;
    RECT 28.05 61.29 28.26 61.36 ;
    RECT 28.05 61.65 28.26 61.72 ;
    RECT 28.05 62.01 28.26 62.08 ;
    RECT 28.51 61.29 28.72 61.36 ;
    RECT 28.51 61.65 28.72 61.72 ;
    RECT 28.51 62.01 28.72 62.08 ;
    RECT 24.73 61.29 24.94 61.36 ;
    RECT 24.73 61.65 24.94 61.72 ;
    RECT 24.73 62.01 24.94 62.08 ;
    RECT 25.19 61.29 25.4 61.36 ;
    RECT 25.19 61.65 25.4 61.72 ;
    RECT 25.19 62.01 25.4 62.08 ;
    RECT 21.41 61.29 21.62 61.36 ;
    RECT 21.41 61.65 21.62 61.72 ;
    RECT 21.41 62.01 21.62 62.08 ;
    RECT 21.87 61.29 22.08 61.36 ;
    RECT 21.87 61.65 22.08 61.72 ;
    RECT 21.87 62.01 22.08 62.08 ;
    RECT 18.09 61.29 18.3 61.36 ;
    RECT 18.09 61.65 18.3 61.72 ;
    RECT 18.09 62.01 18.3 62.08 ;
    RECT 18.55 61.29 18.76 61.36 ;
    RECT 18.55 61.65 18.76 61.72 ;
    RECT 18.55 62.01 18.76 62.08 ;
    RECT 120.825 61.65 120.895 61.72 ;
    RECT 14.77 61.29 14.98 61.36 ;
    RECT 14.77 61.65 14.98 61.72 ;
    RECT 14.77 62.01 14.98 62.08 ;
    RECT 15.23 61.29 15.44 61.36 ;
    RECT 15.23 61.65 15.44 61.72 ;
    RECT 15.23 62.01 15.44 62.08 ;
    RECT 11.45 61.29 11.66 61.36 ;
    RECT 11.45 61.65 11.66 61.72 ;
    RECT 11.45 62.01 11.66 62.08 ;
    RECT 11.91 61.29 12.12 61.36 ;
    RECT 11.91 61.65 12.12 61.72 ;
    RECT 11.91 62.01 12.12 62.08 ;
    RECT 8.13 61.29 8.34 61.36 ;
    RECT 8.13 61.65 8.34 61.72 ;
    RECT 8.13 62.01 8.34 62.08 ;
    RECT 8.59 61.29 8.8 61.36 ;
    RECT 8.59 61.65 8.8 61.72 ;
    RECT 8.59 62.01 8.8 62.08 ;
    RECT 4.81 61.29 5.02 61.36 ;
    RECT 4.81 61.65 5.02 61.72 ;
    RECT 4.81 62.01 5.02 62.08 ;
    RECT 5.27 61.29 5.48 61.36 ;
    RECT 5.27 61.65 5.48 61.72 ;
    RECT 5.27 62.01 5.48 62.08 ;
    RECT 1.49 61.29 1.7 61.36 ;
    RECT 1.49 61.65 1.7 61.72 ;
    RECT 1.49 62.01 1.7 62.08 ;
    RECT 1.95 61.29 2.16 61.36 ;
    RECT 1.95 61.65 2.16 61.72 ;
    RECT 1.95 62.01 2.16 62.08 ;
    RECT 64.57 61.29 64.78 61.36 ;
    RECT 64.57 61.65 64.78 61.72 ;
    RECT 64.57 62.01 64.78 62.08 ;
    RECT 65.03 61.29 65.24 61.36 ;
    RECT 65.03 61.65 65.24 61.72 ;
    RECT 65.03 62.01 65.24 62.08 ;
    RECT 81.63 61.05 81.84 61.12 ;
    RECT 81.17 61.05 81.38 61.12 ;
    RECT 78.8 60.79 79.01 60.86 ;
    RECT 35.15 61.05 35.36 61.12 ;
    RECT 118.15 61.05 118.36 61.12 ;
    RECT 34.69 61.05 34.9 61.12 ;
    RECT 117.69 61.05 117.9 61.12 ;
    RECT 57.93 61.05 58.14 61.12 ;
    RECT 21.87 61.05 22.08 61.12 ;
    RECT 21.41 61.05 21.62 61.12 ;
    RECT 48.92 60.79 49.13 60.86 ;
    RECT 68.84 60.79 69.05 60.86 ;
    RECT 19.04 60.79 19.25 60.86 ;
    RECT 74.99 61.05 75.2 61.12 ;
    RECT 98.23 61.05 98.44 61.12 ;
    RECT 97.77 61.05 97.98 61.12 ;
    RECT 115.32 60.79 115.53 60.86 ;
    RECT 111.51 61.05 111.72 61.12 ;
    RECT 111.05 61.05 111.26 61.12 ;
    RECT 51.75 61.05 51.96 61.12 ;
    RECT 51.29 61.05 51.5 61.12 ;
    RECT 15.23 61.05 15.44 61.12 ;
    RECT 14.77 61.05 14.98 61.12 ;
    RECT 74.53 61.05 74.74 61.12 ;
    RECT 42.28 60.79 42.49 60.86 ;
    RECT 12.4 60.79 12.61 60.86 ;
    RECT 95.4 60.79 95.61 60.86 ;
    RECT 91.59 61.05 91.8 61.12 ;
    RECT 31.83 61.05 32.04 61.12 ;
    RECT 31.37 61.05 31.58 61.12 ;
    RECT 108.68 60.79 108.89 60.86 ;
    RECT 121.035 60.79 121.105 60.86 ;
    RECT 120.825 61.05 120.895 61.12 ;
    RECT 45.11 61.05 45.32 61.12 ;
    RECT 44.65 61.05 44.86 61.12 ;
    RECT 0.19 60.79 0.26 60.86 ;
    RECT 0.4 61.05 0.47 61.12 ;
    RECT 8.59 61.05 8.8 61.12 ;
    RECT 65.52 60.79 65.73 60.86 ;
    RECT 68.35 61.05 68.56 61.12 ;
    RECT 67.89 61.05 68.1 61.12 ;
    RECT 91.13 61.05 91.34 61.12 ;
    RECT 5.76 60.79 5.97 60.86 ;
    RECT 88.76 60.79 88.97 60.86 ;
    RECT 104.87 61.05 105.08 61.12 ;
    RECT 104.41 61.05 104.62 61.12 ;
    RECT 8.13 61.05 8.34 61.12 ;
    RECT 25.19 61.05 25.4 61.12 ;
    RECT 35.64 60.79 35.85 60.86 ;
    RECT 58.88 60.79 59.09 60.86 ;
    RECT 61.71 61.05 61.92 61.12 ;
    RECT 29.0 60.79 29.21 60.86 ;
    RECT 61.25 61.05 61.46 61.12 ;
    RECT 84.95 61.05 85.16 61.12 ;
    RECT 84.49 61.05 84.7 61.12 ;
    RECT 102.04 60.79 102.25 60.86 ;
    RECT 82.12 60.79 82.33 60.86 ;
    RECT 72.16 60.79 72.37 60.86 ;
    RECT 38.47 61.05 38.68 61.12 ;
    RECT 38.01 61.05 38.22 61.12 ;
    RECT 1.95 61.05 2.16 61.12 ;
    RECT 1.49 61.05 1.7 61.12 ;
    RECT 24.73 61.05 24.94 61.12 ;
    RECT 52.24 60.79 52.45 60.86 ;
    RECT 22.36 60.79 22.57 60.86 ;
    RECT 78.31 61.05 78.52 61.12 ;
    RECT 77.85 61.05 78.06 61.12 ;
    RECT 118.64 60.79 118.85 60.86 ;
    RECT 114.83 61.05 115.04 61.12 ;
    RECT 114.37 61.05 114.58 61.12 ;
    RECT 55.07 61.05 55.28 61.12 ;
    RECT 54.61 61.05 54.82 61.12 ;
    RECT 18.55 61.05 18.76 61.12 ;
    RECT 18.09 61.05 18.3 61.12 ;
    RECT 45.6 60.79 45.81 60.86 ;
    RECT 15.72 60.79 15.93 60.86 ;
    RECT 98.72 60.79 98.93 60.86 ;
    RECT 94.91 61.05 95.12 61.12 ;
    RECT 94.45 61.05 94.66 61.12 ;
    RECT 112.0 60.79 112.21 60.86 ;
    RECT 108.19 61.05 108.4 61.12 ;
    RECT 48.43 61.05 48.64 61.12 ;
    RECT 47.97 61.05 48.18 61.12 ;
    RECT 11.91 61.05 12.12 61.12 ;
    RECT 71.67 61.05 71.88 61.12 ;
    RECT 11.45 61.05 11.66 61.12 ;
    RECT 71.21 61.05 71.42 61.12 ;
    RECT 38.96 60.79 39.17 60.86 ;
    RECT 9.08 60.79 9.29 60.86 ;
    RECT 92.08 60.79 92.29 60.86 ;
    RECT 107.73 61.05 107.94 61.12 ;
    RECT 28.51 61.05 28.72 61.12 ;
    RECT 28.05 61.05 28.26 61.12 ;
    RECT 105.36 60.79 105.57 60.86 ;
    RECT 41.79 61.05 42.0 61.12 ;
    RECT 65.03 61.05 65.24 61.12 ;
    RECT 64.57 61.05 64.78 61.12 ;
    RECT 62.2 60.79 62.41 60.86 ;
    RECT 32.32 60.79 32.53 60.86 ;
    RECT 88.27 61.05 88.48 61.12 ;
    RECT 87.81 61.05 88.02 61.12 ;
    RECT 85.44 60.79 85.65 60.86 ;
    RECT 101.55 61.05 101.76 61.12 ;
    RECT 75.48 60.79 75.69 60.86 ;
    RECT 101.09 61.05 101.3 61.12 ;
    RECT 41.33 61.05 41.54 61.12 ;
    RECT 5.27 61.05 5.48 61.12 ;
    RECT 4.81 61.05 5.02 61.12 ;
    RECT 2.44 60.79 2.65 60.86 ;
    RECT 55.56 60.79 55.77 60.86 ;
    RECT 58.39 61.05 58.6 61.12 ;
    RECT 25.68 60.79 25.89 60.86 ;
    RECT 61.25 59.83 61.46 59.9 ;
    RECT 61.25 60.19 61.46 60.26 ;
    RECT 61.25 60.55 61.46 60.62 ;
    RECT 61.71 59.83 61.92 59.9 ;
    RECT 61.71 60.19 61.92 60.26 ;
    RECT 61.71 60.55 61.92 60.62 ;
    RECT 57.93 59.83 58.14 59.9 ;
    RECT 57.93 60.19 58.14 60.26 ;
    RECT 57.93 60.55 58.14 60.62 ;
    RECT 58.39 59.83 58.6 59.9 ;
    RECT 58.39 60.19 58.6 60.26 ;
    RECT 58.39 60.55 58.6 60.62 ;
    RECT 54.61 59.83 54.82 59.9 ;
    RECT 54.61 60.19 54.82 60.26 ;
    RECT 54.61 60.55 54.82 60.62 ;
    RECT 55.07 59.83 55.28 59.9 ;
    RECT 55.07 60.19 55.28 60.26 ;
    RECT 55.07 60.55 55.28 60.62 ;
    RECT 51.29 59.83 51.5 59.9 ;
    RECT 51.29 60.19 51.5 60.26 ;
    RECT 51.29 60.55 51.5 60.62 ;
    RECT 51.75 59.83 51.96 59.9 ;
    RECT 51.75 60.19 51.96 60.26 ;
    RECT 51.75 60.55 51.96 60.62 ;
    RECT 47.97 59.83 48.18 59.9 ;
    RECT 47.97 60.19 48.18 60.26 ;
    RECT 47.97 60.55 48.18 60.62 ;
    RECT 48.43 59.83 48.64 59.9 ;
    RECT 48.43 60.19 48.64 60.26 ;
    RECT 48.43 60.55 48.64 60.62 ;
    RECT 44.65 59.83 44.86 59.9 ;
    RECT 44.65 60.19 44.86 60.26 ;
    RECT 44.65 60.55 44.86 60.62 ;
    RECT 45.11 59.83 45.32 59.9 ;
    RECT 45.11 60.19 45.32 60.26 ;
    RECT 45.11 60.55 45.32 60.62 ;
    RECT 41.33 59.83 41.54 59.9 ;
    RECT 41.33 60.19 41.54 60.26 ;
    RECT 41.33 60.55 41.54 60.62 ;
    RECT 41.79 59.83 42.0 59.9 ;
    RECT 41.79 60.19 42.0 60.26 ;
    RECT 41.79 60.55 42.0 60.62 ;
    RECT 38.01 59.83 38.22 59.9 ;
    RECT 38.01 60.19 38.22 60.26 ;
    RECT 38.01 60.55 38.22 60.62 ;
    RECT 38.47 59.83 38.68 59.9 ;
    RECT 38.47 60.19 38.68 60.26 ;
    RECT 38.47 60.55 38.68 60.62 ;
    RECT 0.4 60.19 0.47 60.26 ;
    RECT 34.69 59.83 34.9 59.9 ;
    RECT 34.69 60.19 34.9 60.26 ;
    RECT 34.69 60.55 34.9 60.62 ;
    RECT 35.15 59.83 35.36 59.9 ;
    RECT 35.15 60.19 35.36 60.26 ;
    RECT 35.15 60.55 35.36 60.62 ;
    RECT 117.69 59.83 117.9 59.9 ;
    RECT 117.69 60.19 117.9 60.26 ;
    RECT 117.69 60.55 117.9 60.62 ;
    RECT 118.15 59.83 118.36 59.9 ;
    RECT 118.15 60.19 118.36 60.26 ;
    RECT 118.15 60.55 118.36 60.62 ;
    RECT 114.37 59.83 114.58 59.9 ;
    RECT 114.37 60.19 114.58 60.26 ;
    RECT 114.37 60.55 114.58 60.62 ;
    RECT 114.83 59.83 115.04 59.9 ;
    RECT 114.83 60.19 115.04 60.26 ;
    RECT 114.83 60.55 115.04 60.62 ;
    RECT 111.05 59.83 111.26 59.9 ;
    RECT 111.05 60.19 111.26 60.26 ;
    RECT 111.05 60.55 111.26 60.62 ;
    RECT 111.51 59.83 111.72 59.9 ;
    RECT 111.51 60.19 111.72 60.26 ;
    RECT 111.51 60.55 111.72 60.62 ;
    RECT 107.73 59.83 107.94 59.9 ;
    RECT 107.73 60.19 107.94 60.26 ;
    RECT 107.73 60.55 107.94 60.62 ;
    RECT 108.19 59.83 108.4 59.9 ;
    RECT 108.19 60.19 108.4 60.26 ;
    RECT 108.19 60.55 108.4 60.62 ;
    RECT 104.41 59.83 104.62 59.9 ;
    RECT 104.41 60.19 104.62 60.26 ;
    RECT 104.41 60.55 104.62 60.62 ;
    RECT 104.87 59.83 105.08 59.9 ;
    RECT 104.87 60.19 105.08 60.26 ;
    RECT 104.87 60.55 105.08 60.62 ;
    RECT 101.09 59.83 101.3 59.9 ;
    RECT 101.09 60.19 101.3 60.26 ;
    RECT 101.09 60.55 101.3 60.62 ;
    RECT 101.55 59.83 101.76 59.9 ;
    RECT 101.55 60.19 101.76 60.26 ;
    RECT 101.55 60.55 101.76 60.62 ;
    RECT 97.77 59.83 97.98 59.9 ;
    RECT 97.77 60.19 97.98 60.26 ;
    RECT 97.77 60.55 97.98 60.62 ;
    RECT 98.23 59.83 98.44 59.9 ;
    RECT 98.23 60.19 98.44 60.26 ;
    RECT 98.23 60.55 98.44 60.62 ;
    RECT 94.45 59.83 94.66 59.9 ;
    RECT 94.45 60.19 94.66 60.26 ;
    RECT 94.45 60.55 94.66 60.62 ;
    RECT 94.91 59.83 95.12 59.9 ;
    RECT 94.91 60.19 95.12 60.26 ;
    RECT 94.91 60.55 95.12 60.62 ;
    RECT 91.13 59.83 91.34 59.9 ;
    RECT 91.13 60.19 91.34 60.26 ;
    RECT 91.13 60.55 91.34 60.62 ;
    RECT 91.59 59.83 91.8 59.9 ;
    RECT 91.59 60.19 91.8 60.26 ;
    RECT 91.59 60.55 91.8 60.62 ;
    RECT 87.81 59.83 88.02 59.9 ;
    RECT 87.81 60.19 88.02 60.26 ;
    RECT 87.81 60.55 88.02 60.62 ;
    RECT 88.27 59.83 88.48 59.9 ;
    RECT 88.27 60.19 88.48 60.26 ;
    RECT 88.27 60.55 88.48 60.62 ;
    RECT 84.49 59.83 84.7 59.9 ;
    RECT 84.49 60.19 84.7 60.26 ;
    RECT 84.49 60.55 84.7 60.62 ;
    RECT 84.95 59.83 85.16 59.9 ;
    RECT 84.95 60.19 85.16 60.26 ;
    RECT 84.95 60.55 85.16 60.62 ;
    RECT 81.17 59.83 81.38 59.9 ;
    RECT 81.17 60.19 81.38 60.26 ;
    RECT 81.17 60.55 81.38 60.62 ;
    RECT 81.63 59.83 81.84 59.9 ;
    RECT 81.63 60.19 81.84 60.26 ;
    RECT 81.63 60.55 81.84 60.62 ;
    RECT 77.85 59.83 78.06 59.9 ;
    RECT 77.85 60.19 78.06 60.26 ;
    RECT 77.85 60.55 78.06 60.62 ;
    RECT 78.31 59.83 78.52 59.9 ;
    RECT 78.31 60.19 78.52 60.26 ;
    RECT 78.31 60.55 78.52 60.62 ;
    RECT 74.53 59.83 74.74 59.9 ;
    RECT 74.53 60.19 74.74 60.26 ;
    RECT 74.53 60.55 74.74 60.62 ;
    RECT 74.99 59.83 75.2 59.9 ;
    RECT 74.99 60.19 75.2 60.26 ;
    RECT 74.99 60.55 75.2 60.62 ;
    RECT 71.21 59.83 71.42 59.9 ;
    RECT 71.21 60.19 71.42 60.26 ;
    RECT 71.21 60.55 71.42 60.62 ;
    RECT 71.67 59.83 71.88 59.9 ;
    RECT 71.67 60.19 71.88 60.26 ;
    RECT 71.67 60.55 71.88 60.62 ;
    RECT 31.37 59.83 31.58 59.9 ;
    RECT 31.37 60.19 31.58 60.26 ;
    RECT 31.37 60.55 31.58 60.62 ;
    RECT 31.83 59.83 32.04 59.9 ;
    RECT 31.83 60.19 32.04 60.26 ;
    RECT 31.83 60.55 32.04 60.62 ;
    RECT 67.89 59.83 68.1 59.9 ;
    RECT 67.89 60.19 68.1 60.26 ;
    RECT 67.89 60.55 68.1 60.62 ;
    RECT 68.35 59.83 68.56 59.9 ;
    RECT 68.35 60.19 68.56 60.26 ;
    RECT 68.35 60.55 68.56 60.62 ;
    RECT 28.05 59.83 28.26 59.9 ;
    RECT 28.05 60.19 28.26 60.26 ;
    RECT 28.05 60.55 28.26 60.62 ;
    RECT 28.51 59.83 28.72 59.9 ;
    RECT 28.51 60.19 28.72 60.26 ;
    RECT 28.51 60.55 28.72 60.62 ;
    RECT 24.73 59.83 24.94 59.9 ;
    RECT 24.73 60.19 24.94 60.26 ;
    RECT 24.73 60.55 24.94 60.62 ;
    RECT 25.19 59.83 25.4 59.9 ;
    RECT 25.19 60.19 25.4 60.26 ;
    RECT 25.19 60.55 25.4 60.62 ;
    RECT 21.41 59.83 21.62 59.9 ;
    RECT 21.41 60.19 21.62 60.26 ;
    RECT 21.41 60.55 21.62 60.62 ;
    RECT 21.87 59.83 22.08 59.9 ;
    RECT 21.87 60.19 22.08 60.26 ;
    RECT 21.87 60.55 22.08 60.62 ;
    RECT 18.09 59.83 18.3 59.9 ;
    RECT 18.09 60.19 18.3 60.26 ;
    RECT 18.09 60.55 18.3 60.62 ;
    RECT 18.55 59.83 18.76 59.9 ;
    RECT 18.55 60.19 18.76 60.26 ;
    RECT 18.55 60.55 18.76 60.62 ;
    RECT 120.825 60.19 120.895 60.26 ;
    RECT 14.77 59.83 14.98 59.9 ;
    RECT 14.77 60.19 14.98 60.26 ;
    RECT 14.77 60.55 14.98 60.62 ;
    RECT 15.23 59.83 15.44 59.9 ;
    RECT 15.23 60.19 15.44 60.26 ;
    RECT 15.23 60.55 15.44 60.62 ;
    RECT 11.45 59.83 11.66 59.9 ;
    RECT 11.45 60.19 11.66 60.26 ;
    RECT 11.45 60.55 11.66 60.62 ;
    RECT 11.91 59.83 12.12 59.9 ;
    RECT 11.91 60.19 12.12 60.26 ;
    RECT 11.91 60.55 12.12 60.62 ;
    RECT 8.13 59.83 8.34 59.9 ;
    RECT 8.13 60.19 8.34 60.26 ;
    RECT 8.13 60.55 8.34 60.62 ;
    RECT 8.59 59.83 8.8 59.9 ;
    RECT 8.59 60.19 8.8 60.26 ;
    RECT 8.59 60.55 8.8 60.62 ;
    RECT 4.81 59.83 5.02 59.9 ;
    RECT 4.81 60.19 5.02 60.26 ;
    RECT 4.81 60.55 5.02 60.62 ;
    RECT 5.27 59.83 5.48 59.9 ;
    RECT 5.27 60.19 5.48 60.26 ;
    RECT 5.27 60.55 5.48 60.62 ;
    RECT 1.49 59.83 1.7 59.9 ;
    RECT 1.49 60.19 1.7 60.26 ;
    RECT 1.49 60.55 1.7 60.62 ;
    RECT 1.95 59.83 2.16 59.9 ;
    RECT 1.95 60.19 2.16 60.26 ;
    RECT 1.95 60.55 2.16 60.62 ;
    RECT 64.57 59.83 64.78 59.9 ;
    RECT 64.57 60.19 64.78 60.26 ;
    RECT 64.57 60.55 64.78 60.62 ;
    RECT 65.03 59.83 65.24 59.9 ;
    RECT 65.03 60.19 65.24 60.26 ;
    RECT 65.03 60.55 65.24 60.62 ;
    RECT 61.25 59.11 61.46 59.18 ;
    RECT 61.25 59.47 61.46 59.54 ;
    RECT 61.25 59.83 61.46 59.9 ;
    RECT 61.71 59.11 61.92 59.18 ;
    RECT 61.71 59.47 61.92 59.54 ;
    RECT 61.71 59.83 61.92 59.9 ;
    RECT 57.93 59.11 58.14 59.18 ;
    RECT 57.93 59.47 58.14 59.54 ;
    RECT 57.93 59.83 58.14 59.9 ;
    RECT 58.39 59.11 58.6 59.18 ;
    RECT 58.39 59.47 58.6 59.54 ;
    RECT 58.39 59.83 58.6 59.9 ;
    RECT 54.61 59.11 54.82 59.18 ;
    RECT 54.61 59.47 54.82 59.54 ;
    RECT 54.61 59.83 54.82 59.9 ;
    RECT 55.07 59.11 55.28 59.18 ;
    RECT 55.07 59.47 55.28 59.54 ;
    RECT 55.07 59.83 55.28 59.9 ;
    RECT 51.29 59.11 51.5 59.18 ;
    RECT 51.29 59.47 51.5 59.54 ;
    RECT 51.29 59.83 51.5 59.9 ;
    RECT 51.75 59.11 51.96 59.18 ;
    RECT 51.75 59.47 51.96 59.54 ;
    RECT 51.75 59.83 51.96 59.9 ;
    RECT 47.97 59.11 48.18 59.18 ;
    RECT 47.97 59.47 48.18 59.54 ;
    RECT 47.97 59.83 48.18 59.9 ;
    RECT 48.43 59.11 48.64 59.18 ;
    RECT 48.43 59.47 48.64 59.54 ;
    RECT 48.43 59.83 48.64 59.9 ;
    RECT 44.65 59.11 44.86 59.18 ;
    RECT 44.65 59.47 44.86 59.54 ;
    RECT 44.65 59.83 44.86 59.9 ;
    RECT 45.11 59.11 45.32 59.18 ;
    RECT 45.11 59.47 45.32 59.54 ;
    RECT 45.11 59.83 45.32 59.9 ;
    RECT 41.33 59.11 41.54 59.18 ;
    RECT 41.33 59.47 41.54 59.54 ;
    RECT 41.33 59.83 41.54 59.9 ;
    RECT 41.79 59.11 42.0 59.18 ;
    RECT 41.79 59.47 42.0 59.54 ;
    RECT 41.79 59.83 42.0 59.9 ;
    RECT 38.01 59.11 38.22 59.18 ;
    RECT 38.01 59.47 38.22 59.54 ;
    RECT 38.01 59.83 38.22 59.9 ;
    RECT 38.47 59.11 38.68 59.18 ;
    RECT 38.47 59.47 38.68 59.54 ;
    RECT 38.47 59.83 38.68 59.9 ;
    RECT 0.4 59.47 0.47 59.54 ;
    RECT 34.69 59.11 34.9 59.18 ;
    RECT 34.69 59.47 34.9 59.54 ;
    RECT 34.69 59.83 34.9 59.9 ;
    RECT 35.15 59.11 35.36 59.18 ;
    RECT 35.15 59.47 35.36 59.54 ;
    RECT 35.15 59.83 35.36 59.9 ;
    RECT 117.69 59.11 117.9 59.18 ;
    RECT 117.69 59.47 117.9 59.54 ;
    RECT 117.69 59.83 117.9 59.9 ;
    RECT 118.15 59.11 118.36 59.18 ;
    RECT 118.15 59.47 118.36 59.54 ;
    RECT 118.15 59.83 118.36 59.9 ;
    RECT 114.37 59.11 114.58 59.18 ;
    RECT 114.37 59.47 114.58 59.54 ;
    RECT 114.37 59.83 114.58 59.9 ;
    RECT 114.83 59.11 115.04 59.18 ;
    RECT 114.83 59.47 115.04 59.54 ;
    RECT 114.83 59.83 115.04 59.9 ;
    RECT 111.05 59.11 111.26 59.18 ;
    RECT 111.05 59.47 111.26 59.54 ;
    RECT 111.05 59.83 111.26 59.9 ;
    RECT 111.51 59.11 111.72 59.18 ;
    RECT 111.51 59.47 111.72 59.54 ;
    RECT 111.51 59.83 111.72 59.9 ;
    RECT 107.73 59.11 107.94 59.18 ;
    RECT 107.73 59.47 107.94 59.54 ;
    RECT 107.73 59.83 107.94 59.9 ;
    RECT 108.19 59.11 108.4 59.18 ;
    RECT 108.19 59.47 108.4 59.54 ;
    RECT 108.19 59.83 108.4 59.9 ;
    RECT 104.41 59.11 104.62 59.18 ;
    RECT 104.41 59.47 104.62 59.54 ;
    RECT 104.41 59.83 104.62 59.9 ;
    RECT 104.87 59.11 105.08 59.18 ;
    RECT 104.87 59.47 105.08 59.54 ;
    RECT 104.87 59.83 105.08 59.9 ;
    RECT 101.09 59.11 101.3 59.18 ;
    RECT 101.09 59.47 101.3 59.54 ;
    RECT 101.09 59.83 101.3 59.9 ;
    RECT 101.55 59.11 101.76 59.18 ;
    RECT 101.55 59.47 101.76 59.54 ;
    RECT 101.55 59.83 101.76 59.9 ;
    RECT 97.77 59.11 97.98 59.18 ;
    RECT 97.77 59.47 97.98 59.54 ;
    RECT 97.77 59.83 97.98 59.9 ;
    RECT 98.23 59.11 98.44 59.18 ;
    RECT 98.23 59.47 98.44 59.54 ;
    RECT 98.23 59.83 98.44 59.9 ;
    RECT 94.45 59.11 94.66 59.18 ;
    RECT 94.45 59.47 94.66 59.54 ;
    RECT 94.45 59.83 94.66 59.9 ;
    RECT 94.91 59.11 95.12 59.18 ;
    RECT 94.91 59.47 95.12 59.54 ;
    RECT 94.91 59.83 95.12 59.9 ;
    RECT 91.13 59.11 91.34 59.18 ;
    RECT 91.13 59.47 91.34 59.54 ;
    RECT 91.13 59.83 91.34 59.9 ;
    RECT 91.59 59.11 91.8 59.18 ;
    RECT 91.59 59.47 91.8 59.54 ;
    RECT 91.59 59.83 91.8 59.9 ;
    RECT 87.81 59.11 88.02 59.18 ;
    RECT 87.81 59.47 88.02 59.54 ;
    RECT 87.81 59.83 88.02 59.9 ;
    RECT 88.27 59.11 88.48 59.18 ;
    RECT 88.27 59.47 88.48 59.54 ;
    RECT 88.27 59.83 88.48 59.9 ;
    RECT 84.49 59.11 84.7 59.18 ;
    RECT 84.49 59.47 84.7 59.54 ;
    RECT 84.49 59.83 84.7 59.9 ;
    RECT 84.95 59.11 85.16 59.18 ;
    RECT 84.95 59.47 85.16 59.54 ;
    RECT 84.95 59.83 85.16 59.9 ;
    RECT 81.17 59.11 81.38 59.18 ;
    RECT 81.17 59.47 81.38 59.54 ;
    RECT 81.17 59.83 81.38 59.9 ;
    RECT 81.63 59.11 81.84 59.18 ;
    RECT 81.63 59.47 81.84 59.54 ;
    RECT 81.63 59.83 81.84 59.9 ;
    RECT 77.85 59.11 78.06 59.18 ;
    RECT 77.85 59.47 78.06 59.54 ;
    RECT 77.85 59.83 78.06 59.9 ;
    RECT 78.31 59.11 78.52 59.18 ;
    RECT 78.31 59.47 78.52 59.54 ;
    RECT 78.31 59.83 78.52 59.9 ;
    RECT 74.53 59.11 74.74 59.18 ;
    RECT 74.53 59.47 74.74 59.54 ;
    RECT 74.53 59.83 74.74 59.9 ;
    RECT 74.99 59.11 75.2 59.18 ;
    RECT 74.99 59.47 75.2 59.54 ;
    RECT 74.99 59.83 75.2 59.9 ;
    RECT 71.21 59.11 71.42 59.18 ;
    RECT 71.21 59.47 71.42 59.54 ;
    RECT 71.21 59.83 71.42 59.9 ;
    RECT 71.67 59.11 71.88 59.18 ;
    RECT 71.67 59.47 71.88 59.54 ;
    RECT 71.67 59.83 71.88 59.9 ;
    RECT 31.37 59.11 31.58 59.18 ;
    RECT 31.37 59.47 31.58 59.54 ;
    RECT 31.37 59.83 31.58 59.9 ;
    RECT 31.83 59.11 32.04 59.18 ;
    RECT 31.83 59.47 32.04 59.54 ;
    RECT 31.83 59.83 32.04 59.9 ;
    RECT 67.89 59.11 68.1 59.18 ;
    RECT 67.89 59.47 68.1 59.54 ;
    RECT 67.89 59.83 68.1 59.9 ;
    RECT 68.35 59.11 68.56 59.18 ;
    RECT 68.35 59.47 68.56 59.54 ;
    RECT 68.35 59.83 68.56 59.9 ;
    RECT 28.05 59.11 28.26 59.18 ;
    RECT 28.05 59.47 28.26 59.54 ;
    RECT 28.05 59.83 28.26 59.9 ;
    RECT 28.51 59.11 28.72 59.18 ;
    RECT 28.51 59.47 28.72 59.54 ;
    RECT 28.51 59.83 28.72 59.9 ;
    RECT 24.73 59.11 24.94 59.18 ;
    RECT 24.73 59.47 24.94 59.54 ;
    RECT 24.73 59.83 24.94 59.9 ;
    RECT 25.19 59.11 25.4 59.18 ;
    RECT 25.19 59.47 25.4 59.54 ;
    RECT 25.19 59.83 25.4 59.9 ;
    RECT 21.41 59.11 21.62 59.18 ;
    RECT 21.41 59.47 21.62 59.54 ;
    RECT 21.41 59.83 21.62 59.9 ;
    RECT 21.87 59.11 22.08 59.18 ;
    RECT 21.87 59.47 22.08 59.54 ;
    RECT 21.87 59.83 22.08 59.9 ;
    RECT 18.09 59.11 18.3 59.18 ;
    RECT 18.09 59.47 18.3 59.54 ;
    RECT 18.09 59.83 18.3 59.9 ;
    RECT 18.55 59.11 18.76 59.18 ;
    RECT 18.55 59.47 18.76 59.54 ;
    RECT 18.55 59.83 18.76 59.9 ;
    RECT 120.825 59.47 120.895 59.54 ;
    RECT 14.77 59.11 14.98 59.18 ;
    RECT 14.77 59.47 14.98 59.54 ;
    RECT 14.77 59.83 14.98 59.9 ;
    RECT 15.23 59.11 15.44 59.18 ;
    RECT 15.23 59.47 15.44 59.54 ;
    RECT 15.23 59.83 15.44 59.9 ;
    RECT 11.45 59.11 11.66 59.18 ;
    RECT 11.45 59.47 11.66 59.54 ;
    RECT 11.45 59.83 11.66 59.9 ;
    RECT 11.91 59.11 12.12 59.18 ;
    RECT 11.91 59.47 12.12 59.54 ;
    RECT 11.91 59.83 12.12 59.9 ;
    RECT 8.13 59.11 8.34 59.18 ;
    RECT 8.13 59.47 8.34 59.54 ;
    RECT 8.13 59.83 8.34 59.9 ;
    RECT 8.59 59.11 8.8 59.18 ;
    RECT 8.59 59.47 8.8 59.54 ;
    RECT 8.59 59.83 8.8 59.9 ;
    RECT 4.81 59.11 5.02 59.18 ;
    RECT 4.81 59.47 5.02 59.54 ;
    RECT 4.81 59.83 5.02 59.9 ;
    RECT 5.27 59.11 5.48 59.18 ;
    RECT 5.27 59.47 5.48 59.54 ;
    RECT 5.27 59.83 5.48 59.9 ;
    RECT 1.49 59.11 1.7 59.18 ;
    RECT 1.49 59.47 1.7 59.54 ;
    RECT 1.49 59.83 1.7 59.9 ;
    RECT 1.95 59.11 2.16 59.18 ;
    RECT 1.95 59.47 2.16 59.54 ;
    RECT 1.95 59.83 2.16 59.9 ;
    RECT 64.57 59.11 64.78 59.18 ;
    RECT 64.57 59.47 64.78 59.54 ;
    RECT 64.57 59.83 64.78 59.9 ;
    RECT 65.03 59.11 65.24 59.18 ;
    RECT 65.03 59.47 65.24 59.54 ;
    RECT 65.03 59.83 65.24 59.9 ;
    RECT 61.25 58.39 61.46 58.46 ;
    RECT 61.25 58.75 61.46 58.82 ;
    RECT 61.25 59.11 61.46 59.18 ;
    RECT 61.71 58.39 61.92 58.46 ;
    RECT 61.71 58.75 61.92 58.82 ;
    RECT 61.71 59.11 61.92 59.18 ;
    RECT 57.93 58.39 58.14 58.46 ;
    RECT 57.93 58.75 58.14 58.82 ;
    RECT 57.93 59.11 58.14 59.18 ;
    RECT 58.39 58.39 58.6 58.46 ;
    RECT 58.39 58.75 58.6 58.82 ;
    RECT 58.39 59.11 58.6 59.18 ;
    RECT 54.61 58.39 54.82 58.46 ;
    RECT 54.61 58.75 54.82 58.82 ;
    RECT 54.61 59.11 54.82 59.18 ;
    RECT 55.07 58.39 55.28 58.46 ;
    RECT 55.07 58.75 55.28 58.82 ;
    RECT 55.07 59.11 55.28 59.18 ;
    RECT 51.29 58.39 51.5 58.46 ;
    RECT 51.29 58.75 51.5 58.82 ;
    RECT 51.29 59.11 51.5 59.18 ;
    RECT 51.75 58.39 51.96 58.46 ;
    RECT 51.75 58.75 51.96 58.82 ;
    RECT 51.75 59.11 51.96 59.18 ;
    RECT 47.97 58.39 48.18 58.46 ;
    RECT 47.97 58.75 48.18 58.82 ;
    RECT 47.97 59.11 48.18 59.18 ;
    RECT 48.43 58.39 48.64 58.46 ;
    RECT 48.43 58.75 48.64 58.82 ;
    RECT 48.43 59.11 48.64 59.18 ;
    RECT 44.65 58.39 44.86 58.46 ;
    RECT 44.65 58.75 44.86 58.82 ;
    RECT 44.65 59.11 44.86 59.18 ;
    RECT 45.11 58.39 45.32 58.46 ;
    RECT 45.11 58.75 45.32 58.82 ;
    RECT 45.11 59.11 45.32 59.18 ;
    RECT 41.33 58.39 41.54 58.46 ;
    RECT 41.33 58.75 41.54 58.82 ;
    RECT 41.33 59.11 41.54 59.18 ;
    RECT 41.79 58.39 42.0 58.46 ;
    RECT 41.79 58.75 42.0 58.82 ;
    RECT 41.79 59.11 42.0 59.18 ;
    RECT 38.01 58.39 38.22 58.46 ;
    RECT 38.01 58.75 38.22 58.82 ;
    RECT 38.01 59.11 38.22 59.18 ;
    RECT 38.47 58.39 38.68 58.46 ;
    RECT 38.47 58.75 38.68 58.82 ;
    RECT 38.47 59.11 38.68 59.18 ;
    RECT 0.4 58.75 0.47 58.82 ;
    RECT 34.69 58.39 34.9 58.46 ;
    RECT 34.69 58.75 34.9 58.82 ;
    RECT 34.69 59.11 34.9 59.18 ;
    RECT 35.15 58.39 35.36 58.46 ;
    RECT 35.15 58.75 35.36 58.82 ;
    RECT 35.15 59.11 35.36 59.18 ;
    RECT 117.69 58.39 117.9 58.46 ;
    RECT 117.69 58.75 117.9 58.82 ;
    RECT 117.69 59.11 117.9 59.18 ;
    RECT 118.15 58.39 118.36 58.46 ;
    RECT 118.15 58.75 118.36 58.82 ;
    RECT 118.15 59.11 118.36 59.18 ;
    RECT 114.37 58.39 114.58 58.46 ;
    RECT 114.37 58.75 114.58 58.82 ;
    RECT 114.37 59.11 114.58 59.18 ;
    RECT 114.83 58.39 115.04 58.46 ;
    RECT 114.83 58.75 115.04 58.82 ;
    RECT 114.83 59.11 115.04 59.18 ;
    RECT 111.05 58.39 111.26 58.46 ;
    RECT 111.05 58.75 111.26 58.82 ;
    RECT 111.05 59.11 111.26 59.18 ;
    RECT 111.51 58.39 111.72 58.46 ;
    RECT 111.51 58.75 111.72 58.82 ;
    RECT 111.51 59.11 111.72 59.18 ;
    RECT 107.73 58.39 107.94 58.46 ;
    RECT 107.73 58.75 107.94 58.82 ;
    RECT 107.73 59.11 107.94 59.18 ;
    RECT 108.19 58.39 108.4 58.46 ;
    RECT 108.19 58.75 108.4 58.82 ;
    RECT 108.19 59.11 108.4 59.18 ;
    RECT 104.41 58.39 104.62 58.46 ;
    RECT 104.41 58.75 104.62 58.82 ;
    RECT 104.41 59.11 104.62 59.18 ;
    RECT 104.87 58.39 105.08 58.46 ;
    RECT 104.87 58.75 105.08 58.82 ;
    RECT 104.87 59.11 105.08 59.18 ;
    RECT 101.09 58.39 101.3 58.46 ;
    RECT 101.09 58.75 101.3 58.82 ;
    RECT 101.09 59.11 101.3 59.18 ;
    RECT 101.55 58.39 101.76 58.46 ;
    RECT 101.55 58.75 101.76 58.82 ;
    RECT 101.55 59.11 101.76 59.18 ;
    RECT 97.77 58.39 97.98 58.46 ;
    RECT 97.77 58.75 97.98 58.82 ;
    RECT 97.77 59.11 97.98 59.18 ;
    RECT 98.23 58.39 98.44 58.46 ;
    RECT 98.23 58.75 98.44 58.82 ;
    RECT 98.23 59.11 98.44 59.18 ;
    RECT 94.45 58.39 94.66 58.46 ;
    RECT 94.45 58.75 94.66 58.82 ;
    RECT 94.45 59.11 94.66 59.18 ;
    RECT 94.91 58.39 95.12 58.46 ;
    RECT 94.91 58.75 95.12 58.82 ;
    RECT 94.91 59.11 95.12 59.18 ;
    RECT 91.13 58.39 91.34 58.46 ;
    RECT 91.13 58.75 91.34 58.82 ;
    RECT 91.13 59.11 91.34 59.18 ;
    RECT 91.59 58.39 91.8 58.46 ;
    RECT 91.59 58.75 91.8 58.82 ;
    RECT 91.59 59.11 91.8 59.18 ;
    RECT 87.81 58.39 88.02 58.46 ;
    RECT 87.81 58.75 88.02 58.82 ;
    RECT 87.81 59.11 88.02 59.18 ;
    RECT 88.27 58.39 88.48 58.46 ;
    RECT 88.27 58.75 88.48 58.82 ;
    RECT 88.27 59.11 88.48 59.18 ;
    RECT 84.49 58.39 84.7 58.46 ;
    RECT 84.49 58.75 84.7 58.82 ;
    RECT 84.49 59.11 84.7 59.18 ;
    RECT 84.95 58.39 85.16 58.46 ;
    RECT 84.95 58.75 85.16 58.82 ;
    RECT 84.95 59.11 85.16 59.18 ;
    RECT 81.17 58.39 81.38 58.46 ;
    RECT 81.17 58.75 81.38 58.82 ;
    RECT 81.17 59.11 81.38 59.18 ;
    RECT 81.63 58.39 81.84 58.46 ;
    RECT 81.63 58.75 81.84 58.82 ;
    RECT 81.63 59.11 81.84 59.18 ;
    RECT 77.85 58.39 78.06 58.46 ;
    RECT 77.85 58.75 78.06 58.82 ;
    RECT 77.85 59.11 78.06 59.18 ;
    RECT 78.31 58.39 78.52 58.46 ;
    RECT 78.31 58.75 78.52 58.82 ;
    RECT 78.31 59.11 78.52 59.18 ;
    RECT 74.53 58.39 74.74 58.46 ;
    RECT 74.53 58.75 74.74 58.82 ;
    RECT 74.53 59.11 74.74 59.18 ;
    RECT 74.99 58.39 75.2 58.46 ;
    RECT 74.99 58.75 75.2 58.82 ;
    RECT 74.99 59.11 75.2 59.18 ;
    RECT 71.21 58.39 71.42 58.46 ;
    RECT 71.21 58.75 71.42 58.82 ;
    RECT 71.21 59.11 71.42 59.18 ;
    RECT 71.67 58.39 71.88 58.46 ;
    RECT 71.67 58.75 71.88 58.82 ;
    RECT 71.67 59.11 71.88 59.18 ;
    RECT 31.37 58.39 31.58 58.46 ;
    RECT 31.37 58.75 31.58 58.82 ;
    RECT 31.37 59.11 31.58 59.18 ;
    RECT 31.83 58.39 32.04 58.46 ;
    RECT 31.83 58.75 32.04 58.82 ;
    RECT 31.83 59.11 32.04 59.18 ;
    RECT 67.89 58.39 68.1 58.46 ;
    RECT 67.89 58.75 68.1 58.82 ;
    RECT 67.89 59.11 68.1 59.18 ;
    RECT 68.35 58.39 68.56 58.46 ;
    RECT 68.35 58.75 68.56 58.82 ;
    RECT 68.35 59.11 68.56 59.18 ;
    RECT 28.05 58.39 28.26 58.46 ;
    RECT 28.05 58.75 28.26 58.82 ;
    RECT 28.05 59.11 28.26 59.18 ;
    RECT 28.51 58.39 28.72 58.46 ;
    RECT 28.51 58.75 28.72 58.82 ;
    RECT 28.51 59.11 28.72 59.18 ;
    RECT 24.73 58.39 24.94 58.46 ;
    RECT 24.73 58.75 24.94 58.82 ;
    RECT 24.73 59.11 24.94 59.18 ;
    RECT 25.19 58.39 25.4 58.46 ;
    RECT 25.19 58.75 25.4 58.82 ;
    RECT 25.19 59.11 25.4 59.18 ;
    RECT 21.41 58.39 21.62 58.46 ;
    RECT 21.41 58.75 21.62 58.82 ;
    RECT 21.41 59.11 21.62 59.18 ;
    RECT 21.87 58.39 22.08 58.46 ;
    RECT 21.87 58.75 22.08 58.82 ;
    RECT 21.87 59.11 22.08 59.18 ;
    RECT 18.09 58.39 18.3 58.46 ;
    RECT 18.09 58.75 18.3 58.82 ;
    RECT 18.09 59.11 18.3 59.18 ;
    RECT 18.55 58.39 18.76 58.46 ;
    RECT 18.55 58.75 18.76 58.82 ;
    RECT 18.55 59.11 18.76 59.18 ;
    RECT 120.825 58.75 120.895 58.82 ;
    RECT 14.77 58.39 14.98 58.46 ;
    RECT 14.77 58.75 14.98 58.82 ;
    RECT 14.77 59.11 14.98 59.18 ;
    RECT 15.23 58.39 15.44 58.46 ;
    RECT 15.23 58.75 15.44 58.82 ;
    RECT 15.23 59.11 15.44 59.18 ;
    RECT 11.45 58.39 11.66 58.46 ;
    RECT 11.45 58.75 11.66 58.82 ;
    RECT 11.45 59.11 11.66 59.18 ;
    RECT 11.91 58.39 12.12 58.46 ;
    RECT 11.91 58.75 12.12 58.82 ;
    RECT 11.91 59.11 12.12 59.18 ;
    RECT 8.13 58.39 8.34 58.46 ;
    RECT 8.13 58.75 8.34 58.82 ;
    RECT 8.13 59.11 8.34 59.18 ;
    RECT 8.59 58.39 8.8 58.46 ;
    RECT 8.59 58.75 8.8 58.82 ;
    RECT 8.59 59.11 8.8 59.18 ;
    RECT 4.81 58.39 5.02 58.46 ;
    RECT 4.81 58.75 5.02 58.82 ;
    RECT 4.81 59.11 5.02 59.18 ;
    RECT 5.27 58.39 5.48 58.46 ;
    RECT 5.27 58.75 5.48 58.82 ;
    RECT 5.27 59.11 5.48 59.18 ;
    RECT 1.49 58.39 1.7 58.46 ;
    RECT 1.49 58.75 1.7 58.82 ;
    RECT 1.49 59.11 1.7 59.18 ;
    RECT 1.95 58.39 2.16 58.46 ;
    RECT 1.95 58.75 2.16 58.82 ;
    RECT 1.95 59.11 2.16 59.18 ;
    RECT 64.57 58.39 64.78 58.46 ;
    RECT 64.57 58.75 64.78 58.82 ;
    RECT 64.57 59.11 64.78 59.18 ;
    RECT 65.03 58.39 65.24 58.46 ;
    RECT 65.03 58.75 65.24 58.82 ;
    RECT 65.03 59.11 65.24 59.18 ;
    RECT 61.25 57.67 61.46 57.74 ;
    RECT 61.25 58.03 61.46 58.1 ;
    RECT 61.25 58.39 61.46 58.46 ;
    RECT 61.71 57.67 61.92 57.74 ;
    RECT 61.71 58.03 61.92 58.1 ;
    RECT 61.71 58.39 61.92 58.46 ;
    RECT 57.93 57.67 58.14 57.74 ;
    RECT 57.93 58.03 58.14 58.1 ;
    RECT 57.93 58.39 58.14 58.46 ;
    RECT 58.39 57.67 58.6 57.74 ;
    RECT 58.39 58.03 58.6 58.1 ;
    RECT 58.39 58.39 58.6 58.46 ;
    RECT 54.61 57.67 54.82 57.74 ;
    RECT 54.61 58.03 54.82 58.1 ;
    RECT 54.61 58.39 54.82 58.46 ;
    RECT 55.07 57.67 55.28 57.74 ;
    RECT 55.07 58.03 55.28 58.1 ;
    RECT 55.07 58.39 55.28 58.46 ;
    RECT 51.29 57.67 51.5 57.74 ;
    RECT 51.29 58.03 51.5 58.1 ;
    RECT 51.29 58.39 51.5 58.46 ;
    RECT 51.75 57.67 51.96 57.74 ;
    RECT 51.75 58.03 51.96 58.1 ;
    RECT 51.75 58.39 51.96 58.46 ;
    RECT 47.97 57.67 48.18 57.74 ;
    RECT 47.97 58.03 48.18 58.1 ;
    RECT 47.97 58.39 48.18 58.46 ;
    RECT 48.43 57.67 48.64 57.74 ;
    RECT 48.43 58.03 48.64 58.1 ;
    RECT 48.43 58.39 48.64 58.46 ;
    RECT 44.65 57.67 44.86 57.74 ;
    RECT 44.65 58.03 44.86 58.1 ;
    RECT 44.65 58.39 44.86 58.46 ;
    RECT 45.11 57.67 45.32 57.74 ;
    RECT 45.11 58.03 45.32 58.1 ;
    RECT 45.11 58.39 45.32 58.46 ;
    RECT 41.33 57.67 41.54 57.74 ;
    RECT 41.33 58.03 41.54 58.1 ;
    RECT 41.33 58.39 41.54 58.46 ;
    RECT 41.79 57.67 42.0 57.74 ;
    RECT 41.79 58.03 42.0 58.1 ;
    RECT 41.79 58.39 42.0 58.46 ;
    RECT 38.01 57.67 38.22 57.74 ;
    RECT 38.01 58.03 38.22 58.1 ;
    RECT 38.01 58.39 38.22 58.46 ;
    RECT 38.47 57.67 38.68 57.74 ;
    RECT 38.47 58.03 38.68 58.1 ;
    RECT 38.47 58.39 38.68 58.46 ;
    RECT 0.4 58.03 0.47 58.1 ;
    RECT 34.69 57.67 34.9 57.74 ;
    RECT 34.69 58.03 34.9 58.1 ;
    RECT 34.69 58.39 34.9 58.46 ;
    RECT 35.15 57.67 35.36 57.74 ;
    RECT 35.15 58.03 35.36 58.1 ;
    RECT 35.15 58.39 35.36 58.46 ;
    RECT 117.69 57.67 117.9 57.74 ;
    RECT 117.69 58.03 117.9 58.1 ;
    RECT 117.69 58.39 117.9 58.46 ;
    RECT 118.15 57.67 118.36 57.74 ;
    RECT 118.15 58.03 118.36 58.1 ;
    RECT 118.15 58.39 118.36 58.46 ;
    RECT 114.37 57.67 114.58 57.74 ;
    RECT 114.37 58.03 114.58 58.1 ;
    RECT 114.37 58.39 114.58 58.46 ;
    RECT 114.83 57.67 115.04 57.74 ;
    RECT 114.83 58.03 115.04 58.1 ;
    RECT 114.83 58.39 115.04 58.46 ;
    RECT 111.05 57.67 111.26 57.74 ;
    RECT 111.05 58.03 111.26 58.1 ;
    RECT 111.05 58.39 111.26 58.46 ;
    RECT 111.51 57.67 111.72 57.74 ;
    RECT 111.51 58.03 111.72 58.1 ;
    RECT 111.51 58.39 111.72 58.46 ;
    RECT 107.73 57.67 107.94 57.74 ;
    RECT 107.73 58.03 107.94 58.1 ;
    RECT 107.73 58.39 107.94 58.46 ;
    RECT 108.19 57.67 108.4 57.74 ;
    RECT 108.19 58.03 108.4 58.1 ;
    RECT 108.19 58.39 108.4 58.46 ;
    RECT 104.41 57.67 104.62 57.74 ;
    RECT 104.41 58.03 104.62 58.1 ;
    RECT 104.41 58.39 104.62 58.46 ;
    RECT 104.87 57.67 105.08 57.74 ;
    RECT 104.87 58.03 105.08 58.1 ;
    RECT 104.87 58.39 105.08 58.46 ;
    RECT 101.09 57.67 101.3 57.74 ;
    RECT 101.09 58.03 101.3 58.1 ;
    RECT 101.09 58.39 101.3 58.46 ;
    RECT 101.55 57.67 101.76 57.74 ;
    RECT 101.55 58.03 101.76 58.1 ;
    RECT 101.55 58.39 101.76 58.46 ;
    RECT 97.77 57.67 97.98 57.74 ;
    RECT 97.77 58.03 97.98 58.1 ;
    RECT 97.77 58.39 97.98 58.46 ;
    RECT 98.23 57.67 98.44 57.74 ;
    RECT 98.23 58.03 98.44 58.1 ;
    RECT 98.23 58.39 98.44 58.46 ;
    RECT 94.45 57.67 94.66 57.74 ;
    RECT 94.45 58.03 94.66 58.1 ;
    RECT 94.45 58.39 94.66 58.46 ;
    RECT 94.91 57.67 95.12 57.74 ;
    RECT 94.91 58.03 95.12 58.1 ;
    RECT 94.91 58.39 95.12 58.46 ;
    RECT 91.13 57.67 91.34 57.74 ;
    RECT 91.13 58.03 91.34 58.1 ;
    RECT 91.13 58.39 91.34 58.46 ;
    RECT 91.59 57.67 91.8 57.74 ;
    RECT 91.59 58.03 91.8 58.1 ;
    RECT 91.59 58.39 91.8 58.46 ;
    RECT 87.81 57.67 88.02 57.74 ;
    RECT 87.81 58.03 88.02 58.1 ;
    RECT 87.81 58.39 88.02 58.46 ;
    RECT 88.27 57.67 88.48 57.74 ;
    RECT 88.27 58.03 88.48 58.1 ;
    RECT 88.27 58.39 88.48 58.46 ;
    RECT 84.49 57.67 84.7 57.74 ;
    RECT 84.49 58.03 84.7 58.1 ;
    RECT 84.49 58.39 84.7 58.46 ;
    RECT 84.95 57.67 85.16 57.74 ;
    RECT 84.95 58.03 85.16 58.1 ;
    RECT 84.95 58.39 85.16 58.46 ;
    RECT 81.17 57.67 81.38 57.74 ;
    RECT 81.17 58.03 81.38 58.1 ;
    RECT 81.17 58.39 81.38 58.46 ;
    RECT 81.63 57.67 81.84 57.74 ;
    RECT 81.63 58.03 81.84 58.1 ;
    RECT 81.63 58.39 81.84 58.46 ;
    RECT 77.85 57.67 78.06 57.74 ;
    RECT 77.85 58.03 78.06 58.1 ;
    RECT 77.85 58.39 78.06 58.46 ;
    RECT 78.31 57.67 78.52 57.74 ;
    RECT 78.31 58.03 78.52 58.1 ;
    RECT 78.31 58.39 78.52 58.46 ;
    RECT 74.53 57.67 74.74 57.74 ;
    RECT 74.53 58.03 74.74 58.1 ;
    RECT 74.53 58.39 74.74 58.46 ;
    RECT 74.99 57.67 75.2 57.74 ;
    RECT 74.99 58.03 75.2 58.1 ;
    RECT 74.99 58.39 75.2 58.46 ;
    RECT 71.21 57.67 71.42 57.74 ;
    RECT 71.21 58.03 71.42 58.1 ;
    RECT 71.21 58.39 71.42 58.46 ;
    RECT 71.67 57.67 71.88 57.74 ;
    RECT 71.67 58.03 71.88 58.1 ;
    RECT 71.67 58.39 71.88 58.46 ;
    RECT 31.37 57.67 31.58 57.74 ;
    RECT 31.37 58.03 31.58 58.1 ;
    RECT 31.37 58.39 31.58 58.46 ;
    RECT 31.83 57.67 32.04 57.74 ;
    RECT 31.83 58.03 32.04 58.1 ;
    RECT 31.83 58.39 32.04 58.46 ;
    RECT 67.89 57.67 68.1 57.74 ;
    RECT 67.89 58.03 68.1 58.1 ;
    RECT 67.89 58.39 68.1 58.46 ;
    RECT 68.35 57.67 68.56 57.74 ;
    RECT 68.35 58.03 68.56 58.1 ;
    RECT 68.35 58.39 68.56 58.46 ;
    RECT 28.05 57.67 28.26 57.74 ;
    RECT 28.05 58.03 28.26 58.1 ;
    RECT 28.05 58.39 28.26 58.46 ;
    RECT 28.51 57.67 28.72 57.74 ;
    RECT 28.51 58.03 28.72 58.1 ;
    RECT 28.51 58.39 28.72 58.46 ;
    RECT 24.73 57.67 24.94 57.74 ;
    RECT 24.73 58.03 24.94 58.1 ;
    RECT 24.73 58.39 24.94 58.46 ;
    RECT 25.19 57.67 25.4 57.74 ;
    RECT 25.19 58.03 25.4 58.1 ;
    RECT 25.19 58.39 25.4 58.46 ;
    RECT 21.41 57.67 21.62 57.74 ;
    RECT 21.41 58.03 21.62 58.1 ;
    RECT 21.41 58.39 21.62 58.46 ;
    RECT 21.87 57.67 22.08 57.74 ;
    RECT 21.87 58.03 22.08 58.1 ;
    RECT 21.87 58.39 22.08 58.46 ;
    RECT 18.09 57.67 18.3 57.74 ;
    RECT 18.09 58.03 18.3 58.1 ;
    RECT 18.09 58.39 18.3 58.46 ;
    RECT 18.55 57.67 18.76 57.74 ;
    RECT 18.55 58.03 18.76 58.1 ;
    RECT 18.55 58.39 18.76 58.46 ;
    RECT 120.825 58.03 120.895 58.1 ;
    RECT 14.77 57.67 14.98 57.74 ;
    RECT 14.77 58.03 14.98 58.1 ;
    RECT 14.77 58.39 14.98 58.46 ;
    RECT 15.23 57.67 15.44 57.74 ;
    RECT 15.23 58.03 15.44 58.1 ;
    RECT 15.23 58.39 15.44 58.46 ;
    RECT 11.45 57.67 11.66 57.74 ;
    RECT 11.45 58.03 11.66 58.1 ;
    RECT 11.45 58.39 11.66 58.46 ;
    RECT 11.91 57.67 12.12 57.74 ;
    RECT 11.91 58.03 12.12 58.1 ;
    RECT 11.91 58.39 12.12 58.46 ;
    RECT 8.13 57.67 8.34 57.74 ;
    RECT 8.13 58.03 8.34 58.1 ;
    RECT 8.13 58.39 8.34 58.46 ;
    RECT 8.59 57.67 8.8 57.74 ;
    RECT 8.59 58.03 8.8 58.1 ;
    RECT 8.59 58.39 8.8 58.46 ;
    RECT 4.81 57.67 5.02 57.74 ;
    RECT 4.81 58.03 5.02 58.1 ;
    RECT 4.81 58.39 5.02 58.46 ;
    RECT 5.27 57.67 5.48 57.74 ;
    RECT 5.27 58.03 5.48 58.1 ;
    RECT 5.27 58.39 5.48 58.46 ;
    RECT 1.49 57.67 1.7 57.74 ;
    RECT 1.49 58.03 1.7 58.1 ;
    RECT 1.49 58.39 1.7 58.46 ;
    RECT 1.95 57.67 2.16 57.74 ;
    RECT 1.95 58.03 2.16 58.1 ;
    RECT 1.95 58.39 2.16 58.46 ;
    RECT 64.57 57.67 64.78 57.74 ;
    RECT 64.57 58.03 64.78 58.1 ;
    RECT 64.57 58.39 64.78 58.46 ;
    RECT 65.03 57.67 65.24 57.74 ;
    RECT 65.03 58.03 65.24 58.1 ;
    RECT 65.03 58.39 65.24 58.46 ;
    RECT 74.99 98.97 75.2 99.04 ;
    RECT 74.53 98.97 74.74 99.04 ;
    RECT 95.4 99.23 95.61 99.3 ;
    RECT 2.44 99.49 2.65 99.56 ;
    RECT 98.23 98.97 98.44 99.04 ;
    RECT 97.77 98.97 97.98 99.04 ;
    RECT 68.84 99.49 69.05 99.56 ;
    RECT 108.68 99.23 108.89 99.3 ;
    RECT 15.23 98.97 15.44 99.04 ;
    RECT 14.77 98.97 14.98 99.04 ;
    RECT 111.51 98.97 111.72 99.04 ;
    RECT 111.05 98.97 111.26 99.04 ;
    RECT 51.75 98.97 51.96 99.04 ;
    RECT 51.29 98.97 51.5 99.04 ;
    RECT 48.92 99.49 49.13 99.56 ;
    RECT 65.52 99.23 65.73 99.3 ;
    RECT 25.68 99.49 25.89 99.56 ;
    RECT 92.08 99.49 92.29 99.56 ;
    RECT 35.64 99.23 35.85 99.3 ;
    RECT 5.76 99.23 5.97 99.3 ;
    RECT 88.76 99.23 88.97 99.3 ;
    RECT 102.04 99.23 102.25 99.3 ;
    RECT 91.59 98.97 91.8 99.04 ;
    RECT 91.13 98.97 91.34 99.04 ;
    RECT 115.32 99.49 115.53 99.56 ;
    RECT 8.59 98.97 8.8 99.04 ;
    RECT 8.13 98.97 8.34 99.04 ;
    RECT 31.83 98.97 32.04 99.04 ;
    RECT 31.37 98.97 31.58 99.04 ;
    RECT 104.87 98.97 105.08 99.04 ;
    RECT 104.41 98.97 104.62 99.04 ;
    RECT 45.11 98.97 45.32 99.04 ;
    RECT 44.65 98.97 44.86 99.04 ;
    RECT 68.35 98.97 68.56 99.04 ;
    RECT 67.89 98.97 68.1 99.04 ;
    RECT 42.28 99.49 42.49 99.56 ;
    RECT 58.88 99.23 59.09 99.3 ;
    RECT 117.225 99.75 117.445 99.82 ;
    RECT 29.0 99.23 29.21 99.3 ;
    RECT 113.905 99.75 114.125 99.82 ;
    RECT 110.585 99.75 110.805 99.82 ;
    RECT 107.265 99.75 107.485 99.82 ;
    RECT 103.945 99.75 104.165 99.82 ;
    RECT 19.04 99.49 19.25 99.56 ;
    RECT 100.625 99.75 100.845 99.82 ;
    RECT 85.44 99.49 85.65 99.56 ;
    RECT 82.12 99.23 82.33 99.3 ;
    RECT 72.16 99.23 72.37 99.3 ;
    RECT 108.68 99.49 108.89 99.56 ;
    RECT 25.19 98.97 25.4 99.04 ;
    RECT 24.73 98.97 24.94 99.04 ;
    RECT 65.52 99.49 65.73 99.56 ;
    RECT 97.305 99.75 97.525 99.82 ;
    RECT 93.985 99.75 94.205 99.82 ;
    RECT 90.665 99.75 90.885 99.82 ;
    RECT 38.47 98.97 38.68 99.04 ;
    RECT 87.345 99.75 87.565 99.82 ;
    RECT 38.01 98.97 38.22 99.04 ;
    RECT 84.025 99.75 84.245 99.82 ;
    RECT 61.71 98.97 61.92 99.04 ;
    RECT 80.705 99.75 80.925 99.82 ;
    RECT 61.25 98.97 61.46 99.04 ;
    RECT 77.385 99.75 77.605 99.82 ;
    RECT 35.64 99.49 35.85 99.56 ;
    RECT 74.065 99.75 74.285 99.82 ;
    RECT 70.745 99.75 70.965 99.82 ;
    RECT 52.24 99.23 52.45 99.3 ;
    RECT 67.425 99.75 67.645 99.82 ;
    RECT 22.36 99.23 22.57 99.3 ;
    RECT 84.95 98.97 85.16 99.04 ;
    RECT 84.49 98.97 84.7 99.04 ;
    RECT 12.4 99.49 12.61 99.56 ;
    RECT 78.8 99.49 79.01 99.56 ;
    RECT 118.64 99.23 118.85 99.3 ;
    RECT 1.95 98.97 2.16 99.04 ;
    RECT 102.04 99.49 102.25 99.56 ;
    RECT 1.49 98.97 1.7 99.04 ;
    RECT 64.105 99.75 64.325 99.82 ;
    RECT 60.785 99.75 61.005 99.82 ;
    RECT 57.465 99.75 57.685 99.82 ;
    RECT 54.145 99.75 54.365 99.82 ;
    RECT 50.825 99.75 51.045 99.82 ;
    RECT 47.505 99.75 47.725 99.82 ;
    RECT 58.88 99.49 59.09 99.56 ;
    RECT 44.185 99.75 44.405 99.82 ;
    RECT 40.865 99.75 41.085 99.82 ;
    RECT 37.545 99.75 37.765 99.82 ;
    RECT 34.225 99.75 34.445 99.82 ;
    RECT 55.07 98.97 55.28 99.04 ;
    RECT 54.61 98.97 54.82 99.04 ;
    RECT 45.6 99.23 45.81 99.3 ;
    RECT 15.72 99.23 15.93 99.3 ;
    RECT 78.31 98.97 78.52 99.04 ;
    RECT 77.85 98.97 78.06 99.04 ;
    RECT 5.76 99.49 5.97 99.56 ;
    RECT 98.72 99.23 98.93 99.3 ;
    RECT 72.16 99.49 72.37 99.56 ;
    RECT 112.0 99.23 112.21 99.3 ;
    RECT 18.55 98.97 18.76 99.04 ;
    RECT 18.09 98.97 18.3 99.04 ;
    RECT 114.83 98.97 115.04 99.04 ;
    RECT 114.37 98.97 114.58 99.04 ;
    RECT 30.905 99.75 31.125 99.82 ;
    RECT 27.585 99.75 27.805 99.82 ;
    RECT 24.265 99.75 24.485 99.82 ;
    RECT 52.24 99.49 52.45 99.56 ;
    RECT 20.945 99.75 21.165 99.82 ;
    RECT 17.625 99.75 17.845 99.82 ;
    RECT 14.305 99.75 14.525 99.82 ;
    RECT 10.985 99.75 11.205 99.82 ;
    RECT 7.665 99.75 7.885 99.82 ;
    RECT 4.345 99.75 4.565 99.82 ;
    RECT 1.025 99.75 1.245 99.82 ;
    RECT 29.0 99.49 29.21 99.56 ;
    RECT 38.96 99.23 39.17 99.3 ;
    RECT 95.4 99.49 95.61 99.56 ;
    RECT 9.08 99.23 9.29 99.3 ;
    RECT 71.67 98.97 71.88 99.04 ;
    RECT 92.08 99.23 92.29 99.3 ;
    RECT 71.21 98.97 71.42 99.04 ;
    RECT 94.91 98.97 95.12 99.04 ;
    RECT 105.36 99.23 105.57 99.3 ;
    RECT 94.45 98.97 94.66 99.04 ;
    RECT 118.64 99.49 118.85 99.56 ;
    RECT 11.91 98.97 12.12 99.04 ;
    RECT 11.45 98.97 11.66 99.04 ;
    RECT 108.19 98.97 108.4 99.04 ;
    RECT 107.73 98.97 107.94 99.04 ;
    RECT 48.43 98.97 48.64 99.04 ;
    RECT 47.97 98.97 48.18 99.04 ;
    RECT 45.6 99.49 45.81 99.56 ;
    RECT 62.2 99.23 62.41 99.3 ;
    RECT 32.32 99.23 32.53 99.3 ;
    RECT 22.36 99.49 22.57 99.56 ;
    RECT 88.76 99.49 88.97 99.56 ;
    RECT 2.44 99.23 2.65 99.3 ;
    RECT 85.44 99.23 85.65 99.3 ;
    RECT 75.48 99.23 75.69 99.3 ;
    RECT 88.27 98.97 88.48 99.04 ;
    RECT 87.81 98.97 88.02 99.04 ;
    RECT 112.0 99.49 112.21 99.56 ;
    RECT 5.27 98.97 5.48 99.04 ;
    RECT 4.81 98.97 5.02 99.04 ;
    RECT 28.51 98.97 28.72 99.04 ;
    RECT 28.05 98.97 28.26 99.04 ;
    RECT 41.79 98.97 42.0 99.04 ;
    RECT 41.33 98.97 41.54 99.04 ;
    RECT 65.03 98.97 65.24 99.04 ;
    RECT 64.57 98.97 64.78 99.04 ;
    RECT 38.96 99.49 39.17 99.56 ;
    RECT 55.56 99.23 55.77 99.3 ;
    RECT 25.68 99.23 25.89 99.3 ;
    RECT 15.72 99.49 15.93 99.56 ;
    RECT 82.12 99.49 82.33 99.56 ;
    RECT 101.55 98.97 101.76 99.04 ;
    RECT 78.8 99.23 79.01 99.3 ;
    RECT 101.09 98.97 101.3 99.04 ;
    RECT 68.84 99.23 69.05 99.3 ;
    RECT 105.36 99.49 105.57 99.56 ;
    RECT 21.87 98.97 22.08 99.04 ;
    RECT 21.41 98.97 21.62 99.04 ;
    RECT 62.2 99.49 62.41 99.56 ;
    RECT 58.39 98.97 58.6 99.04 ;
    RECT 57.93 98.97 58.14 99.04 ;
    RECT 48.92 99.23 49.13 99.3 ;
    RECT 19.04 99.23 19.25 99.3 ;
    RECT 81.63 98.97 81.84 99.04 ;
    RECT 81.17 98.97 81.38 99.04 ;
    RECT 9.08 99.49 9.29 99.56 ;
    RECT 75.48 99.49 75.69 99.56 ;
    RECT 115.32 99.23 115.53 99.3 ;
    RECT 35.15 98.97 35.36 99.04 ;
    RECT 118.15 98.97 118.36 99.04 ;
    RECT 34.69 98.97 34.9 99.04 ;
    RECT 117.69 98.97 117.9 99.04 ;
    RECT 121.035 99.23 121.105 99.3 ;
    RECT 120.825 98.97 120.895 99.04 ;
    RECT 0.19 99.23 0.26 99.3 ;
    RECT 0.4 98.97 0.47 99.04 ;
    RECT 55.56 99.49 55.77 99.56 ;
    RECT 32.32 99.49 32.53 99.56 ;
    RECT 98.72 99.49 98.93 99.56 ;
    RECT 42.28 99.23 42.49 99.3 ;
    RECT 12.4 99.23 12.61 99.3 ;
    RECT 61.25 54.79 61.46 54.86 ;
    RECT 61.25 55.15 61.46 55.22 ;
    RECT 61.25 55.51 61.46 55.58 ;
    RECT 61.71 54.79 61.92 54.86 ;
    RECT 61.71 55.15 61.92 55.22 ;
    RECT 61.71 55.51 61.92 55.58 ;
    RECT 57.93 54.79 58.14 54.86 ;
    RECT 57.93 55.15 58.14 55.22 ;
    RECT 57.93 55.51 58.14 55.58 ;
    RECT 58.39 54.79 58.6 54.86 ;
    RECT 58.39 55.15 58.6 55.22 ;
    RECT 58.39 55.51 58.6 55.58 ;
    RECT 54.61 54.79 54.82 54.86 ;
    RECT 54.61 55.15 54.82 55.22 ;
    RECT 54.61 55.51 54.82 55.58 ;
    RECT 55.07 54.79 55.28 54.86 ;
    RECT 55.07 55.15 55.28 55.22 ;
    RECT 55.07 55.51 55.28 55.58 ;
    RECT 51.29 54.79 51.5 54.86 ;
    RECT 51.29 55.15 51.5 55.22 ;
    RECT 51.29 55.51 51.5 55.58 ;
    RECT 51.75 54.79 51.96 54.86 ;
    RECT 51.75 55.15 51.96 55.22 ;
    RECT 51.75 55.51 51.96 55.58 ;
    RECT 47.97 54.79 48.18 54.86 ;
    RECT 47.97 55.15 48.18 55.22 ;
    RECT 47.97 55.51 48.18 55.58 ;
    RECT 48.43 54.79 48.64 54.86 ;
    RECT 48.43 55.15 48.64 55.22 ;
    RECT 48.43 55.51 48.64 55.58 ;
    RECT 0.4 55.15 0.47 55.22 ;
    RECT 44.65 54.79 44.86 54.86 ;
    RECT 44.65 55.15 44.86 55.22 ;
    RECT 44.65 55.51 44.86 55.58 ;
    RECT 45.11 54.79 45.32 54.86 ;
    RECT 45.11 55.15 45.32 55.22 ;
    RECT 45.11 55.51 45.32 55.58 ;
    RECT 41.33 54.79 41.54 54.86 ;
    RECT 41.33 55.15 41.54 55.22 ;
    RECT 41.33 55.51 41.54 55.58 ;
    RECT 41.79 54.79 42.0 54.86 ;
    RECT 41.79 55.15 42.0 55.22 ;
    RECT 41.79 55.51 42.0 55.58 ;
    RECT 38.01 54.79 38.22 54.86 ;
    RECT 38.01 55.15 38.22 55.22 ;
    RECT 38.01 55.51 38.22 55.58 ;
    RECT 38.47 54.79 38.68 54.86 ;
    RECT 38.47 55.15 38.68 55.22 ;
    RECT 38.47 55.51 38.68 55.58 ;
    RECT 34.69 54.79 34.9 54.86 ;
    RECT 34.69 55.15 34.9 55.22 ;
    RECT 34.69 55.51 34.9 55.58 ;
    RECT 35.15 54.79 35.36 54.86 ;
    RECT 35.15 55.15 35.36 55.22 ;
    RECT 35.15 55.51 35.36 55.58 ;
    RECT 117.69 54.79 117.9 54.86 ;
    RECT 117.69 55.15 117.9 55.22 ;
    RECT 117.69 55.51 117.9 55.58 ;
    RECT 118.15 54.79 118.36 54.86 ;
    RECT 118.15 55.15 118.36 55.22 ;
    RECT 118.15 55.51 118.36 55.58 ;
    RECT 114.37 54.79 114.58 54.86 ;
    RECT 114.37 55.15 114.58 55.22 ;
    RECT 114.37 55.51 114.58 55.58 ;
    RECT 114.83 54.79 115.04 54.86 ;
    RECT 114.83 55.15 115.04 55.22 ;
    RECT 114.83 55.51 115.04 55.58 ;
    RECT 111.05 54.79 111.26 54.86 ;
    RECT 111.05 55.15 111.26 55.22 ;
    RECT 111.05 55.51 111.26 55.58 ;
    RECT 111.51 54.79 111.72 54.86 ;
    RECT 111.51 55.15 111.72 55.22 ;
    RECT 111.51 55.51 111.72 55.58 ;
    RECT 107.73 54.79 107.94 54.86 ;
    RECT 107.73 55.15 107.94 55.22 ;
    RECT 107.73 55.51 107.94 55.58 ;
    RECT 108.19 54.79 108.4 54.86 ;
    RECT 108.19 55.15 108.4 55.22 ;
    RECT 108.19 55.51 108.4 55.58 ;
    RECT 104.41 54.79 104.62 54.86 ;
    RECT 104.41 55.15 104.62 55.22 ;
    RECT 104.41 55.51 104.62 55.58 ;
    RECT 104.87 54.79 105.08 54.86 ;
    RECT 104.87 55.15 105.08 55.22 ;
    RECT 104.87 55.51 105.08 55.58 ;
    RECT 101.09 54.79 101.3 54.86 ;
    RECT 101.09 55.15 101.3 55.22 ;
    RECT 101.09 55.51 101.3 55.58 ;
    RECT 101.55 54.79 101.76 54.86 ;
    RECT 101.55 55.15 101.76 55.22 ;
    RECT 101.55 55.51 101.76 55.58 ;
    RECT 120.825 55.15 120.895 55.22 ;
    RECT 97.77 54.79 97.98 54.86 ;
    RECT 97.77 55.15 97.98 55.22 ;
    RECT 97.77 55.51 97.98 55.58 ;
    RECT 98.23 54.79 98.44 54.86 ;
    RECT 98.23 55.15 98.44 55.22 ;
    RECT 98.23 55.51 98.44 55.58 ;
    RECT 94.45 54.79 94.66 54.86 ;
    RECT 94.45 55.15 94.66 55.22 ;
    RECT 94.45 55.51 94.66 55.58 ;
    RECT 94.91 54.79 95.12 54.86 ;
    RECT 94.91 55.15 95.12 55.22 ;
    RECT 94.91 55.51 95.12 55.58 ;
    RECT 91.13 54.79 91.34 54.86 ;
    RECT 91.13 55.15 91.34 55.22 ;
    RECT 91.13 55.51 91.34 55.58 ;
    RECT 91.59 54.79 91.8 54.86 ;
    RECT 91.59 55.15 91.8 55.22 ;
    RECT 91.59 55.51 91.8 55.58 ;
    RECT 87.81 54.79 88.02 54.86 ;
    RECT 87.81 55.15 88.02 55.22 ;
    RECT 87.81 55.51 88.02 55.58 ;
    RECT 88.27 54.79 88.48 54.86 ;
    RECT 88.27 55.15 88.48 55.22 ;
    RECT 88.27 55.51 88.48 55.58 ;
    RECT 84.49 54.79 84.7 54.86 ;
    RECT 84.49 55.15 84.7 55.22 ;
    RECT 84.49 55.51 84.7 55.58 ;
    RECT 84.95 54.79 85.16 54.86 ;
    RECT 84.95 55.15 85.16 55.22 ;
    RECT 84.95 55.51 85.16 55.58 ;
    RECT 81.17 54.79 81.38 54.86 ;
    RECT 81.17 55.15 81.38 55.22 ;
    RECT 81.17 55.51 81.38 55.58 ;
    RECT 81.63 54.79 81.84 54.86 ;
    RECT 81.63 55.15 81.84 55.22 ;
    RECT 81.63 55.51 81.84 55.58 ;
    RECT 77.85 54.79 78.06 54.86 ;
    RECT 77.85 55.15 78.06 55.22 ;
    RECT 77.85 55.51 78.06 55.58 ;
    RECT 78.31 54.79 78.52 54.86 ;
    RECT 78.31 55.15 78.52 55.22 ;
    RECT 78.31 55.51 78.52 55.58 ;
    RECT 74.53 54.79 74.74 54.86 ;
    RECT 74.53 55.15 74.74 55.22 ;
    RECT 74.53 55.51 74.74 55.58 ;
    RECT 74.99 54.79 75.2 54.86 ;
    RECT 74.99 55.15 75.2 55.22 ;
    RECT 74.99 55.51 75.2 55.58 ;
    RECT 71.21 54.79 71.42 54.86 ;
    RECT 71.21 55.15 71.42 55.22 ;
    RECT 71.21 55.51 71.42 55.58 ;
    RECT 71.67 54.79 71.88 54.86 ;
    RECT 71.67 55.15 71.88 55.22 ;
    RECT 71.67 55.51 71.88 55.58 ;
    RECT 31.37 54.79 31.58 54.86 ;
    RECT 31.37 55.15 31.58 55.22 ;
    RECT 31.37 55.51 31.58 55.58 ;
    RECT 31.83 54.79 32.04 54.86 ;
    RECT 31.83 55.15 32.04 55.22 ;
    RECT 31.83 55.51 32.04 55.58 ;
    RECT 67.89 54.79 68.1 54.86 ;
    RECT 67.89 55.15 68.1 55.22 ;
    RECT 67.89 55.51 68.1 55.58 ;
    RECT 68.35 54.79 68.56 54.86 ;
    RECT 68.35 55.15 68.56 55.22 ;
    RECT 68.35 55.51 68.56 55.58 ;
    RECT 28.05 54.79 28.26 54.86 ;
    RECT 28.05 55.15 28.26 55.22 ;
    RECT 28.05 55.51 28.26 55.58 ;
    RECT 28.51 54.79 28.72 54.86 ;
    RECT 28.51 55.15 28.72 55.22 ;
    RECT 28.51 55.51 28.72 55.58 ;
    RECT 24.73 54.79 24.94 54.86 ;
    RECT 24.73 55.15 24.94 55.22 ;
    RECT 24.73 55.51 24.94 55.58 ;
    RECT 25.19 54.79 25.4 54.86 ;
    RECT 25.19 55.15 25.4 55.22 ;
    RECT 25.19 55.51 25.4 55.58 ;
    RECT 21.41 54.79 21.62 54.86 ;
    RECT 21.41 55.15 21.62 55.22 ;
    RECT 21.41 55.51 21.62 55.58 ;
    RECT 21.87 54.79 22.08 54.86 ;
    RECT 21.87 55.15 22.08 55.22 ;
    RECT 21.87 55.51 22.08 55.58 ;
    RECT 18.09 54.79 18.3 54.86 ;
    RECT 18.09 55.15 18.3 55.22 ;
    RECT 18.09 55.51 18.3 55.58 ;
    RECT 18.55 54.79 18.76 54.86 ;
    RECT 18.55 55.15 18.76 55.22 ;
    RECT 18.55 55.51 18.76 55.58 ;
    RECT 14.77 54.79 14.98 54.86 ;
    RECT 14.77 55.15 14.98 55.22 ;
    RECT 14.77 55.51 14.98 55.58 ;
    RECT 15.23 54.79 15.44 54.86 ;
    RECT 15.23 55.15 15.44 55.22 ;
    RECT 15.23 55.51 15.44 55.58 ;
    RECT 11.45 54.79 11.66 54.86 ;
    RECT 11.45 55.15 11.66 55.22 ;
    RECT 11.45 55.51 11.66 55.58 ;
    RECT 11.91 54.79 12.12 54.86 ;
    RECT 11.91 55.15 12.12 55.22 ;
    RECT 11.91 55.51 12.12 55.58 ;
    RECT 8.13 54.79 8.34 54.86 ;
    RECT 8.13 55.15 8.34 55.22 ;
    RECT 8.13 55.51 8.34 55.58 ;
    RECT 8.59 54.79 8.8 54.86 ;
    RECT 8.59 55.15 8.8 55.22 ;
    RECT 8.59 55.51 8.8 55.58 ;
    RECT 4.81 54.79 5.02 54.86 ;
    RECT 4.81 55.15 5.02 55.22 ;
    RECT 4.81 55.51 5.02 55.58 ;
    RECT 5.27 54.79 5.48 54.86 ;
    RECT 5.27 55.15 5.48 55.22 ;
    RECT 5.27 55.51 5.48 55.58 ;
    RECT 1.49 54.79 1.7 54.86 ;
    RECT 1.49 55.15 1.7 55.22 ;
    RECT 1.49 55.51 1.7 55.58 ;
    RECT 1.95 54.79 2.16 54.86 ;
    RECT 1.95 55.15 2.16 55.22 ;
    RECT 1.95 55.51 2.16 55.58 ;
    RECT 64.57 54.79 64.78 54.86 ;
    RECT 64.57 55.15 64.78 55.22 ;
    RECT 64.57 55.51 64.78 55.58 ;
    RECT 65.03 54.79 65.24 54.86 ;
    RECT 65.03 55.15 65.24 55.22 ;
    RECT 65.03 55.51 65.24 55.58 ;
    RECT 61.25 55.51 61.46 55.58 ;
    RECT 61.25 55.87 61.46 55.94 ;
    RECT 61.25 56.23 61.46 56.3 ;
    RECT 61.71 55.51 61.92 55.58 ;
    RECT 61.71 55.87 61.92 55.94 ;
    RECT 61.71 56.23 61.92 56.3 ;
    RECT 57.93 55.51 58.14 55.58 ;
    RECT 57.93 55.87 58.14 55.94 ;
    RECT 57.93 56.23 58.14 56.3 ;
    RECT 58.39 55.51 58.6 55.58 ;
    RECT 58.39 55.87 58.6 55.94 ;
    RECT 58.39 56.23 58.6 56.3 ;
    RECT 54.61 55.51 54.82 55.58 ;
    RECT 54.61 55.87 54.82 55.94 ;
    RECT 54.61 56.23 54.82 56.3 ;
    RECT 55.07 55.51 55.28 55.58 ;
    RECT 55.07 55.87 55.28 55.94 ;
    RECT 55.07 56.23 55.28 56.3 ;
    RECT 51.29 55.51 51.5 55.58 ;
    RECT 51.29 55.87 51.5 55.94 ;
    RECT 51.29 56.23 51.5 56.3 ;
    RECT 51.75 55.51 51.96 55.58 ;
    RECT 51.75 55.87 51.96 55.94 ;
    RECT 51.75 56.23 51.96 56.3 ;
    RECT 47.97 55.51 48.18 55.58 ;
    RECT 47.97 55.87 48.18 55.94 ;
    RECT 47.97 56.23 48.18 56.3 ;
    RECT 48.43 55.51 48.64 55.58 ;
    RECT 48.43 55.87 48.64 55.94 ;
    RECT 48.43 56.23 48.64 56.3 ;
    RECT 44.65 55.51 44.86 55.58 ;
    RECT 44.65 55.87 44.86 55.94 ;
    RECT 44.65 56.23 44.86 56.3 ;
    RECT 45.11 55.51 45.32 55.58 ;
    RECT 45.11 55.87 45.32 55.94 ;
    RECT 45.11 56.23 45.32 56.3 ;
    RECT 41.33 55.51 41.54 55.58 ;
    RECT 41.33 55.87 41.54 55.94 ;
    RECT 41.33 56.23 41.54 56.3 ;
    RECT 41.79 55.51 42.0 55.58 ;
    RECT 41.79 55.87 42.0 55.94 ;
    RECT 41.79 56.23 42.0 56.3 ;
    RECT 38.01 55.51 38.22 55.58 ;
    RECT 38.01 55.87 38.22 55.94 ;
    RECT 38.01 56.23 38.22 56.3 ;
    RECT 38.47 55.51 38.68 55.58 ;
    RECT 38.47 55.87 38.68 55.94 ;
    RECT 38.47 56.23 38.68 56.3 ;
    RECT 34.69 55.51 34.9 55.58 ;
    RECT 34.69 55.87 34.9 55.94 ;
    RECT 34.69 56.23 34.9 56.3 ;
    RECT 35.15 55.51 35.36 55.58 ;
    RECT 35.15 55.87 35.36 55.94 ;
    RECT 35.15 56.23 35.36 56.3 ;
    RECT 117.69 55.51 117.9 55.58 ;
    RECT 117.69 55.87 117.9 55.94 ;
    RECT 117.69 56.23 117.9 56.3 ;
    RECT 118.15 55.51 118.36 55.58 ;
    RECT 118.15 55.87 118.36 55.94 ;
    RECT 118.15 56.23 118.36 56.3 ;
    RECT 114.37 55.51 114.58 55.58 ;
    RECT 114.37 55.87 114.58 55.94 ;
    RECT 114.37 56.23 114.58 56.3 ;
    RECT 114.83 55.51 115.04 55.58 ;
    RECT 114.83 55.87 115.04 55.94 ;
    RECT 114.83 56.23 115.04 56.3 ;
    RECT 111.05 55.51 111.26 55.58 ;
    RECT 111.05 55.87 111.26 55.94 ;
    RECT 111.05 56.23 111.26 56.3 ;
    RECT 111.51 55.51 111.72 55.58 ;
    RECT 111.51 55.87 111.72 55.94 ;
    RECT 111.51 56.23 111.72 56.3 ;
    RECT 107.73 55.51 107.94 55.58 ;
    RECT 107.73 55.87 107.94 55.94 ;
    RECT 107.73 56.23 107.94 56.3 ;
    RECT 108.19 55.51 108.4 55.58 ;
    RECT 108.19 55.87 108.4 55.94 ;
    RECT 108.19 56.23 108.4 56.3 ;
    RECT 104.41 55.51 104.62 55.58 ;
    RECT 104.41 55.87 104.62 55.94 ;
    RECT 104.41 56.23 104.62 56.3 ;
    RECT 104.87 55.51 105.08 55.58 ;
    RECT 104.87 55.87 105.08 55.94 ;
    RECT 104.87 56.23 105.08 56.3 ;
    RECT 101.09 55.51 101.3 55.58 ;
    RECT 101.09 55.87 101.3 55.94 ;
    RECT 101.09 56.23 101.3 56.3 ;
    RECT 101.55 55.51 101.76 55.58 ;
    RECT 101.55 55.87 101.76 55.94 ;
    RECT 101.55 56.23 101.76 56.3 ;
    RECT 120.825 55.87 120.895 55.94 ;
    RECT 97.77 55.51 97.98 55.58 ;
    RECT 97.77 55.87 97.98 55.94 ;
    RECT 97.77 56.23 97.98 56.3 ;
    RECT 98.23 55.51 98.44 55.58 ;
    RECT 98.23 55.87 98.44 55.94 ;
    RECT 98.23 56.23 98.44 56.3 ;
    RECT 94.45 55.51 94.66 55.58 ;
    RECT 94.45 55.87 94.66 55.94 ;
    RECT 94.45 56.23 94.66 56.3 ;
    RECT 94.91 55.51 95.12 55.58 ;
    RECT 94.91 55.87 95.12 55.94 ;
    RECT 94.91 56.23 95.12 56.3 ;
    RECT 91.13 55.51 91.34 55.58 ;
    RECT 91.13 55.87 91.34 55.94 ;
    RECT 91.13 56.23 91.34 56.3 ;
    RECT 91.59 55.51 91.8 55.58 ;
    RECT 91.59 55.87 91.8 55.94 ;
    RECT 91.59 56.23 91.8 56.3 ;
    RECT 87.81 55.51 88.02 55.58 ;
    RECT 87.81 55.87 88.02 55.94 ;
    RECT 87.81 56.23 88.02 56.3 ;
    RECT 88.27 55.51 88.48 55.58 ;
    RECT 88.27 55.87 88.48 55.94 ;
    RECT 88.27 56.23 88.48 56.3 ;
    RECT 84.49 55.51 84.7 55.58 ;
    RECT 84.49 55.87 84.7 55.94 ;
    RECT 84.49 56.23 84.7 56.3 ;
    RECT 84.95 55.51 85.16 55.58 ;
    RECT 84.95 55.87 85.16 55.94 ;
    RECT 84.95 56.23 85.16 56.3 ;
    RECT 81.17 55.51 81.38 55.58 ;
    RECT 81.17 55.87 81.38 55.94 ;
    RECT 81.17 56.23 81.38 56.3 ;
    RECT 81.63 55.51 81.84 55.58 ;
    RECT 81.63 55.87 81.84 55.94 ;
    RECT 81.63 56.23 81.84 56.3 ;
    RECT 77.85 55.51 78.06 55.58 ;
    RECT 77.85 55.87 78.06 55.94 ;
    RECT 77.85 56.23 78.06 56.3 ;
    RECT 78.31 55.51 78.52 55.58 ;
    RECT 78.31 55.87 78.52 55.94 ;
    RECT 78.31 56.23 78.52 56.3 ;
    RECT 74.53 55.51 74.74 55.58 ;
    RECT 74.53 55.87 74.74 55.94 ;
    RECT 74.53 56.23 74.74 56.3 ;
    RECT 74.99 55.51 75.2 55.58 ;
    RECT 74.99 55.87 75.2 55.94 ;
    RECT 74.99 56.23 75.2 56.3 ;
    RECT 71.21 55.51 71.42 55.58 ;
    RECT 71.21 55.87 71.42 55.94 ;
    RECT 71.21 56.23 71.42 56.3 ;
    RECT 71.67 55.51 71.88 55.58 ;
    RECT 71.67 55.87 71.88 55.94 ;
    RECT 71.67 56.23 71.88 56.3 ;
    RECT 31.37 55.51 31.58 55.58 ;
    RECT 31.37 55.87 31.58 55.94 ;
    RECT 31.37 56.23 31.58 56.3 ;
    RECT 31.83 55.51 32.04 55.58 ;
    RECT 31.83 55.87 32.04 55.94 ;
    RECT 31.83 56.23 32.04 56.3 ;
    RECT 67.89 55.51 68.1 55.58 ;
    RECT 67.89 55.87 68.1 55.94 ;
    RECT 67.89 56.23 68.1 56.3 ;
    RECT 68.35 55.51 68.56 55.58 ;
    RECT 68.35 55.87 68.56 55.94 ;
    RECT 68.35 56.23 68.56 56.3 ;
    RECT 28.05 55.51 28.26 55.58 ;
    RECT 28.05 55.87 28.26 55.94 ;
    RECT 28.05 56.23 28.26 56.3 ;
    RECT 28.51 55.51 28.72 55.58 ;
    RECT 28.51 55.87 28.72 55.94 ;
    RECT 28.51 56.23 28.72 56.3 ;
    RECT 24.73 55.51 24.94 55.58 ;
    RECT 24.73 55.87 24.94 55.94 ;
    RECT 24.73 56.23 24.94 56.3 ;
    RECT 25.19 55.51 25.4 55.58 ;
    RECT 25.19 55.87 25.4 55.94 ;
    RECT 25.19 56.23 25.4 56.3 ;
    RECT 21.41 55.51 21.62 55.58 ;
    RECT 21.41 55.87 21.62 55.94 ;
    RECT 21.41 56.23 21.62 56.3 ;
    RECT 21.87 55.51 22.08 55.58 ;
    RECT 21.87 55.87 22.08 55.94 ;
    RECT 21.87 56.23 22.08 56.3 ;
    RECT 0.4 55.87 0.47 55.94 ;
    RECT 18.09 55.51 18.3 55.58 ;
    RECT 18.09 55.87 18.3 55.94 ;
    RECT 18.09 56.23 18.3 56.3 ;
    RECT 18.55 55.51 18.76 55.58 ;
    RECT 18.55 55.87 18.76 55.94 ;
    RECT 18.55 56.23 18.76 56.3 ;
    RECT 14.77 55.51 14.98 55.58 ;
    RECT 14.77 55.87 14.98 55.94 ;
    RECT 14.77 56.23 14.98 56.3 ;
    RECT 15.23 55.51 15.44 55.58 ;
    RECT 15.23 55.87 15.44 55.94 ;
    RECT 15.23 56.23 15.44 56.3 ;
    RECT 11.45 55.51 11.66 55.58 ;
    RECT 11.45 55.87 11.66 55.94 ;
    RECT 11.45 56.23 11.66 56.3 ;
    RECT 11.91 55.51 12.12 55.58 ;
    RECT 11.91 55.87 12.12 55.94 ;
    RECT 11.91 56.23 12.12 56.3 ;
    RECT 8.13 55.51 8.34 55.58 ;
    RECT 8.13 55.87 8.34 55.94 ;
    RECT 8.13 56.23 8.34 56.3 ;
    RECT 8.59 55.51 8.8 55.58 ;
    RECT 8.59 55.87 8.8 55.94 ;
    RECT 8.59 56.23 8.8 56.3 ;
    RECT 4.81 55.51 5.02 55.58 ;
    RECT 4.81 55.87 5.02 55.94 ;
    RECT 4.81 56.23 5.02 56.3 ;
    RECT 5.27 55.51 5.48 55.58 ;
    RECT 5.27 55.87 5.48 55.94 ;
    RECT 5.27 56.23 5.48 56.3 ;
    RECT 1.49 55.51 1.7 55.58 ;
    RECT 1.49 55.87 1.7 55.94 ;
    RECT 1.49 56.23 1.7 56.3 ;
    RECT 1.95 55.51 2.16 55.58 ;
    RECT 1.95 55.87 2.16 55.94 ;
    RECT 1.95 56.23 2.16 56.3 ;
    RECT 64.57 55.51 64.78 55.58 ;
    RECT 64.57 55.87 64.78 55.94 ;
    RECT 64.57 56.23 64.78 56.3 ;
    RECT 65.03 55.51 65.24 55.58 ;
    RECT 65.03 55.87 65.24 55.94 ;
    RECT 65.03 56.23 65.24 56.3 ;
    RECT 61.25 97.29 61.46 97.36 ;
    RECT 61.25 97.65 61.46 97.72 ;
    RECT 61.25 98.01 61.46 98.08 ;
    RECT 61.71 97.29 61.92 97.36 ;
    RECT 61.71 97.65 61.92 97.72 ;
    RECT 61.71 98.01 61.92 98.08 ;
    RECT 57.93 97.29 58.14 97.36 ;
    RECT 57.93 97.65 58.14 97.72 ;
    RECT 57.93 98.01 58.14 98.08 ;
    RECT 58.39 97.29 58.6 97.36 ;
    RECT 58.39 97.65 58.6 97.72 ;
    RECT 58.39 98.01 58.6 98.08 ;
    RECT 54.61 97.29 54.82 97.36 ;
    RECT 54.61 97.65 54.82 97.72 ;
    RECT 54.61 98.01 54.82 98.08 ;
    RECT 55.07 97.29 55.28 97.36 ;
    RECT 55.07 97.65 55.28 97.72 ;
    RECT 55.07 98.01 55.28 98.08 ;
    RECT 51.29 97.29 51.5 97.36 ;
    RECT 51.29 97.65 51.5 97.72 ;
    RECT 51.29 98.01 51.5 98.08 ;
    RECT 51.75 97.29 51.96 97.36 ;
    RECT 51.75 97.65 51.96 97.72 ;
    RECT 51.75 98.01 51.96 98.08 ;
    RECT 47.97 97.29 48.18 97.36 ;
    RECT 47.97 97.65 48.18 97.72 ;
    RECT 47.97 98.01 48.18 98.08 ;
    RECT 48.43 97.29 48.64 97.36 ;
    RECT 48.43 97.65 48.64 97.72 ;
    RECT 48.43 98.01 48.64 98.08 ;
    RECT 44.65 97.29 44.86 97.36 ;
    RECT 44.65 97.65 44.86 97.72 ;
    RECT 44.65 98.01 44.86 98.08 ;
    RECT 45.11 97.29 45.32 97.36 ;
    RECT 45.11 97.65 45.32 97.72 ;
    RECT 45.11 98.01 45.32 98.08 ;
    RECT 41.33 97.29 41.54 97.36 ;
    RECT 41.33 97.65 41.54 97.72 ;
    RECT 41.33 98.01 41.54 98.08 ;
    RECT 41.79 97.29 42.0 97.36 ;
    RECT 41.79 97.65 42.0 97.72 ;
    RECT 41.79 98.01 42.0 98.08 ;
    RECT 38.01 97.29 38.22 97.36 ;
    RECT 38.01 97.65 38.22 97.72 ;
    RECT 38.01 98.01 38.22 98.08 ;
    RECT 38.47 97.29 38.68 97.36 ;
    RECT 38.47 97.65 38.68 97.72 ;
    RECT 38.47 98.01 38.68 98.08 ;
    RECT 0.4 97.65 0.47 97.72 ;
    RECT 34.69 97.29 34.9 97.36 ;
    RECT 34.69 97.65 34.9 97.72 ;
    RECT 34.69 98.01 34.9 98.08 ;
    RECT 35.15 97.29 35.36 97.36 ;
    RECT 35.15 97.65 35.36 97.72 ;
    RECT 35.15 98.01 35.36 98.08 ;
    RECT 117.69 97.29 117.9 97.36 ;
    RECT 117.69 97.65 117.9 97.72 ;
    RECT 117.69 98.01 117.9 98.08 ;
    RECT 118.15 97.29 118.36 97.36 ;
    RECT 118.15 97.65 118.36 97.72 ;
    RECT 118.15 98.01 118.36 98.08 ;
    RECT 114.37 97.29 114.58 97.36 ;
    RECT 114.37 97.65 114.58 97.72 ;
    RECT 114.37 98.01 114.58 98.08 ;
    RECT 114.83 97.29 115.04 97.36 ;
    RECT 114.83 97.65 115.04 97.72 ;
    RECT 114.83 98.01 115.04 98.08 ;
    RECT 111.05 97.29 111.26 97.36 ;
    RECT 111.05 97.65 111.26 97.72 ;
    RECT 111.05 98.01 111.26 98.08 ;
    RECT 111.51 97.29 111.72 97.36 ;
    RECT 111.51 97.65 111.72 97.72 ;
    RECT 111.51 98.01 111.72 98.08 ;
    RECT 107.73 97.29 107.94 97.36 ;
    RECT 107.73 97.65 107.94 97.72 ;
    RECT 107.73 98.01 107.94 98.08 ;
    RECT 108.19 97.29 108.4 97.36 ;
    RECT 108.19 97.65 108.4 97.72 ;
    RECT 108.19 98.01 108.4 98.08 ;
    RECT 104.41 97.29 104.62 97.36 ;
    RECT 104.41 97.65 104.62 97.72 ;
    RECT 104.41 98.01 104.62 98.08 ;
    RECT 104.87 97.29 105.08 97.36 ;
    RECT 104.87 97.65 105.08 97.72 ;
    RECT 104.87 98.01 105.08 98.08 ;
    RECT 101.09 97.29 101.3 97.36 ;
    RECT 101.09 97.65 101.3 97.72 ;
    RECT 101.09 98.01 101.3 98.08 ;
    RECT 101.55 97.29 101.76 97.36 ;
    RECT 101.55 97.65 101.76 97.72 ;
    RECT 101.55 98.01 101.76 98.08 ;
    RECT 97.77 97.29 97.98 97.36 ;
    RECT 97.77 97.65 97.98 97.72 ;
    RECT 97.77 98.01 97.98 98.08 ;
    RECT 98.23 97.29 98.44 97.36 ;
    RECT 98.23 97.65 98.44 97.72 ;
    RECT 98.23 98.01 98.44 98.08 ;
    RECT 94.45 97.29 94.66 97.36 ;
    RECT 94.45 97.65 94.66 97.72 ;
    RECT 94.45 98.01 94.66 98.08 ;
    RECT 94.91 97.29 95.12 97.36 ;
    RECT 94.91 97.65 95.12 97.72 ;
    RECT 94.91 98.01 95.12 98.08 ;
    RECT 91.13 97.29 91.34 97.36 ;
    RECT 91.13 97.65 91.34 97.72 ;
    RECT 91.13 98.01 91.34 98.08 ;
    RECT 91.59 97.29 91.8 97.36 ;
    RECT 91.59 97.65 91.8 97.72 ;
    RECT 91.59 98.01 91.8 98.08 ;
    RECT 87.81 97.29 88.02 97.36 ;
    RECT 87.81 97.65 88.02 97.72 ;
    RECT 87.81 98.01 88.02 98.08 ;
    RECT 88.27 97.29 88.48 97.36 ;
    RECT 88.27 97.65 88.48 97.72 ;
    RECT 88.27 98.01 88.48 98.08 ;
    RECT 84.49 97.29 84.7 97.36 ;
    RECT 84.49 97.65 84.7 97.72 ;
    RECT 84.49 98.01 84.7 98.08 ;
    RECT 84.95 97.29 85.16 97.36 ;
    RECT 84.95 97.65 85.16 97.72 ;
    RECT 84.95 98.01 85.16 98.08 ;
    RECT 81.17 97.29 81.38 97.36 ;
    RECT 81.17 97.65 81.38 97.72 ;
    RECT 81.17 98.01 81.38 98.08 ;
    RECT 81.63 97.29 81.84 97.36 ;
    RECT 81.63 97.65 81.84 97.72 ;
    RECT 81.63 98.01 81.84 98.08 ;
    RECT 77.85 97.29 78.06 97.36 ;
    RECT 77.85 97.65 78.06 97.72 ;
    RECT 77.85 98.01 78.06 98.08 ;
    RECT 78.31 97.29 78.52 97.36 ;
    RECT 78.31 97.65 78.52 97.72 ;
    RECT 78.31 98.01 78.52 98.08 ;
    RECT 74.53 97.29 74.74 97.36 ;
    RECT 74.53 97.65 74.74 97.72 ;
    RECT 74.53 98.01 74.74 98.08 ;
    RECT 74.99 97.29 75.2 97.36 ;
    RECT 74.99 97.65 75.2 97.72 ;
    RECT 74.99 98.01 75.2 98.08 ;
    RECT 71.21 97.29 71.42 97.36 ;
    RECT 71.21 97.65 71.42 97.72 ;
    RECT 71.21 98.01 71.42 98.08 ;
    RECT 71.67 97.29 71.88 97.36 ;
    RECT 71.67 97.65 71.88 97.72 ;
    RECT 71.67 98.01 71.88 98.08 ;
    RECT 31.37 97.29 31.58 97.36 ;
    RECT 31.37 97.65 31.58 97.72 ;
    RECT 31.37 98.01 31.58 98.08 ;
    RECT 31.83 97.29 32.04 97.36 ;
    RECT 31.83 97.65 32.04 97.72 ;
    RECT 31.83 98.01 32.04 98.08 ;
    RECT 67.89 97.29 68.1 97.36 ;
    RECT 67.89 97.65 68.1 97.72 ;
    RECT 67.89 98.01 68.1 98.08 ;
    RECT 68.35 97.29 68.56 97.36 ;
    RECT 68.35 97.65 68.56 97.72 ;
    RECT 68.35 98.01 68.56 98.08 ;
    RECT 28.05 97.29 28.26 97.36 ;
    RECT 28.05 97.65 28.26 97.72 ;
    RECT 28.05 98.01 28.26 98.08 ;
    RECT 28.51 97.29 28.72 97.36 ;
    RECT 28.51 97.65 28.72 97.72 ;
    RECT 28.51 98.01 28.72 98.08 ;
    RECT 24.73 97.29 24.94 97.36 ;
    RECT 24.73 97.65 24.94 97.72 ;
    RECT 24.73 98.01 24.94 98.08 ;
    RECT 25.19 97.29 25.4 97.36 ;
    RECT 25.19 97.65 25.4 97.72 ;
    RECT 25.19 98.01 25.4 98.08 ;
    RECT 21.41 97.29 21.62 97.36 ;
    RECT 21.41 97.65 21.62 97.72 ;
    RECT 21.41 98.01 21.62 98.08 ;
    RECT 21.87 97.29 22.08 97.36 ;
    RECT 21.87 97.65 22.08 97.72 ;
    RECT 21.87 98.01 22.08 98.08 ;
    RECT 18.09 97.29 18.3 97.36 ;
    RECT 18.09 97.65 18.3 97.72 ;
    RECT 18.09 98.01 18.3 98.08 ;
    RECT 18.55 97.29 18.76 97.36 ;
    RECT 18.55 97.65 18.76 97.72 ;
    RECT 18.55 98.01 18.76 98.08 ;
    RECT 120.825 97.65 120.895 97.72 ;
    RECT 14.77 97.29 14.98 97.36 ;
    RECT 14.77 97.65 14.98 97.72 ;
    RECT 14.77 98.01 14.98 98.08 ;
    RECT 15.23 97.29 15.44 97.36 ;
    RECT 15.23 97.65 15.44 97.72 ;
    RECT 15.23 98.01 15.44 98.08 ;
    RECT 11.45 97.29 11.66 97.36 ;
    RECT 11.45 97.65 11.66 97.72 ;
    RECT 11.45 98.01 11.66 98.08 ;
    RECT 11.91 97.29 12.12 97.36 ;
    RECT 11.91 97.65 12.12 97.72 ;
    RECT 11.91 98.01 12.12 98.08 ;
    RECT 8.13 97.29 8.34 97.36 ;
    RECT 8.13 97.65 8.34 97.72 ;
    RECT 8.13 98.01 8.34 98.08 ;
    RECT 8.59 97.29 8.8 97.36 ;
    RECT 8.59 97.65 8.8 97.72 ;
    RECT 8.59 98.01 8.8 98.08 ;
    RECT 4.81 97.29 5.02 97.36 ;
    RECT 4.81 97.65 5.02 97.72 ;
    RECT 4.81 98.01 5.02 98.08 ;
    RECT 5.27 97.29 5.48 97.36 ;
    RECT 5.27 97.65 5.48 97.72 ;
    RECT 5.27 98.01 5.48 98.08 ;
    RECT 1.49 97.29 1.7 97.36 ;
    RECT 1.49 97.65 1.7 97.72 ;
    RECT 1.49 98.01 1.7 98.08 ;
    RECT 1.95 97.29 2.16 97.36 ;
    RECT 1.95 97.65 2.16 97.72 ;
    RECT 1.95 98.01 2.16 98.08 ;
    RECT 64.57 97.29 64.78 97.36 ;
    RECT 64.57 97.65 64.78 97.72 ;
    RECT 64.57 98.01 64.78 98.08 ;
    RECT 65.03 97.29 65.24 97.36 ;
    RECT 65.03 97.65 65.24 97.72 ;
    RECT 65.03 98.01 65.24 98.08 ;
    RECT 61.25 96.57 61.46 96.64 ;
    RECT 61.25 96.93 61.46 97.0 ;
    RECT 61.25 97.29 61.46 97.36 ;
    RECT 61.71 96.57 61.92 96.64 ;
    RECT 61.71 96.93 61.92 97.0 ;
    RECT 61.71 97.29 61.92 97.36 ;
    RECT 57.93 96.57 58.14 96.64 ;
    RECT 57.93 96.93 58.14 97.0 ;
    RECT 57.93 97.29 58.14 97.36 ;
    RECT 58.39 96.57 58.6 96.64 ;
    RECT 58.39 96.93 58.6 97.0 ;
    RECT 58.39 97.29 58.6 97.36 ;
    RECT 54.61 96.57 54.82 96.64 ;
    RECT 54.61 96.93 54.82 97.0 ;
    RECT 54.61 97.29 54.82 97.36 ;
    RECT 55.07 96.57 55.28 96.64 ;
    RECT 55.07 96.93 55.28 97.0 ;
    RECT 55.07 97.29 55.28 97.36 ;
    RECT 51.29 96.57 51.5 96.64 ;
    RECT 51.29 96.93 51.5 97.0 ;
    RECT 51.29 97.29 51.5 97.36 ;
    RECT 51.75 96.57 51.96 96.64 ;
    RECT 51.75 96.93 51.96 97.0 ;
    RECT 51.75 97.29 51.96 97.36 ;
    RECT 47.97 96.57 48.18 96.64 ;
    RECT 47.97 96.93 48.18 97.0 ;
    RECT 47.97 97.29 48.18 97.36 ;
    RECT 48.43 96.57 48.64 96.64 ;
    RECT 48.43 96.93 48.64 97.0 ;
    RECT 48.43 97.29 48.64 97.36 ;
    RECT 44.65 96.57 44.86 96.64 ;
    RECT 44.65 96.93 44.86 97.0 ;
    RECT 44.65 97.29 44.86 97.36 ;
    RECT 45.11 96.57 45.32 96.64 ;
    RECT 45.11 96.93 45.32 97.0 ;
    RECT 45.11 97.29 45.32 97.36 ;
    RECT 41.33 96.57 41.54 96.64 ;
    RECT 41.33 96.93 41.54 97.0 ;
    RECT 41.33 97.29 41.54 97.36 ;
    RECT 41.79 96.57 42.0 96.64 ;
    RECT 41.79 96.93 42.0 97.0 ;
    RECT 41.79 97.29 42.0 97.36 ;
    RECT 38.01 96.57 38.22 96.64 ;
    RECT 38.01 96.93 38.22 97.0 ;
    RECT 38.01 97.29 38.22 97.36 ;
    RECT 38.47 96.57 38.68 96.64 ;
    RECT 38.47 96.93 38.68 97.0 ;
    RECT 38.47 97.29 38.68 97.36 ;
    RECT 0.4 96.93 0.47 97.0 ;
    RECT 34.69 96.57 34.9 96.64 ;
    RECT 34.69 96.93 34.9 97.0 ;
    RECT 34.69 97.29 34.9 97.36 ;
    RECT 35.15 96.57 35.36 96.64 ;
    RECT 35.15 96.93 35.36 97.0 ;
    RECT 35.15 97.29 35.36 97.36 ;
    RECT 117.69 96.57 117.9 96.64 ;
    RECT 117.69 96.93 117.9 97.0 ;
    RECT 117.69 97.29 117.9 97.36 ;
    RECT 118.15 96.57 118.36 96.64 ;
    RECT 118.15 96.93 118.36 97.0 ;
    RECT 118.15 97.29 118.36 97.36 ;
    RECT 114.37 96.57 114.58 96.64 ;
    RECT 114.37 96.93 114.58 97.0 ;
    RECT 114.37 97.29 114.58 97.36 ;
    RECT 114.83 96.57 115.04 96.64 ;
    RECT 114.83 96.93 115.04 97.0 ;
    RECT 114.83 97.29 115.04 97.36 ;
    RECT 111.05 96.57 111.26 96.64 ;
    RECT 111.05 96.93 111.26 97.0 ;
    RECT 111.05 97.29 111.26 97.36 ;
    RECT 111.51 96.57 111.72 96.64 ;
    RECT 111.51 96.93 111.72 97.0 ;
    RECT 111.51 97.29 111.72 97.36 ;
    RECT 107.73 96.57 107.94 96.64 ;
    RECT 107.73 96.93 107.94 97.0 ;
    RECT 107.73 97.29 107.94 97.36 ;
    RECT 108.19 96.57 108.4 96.64 ;
    RECT 108.19 96.93 108.4 97.0 ;
    RECT 108.19 97.29 108.4 97.36 ;
    RECT 104.41 96.57 104.62 96.64 ;
    RECT 104.41 96.93 104.62 97.0 ;
    RECT 104.41 97.29 104.62 97.36 ;
    RECT 104.87 96.57 105.08 96.64 ;
    RECT 104.87 96.93 105.08 97.0 ;
    RECT 104.87 97.29 105.08 97.36 ;
    RECT 101.09 96.57 101.3 96.64 ;
    RECT 101.09 96.93 101.3 97.0 ;
    RECT 101.09 97.29 101.3 97.36 ;
    RECT 101.55 96.57 101.76 96.64 ;
    RECT 101.55 96.93 101.76 97.0 ;
    RECT 101.55 97.29 101.76 97.36 ;
    RECT 97.77 96.57 97.98 96.64 ;
    RECT 97.77 96.93 97.98 97.0 ;
    RECT 97.77 97.29 97.98 97.36 ;
    RECT 98.23 96.57 98.44 96.64 ;
    RECT 98.23 96.93 98.44 97.0 ;
    RECT 98.23 97.29 98.44 97.36 ;
    RECT 94.45 96.57 94.66 96.64 ;
    RECT 94.45 96.93 94.66 97.0 ;
    RECT 94.45 97.29 94.66 97.36 ;
    RECT 94.91 96.57 95.12 96.64 ;
    RECT 94.91 96.93 95.12 97.0 ;
    RECT 94.91 97.29 95.12 97.36 ;
    RECT 91.13 96.57 91.34 96.64 ;
    RECT 91.13 96.93 91.34 97.0 ;
    RECT 91.13 97.29 91.34 97.36 ;
    RECT 91.59 96.57 91.8 96.64 ;
    RECT 91.59 96.93 91.8 97.0 ;
    RECT 91.59 97.29 91.8 97.36 ;
    RECT 87.81 96.57 88.02 96.64 ;
    RECT 87.81 96.93 88.02 97.0 ;
    RECT 87.81 97.29 88.02 97.36 ;
    RECT 88.27 96.57 88.48 96.64 ;
    RECT 88.27 96.93 88.48 97.0 ;
    RECT 88.27 97.29 88.48 97.36 ;
    RECT 84.49 96.57 84.7 96.64 ;
    RECT 84.49 96.93 84.7 97.0 ;
    RECT 84.49 97.29 84.7 97.36 ;
    RECT 84.95 96.57 85.16 96.64 ;
    RECT 84.95 96.93 85.16 97.0 ;
    RECT 84.95 97.29 85.16 97.36 ;
    RECT 81.17 96.57 81.38 96.64 ;
    RECT 81.17 96.93 81.38 97.0 ;
    RECT 81.17 97.29 81.38 97.36 ;
    RECT 81.63 96.57 81.84 96.64 ;
    RECT 81.63 96.93 81.84 97.0 ;
    RECT 81.63 97.29 81.84 97.36 ;
    RECT 77.85 96.57 78.06 96.64 ;
    RECT 77.85 96.93 78.06 97.0 ;
    RECT 77.85 97.29 78.06 97.36 ;
    RECT 78.31 96.57 78.52 96.64 ;
    RECT 78.31 96.93 78.52 97.0 ;
    RECT 78.31 97.29 78.52 97.36 ;
    RECT 74.53 96.57 74.74 96.64 ;
    RECT 74.53 96.93 74.74 97.0 ;
    RECT 74.53 97.29 74.74 97.36 ;
    RECT 74.99 96.57 75.2 96.64 ;
    RECT 74.99 96.93 75.2 97.0 ;
    RECT 74.99 97.29 75.2 97.36 ;
    RECT 71.21 96.57 71.42 96.64 ;
    RECT 71.21 96.93 71.42 97.0 ;
    RECT 71.21 97.29 71.42 97.36 ;
    RECT 71.67 96.57 71.88 96.64 ;
    RECT 71.67 96.93 71.88 97.0 ;
    RECT 71.67 97.29 71.88 97.36 ;
    RECT 31.37 96.57 31.58 96.64 ;
    RECT 31.37 96.93 31.58 97.0 ;
    RECT 31.37 97.29 31.58 97.36 ;
    RECT 31.83 96.57 32.04 96.64 ;
    RECT 31.83 96.93 32.04 97.0 ;
    RECT 31.83 97.29 32.04 97.36 ;
    RECT 67.89 96.57 68.1 96.64 ;
    RECT 67.89 96.93 68.1 97.0 ;
    RECT 67.89 97.29 68.1 97.36 ;
    RECT 68.35 96.57 68.56 96.64 ;
    RECT 68.35 96.93 68.56 97.0 ;
    RECT 68.35 97.29 68.56 97.36 ;
    RECT 28.05 96.57 28.26 96.64 ;
    RECT 28.05 96.93 28.26 97.0 ;
    RECT 28.05 97.29 28.26 97.36 ;
    RECT 28.51 96.57 28.72 96.64 ;
    RECT 28.51 96.93 28.72 97.0 ;
    RECT 28.51 97.29 28.72 97.36 ;
    RECT 24.73 96.57 24.94 96.64 ;
    RECT 24.73 96.93 24.94 97.0 ;
    RECT 24.73 97.29 24.94 97.36 ;
    RECT 25.19 96.57 25.4 96.64 ;
    RECT 25.19 96.93 25.4 97.0 ;
    RECT 25.19 97.29 25.4 97.36 ;
    RECT 21.41 96.57 21.62 96.64 ;
    RECT 21.41 96.93 21.62 97.0 ;
    RECT 21.41 97.29 21.62 97.36 ;
    RECT 21.87 96.57 22.08 96.64 ;
    RECT 21.87 96.93 22.08 97.0 ;
    RECT 21.87 97.29 22.08 97.36 ;
    RECT 18.09 96.57 18.3 96.64 ;
    RECT 18.09 96.93 18.3 97.0 ;
    RECT 18.09 97.29 18.3 97.36 ;
    RECT 18.55 96.57 18.76 96.64 ;
    RECT 18.55 96.93 18.76 97.0 ;
    RECT 18.55 97.29 18.76 97.36 ;
    RECT 120.825 96.93 120.895 97.0 ;
    RECT 14.77 96.57 14.98 96.64 ;
    RECT 14.77 96.93 14.98 97.0 ;
    RECT 14.77 97.29 14.98 97.36 ;
    RECT 15.23 96.57 15.44 96.64 ;
    RECT 15.23 96.93 15.44 97.0 ;
    RECT 15.23 97.29 15.44 97.36 ;
    RECT 11.45 96.57 11.66 96.64 ;
    RECT 11.45 96.93 11.66 97.0 ;
    RECT 11.45 97.29 11.66 97.36 ;
    RECT 11.91 96.57 12.12 96.64 ;
    RECT 11.91 96.93 12.12 97.0 ;
    RECT 11.91 97.29 12.12 97.36 ;
    RECT 8.13 96.57 8.34 96.64 ;
    RECT 8.13 96.93 8.34 97.0 ;
    RECT 8.13 97.29 8.34 97.36 ;
    RECT 8.59 96.57 8.8 96.64 ;
    RECT 8.59 96.93 8.8 97.0 ;
    RECT 8.59 97.29 8.8 97.36 ;
    RECT 4.81 96.57 5.02 96.64 ;
    RECT 4.81 96.93 5.02 97.0 ;
    RECT 4.81 97.29 5.02 97.36 ;
    RECT 5.27 96.57 5.48 96.64 ;
    RECT 5.27 96.93 5.48 97.0 ;
    RECT 5.27 97.29 5.48 97.36 ;
    RECT 1.49 96.57 1.7 96.64 ;
    RECT 1.49 96.93 1.7 97.0 ;
    RECT 1.49 97.29 1.7 97.36 ;
    RECT 1.95 96.57 2.16 96.64 ;
    RECT 1.95 96.93 2.16 97.0 ;
    RECT 1.95 97.29 2.16 97.36 ;
    RECT 64.57 96.57 64.78 96.64 ;
    RECT 64.57 96.93 64.78 97.0 ;
    RECT 64.57 97.29 64.78 97.36 ;
    RECT 65.03 96.57 65.24 96.64 ;
    RECT 65.03 96.93 65.24 97.0 ;
    RECT 65.03 97.29 65.24 97.36 ;
    RECT 61.25 95.85 61.46 95.92 ;
    RECT 61.25 96.21 61.46 96.28 ;
    RECT 61.25 96.57 61.46 96.64 ;
    RECT 61.71 95.85 61.92 95.92 ;
    RECT 61.71 96.21 61.92 96.28 ;
    RECT 61.71 96.57 61.92 96.64 ;
    RECT 57.93 95.85 58.14 95.92 ;
    RECT 57.93 96.21 58.14 96.28 ;
    RECT 57.93 96.57 58.14 96.64 ;
    RECT 58.39 95.85 58.6 95.92 ;
    RECT 58.39 96.21 58.6 96.28 ;
    RECT 58.39 96.57 58.6 96.64 ;
    RECT 54.61 95.85 54.82 95.92 ;
    RECT 54.61 96.21 54.82 96.28 ;
    RECT 54.61 96.57 54.82 96.64 ;
    RECT 55.07 95.85 55.28 95.92 ;
    RECT 55.07 96.21 55.28 96.28 ;
    RECT 55.07 96.57 55.28 96.64 ;
    RECT 51.29 95.85 51.5 95.92 ;
    RECT 51.29 96.21 51.5 96.28 ;
    RECT 51.29 96.57 51.5 96.64 ;
    RECT 51.75 95.85 51.96 95.92 ;
    RECT 51.75 96.21 51.96 96.28 ;
    RECT 51.75 96.57 51.96 96.64 ;
    RECT 47.97 95.85 48.18 95.92 ;
    RECT 47.97 96.21 48.18 96.28 ;
    RECT 47.97 96.57 48.18 96.64 ;
    RECT 48.43 95.85 48.64 95.92 ;
    RECT 48.43 96.21 48.64 96.28 ;
    RECT 48.43 96.57 48.64 96.64 ;
    RECT 44.65 95.85 44.86 95.92 ;
    RECT 44.65 96.21 44.86 96.28 ;
    RECT 44.65 96.57 44.86 96.64 ;
    RECT 45.11 95.85 45.32 95.92 ;
    RECT 45.11 96.21 45.32 96.28 ;
    RECT 45.11 96.57 45.32 96.64 ;
    RECT 41.33 95.85 41.54 95.92 ;
    RECT 41.33 96.21 41.54 96.28 ;
    RECT 41.33 96.57 41.54 96.64 ;
    RECT 41.79 95.85 42.0 95.92 ;
    RECT 41.79 96.21 42.0 96.28 ;
    RECT 41.79 96.57 42.0 96.64 ;
    RECT 38.01 95.85 38.22 95.92 ;
    RECT 38.01 96.21 38.22 96.28 ;
    RECT 38.01 96.57 38.22 96.64 ;
    RECT 38.47 95.85 38.68 95.92 ;
    RECT 38.47 96.21 38.68 96.28 ;
    RECT 38.47 96.57 38.68 96.64 ;
    RECT 0.4 96.21 0.47 96.28 ;
    RECT 34.69 95.85 34.9 95.92 ;
    RECT 34.69 96.21 34.9 96.28 ;
    RECT 34.69 96.57 34.9 96.64 ;
    RECT 35.15 95.85 35.36 95.92 ;
    RECT 35.15 96.21 35.36 96.28 ;
    RECT 35.15 96.57 35.36 96.64 ;
    RECT 117.69 95.85 117.9 95.92 ;
    RECT 117.69 96.21 117.9 96.28 ;
    RECT 117.69 96.57 117.9 96.64 ;
    RECT 118.15 95.85 118.36 95.92 ;
    RECT 118.15 96.21 118.36 96.28 ;
    RECT 118.15 96.57 118.36 96.64 ;
    RECT 114.37 95.85 114.58 95.92 ;
    RECT 114.37 96.21 114.58 96.28 ;
    RECT 114.37 96.57 114.58 96.64 ;
    RECT 114.83 95.85 115.04 95.92 ;
    RECT 114.83 96.21 115.04 96.28 ;
    RECT 114.83 96.57 115.04 96.64 ;
    RECT 111.05 95.85 111.26 95.92 ;
    RECT 111.05 96.21 111.26 96.28 ;
    RECT 111.05 96.57 111.26 96.64 ;
    RECT 111.51 95.85 111.72 95.92 ;
    RECT 111.51 96.21 111.72 96.28 ;
    RECT 111.51 96.57 111.72 96.64 ;
    RECT 107.73 95.85 107.94 95.92 ;
    RECT 107.73 96.21 107.94 96.28 ;
    RECT 107.73 96.57 107.94 96.64 ;
    RECT 108.19 95.85 108.4 95.92 ;
    RECT 108.19 96.21 108.4 96.28 ;
    RECT 108.19 96.57 108.4 96.64 ;
    RECT 104.41 95.85 104.62 95.92 ;
    RECT 104.41 96.21 104.62 96.28 ;
    RECT 104.41 96.57 104.62 96.64 ;
    RECT 104.87 95.85 105.08 95.92 ;
    RECT 104.87 96.21 105.08 96.28 ;
    RECT 104.87 96.57 105.08 96.64 ;
    RECT 101.09 95.85 101.3 95.92 ;
    RECT 101.09 96.21 101.3 96.28 ;
    RECT 101.09 96.57 101.3 96.64 ;
    RECT 101.55 95.85 101.76 95.92 ;
    RECT 101.55 96.21 101.76 96.28 ;
    RECT 101.55 96.57 101.76 96.64 ;
    RECT 97.77 95.85 97.98 95.92 ;
    RECT 97.77 96.21 97.98 96.28 ;
    RECT 97.77 96.57 97.98 96.64 ;
    RECT 98.23 95.85 98.44 95.92 ;
    RECT 98.23 96.21 98.44 96.28 ;
    RECT 98.23 96.57 98.44 96.64 ;
    RECT 94.45 95.85 94.66 95.92 ;
    RECT 94.45 96.21 94.66 96.28 ;
    RECT 94.45 96.57 94.66 96.64 ;
    RECT 94.91 95.85 95.12 95.92 ;
    RECT 94.91 96.21 95.12 96.28 ;
    RECT 94.91 96.57 95.12 96.64 ;
    RECT 91.13 95.85 91.34 95.92 ;
    RECT 91.13 96.21 91.34 96.28 ;
    RECT 91.13 96.57 91.34 96.64 ;
    RECT 91.59 95.85 91.8 95.92 ;
    RECT 91.59 96.21 91.8 96.28 ;
    RECT 91.59 96.57 91.8 96.64 ;
    RECT 87.81 95.85 88.02 95.92 ;
    RECT 87.81 96.21 88.02 96.28 ;
    RECT 87.81 96.57 88.02 96.64 ;
    RECT 88.27 95.85 88.48 95.92 ;
    RECT 88.27 96.21 88.48 96.28 ;
    RECT 88.27 96.57 88.48 96.64 ;
    RECT 84.49 95.85 84.7 95.92 ;
    RECT 84.49 96.21 84.7 96.28 ;
    RECT 84.49 96.57 84.7 96.64 ;
    RECT 84.95 95.85 85.16 95.92 ;
    RECT 84.95 96.21 85.16 96.28 ;
    RECT 84.95 96.57 85.16 96.64 ;
    RECT 81.17 95.85 81.38 95.92 ;
    RECT 81.17 96.21 81.38 96.28 ;
    RECT 81.17 96.57 81.38 96.64 ;
    RECT 81.63 95.85 81.84 95.92 ;
    RECT 81.63 96.21 81.84 96.28 ;
    RECT 81.63 96.57 81.84 96.64 ;
    RECT 77.85 95.85 78.06 95.92 ;
    RECT 77.85 96.21 78.06 96.28 ;
    RECT 77.85 96.57 78.06 96.64 ;
    RECT 78.31 95.85 78.52 95.92 ;
    RECT 78.31 96.21 78.52 96.28 ;
    RECT 78.31 96.57 78.52 96.64 ;
    RECT 74.53 95.85 74.74 95.92 ;
    RECT 74.53 96.21 74.74 96.28 ;
    RECT 74.53 96.57 74.74 96.64 ;
    RECT 74.99 95.85 75.2 95.92 ;
    RECT 74.99 96.21 75.2 96.28 ;
    RECT 74.99 96.57 75.2 96.64 ;
    RECT 71.21 95.85 71.42 95.92 ;
    RECT 71.21 96.21 71.42 96.28 ;
    RECT 71.21 96.57 71.42 96.64 ;
    RECT 71.67 95.85 71.88 95.92 ;
    RECT 71.67 96.21 71.88 96.28 ;
    RECT 71.67 96.57 71.88 96.64 ;
    RECT 31.37 95.85 31.58 95.92 ;
    RECT 31.37 96.21 31.58 96.28 ;
    RECT 31.37 96.57 31.58 96.64 ;
    RECT 31.83 95.85 32.04 95.92 ;
    RECT 31.83 96.21 32.04 96.28 ;
    RECT 31.83 96.57 32.04 96.64 ;
    RECT 67.89 95.85 68.1 95.92 ;
    RECT 67.89 96.21 68.1 96.28 ;
    RECT 67.89 96.57 68.1 96.64 ;
    RECT 68.35 95.85 68.56 95.92 ;
    RECT 68.35 96.21 68.56 96.28 ;
    RECT 68.35 96.57 68.56 96.64 ;
    RECT 28.05 95.85 28.26 95.92 ;
    RECT 28.05 96.21 28.26 96.28 ;
    RECT 28.05 96.57 28.26 96.64 ;
    RECT 28.51 95.85 28.72 95.92 ;
    RECT 28.51 96.21 28.72 96.28 ;
    RECT 28.51 96.57 28.72 96.64 ;
    RECT 24.73 95.85 24.94 95.92 ;
    RECT 24.73 96.21 24.94 96.28 ;
    RECT 24.73 96.57 24.94 96.64 ;
    RECT 25.19 95.85 25.4 95.92 ;
    RECT 25.19 96.21 25.4 96.28 ;
    RECT 25.19 96.57 25.4 96.64 ;
    RECT 21.41 95.85 21.62 95.92 ;
    RECT 21.41 96.21 21.62 96.28 ;
    RECT 21.41 96.57 21.62 96.64 ;
    RECT 21.87 95.85 22.08 95.92 ;
    RECT 21.87 96.21 22.08 96.28 ;
    RECT 21.87 96.57 22.08 96.64 ;
    RECT 18.09 95.85 18.3 95.92 ;
    RECT 18.09 96.21 18.3 96.28 ;
    RECT 18.09 96.57 18.3 96.64 ;
    RECT 18.55 95.85 18.76 95.92 ;
    RECT 18.55 96.21 18.76 96.28 ;
    RECT 18.55 96.57 18.76 96.64 ;
    RECT 120.825 96.21 120.895 96.28 ;
    RECT 14.77 95.85 14.98 95.92 ;
    RECT 14.77 96.21 14.98 96.28 ;
    RECT 14.77 96.57 14.98 96.64 ;
    RECT 15.23 95.85 15.44 95.92 ;
    RECT 15.23 96.21 15.44 96.28 ;
    RECT 15.23 96.57 15.44 96.64 ;
    RECT 11.45 95.85 11.66 95.92 ;
    RECT 11.45 96.21 11.66 96.28 ;
    RECT 11.45 96.57 11.66 96.64 ;
    RECT 11.91 95.85 12.12 95.92 ;
    RECT 11.91 96.21 12.12 96.28 ;
    RECT 11.91 96.57 12.12 96.64 ;
    RECT 8.13 95.85 8.34 95.92 ;
    RECT 8.13 96.21 8.34 96.28 ;
    RECT 8.13 96.57 8.34 96.64 ;
    RECT 8.59 95.85 8.8 95.92 ;
    RECT 8.59 96.21 8.8 96.28 ;
    RECT 8.59 96.57 8.8 96.64 ;
    RECT 4.81 95.85 5.02 95.92 ;
    RECT 4.81 96.21 5.02 96.28 ;
    RECT 4.81 96.57 5.02 96.64 ;
    RECT 5.27 95.85 5.48 95.92 ;
    RECT 5.27 96.21 5.48 96.28 ;
    RECT 5.27 96.57 5.48 96.64 ;
    RECT 1.49 95.85 1.7 95.92 ;
    RECT 1.49 96.21 1.7 96.28 ;
    RECT 1.49 96.57 1.7 96.64 ;
    RECT 1.95 95.85 2.16 95.92 ;
    RECT 1.95 96.21 2.16 96.28 ;
    RECT 1.95 96.57 2.16 96.64 ;
    RECT 64.57 95.85 64.78 95.92 ;
    RECT 64.57 96.21 64.78 96.28 ;
    RECT 64.57 96.57 64.78 96.64 ;
    RECT 65.03 95.85 65.24 95.92 ;
    RECT 65.03 96.21 65.24 96.28 ;
    RECT 65.03 96.57 65.24 96.64 ;
    RECT 61.25 95.13 61.46 95.2 ;
    RECT 61.25 95.49 61.46 95.56 ;
    RECT 61.25 95.85 61.46 95.92 ;
    RECT 61.71 95.13 61.92 95.2 ;
    RECT 61.71 95.49 61.92 95.56 ;
    RECT 61.71 95.85 61.92 95.92 ;
    RECT 57.93 95.13 58.14 95.2 ;
    RECT 57.93 95.49 58.14 95.56 ;
    RECT 57.93 95.85 58.14 95.92 ;
    RECT 58.39 95.13 58.6 95.2 ;
    RECT 58.39 95.49 58.6 95.56 ;
    RECT 58.39 95.85 58.6 95.92 ;
    RECT 54.61 95.13 54.82 95.2 ;
    RECT 54.61 95.49 54.82 95.56 ;
    RECT 54.61 95.85 54.82 95.92 ;
    RECT 55.07 95.13 55.28 95.2 ;
    RECT 55.07 95.49 55.28 95.56 ;
    RECT 55.07 95.85 55.28 95.92 ;
    RECT 51.29 95.13 51.5 95.2 ;
    RECT 51.29 95.49 51.5 95.56 ;
    RECT 51.29 95.85 51.5 95.92 ;
    RECT 51.75 95.13 51.96 95.2 ;
    RECT 51.75 95.49 51.96 95.56 ;
    RECT 51.75 95.85 51.96 95.92 ;
    RECT 47.97 95.13 48.18 95.2 ;
    RECT 47.97 95.49 48.18 95.56 ;
    RECT 47.97 95.85 48.18 95.92 ;
    RECT 48.43 95.13 48.64 95.2 ;
    RECT 48.43 95.49 48.64 95.56 ;
    RECT 48.43 95.85 48.64 95.92 ;
    RECT 44.65 95.13 44.86 95.2 ;
    RECT 44.65 95.49 44.86 95.56 ;
    RECT 44.65 95.85 44.86 95.92 ;
    RECT 45.11 95.13 45.32 95.2 ;
    RECT 45.11 95.49 45.32 95.56 ;
    RECT 45.11 95.85 45.32 95.92 ;
    RECT 41.33 95.13 41.54 95.2 ;
    RECT 41.33 95.49 41.54 95.56 ;
    RECT 41.33 95.85 41.54 95.92 ;
    RECT 41.79 95.13 42.0 95.2 ;
    RECT 41.79 95.49 42.0 95.56 ;
    RECT 41.79 95.85 42.0 95.92 ;
    RECT 38.01 95.13 38.22 95.2 ;
    RECT 38.01 95.49 38.22 95.56 ;
    RECT 38.01 95.85 38.22 95.92 ;
    RECT 38.47 95.13 38.68 95.2 ;
    RECT 38.47 95.49 38.68 95.56 ;
    RECT 38.47 95.85 38.68 95.92 ;
    RECT 0.4 95.49 0.47 95.56 ;
    RECT 34.69 95.13 34.9 95.2 ;
    RECT 34.69 95.49 34.9 95.56 ;
    RECT 34.69 95.85 34.9 95.92 ;
    RECT 35.15 95.13 35.36 95.2 ;
    RECT 35.15 95.49 35.36 95.56 ;
    RECT 35.15 95.85 35.36 95.92 ;
    RECT 117.69 95.13 117.9 95.2 ;
    RECT 117.69 95.49 117.9 95.56 ;
    RECT 117.69 95.85 117.9 95.92 ;
    RECT 118.15 95.13 118.36 95.2 ;
    RECT 118.15 95.49 118.36 95.56 ;
    RECT 118.15 95.85 118.36 95.92 ;
    RECT 114.37 95.13 114.58 95.2 ;
    RECT 114.37 95.49 114.58 95.56 ;
    RECT 114.37 95.85 114.58 95.92 ;
    RECT 114.83 95.13 115.04 95.2 ;
    RECT 114.83 95.49 115.04 95.56 ;
    RECT 114.83 95.85 115.04 95.92 ;
    RECT 111.05 95.13 111.26 95.2 ;
    RECT 111.05 95.49 111.26 95.56 ;
    RECT 111.05 95.85 111.26 95.92 ;
    RECT 111.51 95.13 111.72 95.2 ;
    RECT 111.51 95.49 111.72 95.56 ;
    RECT 111.51 95.85 111.72 95.92 ;
    RECT 107.73 95.13 107.94 95.2 ;
    RECT 107.73 95.49 107.94 95.56 ;
    RECT 107.73 95.85 107.94 95.92 ;
    RECT 108.19 95.13 108.4 95.2 ;
    RECT 108.19 95.49 108.4 95.56 ;
    RECT 108.19 95.85 108.4 95.92 ;
    RECT 104.41 95.13 104.62 95.2 ;
    RECT 104.41 95.49 104.62 95.56 ;
    RECT 104.41 95.85 104.62 95.92 ;
    RECT 104.87 95.13 105.08 95.2 ;
    RECT 104.87 95.49 105.08 95.56 ;
    RECT 104.87 95.85 105.08 95.92 ;
    RECT 101.09 95.13 101.3 95.2 ;
    RECT 101.09 95.49 101.3 95.56 ;
    RECT 101.09 95.85 101.3 95.92 ;
    RECT 101.55 95.13 101.76 95.2 ;
    RECT 101.55 95.49 101.76 95.56 ;
    RECT 101.55 95.85 101.76 95.92 ;
    RECT 97.77 95.13 97.98 95.2 ;
    RECT 97.77 95.49 97.98 95.56 ;
    RECT 97.77 95.85 97.98 95.92 ;
    RECT 98.23 95.13 98.44 95.2 ;
    RECT 98.23 95.49 98.44 95.56 ;
    RECT 98.23 95.85 98.44 95.92 ;
    RECT 94.45 95.13 94.66 95.2 ;
    RECT 94.45 95.49 94.66 95.56 ;
    RECT 94.45 95.85 94.66 95.92 ;
    RECT 94.91 95.13 95.12 95.2 ;
    RECT 94.91 95.49 95.12 95.56 ;
    RECT 94.91 95.85 95.12 95.92 ;
    RECT 91.13 95.13 91.34 95.2 ;
    RECT 91.13 95.49 91.34 95.56 ;
    RECT 91.13 95.85 91.34 95.92 ;
    RECT 91.59 95.13 91.8 95.2 ;
    RECT 91.59 95.49 91.8 95.56 ;
    RECT 91.59 95.85 91.8 95.92 ;
    RECT 87.81 95.13 88.02 95.2 ;
    RECT 87.81 95.49 88.02 95.56 ;
    RECT 87.81 95.85 88.02 95.92 ;
    RECT 88.27 95.13 88.48 95.2 ;
    RECT 88.27 95.49 88.48 95.56 ;
    RECT 88.27 95.85 88.48 95.92 ;
    RECT 84.49 95.13 84.7 95.2 ;
    RECT 84.49 95.49 84.7 95.56 ;
    RECT 84.49 95.85 84.7 95.92 ;
    RECT 84.95 95.13 85.16 95.2 ;
    RECT 84.95 95.49 85.16 95.56 ;
    RECT 84.95 95.85 85.16 95.92 ;
    RECT 81.17 95.13 81.38 95.2 ;
    RECT 81.17 95.49 81.38 95.56 ;
    RECT 81.17 95.85 81.38 95.92 ;
    RECT 81.63 95.13 81.84 95.2 ;
    RECT 81.63 95.49 81.84 95.56 ;
    RECT 81.63 95.85 81.84 95.92 ;
    RECT 77.85 95.13 78.06 95.2 ;
    RECT 77.85 95.49 78.06 95.56 ;
    RECT 77.85 95.85 78.06 95.92 ;
    RECT 78.31 95.13 78.52 95.2 ;
    RECT 78.31 95.49 78.52 95.56 ;
    RECT 78.31 95.85 78.52 95.92 ;
    RECT 74.53 95.13 74.74 95.2 ;
    RECT 74.53 95.49 74.74 95.56 ;
    RECT 74.53 95.85 74.74 95.92 ;
    RECT 74.99 95.13 75.2 95.2 ;
    RECT 74.99 95.49 75.2 95.56 ;
    RECT 74.99 95.85 75.2 95.92 ;
    RECT 71.21 95.13 71.42 95.2 ;
    RECT 71.21 95.49 71.42 95.56 ;
    RECT 71.21 95.85 71.42 95.92 ;
    RECT 71.67 95.13 71.88 95.2 ;
    RECT 71.67 95.49 71.88 95.56 ;
    RECT 71.67 95.85 71.88 95.92 ;
    RECT 31.37 95.13 31.58 95.2 ;
    RECT 31.37 95.49 31.58 95.56 ;
    RECT 31.37 95.85 31.58 95.92 ;
    RECT 31.83 95.13 32.04 95.2 ;
    RECT 31.83 95.49 32.04 95.56 ;
    RECT 31.83 95.85 32.04 95.92 ;
    RECT 67.89 95.13 68.1 95.2 ;
    RECT 67.89 95.49 68.1 95.56 ;
    RECT 67.89 95.85 68.1 95.92 ;
    RECT 68.35 95.13 68.56 95.2 ;
    RECT 68.35 95.49 68.56 95.56 ;
    RECT 68.35 95.85 68.56 95.92 ;
    RECT 28.05 95.13 28.26 95.2 ;
    RECT 28.05 95.49 28.26 95.56 ;
    RECT 28.05 95.85 28.26 95.92 ;
    RECT 28.51 95.13 28.72 95.2 ;
    RECT 28.51 95.49 28.72 95.56 ;
    RECT 28.51 95.85 28.72 95.92 ;
    RECT 24.73 95.13 24.94 95.2 ;
    RECT 24.73 95.49 24.94 95.56 ;
    RECT 24.73 95.85 24.94 95.92 ;
    RECT 25.19 95.13 25.4 95.2 ;
    RECT 25.19 95.49 25.4 95.56 ;
    RECT 25.19 95.85 25.4 95.92 ;
    RECT 21.41 95.13 21.62 95.2 ;
    RECT 21.41 95.49 21.62 95.56 ;
    RECT 21.41 95.85 21.62 95.92 ;
    RECT 21.87 95.13 22.08 95.2 ;
    RECT 21.87 95.49 22.08 95.56 ;
    RECT 21.87 95.85 22.08 95.92 ;
    RECT 18.09 95.13 18.3 95.2 ;
    RECT 18.09 95.49 18.3 95.56 ;
    RECT 18.09 95.85 18.3 95.92 ;
    RECT 18.55 95.13 18.76 95.2 ;
    RECT 18.55 95.49 18.76 95.56 ;
    RECT 18.55 95.85 18.76 95.92 ;
    RECT 120.825 95.49 120.895 95.56 ;
    RECT 14.77 95.13 14.98 95.2 ;
    RECT 14.77 95.49 14.98 95.56 ;
    RECT 14.77 95.85 14.98 95.92 ;
    RECT 15.23 95.13 15.44 95.2 ;
    RECT 15.23 95.49 15.44 95.56 ;
    RECT 15.23 95.85 15.44 95.92 ;
    RECT 11.45 95.13 11.66 95.2 ;
    RECT 11.45 95.49 11.66 95.56 ;
    RECT 11.45 95.85 11.66 95.92 ;
    RECT 11.91 95.13 12.12 95.2 ;
    RECT 11.91 95.49 12.12 95.56 ;
    RECT 11.91 95.85 12.12 95.92 ;
    RECT 8.13 95.13 8.34 95.2 ;
    RECT 8.13 95.49 8.34 95.56 ;
    RECT 8.13 95.85 8.34 95.92 ;
    RECT 8.59 95.13 8.8 95.2 ;
    RECT 8.59 95.49 8.8 95.56 ;
    RECT 8.59 95.85 8.8 95.92 ;
    RECT 4.81 95.13 5.02 95.2 ;
    RECT 4.81 95.49 5.02 95.56 ;
    RECT 4.81 95.85 5.02 95.92 ;
    RECT 5.27 95.13 5.48 95.2 ;
    RECT 5.27 95.49 5.48 95.56 ;
    RECT 5.27 95.85 5.48 95.92 ;
    RECT 1.49 95.13 1.7 95.2 ;
    RECT 1.49 95.49 1.7 95.56 ;
    RECT 1.49 95.85 1.7 95.92 ;
    RECT 1.95 95.13 2.16 95.2 ;
    RECT 1.95 95.49 2.16 95.56 ;
    RECT 1.95 95.85 2.16 95.92 ;
    RECT 64.57 95.13 64.78 95.2 ;
    RECT 64.57 95.49 64.78 95.56 ;
    RECT 64.57 95.85 64.78 95.92 ;
    RECT 65.03 95.13 65.24 95.2 ;
    RECT 65.03 95.49 65.24 95.56 ;
    RECT 65.03 95.85 65.24 95.92 ;
    RECT 61.25 94.41 61.46 94.48 ;
    RECT 61.25 94.77 61.46 94.84 ;
    RECT 61.25 95.13 61.46 95.2 ;
    RECT 61.71 94.41 61.92 94.48 ;
    RECT 61.71 94.77 61.92 94.84 ;
    RECT 61.71 95.13 61.92 95.2 ;
    RECT 57.93 94.41 58.14 94.48 ;
    RECT 57.93 94.77 58.14 94.84 ;
    RECT 57.93 95.13 58.14 95.2 ;
    RECT 58.39 94.41 58.6 94.48 ;
    RECT 58.39 94.77 58.6 94.84 ;
    RECT 58.39 95.13 58.6 95.2 ;
    RECT 54.61 94.41 54.82 94.48 ;
    RECT 54.61 94.77 54.82 94.84 ;
    RECT 54.61 95.13 54.82 95.2 ;
    RECT 55.07 94.41 55.28 94.48 ;
    RECT 55.07 94.77 55.28 94.84 ;
    RECT 55.07 95.13 55.28 95.2 ;
    RECT 51.29 94.41 51.5 94.48 ;
    RECT 51.29 94.77 51.5 94.84 ;
    RECT 51.29 95.13 51.5 95.2 ;
    RECT 51.75 94.41 51.96 94.48 ;
    RECT 51.75 94.77 51.96 94.84 ;
    RECT 51.75 95.13 51.96 95.2 ;
    RECT 47.97 94.41 48.18 94.48 ;
    RECT 47.97 94.77 48.18 94.84 ;
    RECT 47.97 95.13 48.18 95.2 ;
    RECT 48.43 94.41 48.64 94.48 ;
    RECT 48.43 94.77 48.64 94.84 ;
    RECT 48.43 95.13 48.64 95.2 ;
    RECT 44.65 94.41 44.86 94.48 ;
    RECT 44.65 94.77 44.86 94.84 ;
    RECT 44.65 95.13 44.86 95.2 ;
    RECT 45.11 94.41 45.32 94.48 ;
    RECT 45.11 94.77 45.32 94.84 ;
    RECT 45.11 95.13 45.32 95.2 ;
    RECT 41.33 94.41 41.54 94.48 ;
    RECT 41.33 94.77 41.54 94.84 ;
    RECT 41.33 95.13 41.54 95.2 ;
    RECT 41.79 94.41 42.0 94.48 ;
    RECT 41.79 94.77 42.0 94.84 ;
    RECT 41.79 95.13 42.0 95.2 ;
    RECT 38.01 94.41 38.22 94.48 ;
    RECT 38.01 94.77 38.22 94.84 ;
    RECT 38.01 95.13 38.22 95.2 ;
    RECT 38.47 94.41 38.68 94.48 ;
    RECT 38.47 94.77 38.68 94.84 ;
    RECT 38.47 95.13 38.68 95.2 ;
    RECT 0.4 94.77 0.47 94.84 ;
    RECT 34.69 94.41 34.9 94.48 ;
    RECT 34.69 94.77 34.9 94.84 ;
    RECT 34.69 95.13 34.9 95.2 ;
    RECT 35.15 94.41 35.36 94.48 ;
    RECT 35.15 94.77 35.36 94.84 ;
    RECT 35.15 95.13 35.36 95.2 ;
    RECT 117.69 94.41 117.9 94.48 ;
    RECT 117.69 94.77 117.9 94.84 ;
    RECT 117.69 95.13 117.9 95.2 ;
    RECT 118.15 94.41 118.36 94.48 ;
    RECT 118.15 94.77 118.36 94.84 ;
    RECT 118.15 95.13 118.36 95.2 ;
    RECT 114.37 94.41 114.58 94.48 ;
    RECT 114.37 94.77 114.58 94.84 ;
    RECT 114.37 95.13 114.58 95.2 ;
    RECT 114.83 94.41 115.04 94.48 ;
    RECT 114.83 94.77 115.04 94.84 ;
    RECT 114.83 95.13 115.04 95.2 ;
    RECT 111.05 94.41 111.26 94.48 ;
    RECT 111.05 94.77 111.26 94.84 ;
    RECT 111.05 95.13 111.26 95.2 ;
    RECT 111.51 94.41 111.72 94.48 ;
    RECT 111.51 94.77 111.72 94.84 ;
    RECT 111.51 95.13 111.72 95.2 ;
    RECT 107.73 94.41 107.94 94.48 ;
    RECT 107.73 94.77 107.94 94.84 ;
    RECT 107.73 95.13 107.94 95.2 ;
    RECT 108.19 94.41 108.4 94.48 ;
    RECT 108.19 94.77 108.4 94.84 ;
    RECT 108.19 95.13 108.4 95.2 ;
    RECT 104.41 94.41 104.62 94.48 ;
    RECT 104.41 94.77 104.62 94.84 ;
    RECT 104.41 95.13 104.62 95.2 ;
    RECT 104.87 94.41 105.08 94.48 ;
    RECT 104.87 94.77 105.08 94.84 ;
    RECT 104.87 95.13 105.08 95.2 ;
    RECT 101.09 94.41 101.3 94.48 ;
    RECT 101.09 94.77 101.3 94.84 ;
    RECT 101.09 95.13 101.3 95.2 ;
    RECT 101.55 94.41 101.76 94.48 ;
    RECT 101.55 94.77 101.76 94.84 ;
    RECT 101.55 95.13 101.76 95.2 ;
    RECT 97.77 94.41 97.98 94.48 ;
    RECT 97.77 94.77 97.98 94.84 ;
    RECT 97.77 95.13 97.98 95.2 ;
    RECT 98.23 94.41 98.44 94.48 ;
    RECT 98.23 94.77 98.44 94.84 ;
    RECT 98.23 95.13 98.44 95.2 ;
    RECT 94.45 94.41 94.66 94.48 ;
    RECT 94.45 94.77 94.66 94.84 ;
    RECT 94.45 95.13 94.66 95.2 ;
    RECT 94.91 94.41 95.12 94.48 ;
    RECT 94.91 94.77 95.12 94.84 ;
    RECT 94.91 95.13 95.12 95.2 ;
    RECT 91.13 94.41 91.34 94.48 ;
    RECT 91.13 94.77 91.34 94.84 ;
    RECT 91.13 95.13 91.34 95.2 ;
    RECT 91.59 94.41 91.8 94.48 ;
    RECT 91.59 94.77 91.8 94.84 ;
    RECT 91.59 95.13 91.8 95.2 ;
    RECT 87.81 94.41 88.02 94.48 ;
    RECT 87.81 94.77 88.02 94.84 ;
    RECT 87.81 95.13 88.02 95.2 ;
    RECT 88.27 94.41 88.48 94.48 ;
    RECT 88.27 94.77 88.48 94.84 ;
    RECT 88.27 95.13 88.48 95.2 ;
    RECT 84.49 94.41 84.7 94.48 ;
    RECT 84.49 94.77 84.7 94.84 ;
    RECT 84.49 95.13 84.7 95.2 ;
    RECT 84.95 94.41 85.16 94.48 ;
    RECT 84.95 94.77 85.16 94.84 ;
    RECT 84.95 95.13 85.16 95.2 ;
    RECT 81.17 94.41 81.38 94.48 ;
    RECT 81.17 94.77 81.38 94.84 ;
    RECT 81.17 95.13 81.38 95.2 ;
    RECT 81.63 94.41 81.84 94.48 ;
    RECT 81.63 94.77 81.84 94.84 ;
    RECT 81.63 95.13 81.84 95.2 ;
    RECT 77.85 94.41 78.06 94.48 ;
    RECT 77.85 94.77 78.06 94.84 ;
    RECT 77.85 95.13 78.06 95.2 ;
    RECT 78.31 94.41 78.52 94.48 ;
    RECT 78.31 94.77 78.52 94.84 ;
    RECT 78.31 95.13 78.52 95.2 ;
    RECT 74.53 94.41 74.74 94.48 ;
    RECT 74.53 94.77 74.74 94.84 ;
    RECT 74.53 95.13 74.74 95.2 ;
    RECT 74.99 94.41 75.2 94.48 ;
    RECT 74.99 94.77 75.2 94.84 ;
    RECT 74.99 95.13 75.2 95.2 ;
    RECT 71.21 94.41 71.42 94.48 ;
    RECT 71.21 94.77 71.42 94.84 ;
    RECT 71.21 95.13 71.42 95.2 ;
    RECT 71.67 94.41 71.88 94.48 ;
    RECT 71.67 94.77 71.88 94.84 ;
    RECT 71.67 95.13 71.88 95.2 ;
    RECT 31.37 94.41 31.58 94.48 ;
    RECT 31.37 94.77 31.58 94.84 ;
    RECT 31.37 95.13 31.58 95.2 ;
    RECT 31.83 94.41 32.04 94.48 ;
    RECT 31.83 94.77 32.04 94.84 ;
    RECT 31.83 95.13 32.04 95.2 ;
    RECT 67.89 94.41 68.1 94.48 ;
    RECT 67.89 94.77 68.1 94.84 ;
    RECT 67.89 95.13 68.1 95.2 ;
    RECT 68.35 94.41 68.56 94.48 ;
    RECT 68.35 94.77 68.56 94.84 ;
    RECT 68.35 95.13 68.56 95.2 ;
    RECT 28.05 94.41 28.26 94.48 ;
    RECT 28.05 94.77 28.26 94.84 ;
    RECT 28.05 95.13 28.26 95.2 ;
    RECT 28.51 94.41 28.72 94.48 ;
    RECT 28.51 94.77 28.72 94.84 ;
    RECT 28.51 95.13 28.72 95.2 ;
    RECT 24.73 94.41 24.94 94.48 ;
    RECT 24.73 94.77 24.94 94.84 ;
    RECT 24.73 95.13 24.94 95.2 ;
    RECT 25.19 94.41 25.4 94.48 ;
    RECT 25.19 94.77 25.4 94.84 ;
    RECT 25.19 95.13 25.4 95.2 ;
    RECT 21.41 94.41 21.62 94.48 ;
    RECT 21.41 94.77 21.62 94.84 ;
    RECT 21.41 95.13 21.62 95.2 ;
    RECT 21.87 94.41 22.08 94.48 ;
    RECT 21.87 94.77 22.08 94.84 ;
    RECT 21.87 95.13 22.08 95.2 ;
    RECT 18.09 94.41 18.3 94.48 ;
    RECT 18.09 94.77 18.3 94.84 ;
    RECT 18.09 95.13 18.3 95.2 ;
    RECT 18.55 94.41 18.76 94.48 ;
    RECT 18.55 94.77 18.76 94.84 ;
    RECT 18.55 95.13 18.76 95.2 ;
    RECT 120.825 94.77 120.895 94.84 ;
    RECT 14.77 94.41 14.98 94.48 ;
    RECT 14.77 94.77 14.98 94.84 ;
    RECT 14.77 95.13 14.98 95.2 ;
    RECT 15.23 94.41 15.44 94.48 ;
    RECT 15.23 94.77 15.44 94.84 ;
    RECT 15.23 95.13 15.44 95.2 ;
    RECT 11.45 94.41 11.66 94.48 ;
    RECT 11.45 94.77 11.66 94.84 ;
    RECT 11.45 95.13 11.66 95.2 ;
    RECT 11.91 94.41 12.12 94.48 ;
    RECT 11.91 94.77 12.12 94.84 ;
    RECT 11.91 95.13 12.12 95.2 ;
    RECT 8.13 94.41 8.34 94.48 ;
    RECT 8.13 94.77 8.34 94.84 ;
    RECT 8.13 95.13 8.34 95.2 ;
    RECT 8.59 94.41 8.8 94.48 ;
    RECT 8.59 94.77 8.8 94.84 ;
    RECT 8.59 95.13 8.8 95.2 ;
    RECT 4.81 94.41 5.02 94.48 ;
    RECT 4.81 94.77 5.02 94.84 ;
    RECT 4.81 95.13 5.02 95.2 ;
    RECT 5.27 94.41 5.48 94.48 ;
    RECT 5.27 94.77 5.48 94.84 ;
    RECT 5.27 95.13 5.48 95.2 ;
    RECT 1.49 94.41 1.7 94.48 ;
    RECT 1.49 94.77 1.7 94.84 ;
    RECT 1.49 95.13 1.7 95.2 ;
    RECT 1.95 94.41 2.16 94.48 ;
    RECT 1.95 94.77 2.16 94.84 ;
    RECT 1.95 95.13 2.16 95.2 ;
    RECT 64.57 94.41 64.78 94.48 ;
    RECT 64.57 94.77 64.78 94.84 ;
    RECT 64.57 95.13 64.78 95.2 ;
    RECT 65.03 94.41 65.24 94.48 ;
    RECT 65.03 94.77 65.24 94.84 ;
    RECT 65.03 95.13 65.24 95.2 ;
    RECT 61.25 56.95 61.46 57.02 ;
    RECT 61.25 57.31 61.46 57.38 ;
    RECT 61.25 57.67 61.46 57.74 ;
    RECT 61.71 56.95 61.92 57.02 ;
    RECT 61.71 57.31 61.92 57.38 ;
    RECT 61.71 57.67 61.92 57.74 ;
    RECT 57.93 56.95 58.14 57.02 ;
    RECT 57.93 57.31 58.14 57.38 ;
    RECT 57.93 57.67 58.14 57.74 ;
    RECT 58.39 56.95 58.6 57.02 ;
    RECT 58.39 57.31 58.6 57.38 ;
    RECT 58.39 57.67 58.6 57.74 ;
    RECT 54.61 56.95 54.82 57.02 ;
    RECT 54.61 57.31 54.82 57.38 ;
    RECT 54.61 57.67 54.82 57.74 ;
    RECT 55.07 56.95 55.28 57.02 ;
    RECT 55.07 57.31 55.28 57.38 ;
    RECT 55.07 57.67 55.28 57.74 ;
    RECT 51.29 56.95 51.5 57.02 ;
    RECT 51.29 57.31 51.5 57.38 ;
    RECT 51.29 57.67 51.5 57.74 ;
    RECT 51.75 56.95 51.96 57.02 ;
    RECT 51.75 57.31 51.96 57.38 ;
    RECT 51.75 57.67 51.96 57.74 ;
    RECT 47.97 56.95 48.18 57.02 ;
    RECT 47.97 57.31 48.18 57.38 ;
    RECT 47.97 57.67 48.18 57.74 ;
    RECT 48.43 56.95 48.64 57.02 ;
    RECT 48.43 57.31 48.64 57.38 ;
    RECT 48.43 57.67 48.64 57.74 ;
    RECT 44.65 56.95 44.86 57.02 ;
    RECT 44.65 57.31 44.86 57.38 ;
    RECT 44.65 57.67 44.86 57.74 ;
    RECT 45.11 56.95 45.32 57.02 ;
    RECT 45.11 57.31 45.32 57.38 ;
    RECT 45.11 57.67 45.32 57.74 ;
    RECT 41.33 56.95 41.54 57.02 ;
    RECT 41.33 57.31 41.54 57.38 ;
    RECT 41.33 57.67 41.54 57.74 ;
    RECT 41.79 56.95 42.0 57.02 ;
    RECT 41.79 57.31 42.0 57.38 ;
    RECT 41.79 57.67 42.0 57.74 ;
    RECT 38.01 56.95 38.22 57.02 ;
    RECT 38.01 57.31 38.22 57.38 ;
    RECT 38.01 57.67 38.22 57.74 ;
    RECT 38.47 56.95 38.68 57.02 ;
    RECT 38.47 57.31 38.68 57.38 ;
    RECT 38.47 57.67 38.68 57.74 ;
    RECT 0.4 57.31 0.47 57.38 ;
    RECT 34.69 56.95 34.9 57.02 ;
    RECT 34.69 57.31 34.9 57.38 ;
    RECT 34.69 57.67 34.9 57.74 ;
    RECT 35.15 56.95 35.36 57.02 ;
    RECT 35.15 57.31 35.36 57.38 ;
    RECT 35.15 57.67 35.36 57.74 ;
    RECT 117.69 56.95 117.9 57.02 ;
    RECT 117.69 57.31 117.9 57.38 ;
    RECT 117.69 57.67 117.9 57.74 ;
    RECT 118.15 56.95 118.36 57.02 ;
    RECT 118.15 57.31 118.36 57.38 ;
    RECT 118.15 57.67 118.36 57.74 ;
    RECT 114.37 56.95 114.58 57.02 ;
    RECT 114.37 57.31 114.58 57.38 ;
    RECT 114.37 57.67 114.58 57.74 ;
    RECT 114.83 56.95 115.04 57.02 ;
    RECT 114.83 57.31 115.04 57.38 ;
    RECT 114.83 57.67 115.04 57.74 ;
    RECT 111.05 56.95 111.26 57.02 ;
    RECT 111.05 57.31 111.26 57.38 ;
    RECT 111.05 57.67 111.26 57.74 ;
    RECT 111.51 56.95 111.72 57.02 ;
    RECT 111.51 57.31 111.72 57.38 ;
    RECT 111.51 57.67 111.72 57.74 ;
    RECT 107.73 56.95 107.94 57.02 ;
    RECT 107.73 57.31 107.94 57.38 ;
    RECT 107.73 57.67 107.94 57.74 ;
    RECT 108.19 56.95 108.4 57.02 ;
    RECT 108.19 57.31 108.4 57.38 ;
    RECT 108.19 57.67 108.4 57.74 ;
    RECT 104.41 56.95 104.62 57.02 ;
    RECT 104.41 57.31 104.62 57.38 ;
    RECT 104.41 57.67 104.62 57.74 ;
    RECT 104.87 56.95 105.08 57.02 ;
    RECT 104.87 57.31 105.08 57.38 ;
    RECT 104.87 57.67 105.08 57.74 ;
    RECT 101.09 56.95 101.3 57.02 ;
    RECT 101.09 57.31 101.3 57.38 ;
    RECT 101.09 57.67 101.3 57.74 ;
    RECT 101.55 56.95 101.76 57.02 ;
    RECT 101.55 57.31 101.76 57.38 ;
    RECT 101.55 57.67 101.76 57.74 ;
    RECT 97.77 56.95 97.98 57.02 ;
    RECT 97.77 57.31 97.98 57.38 ;
    RECT 97.77 57.67 97.98 57.74 ;
    RECT 98.23 56.95 98.44 57.02 ;
    RECT 98.23 57.31 98.44 57.38 ;
    RECT 98.23 57.67 98.44 57.74 ;
    RECT 94.45 56.95 94.66 57.02 ;
    RECT 94.45 57.31 94.66 57.38 ;
    RECT 94.45 57.67 94.66 57.74 ;
    RECT 94.91 56.95 95.12 57.02 ;
    RECT 94.91 57.31 95.12 57.38 ;
    RECT 94.91 57.67 95.12 57.74 ;
    RECT 91.13 56.95 91.34 57.02 ;
    RECT 91.13 57.31 91.34 57.38 ;
    RECT 91.13 57.67 91.34 57.74 ;
    RECT 91.59 56.95 91.8 57.02 ;
    RECT 91.59 57.31 91.8 57.38 ;
    RECT 91.59 57.67 91.8 57.74 ;
    RECT 87.81 56.95 88.02 57.02 ;
    RECT 87.81 57.31 88.02 57.38 ;
    RECT 87.81 57.67 88.02 57.74 ;
    RECT 88.27 56.95 88.48 57.02 ;
    RECT 88.27 57.31 88.48 57.38 ;
    RECT 88.27 57.67 88.48 57.74 ;
    RECT 84.49 56.95 84.7 57.02 ;
    RECT 84.49 57.31 84.7 57.38 ;
    RECT 84.49 57.67 84.7 57.74 ;
    RECT 84.95 56.95 85.16 57.02 ;
    RECT 84.95 57.31 85.16 57.38 ;
    RECT 84.95 57.67 85.16 57.74 ;
    RECT 81.17 56.95 81.38 57.02 ;
    RECT 81.17 57.31 81.38 57.38 ;
    RECT 81.17 57.67 81.38 57.74 ;
    RECT 81.63 56.95 81.84 57.02 ;
    RECT 81.63 57.31 81.84 57.38 ;
    RECT 81.63 57.67 81.84 57.74 ;
    RECT 77.85 56.95 78.06 57.02 ;
    RECT 77.85 57.31 78.06 57.38 ;
    RECT 77.85 57.67 78.06 57.74 ;
    RECT 78.31 56.95 78.52 57.02 ;
    RECT 78.31 57.31 78.52 57.38 ;
    RECT 78.31 57.67 78.52 57.74 ;
    RECT 74.53 56.95 74.74 57.02 ;
    RECT 74.53 57.31 74.74 57.38 ;
    RECT 74.53 57.67 74.74 57.74 ;
    RECT 74.99 56.95 75.2 57.02 ;
    RECT 74.99 57.31 75.2 57.38 ;
    RECT 74.99 57.67 75.2 57.74 ;
    RECT 71.21 56.95 71.42 57.02 ;
    RECT 71.21 57.31 71.42 57.38 ;
    RECT 71.21 57.67 71.42 57.74 ;
    RECT 71.67 56.95 71.88 57.02 ;
    RECT 71.67 57.31 71.88 57.38 ;
    RECT 71.67 57.67 71.88 57.74 ;
    RECT 31.37 56.95 31.58 57.02 ;
    RECT 31.37 57.31 31.58 57.38 ;
    RECT 31.37 57.67 31.58 57.74 ;
    RECT 31.83 56.95 32.04 57.02 ;
    RECT 31.83 57.31 32.04 57.38 ;
    RECT 31.83 57.67 32.04 57.74 ;
    RECT 67.89 56.95 68.1 57.02 ;
    RECT 67.89 57.31 68.1 57.38 ;
    RECT 67.89 57.67 68.1 57.74 ;
    RECT 68.35 56.95 68.56 57.02 ;
    RECT 68.35 57.31 68.56 57.38 ;
    RECT 68.35 57.67 68.56 57.74 ;
    RECT 28.05 56.95 28.26 57.02 ;
    RECT 28.05 57.31 28.26 57.38 ;
    RECT 28.05 57.67 28.26 57.74 ;
    RECT 28.51 56.95 28.72 57.02 ;
    RECT 28.51 57.31 28.72 57.38 ;
    RECT 28.51 57.67 28.72 57.74 ;
    RECT 24.73 56.95 24.94 57.02 ;
    RECT 24.73 57.31 24.94 57.38 ;
    RECT 24.73 57.67 24.94 57.74 ;
    RECT 25.19 56.95 25.4 57.02 ;
    RECT 25.19 57.31 25.4 57.38 ;
    RECT 25.19 57.67 25.4 57.74 ;
    RECT 21.41 56.95 21.62 57.02 ;
    RECT 21.41 57.31 21.62 57.38 ;
    RECT 21.41 57.67 21.62 57.74 ;
    RECT 21.87 56.95 22.08 57.02 ;
    RECT 21.87 57.31 22.08 57.38 ;
    RECT 21.87 57.67 22.08 57.74 ;
    RECT 18.09 56.95 18.3 57.02 ;
    RECT 18.09 57.31 18.3 57.38 ;
    RECT 18.09 57.67 18.3 57.74 ;
    RECT 18.55 56.95 18.76 57.02 ;
    RECT 18.55 57.31 18.76 57.38 ;
    RECT 18.55 57.67 18.76 57.74 ;
    RECT 120.825 57.31 120.895 57.38 ;
    RECT 14.77 56.95 14.98 57.02 ;
    RECT 14.77 57.31 14.98 57.38 ;
    RECT 14.77 57.67 14.98 57.74 ;
    RECT 15.23 56.95 15.44 57.02 ;
    RECT 15.23 57.31 15.44 57.38 ;
    RECT 15.23 57.67 15.44 57.74 ;
    RECT 11.45 56.95 11.66 57.02 ;
    RECT 11.45 57.31 11.66 57.38 ;
    RECT 11.45 57.67 11.66 57.74 ;
    RECT 11.91 56.95 12.12 57.02 ;
    RECT 11.91 57.31 12.12 57.38 ;
    RECT 11.91 57.67 12.12 57.74 ;
    RECT 8.13 56.95 8.34 57.02 ;
    RECT 8.13 57.31 8.34 57.38 ;
    RECT 8.13 57.67 8.34 57.74 ;
    RECT 8.59 56.95 8.8 57.02 ;
    RECT 8.59 57.31 8.8 57.38 ;
    RECT 8.59 57.67 8.8 57.74 ;
    RECT 4.81 56.95 5.02 57.02 ;
    RECT 4.81 57.31 5.02 57.38 ;
    RECT 4.81 57.67 5.02 57.74 ;
    RECT 5.27 56.95 5.48 57.02 ;
    RECT 5.27 57.31 5.48 57.38 ;
    RECT 5.27 57.67 5.48 57.74 ;
    RECT 1.49 56.95 1.7 57.02 ;
    RECT 1.49 57.31 1.7 57.38 ;
    RECT 1.49 57.67 1.7 57.74 ;
    RECT 1.95 56.95 2.16 57.02 ;
    RECT 1.95 57.31 2.16 57.38 ;
    RECT 1.95 57.67 2.16 57.74 ;
    RECT 64.57 56.95 64.78 57.02 ;
    RECT 64.57 57.31 64.78 57.38 ;
    RECT 64.57 57.67 64.78 57.74 ;
    RECT 65.03 56.95 65.24 57.02 ;
    RECT 65.03 57.31 65.24 57.38 ;
    RECT 65.03 57.67 65.24 57.74 ;
    RECT 61.25 54.07 61.46 54.14 ;
    RECT 61.25 54.43 61.46 54.5 ;
    RECT 61.25 54.79 61.46 54.86 ;
    RECT 61.71 54.07 61.92 54.14 ;
    RECT 61.71 54.43 61.92 54.5 ;
    RECT 61.71 54.79 61.92 54.86 ;
    RECT 57.93 54.07 58.14 54.14 ;
    RECT 57.93 54.43 58.14 54.5 ;
    RECT 57.93 54.79 58.14 54.86 ;
    RECT 58.39 54.07 58.6 54.14 ;
    RECT 58.39 54.43 58.6 54.5 ;
    RECT 58.39 54.79 58.6 54.86 ;
    RECT 54.61 54.07 54.82 54.14 ;
    RECT 54.61 54.43 54.82 54.5 ;
    RECT 54.61 54.79 54.82 54.86 ;
    RECT 55.07 54.07 55.28 54.14 ;
    RECT 55.07 54.43 55.28 54.5 ;
    RECT 55.07 54.79 55.28 54.86 ;
    RECT 51.29 54.07 51.5 54.14 ;
    RECT 51.29 54.43 51.5 54.5 ;
    RECT 51.29 54.79 51.5 54.86 ;
    RECT 51.75 54.07 51.96 54.14 ;
    RECT 51.75 54.43 51.96 54.5 ;
    RECT 51.75 54.79 51.96 54.86 ;
    RECT 47.97 54.07 48.18 54.14 ;
    RECT 47.97 54.43 48.18 54.5 ;
    RECT 47.97 54.79 48.18 54.86 ;
    RECT 48.43 54.07 48.64 54.14 ;
    RECT 48.43 54.43 48.64 54.5 ;
    RECT 48.43 54.79 48.64 54.86 ;
    RECT 44.65 54.07 44.86 54.14 ;
    RECT 44.65 54.43 44.86 54.5 ;
    RECT 44.65 54.79 44.86 54.86 ;
    RECT 45.11 54.07 45.32 54.14 ;
    RECT 45.11 54.43 45.32 54.5 ;
    RECT 45.11 54.79 45.32 54.86 ;
    RECT 41.33 54.07 41.54 54.14 ;
    RECT 41.33 54.43 41.54 54.5 ;
    RECT 41.33 54.79 41.54 54.86 ;
    RECT 41.79 54.07 42.0 54.14 ;
    RECT 41.79 54.43 42.0 54.5 ;
    RECT 41.79 54.79 42.0 54.86 ;
    RECT 38.01 54.07 38.22 54.14 ;
    RECT 38.01 54.43 38.22 54.5 ;
    RECT 38.01 54.79 38.22 54.86 ;
    RECT 38.47 54.07 38.68 54.14 ;
    RECT 38.47 54.43 38.68 54.5 ;
    RECT 38.47 54.79 38.68 54.86 ;
    RECT 0.4 54.43 0.47 54.5 ;
    RECT 34.69 54.07 34.9 54.14 ;
    RECT 34.69 54.43 34.9 54.5 ;
    RECT 34.69 54.79 34.9 54.86 ;
    RECT 35.15 54.07 35.36 54.14 ;
    RECT 35.15 54.43 35.36 54.5 ;
    RECT 35.15 54.79 35.36 54.86 ;
    RECT 117.69 54.07 117.9 54.14 ;
    RECT 117.69 54.43 117.9 54.5 ;
    RECT 117.69 54.79 117.9 54.86 ;
    RECT 118.15 54.07 118.36 54.14 ;
    RECT 118.15 54.43 118.36 54.5 ;
    RECT 118.15 54.79 118.36 54.86 ;
    RECT 114.37 54.07 114.58 54.14 ;
    RECT 114.37 54.43 114.58 54.5 ;
    RECT 114.37 54.79 114.58 54.86 ;
    RECT 114.83 54.07 115.04 54.14 ;
    RECT 114.83 54.43 115.04 54.5 ;
    RECT 114.83 54.79 115.04 54.86 ;
    RECT 111.05 54.07 111.26 54.14 ;
    RECT 111.05 54.43 111.26 54.5 ;
    RECT 111.05 54.79 111.26 54.86 ;
    RECT 111.51 54.07 111.72 54.14 ;
    RECT 111.51 54.43 111.72 54.5 ;
    RECT 111.51 54.79 111.72 54.86 ;
    RECT 107.73 54.07 107.94 54.14 ;
    RECT 107.73 54.43 107.94 54.5 ;
    RECT 107.73 54.79 107.94 54.86 ;
    RECT 108.19 54.07 108.4 54.14 ;
    RECT 108.19 54.43 108.4 54.5 ;
    RECT 108.19 54.79 108.4 54.86 ;
    RECT 104.41 54.07 104.62 54.14 ;
    RECT 104.41 54.43 104.62 54.5 ;
    RECT 104.41 54.79 104.62 54.86 ;
    RECT 104.87 54.07 105.08 54.14 ;
    RECT 104.87 54.43 105.08 54.5 ;
    RECT 104.87 54.79 105.08 54.86 ;
    RECT 101.09 54.07 101.3 54.14 ;
    RECT 101.09 54.43 101.3 54.5 ;
    RECT 101.09 54.79 101.3 54.86 ;
    RECT 101.55 54.07 101.76 54.14 ;
    RECT 101.55 54.43 101.76 54.5 ;
    RECT 101.55 54.79 101.76 54.86 ;
    RECT 97.77 54.07 97.98 54.14 ;
    RECT 97.77 54.43 97.98 54.5 ;
    RECT 97.77 54.79 97.98 54.86 ;
    RECT 98.23 54.07 98.44 54.14 ;
    RECT 98.23 54.43 98.44 54.5 ;
    RECT 98.23 54.79 98.44 54.86 ;
    RECT 94.45 54.07 94.66 54.14 ;
    RECT 94.45 54.43 94.66 54.5 ;
    RECT 94.45 54.79 94.66 54.86 ;
    RECT 94.91 54.07 95.12 54.14 ;
    RECT 94.91 54.43 95.12 54.5 ;
    RECT 94.91 54.79 95.12 54.86 ;
    RECT 91.13 54.07 91.34 54.14 ;
    RECT 91.13 54.43 91.34 54.5 ;
    RECT 91.13 54.79 91.34 54.86 ;
    RECT 91.59 54.07 91.8 54.14 ;
    RECT 91.59 54.43 91.8 54.5 ;
    RECT 91.59 54.79 91.8 54.86 ;
    RECT 87.81 54.07 88.02 54.14 ;
    RECT 87.81 54.43 88.02 54.5 ;
    RECT 87.81 54.79 88.02 54.86 ;
    RECT 88.27 54.07 88.48 54.14 ;
    RECT 88.27 54.43 88.48 54.5 ;
    RECT 88.27 54.79 88.48 54.86 ;
    RECT 84.49 54.07 84.7 54.14 ;
    RECT 84.49 54.43 84.7 54.5 ;
    RECT 84.49 54.79 84.7 54.86 ;
    RECT 84.95 54.07 85.16 54.14 ;
    RECT 84.95 54.43 85.16 54.5 ;
    RECT 84.95 54.79 85.16 54.86 ;
    RECT 81.17 54.07 81.38 54.14 ;
    RECT 81.17 54.43 81.38 54.5 ;
    RECT 81.17 54.79 81.38 54.86 ;
    RECT 81.63 54.07 81.84 54.14 ;
    RECT 81.63 54.43 81.84 54.5 ;
    RECT 81.63 54.79 81.84 54.86 ;
    RECT 77.85 54.07 78.06 54.14 ;
    RECT 77.85 54.43 78.06 54.5 ;
    RECT 77.85 54.79 78.06 54.86 ;
    RECT 78.31 54.07 78.52 54.14 ;
    RECT 78.31 54.43 78.52 54.5 ;
    RECT 78.31 54.79 78.52 54.86 ;
    RECT 74.53 54.07 74.74 54.14 ;
    RECT 74.53 54.43 74.74 54.5 ;
    RECT 74.53 54.79 74.74 54.86 ;
    RECT 74.99 54.07 75.2 54.14 ;
    RECT 74.99 54.43 75.2 54.5 ;
    RECT 74.99 54.79 75.2 54.86 ;
    RECT 71.21 54.07 71.42 54.14 ;
    RECT 71.21 54.43 71.42 54.5 ;
    RECT 71.21 54.79 71.42 54.86 ;
    RECT 71.67 54.07 71.88 54.14 ;
    RECT 71.67 54.43 71.88 54.5 ;
    RECT 71.67 54.79 71.88 54.86 ;
    RECT 31.37 54.07 31.58 54.14 ;
    RECT 31.37 54.43 31.58 54.5 ;
    RECT 31.37 54.79 31.58 54.86 ;
    RECT 31.83 54.07 32.04 54.14 ;
    RECT 31.83 54.43 32.04 54.5 ;
    RECT 31.83 54.79 32.04 54.86 ;
    RECT 67.89 54.07 68.1 54.14 ;
    RECT 67.89 54.43 68.1 54.5 ;
    RECT 67.89 54.79 68.1 54.86 ;
    RECT 68.35 54.07 68.56 54.14 ;
    RECT 68.35 54.43 68.56 54.5 ;
    RECT 68.35 54.79 68.56 54.86 ;
    RECT 28.05 54.07 28.26 54.14 ;
    RECT 28.05 54.43 28.26 54.5 ;
    RECT 28.05 54.79 28.26 54.86 ;
    RECT 28.51 54.07 28.72 54.14 ;
    RECT 28.51 54.43 28.72 54.5 ;
    RECT 28.51 54.79 28.72 54.86 ;
    RECT 24.73 54.07 24.94 54.14 ;
    RECT 24.73 54.43 24.94 54.5 ;
    RECT 24.73 54.79 24.94 54.86 ;
    RECT 25.19 54.07 25.4 54.14 ;
    RECT 25.19 54.43 25.4 54.5 ;
    RECT 25.19 54.79 25.4 54.86 ;
    RECT 21.41 54.07 21.62 54.14 ;
    RECT 21.41 54.43 21.62 54.5 ;
    RECT 21.41 54.79 21.62 54.86 ;
    RECT 21.87 54.07 22.08 54.14 ;
    RECT 21.87 54.43 22.08 54.5 ;
    RECT 21.87 54.79 22.08 54.86 ;
    RECT 18.09 54.07 18.3 54.14 ;
    RECT 18.09 54.43 18.3 54.5 ;
    RECT 18.09 54.79 18.3 54.86 ;
    RECT 18.55 54.07 18.76 54.14 ;
    RECT 18.55 54.43 18.76 54.5 ;
    RECT 18.55 54.79 18.76 54.86 ;
    RECT 120.825 54.43 120.895 54.5 ;
    RECT 14.77 54.07 14.98 54.14 ;
    RECT 14.77 54.43 14.98 54.5 ;
    RECT 14.77 54.79 14.98 54.86 ;
    RECT 15.23 54.07 15.44 54.14 ;
    RECT 15.23 54.43 15.44 54.5 ;
    RECT 15.23 54.79 15.44 54.86 ;
    RECT 11.45 54.07 11.66 54.14 ;
    RECT 11.45 54.43 11.66 54.5 ;
    RECT 11.45 54.79 11.66 54.86 ;
    RECT 11.91 54.07 12.12 54.14 ;
    RECT 11.91 54.43 12.12 54.5 ;
    RECT 11.91 54.79 12.12 54.86 ;
    RECT 8.13 54.07 8.34 54.14 ;
    RECT 8.13 54.43 8.34 54.5 ;
    RECT 8.13 54.79 8.34 54.86 ;
    RECT 8.59 54.07 8.8 54.14 ;
    RECT 8.59 54.43 8.8 54.5 ;
    RECT 8.59 54.79 8.8 54.86 ;
    RECT 4.81 54.07 5.02 54.14 ;
    RECT 4.81 54.43 5.02 54.5 ;
    RECT 4.81 54.79 5.02 54.86 ;
    RECT 5.27 54.07 5.48 54.14 ;
    RECT 5.27 54.43 5.48 54.5 ;
    RECT 5.27 54.79 5.48 54.86 ;
    RECT 1.49 54.07 1.7 54.14 ;
    RECT 1.49 54.43 1.7 54.5 ;
    RECT 1.49 54.79 1.7 54.86 ;
    RECT 1.95 54.07 2.16 54.14 ;
    RECT 1.95 54.43 2.16 54.5 ;
    RECT 1.95 54.79 2.16 54.86 ;
    RECT 64.57 54.07 64.78 54.14 ;
    RECT 64.57 54.43 64.78 54.5 ;
    RECT 64.57 54.79 64.78 54.86 ;
    RECT 65.03 54.07 65.24 54.14 ;
    RECT 65.03 54.43 65.24 54.5 ;
    RECT 65.03 54.79 65.24 54.86 ;
    RECT 61.25 53.35 61.46 53.42 ;
    RECT 61.25 53.71 61.46 53.78 ;
    RECT 61.25 54.07 61.46 54.14 ;
    RECT 61.71 53.35 61.92 53.42 ;
    RECT 61.71 53.71 61.92 53.78 ;
    RECT 61.71 54.07 61.92 54.14 ;
    RECT 57.93 53.35 58.14 53.42 ;
    RECT 57.93 53.71 58.14 53.78 ;
    RECT 57.93 54.07 58.14 54.14 ;
    RECT 58.39 53.35 58.6 53.42 ;
    RECT 58.39 53.71 58.6 53.78 ;
    RECT 58.39 54.07 58.6 54.14 ;
    RECT 54.61 53.35 54.82 53.42 ;
    RECT 54.61 53.71 54.82 53.78 ;
    RECT 54.61 54.07 54.82 54.14 ;
    RECT 55.07 53.35 55.28 53.42 ;
    RECT 55.07 53.71 55.28 53.78 ;
    RECT 55.07 54.07 55.28 54.14 ;
    RECT 51.29 53.35 51.5 53.42 ;
    RECT 51.29 53.71 51.5 53.78 ;
    RECT 51.29 54.07 51.5 54.14 ;
    RECT 51.75 53.35 51.96 53.42 ;
    RECT 51.75 53.71 51.96 53.78 ;
    RECT 51.75 54.07 51.96 54.14 ;
    RECT 47.97 53.35 48.18 53.42 ;
    RECT 47.97 53.71 48.18 53.78 ;
    RECT 47.97 54.07 48.18 54.14 ;
    RECT 48.43 53.35 48.64 53.42 ;
    RECT 48.43 53.71 48.64 53.78 ;
    RECT 48.43 54.07 48.64 54.14 ;
    RECT 44.65 53.35 44.86 53.42 ;
    RECT 44.65 53.71 44.86 53.78 ;
    RECT 44.65 54.07 44.86 54.14 ;
    RECT 45.11 53.35 45.32 53.42 ;
    RECT 45.11 53.71 45.32 53.78 ;
    RECT 45.11 54.07 45.32 54.14 ;
    RECT 41.33 53.35 41.54 53.42 ;
    RECT 41.33 53.71 41.54 53.78 ;
    RECT 41.33 54.07 41.54 54.14 ;
    RECT 41.79 53.35 42.0 53.42 ;
    RECT 41.79 53.71 42.0 53.78 ;
    RECT 41.79 54.07 42.0 54.14 ;
    RECT 38.01 53.35 38.22 53.42 ;
    RECT 38.01 53.71 38.22 53.78 ;
    RECT 38.01 54.07 38.22 54.14 ;
    RECT 38.47 53.35 38.68 53.42 ;
    RECT 38.47 53.71 38.68 53.78 ;
    RECT 38.47 54.07 38.68 54.14 ;
    RECT 0.4 53.71 0.47 53.78 ;
    RECT 34.69 53.35 34.9 53.42 ;
    RECT 34.69 53.71 34.9 53.78 ;
    RECT 34.69 54.07 34.9 54.14 ;
    RECT 35.15 53.35 35.36 53.42 ;
    RECT 35.15 53.71 35.36 53.78 ;
    RECT 35.15 54.07 35.36 54.14 ;
    RECT 117.69 53.35 117.9 53.42 ;
    RECT 117.69 53.71 117.9 53.78 ;
    RECT 117.69 54.07 117.9 54.14 ;
    RECT 118.15 53.35 118.36 53.42 ;
    RECT 118.15 53.71 118.36 53.78 ;
    RECT 118.15 54.07 118.36 54.14 ;
    RECT 114.37 53.35 114.58 53.42 ;
    RECT 114.37 53.71 114.58 53.78 ;
    RECT 114.37 54.07 114.58 54.14 ;
    RECT 114.83 53.35 115.04 53.42 ;
    RECT 114.83 53.71 115.04 53.78 ;
    RECT 114.83 54.07 115.04 54.14 ;
    RECT 111.05 53.35 111.26 53.42 ;
    RECT 111.05 53.71 111.26 53.78 ;
    RECT 111.05 54.07 111.26 54.14 ;
    RECT 111.51 53.35 111.72 53.42 ;
    RECT 111.51 53.71 111.72 53.78 ;
    RECT 111.51 54.07 111.72 54.14 ;
    RECT 107.73 53.35 107.94 53.42 ;
    RECT 107.73 53.71 107.94 53.78 ;
    RECT 107.73 54.07 107.94 54.14 ;
    RECT 108.19 53.35 108.4 53.42 ;
    RECT 108.19 53.71 108.4 53.78 ;
    RECT 108.19 54.07 108.4 54.14 ;
    RECT 104.41 53.35 104.62 53.42 ;
    RECT 104.41 53.71 104.62 53.78 ;
    RECT 104.41 54.07 104.62 54.14 ;
    RECT 104.87 53.35 105.08 53.42 ;
    RECT 104.87 53.71 105.08 53.78 ;
    RECT 104.87 54.07 105.08 54.14 ;
    RECT 101.09 53.35 101.3 53.42 ;
    RECT 101.09 53.71 101.3 53.78 ;
    RECT 101.09 54.07 101.3 54.14 ;
    RECT 101.55 53.35 101.76 53.42 ;
    RECT 101.55 53.71 101.76 53.78 ;
    RECT 101.55 54.07 101.76 54.14 ;
    RECT 97.77 53.35 97.98 53.42 ;
    RECT 97.77 53.71 97.98 53.78 ;
    RECT 97.77 54.07 97.98 54.14 ;
    RECT 98.23 53.35 98.44 53.42 ;
    RECT 98.23 53.71 98.44 53.78 ;
    RECT 98.23 54.07 98.44 54.14 ;
    RECT 94.45 53.35 94.66 53.42 ;
    RECT 94.45 53.71 94.66 53.78 ;
    RECT 94.45 54.07 94.66 54.14 ;
    RECT 94.91 53.35 95.12 53.42 ;
    RECT 94.91 53.71 95.12 53.78 ;
    RECT 94.91 54.07 95.12 54.14 ;
    RECT 91.13 53.35 91.34 53.42 ;
    RECT 91.13 53.71 91.34 53.78 ;
    RECT 91.13 54.07 91.34 54.14 ;
    RECT 91.59 53.35 91.8 53.42 ;
    RECT 91.59 53.71 91.8 53.78 ;
    RECT 91.59 54.07 91.8 54.14 ;
    RECT 87.81 53.35 88.02 53.42 ;
    RECT 87.81 53.71 88.02 53.78 ;
    RECT 87.81 54.07 88.02 54.14 ;
    RECT 88.27 53.35 88.48 53.42 ;
    RECT 88.27 53.71 88.48 53.78 ;
    RECT 88.27 54.07 88.48 54.14 ;
    RECT 84.49 53.35 84.7 53.42 ;
    RECT 84.49 53.71 84.7 53.78 ;
    RECT 84.49 54.07 84.7 54.14 ;
    RECT 84.95 53.35 85.16 53.42 ;
    RECT 84.95 53.71 85.16 53.78 ;
    RECT 84.95 54.07 85.16 54.14 ;
    RECT 81.17 53.35 81.38 53.42 ;
    RECT 81.17 53.71 81.38 53.78 ;
    RECT 81.17 54.07 81.38 54.14 ;
    RECT 81.63 53.35 81.84 53.42 ;
    RECT 81.63 53.71 81.84 53.78 ;
    RECT 81.63 54.07 81.84 54.14 ;
    RECT 77.85 53.35 78.06 53.42 ;
    RECT 77.85 53.71 78.06 53.78 ;
    RECT 77.85 54.07 78.06 54.14 ;
    RECT 78.31 53.35 78.52 53.42 ;
    RECT 78.31 53.71 78.52 53.78 ;
    RECT 78.31 54.07 78.52 54.14 ;
    RECT 74.53 53.35 74.74 53.42 ;
    RECT 74.53 53.71 74.74 53.78 ;
    RECT 74.53 54.07 74.74 54.14 ;
    RECT 74.99 53.35 75.2 53.42 ;
    RECT 74.99 53.71 75.2 53.78 ;
    RECT 74.99 54.07 75.2 54.14 ;
    RECT 71.21 53.35 71.42 53.42 ;
    RECT 71.21 53.71 71.42 53.78 ;
    RECT 71.21 54.07 71.42 54.14 ;
    RECT 71.67 53.35 71.88 53.42 ;
    RECT 71.67 53.71 71.88 53.78 ;
    RECT 71.67 54.07 71.88 54.14 ;
    RECT 31.37 53.35 31.58 53.42 ;
    RECT 31.37 53.71 31.58 53.78 ;
    RECT 31.37 54.07 31.58 54.14 ;
    RECT 31.83 53.35 32.04 53.42 ;
    RECT 31.83 53.71 32.04 53.78 ;
    RECT 31.83 54.07 32.04 54.14 ;
    RECT 67.89 53.35 68.1 53.42 ;
    RECT 67.89 53.71 68.1 53.78 ;
    RECT 67.89 54.07 68.1 54.14 ;
    RECT 68.35 53.35 68.56 53.42 ;
    RECT 68.35 53.71 68.56 53.78 ;
    RECT 68.35 54.07 68.56 54.14 ;
    RECT 28.05 53.35 28.26 53.42 ;
    RECT 28.05 53.71 28.26 53.78 ;
    RECT 28.05 54.07 28.26 54.14 ;
    RECT 28.51 53.35 28.72 53.42 ;
    RECT 28.51 53.71 28.72 53.78 ;
    RECT 28.51 54.07 28.72 54.14 ;
    RECT 24.73 53.35 24.94 53.42 ;
    RECT 24.73 53.71 24.94 53.78 ;
    RECT 24.73 54.07 24.94 54.14 ;
    RECT 25.19 53.35 25.4 53.42 ;
    RECT 25.19 53.71 25.4 53.78 ;
    RECT 25.19 54.07 25.4 54.14 ;
    RECT 21.41 53.35 21.62 53.42 ;
    RECT 21.41 53.71 21.62 53.78 ;
    RECT 21.41 54.07 21.62 54.14 ;
    RECT 21.87 53.35 22.08 53.42 ;
    RECT 21.87 53.71 22.08 53.78 ;
    RECT 21.87 54.07 22.08 54.14 ;
    RECT 18.09 53.35 18.3 53.42 ;
    RECT 18.09 53.71 18.3 53.78 ;
    RECT 18.09 54.07 18.3 54.14 ;
    RECT 18.55 53.35 18.76 53.42 ;
    RECT 18.55 53.71 18.76 53.78 ;
    RECT 18.55 54.07 18.76 54.14 ;
    RECT 120.825 53.71 120.895 53.78 ;
    RECT 14.77 53.35 14.98 53.42 ;
    RECT 14.77 53.71 14.98 53.78 ;
    RECT 14.77 54.07 14.98 54.14 ;
    RECT 15.23 53.35 15.44 53.42 ;
    RECT 15.23 53.71 15.44 53.78 ;
    RECT 15.23 54.07 15.44 54.14 ;
    RECT 11.45 53.35 11.66 53.42 ;
    RECT 11.45 53.71 11.66 53.78 ;
    RECT 11.45 54.07 11.66 54.14 ;
    RECT 11.91 53.35 12.12 53.42 ;
    RECT 11.91 53.71 12.12 53.78 ;
    RECT 11.91 54.07 12.12 54.14 ;
    RECT 8.13 53.35 8.34 53.42 ;
    RECT 8.13 53.71 8.34 53.78 ;
    RECT 8.13 54.07 8.34 54.14 ;
    RECT 8.59 53.35 8.8 53.42 ;
    RECT 8.59 53.71 8.8 53.78 ;
    RECT 8.59 54.07 8.8 54.14 ;
    RECT 4.81 53.35 5.02 53.42 ;
    RECT 4.81 53.71 5.02 53.78 ;
    RECT 4.81 54.07 5.02 54.14 ;
    RECT 5.27 53.35 5.48 53.42 ;
    RECT 5.27 53.71 5.48 53.78 ;
    RECT 5.27 54.07 5.48 54.14 ;
    RECT 1.49 53.35 1.7 53.42 ;
    RECT 1.49 53.71 1.7 53.78 ;
    RECT 1.49 54.07 1.7 54.14 ;
    RECT 1.95 53.35 2.16 53.42 ;
    RECT 1.95 53.71 2.16 53.78 ;
    RECT 1.95 54.07 2.16 54.14 ;
    RECT 64.57 53.35 64.78 53.42 ;
    RECT 64.57 53.71 64.78 53.78 ;
    RECT 64.57 54.07 64.78 54.14 ;
    RECT 65.03 53.35 65.24 53.42 ;
    RECT 65.03 53.71 65.24 53.78 ;
    RECT 65.03 54.07 65.24 54.14 ;
    RECT 121.44 49.75 121.51 50.54 ;
    RECT 122.04 49.75 122.25 49.82 ;
    RECT 122.04 50.105 122.25 50.175 ;
    RECT 122.04 50.47 122.25 50.54 ;
    RECT 123.205 50.195 124.005 50.265 ;
    RECT 125.67 50.02 125.905 50.09 ;
    RECT 126.73 50.02 126.99 50.09 ;
    RECT 128.705 50.02 128.935 50.09 ;
    RECT 129.42 50.02 129.68 50.09 ;
    RECT 130.59 50.02 130.66 50.09 ;
    RECT 133.925 50.02 134.135 50.09 ;
    RECT 134.31 50.02 134.58 50.09 ;
    RECT 138.365 50.02 138.435 50.09 ;
    RECT 138.695 50.02 138.96 50.09 ;
    RECT 140.45 50.02 140.71 50.09 ;
    RECT 140.895 50.02 140.965 50.09 ;
    RECT 141.385 50.02 141.645 50.09 ;
    RECT 142.51 50.02 142.72 50.09 ;
    RECT 144.32 50.195 145.135 50.265 ;
    RECT 146.125 49.75 146.395 49.82 ;
    RECT 146.125 50.105 146.395 50.175 ;
    RECT 146.125 50.47 146.395 50.54 ;
    RECT 121.44 49.03 121.51 49.82 ;
    RECT 122.04 49.03 122.25 49.1 ;
    RECT 122.04 49.385 122.25 49.455 ;
    RECT 122.04 49.75 122.25 49.82 ;
    RECT 123.205 49.475 124.005 49.545 ;
    RECT 125.67 49.3 125.905 49.37 ;
    RECT 126.73 49.3 126.99 49.37 ;
    RECT 128.705 49.3 128.935 49.37 ;
    RECT 129.42 49.3 129.68 49.37 ;
    RECT 130.59 49.3 130.66 49.37 ;
    RECT 133.925 49.3 134.135 49.37 ;
    RECT 134.31 49.3 134.58 49.37 ;
    RECT 138.365 49.3 138.435 49.37 ;
    RECT 138.695 49.3 138.96 49.37 ;
    RECT 140.45 49.3 140.71 49.37 ;
    RECT 140.895 49.3 140.965 49.37 ;
    RECT 141.385 49.3 141.645 49.37 ;
    RECT 142.51 49.3 142.72 49.37 ;
    RECT 144.32 49.475 145.135 49.545 ;
    RECT 146.125 49.03 146.395 49.1 ;
    RECT 146.125 49.385 146.395 49.455 ;
    RECT 146.125 49.75 146.395 49.82 ;
    RECT 121.44 48.31 121.51 49.1 ;
    RECT 122.04 48.31 122.25 48.38 ;
    RECT 122.04 48.665 122.25 48.735 ;
    RECT 122.04 49.03 122.25 49.1 ;
    RECT 123.205 48.755 124.005 48.825 ;
    RECT 125.67 48.58 125.905 48.65 ;
    RECT 126.73 48.58 126.99 48.65 ;
    RECT 128.705 48.58 128.935 48.65 ;
    RECT 129.42 48.58 129.68 48.65 ;
    RECT 130.59 48.58 130.66 48.65 ;
    RECT 133.925 48.58 134.135 48.65 ;
    RECT 134.31 48.58 134.58 48.65 ;
    RECT 138.365 48.58 138.435 48.65 ;
    RECT 138.695 48.58 138.96 48.65 ;
    RECT 140.45 48.58 140.71 48.65 ;
    RECT 140.895 48.58 140.965 48.65 ;
    RECT 141.385 48.58 141.645 48.65 ;
    RECT 142.51 48.58 142.72 48.65 ;
    RECT 144.32 48.755 145.135 48.825 ;
    RECT 146.125 48.31 146.395 48.38 ;
    RECT 146.125 48.665 146.395 48.735 ;
    RECT 146.125 49.03 146.395 49.1 ;
    RECT 121.44 47.59 121.51 48.38 ;
    RECT 122.04 47.59 122.25 47.66 ;
    RECT 122.04 47.945 122.25 48.015 ;
    RECT 122.04 48.31 122.25 48.38 ;
    RECT 123.205 48.035 124.005 48.105 ;
    RECT 125.67 47.86 125.905 47.93 ;
    RECT 126.73 47.86 126.99 47.93 ;
    RECT 128.705 47.86 128.935 47.93 ;
    RECT 129.42 47.86 129.68 47.93 ;
    RECT 130.59 47.86 130.66 47.93 ;
    RECT 133.925 47.86 134.135 47.93 ;
    RECT 134.31 47.86 134.58 47.93 ;
    RECT 138.365 47.86 138.435 47.93 ;
    RECT 138.695 47.86 138.96 47.93 ;
    RECT 140.45 47.86 140.71 47.93 ;
    RECT 140.895 47.86 140.965 47.93 ;
    RECT 141.385 47.86 141.645 47.93 ;
    RECT 142.51 47.86 142.72 47.93 ;
    RECT 144.32 48.035 145.135 48.105 ;
    RECT 146.125 47.59 146.395 47.66 ;
    RECT 146.125 47.945 146.395 48.015 ;
    RECT 146.125 48.31 146.395 48.38 ;
    RECT 121.44 46.87 121.51 47.66 ;
    RECT 122.04 46.87 122.25 46.94 ;
    RECT 122.04 47.225 122.25 47.295 ;
    RECT 122.04 47.59 122.25 47.66 ;
    RECT 123.205 47.315 124.005 47.385 ;
    RECT 125.67 47.14 125.905 47.21 ;
    RECT 126.73 47.14 126.99 47.21 ;
    RECT 128.705 47.14 128.935 47.21 ;
    RECT 129.42 47.14 129.68 47.21 ;
    RECT 130.59 47.14 130.66 47.21 ;
    RECT 133.925 47.14 134.135 47.21 ;
    RECT 134.31 47.14 134.58 47.21 ;
    RECT 138.365 47.14 138.435 47.21 ;
    RECT 138.695 47.14 138.96 47.21 ;
    RECT 140.45 47.14 140.71 47.21 ;
    RECT 140.895 47.14 140.965 47.21 ;
    RECT 141.385 47.14 141.645 47.21 ;
    RECT 142.51 47.14 142.72 47.21 ;
    RECT 144.32 47.315 145.135 47.385 ;
    RECT 146.125 46.87 146.395 46.94 ;
    RECT 146.125 47.225 146.395 47.295 ;
    RECT 146.125 47.59 146.395 47.66 ;
    RECT 135.305 65.877 135.375 65.947 ;
    RECT 121.44 46.15 121.51 46.94 ;
    RECT 122.04 46.15 122.25 46.22 ;
    RECT 122.04 46.505 122.25 46.575 ;
    RECT 122.04 46.87 122.25 46.94 ;
    RECT 123.205 46.595 124.005 46.665 ;
    RECT 125.67 46.42 125.905 46.49 ;
    RECT 126.73 46.42 126.99 46.49 ;
    RECT 128.705 46.42 128.935 46.49 ;
    RECT 129.42 46.42 129.68 46.49 ;
    RECT 130.59 46.42 130.66 46.49 ;
    RECT 133.925 46.42 134.135 46.49 ;
    RECT 134.31 46.42 134.58 46.49 ;
    RECT 138.365 46.42 138.435 46.49 ;
    RECT 138.695 46.42 138.96 46.49 ;
    RECT 140.45 46.42 140.71 46.49 ;
    RECT 140.895 46.42 140.965 46.49 ;
    RECT 141.385 46.42 141.645 46.49 ;
    RECT 142.51 46.42 142.72 46.49 ;
    RECT 144.32 46.595 145.135 46.665 ;
    RECT 146.125 46.15 146.395 46.22 ;
    RECT 146.125 46.505 146.395 46.575 ;
    RECT 146.125 46.87 146.395 46.94 ;
    RECT 121.44 45.43 121.51 46.22 ;
    RECT 122.04 45.43 122.25 45.5 ;
    RECT 122.04 45.785 122.25 45.855 ;
    RECT 122.04 46.15 122.25 46.22 ;
    RECT 123.205 45.875 124.005 45.945 ;
    RECT 125.67 45.7 125.905 45.77 ;
    RECT 126.73 45.7 126.99 45.77 ;
    RECT 128.705 45.7 128.935 45.77 ;
    RECT 129.42 45.7 129.68 45.77 ;
    RECT 130.59 45.7 130.66 45.77 ;
    RECT 133.925 45.7 134.135 45.77 ;
    RECT 134.31 45.7 134.58 45.77 ;
    RECT 138.365 45.7 138.435 45.77 ;
    RECT 138.695 45.7 138.96 45.77 ;
    RECT 140.45 45.7 140.71 45.77 ;
    RECT 140.895 45.7 140.965 45.77 ;
    RECT 141.385 45.7 141.645 45.77 ;
    RECT 142.51 45.7 142.72 45.77 ;
    RECT 144.32 45.875 145.135 45.945 ;
    RECT 146.125 45.43 146.395 45.5 ;
    RECT 146.125 45.785 146.395 45.855 ;
    RECT 146.125 46.15 146.395 46.22 ;
    RECT 121.44 44.71 121.51 45.5 ;
    RECT 122.04 44.71 122.25 44.78 ;
    RECT 122.04 45.065 122.25 45.135 ;
    RECT 122.04 45.43 122.25 45.5 ;
    RECT 123.205 45.155 124.005 45.225 ;
    RECT 125.67 44.98 125.905 45.05 ;
    RECT 126.73 44.98 126.99 45.05 ;
    RECT 128.705 44.98 128.935 45.05 ;
    RECT 129.42 44.98 129.68 45.05 ;
    RECT 130.59 44.98 130.66 45.05 ;
    RECT 133.925 44.98 134.135 45.05 ;
    RECT 134.31 44.98 134.58 45.05 ;
    RECT 138.365 44.98 138.435 45.05 ;
    RECT 138.695 44.98 138.96 45.05 ;
    RECT 140.45 44.98 140.71 45.05 ;
    RECT 140.895 44.98 140.965 45.05 ;
    RECT 141.385 44.98 141.645 45.05 ;
    RECT 142.51 44.98 142.72 45.05 ;
    RECT 144.32 45.155 145.135 45.225 ;
    RECT 146.125 44.71 146.395 44.78 ;
    RECT 146.125 45.065 146.395 45.135 ;
    RECT 146.125 45.43 146.395 45.5 ;
    RECT 135.5 93.237 135.57 93.307 ;
    RECT 127.69 37.057 127.9 37.127 ;
    RECT 127.69 32.022 127.9 32.092 ;
    RECT 135.105 50.737 135.175 50.807 ;
    RECT 122.63 82.53 122.84 82.6 ;
    RECT 133.19 66.597 133.26 66.667 ;
    RECT 145.485 67.41 145.695 67.48 ;
    RECT 139.73 67.32 139.94 67.39 ;
    RECT 132.79 93.957 132.86 94.027 ;
    RECT 127.69 67.317 127.9 67.387 ;
    RECT 132.595 51.457 132.665 51.527 ;
    RECT 133.19 40.657 133.26 40.727 ;
    RECT 127.69 21.937 127.9 22.007 ;
    RECT 145.485 92.61 145.695 92.68 ;
    RECT 145.485 70.29 145.695 70.36 ;
    RECT 132.99 44.977 133.06 45.047 ;
    RECT 127.69 21.217 127.9 21.287 ;
    RECT 127.69 17.602 127.9 17.672 ;
    RECT 139.73 92.52 139.94 92.59 ;
    RECT 127.69 16.887 127.9 16.957 ;
    RECT 139.73 70.2 139.94 70.27 ;
    RECT 127.69 92.517 127.9 92.587 ;
    RECT 122.63 37.15 122.84 37.22 ;
    RECT 127.69 70.197 127.9 70.267 ;
    RECT 122.63 92.61 122.84 92.68 ;
    RECT 142.51 99.182 142.72 99.252 ;
    RECT 135.105 58.657 135.175 58.727 ;
    RECT 145.485 77.49 145.695 77.56 ;
    RECT 122.63 70.29 122.84 70.36 ;
    RECT 125.67 99.182 125.88 99.252 ;
    RECT 122.63 36.43 122.84 36.5 ;
    RECT 122.63 35.71 122.84 35.78 ;
    RECT 139.73 77.4 139.94 77.47 ;
    RECT 145.485 54.43 145.695 54.5 ;
    RECT 122.63 34.99 122.84 35.06 ;
    RECT 122.63 34.27 122.84 34.34 ;
    RECT 127.69 77.397 127.9 77.467 ;
    RECT 139.73 54.34 139.94 54.41 ;
    RECT 145.485 84.69 145.695 84.76 ;
    RECT 122.63 77.49 122.84 77.56 ;
    RECT 127.69 54.337 127.9 54.407 ;
    RECT 135.5 87.477 135.57 87.547 ;
    RECT 122.63 33.55 122.84 33.62 ;
    RECT 135.305 73.077 135.375 73.147 ;
    RECT 139.73 84.6 139.94 84.67 ;
    RECT 145.485 62.37 145.695 62.44 ;
    RECT 122.63 32.83 122.84 32.9 ;
    RECT 122.63 54.43 122.84 54.5 ;
    RECT 133.19 88.197 133.26 88.267 ;
    RECT 139.73 62.28 139.94 62.35 ;
    RECT 127.69 84.597 127.9 84.667 ;
    RECT 127.69 62.277 127.9 62.347 ;
    RECT 122.63 84.69 122.84 84.76 ;
    RECT 132.595 73.797 132.665 73.867 ;
    RECT 122.63 32.11 122.84 32.18 ;
    RECT 145.485 39.31 145.695 39.38 ;
    RECT 145.485 69.57 145.695 69.64 ;
    RECT 122.63 31.39 122.84 31.46 ;
    RECT 139.73 39.22 139.94 39.29 ;
    RECT 122.63 62.37 122.84 62.44 ;
    RECT 139.73 69.48 139.94 69.55 ;
    RECT 122.63 30.67 122.84 30.74 ;
    RECT 127.69 39.217 127.9 39.287 ;
    RECT 127.69 69.477 127.9 69.547 ;
    RECT 135.5 95.397 135.57 95.467 ;
    RECT 122.63 39.31 122.84 39.38 ;
    RECT 122.63 69.57 122.84 69.64 ;
    RECT 133.19 42.817 133.26 42.887 ;
    RECT 132.99 67.317 133.06 67.387 ;
    RECT 140.895 60.812 140.965 60.882 ;
    RECT 139.73 61.177 139.94 61.247 ;
    RECT 145.485 72.45 145.695 72.52 ;
    RECT 135.305 80.997 135.375 81.067 ;
    RECT 136.92 61.177 137.13 61.247 ;
    RECT 139.73 72.36 139.94 72.43 ;
    RECT 145.485 97.65 145.695 97.72 ;
    RECT 139.73 97.56 139.94 97.63 ;
    RECT 134.34 61.177 134.55 61.247 ;
    RECT 130.595 60.812 130.665 60.882 ;
    RECT 135.5 88.917 135.57 88.987 ;
    RECT 127.69 97.557 127.9 97.627 ;
    RECT 135.105 39.217 135.175 39.287 ;
    RECT 132.395 52.177 132.465 52.247 ;
    RECT 127.69 72.357 127.9 72.427 ;
    RECT 145.485 79.65 145.695 79.72 ;
    RECT 126.76 61.177 126.97 61.247 ;
    RECT 122.63 72.45 122.84 72.52 ;
    RECT 125.11 61.177 125.32 61.247 ;
    RECT 139.73 79.56 139.94 79.63 ;
    RECT 124.255 61.177 124.465 61.247 ;
    RECT 122.63 97.65 122.84 97.72 ;
    RECT 121.44 61.05 121.51 61.12 ;
    RECT 145.485 56.59 145.695 56.66 ;
    RECT 139.73 56.5 139.94 56.57 ;
    RECT 135.105 46.417 135.175 46.487 ;
    RECT 135.305 74.517 135.375 74.587 ;
    RECT 127.69 79.557 127.9 79.627 ;
    RECT 122.63 79.65 122.84 79.72 ;
    RECT 127.69 56.497 127.9 56.567 ;
    RECT 145.485 64.53 145.695 64.6 ;
    RECT 135.105 59.377 135.175 59.447 ;
    RECT 122.63 56.59 122.84 56.66 ;
    RECT 139.73 64.44 139.94 64.51 ;
    RECT 132.79 47.137 132.86 47.207 ;
    RECT 132.595 75.237 132.665 75.307 ;
    RECT 131.995 60.097 132.065 60.167 ;
    RECT 127.69 86.757 127.9 86.827 ;
    RECT 127.69 64.437 127.9 64.507 ;
    RECT 122.63 86.85 122.84 86.92 ;
    RECT 122.63 64.53 122.84 64.6 ;
    RECT 145.485 48.67 145.695 48.74 ;
    RECT 135.105 54.337 135.175 54.407 ;
    RECT 133.19 88.917 133.26 88.987 ;
    RECT 139.73 48.58 139.94 48.65 ;
    RECT 127.69 48.577 127.9 48.647 ;
    RECT 122.63 48.67 122.84 48.74 ;
    RECT 135.5 96.117 135.57 96.187 ;
    RECT 135.105 53.617 135.175 53.687 ;
    RECT 145.485 58.75 145.695 58.82 ;
    RECT 139.73 58.66 139.94 58.73 ;
    RECT 135.305 81.717 135.375 81.787 ;
    RECT 132.595 96.837 132.665 96.907 ;
    RECT 135.105 41.377 135.175 41.447 ;
    RECT 132.395 54.337 132.465 54.407 ;
    RECT 131.995 82.437 132.065 82.507 ;
    RECT 127.69 58.657 127.9 58.727 ;
    RECT 145.485 66.69 145.695 66.76 ;
    RECT 122.63 58.75 122.84 58.82 ;
    RECT 139.73 66.6 139.94 66.67 ;
    RECT 135.305 76.677 135.375 76.747 ;
    RECT 127.69 66.597 127.9 66.667 ;
    RECT 122.63 66.69 122.84 66.76 ;
    RECT 135.305 62.277 135.375 62.347 ;
    RECT 145.485 50.83 145.695 50.9 ;
    RECT 139.73 50.74 139.94 50.81 ;
    RECT 132.395 77.397 132.465 77.467 ;
    RECT 133.39 62.997 133.46 63.067 ;
    RECT 145.485 80.37 145.695 80.44 ;
    RECT 139.73 80.28 139.94 80.35 ;
    RECT 127.69 50.737 127.9 50.807 ;
    RECT 122.63 50.83 122.84 50.9 ;
    RECT 135.105 47.137 135.175 47.207 ;
    RECT 135.105 56.497 135.175 56.567 ;
    RECT 145.485 87.57 145.695 87.64 ;
    RECT 139.73 87.48 139.94 87.55 ;
    RECT 132.79 47.857 132.86 47.927 ;
    RECT 127.69 87.477 127.9 87.547 ;
    RECT 142.51 60.992 142.72 61.062 ;
    RECT 122.63 87.57 122.84 87.64 ;
    RECT 145.485 42.19 145.695 42.26 ;
    RECT 139.73 42.1 139.94 42.17 ;
    RECT 121.44 43.99 121.51 44.78 ;
    RECT 122.04 43.99 122.25 44.06 ;
    RECT 122.04 44.345 122.25 44.415 ;
    RECT 122.04 44.71 122.25 44.78 ;
    RECT 123.205 44.435 124.005 44.505 ;
    RECT 125.67 44.26 125.905 44.33 ;
    RECT 126.73 44.26 126.99 44.33 ;
    RECT 128.705 44.26 128.935 44.33 ;
    RECT 129.42 44.26 129.68 44.33 ;
    RECT 130.59 44.26 130.66 44.33 ;
    RECT 133.925 44.26 134.135 44.33 ;
    RECT 134.31 44.26 134.58 44.33 ;
    RECT 138.365 44.26 138.435 44.33 ;
    RECT 138.695 44.26 138.96 44.33 ;
    RECT 140.45 44.26 140.71 44.33 ;
    RECT 140.895 44.26 140.965 44.33 ;
    RECT 141.385 44.26 141.645 44.33 ;
    RECT 142.51 44.26 142.72 44.33 ;
    RECT 144.32 44.435 145.135 44.505 ;
    RECT 146.125 43.99 146.395 44.06 ;
    RECT 146.125 44.345 146.395 44.415 ;
    RECT 146.125 44.71 146.395 44.78 ;
    RECT 121.44 43.27 121.51 44.06 ;
    RECT 122.04 43.27 122.25 43.34 ;
    RECT 122.04 43.625 122.25 43.695 ;
    RECT 122.04 43.99 122.25 44.06 ;
    RECT 123.205 43.715 124.005 43.785 ;
    RECT 125.67 43.54 125.905 43.61 ;
    RECT 126.73 43.54 126.99 43.61 ;
    RECT 128.705 43.54 128.935 43.61 ;
    RECT 129.42 43.54 129.68 43.61 ;
    RECT 130.59 43.54 130.66 43.61 ;
    RECT 133.925 43.54 134.135 43.61 ;
    RECT 134.31 43.54 134.58 43.61 ;
    RECT 138.365 43.54 138.435 43.61 ;
    RECT 138.695 43.54 138.96 43.61 ;
    RECT 140.45 43.54 140.71 43.61 ;
    RECT 140.895 43.54 140.965 43.61 ;
    RECT 141.385 43.54 141.645 43.61 ;
    RECT 142.51 43.54 142.72 43.61 ;
    RECT 144.32 43.715 145.135 43.785 ;
    RECT 146.125 43.27 146.395 43.34 ;
    RECT 146.125 43.625 146.395 43.695 ;
    RECT 146.125 43.99 146.395 44.06 ;
    RECT 121.44 42.55 121.51 43.34 ;
    RECT 122.04 42.55 122.25 42.62 ;
    RECT 122.04 42.905 122.25 42.975 ;
    RECT 122.04 43.27 122.25 43.34 ;
    RECT 123.205 42.995 124.005 43.065 ;
    RECT 125.67 42.82 125.905 42.89 ;
    RECT 126.73 42.82 126.99 42.89 ;
    RECT 128.705 42.82 128.935 42.89 ;
    RECT 129.42 42.82 129.68 42.89 ;
    RECT 130.59 42.82 130.66 42.89 ;
    RECT 133.925 42.82 134.135 42.89 ;
    RECT 134.31 42.82 134.58 42.89 ;
    RECT 138.365 42.82 138.435 42.89 ;
    RECT 138.695 42.82 138.96 42.89 ;
    RECT 140.45 42.82 140.71 42.89 ;
    RECT 140.895 42.82 140.965 42.89 ;
    RECT 141.385 42.82 141.645 42.89 ;
    RECT 142.51 42.82 142.72 42.89 ;
    RECT 144.32 42.995 145.135 43.065 ;
    RECT 146.125 42.55 146.395 42.62 ;
    RECT 146.125 42.905 146.395 42.975 ;
    RECT 146.125 43.27 146.395 43.34 ;
    RECT 121.44 41.83 121.51 42.62 ;
    RECT 122.04 41.83 122.25 41.9 ;
    RECT 122.04 42.185 122.25 42.255 ;
    RECT 122.04 42.55 122.25 42.62 ;
    RECT 123.205 42.275 124.005 42.345 ;
    RECT 125.67 42.1 125.905 42.17 ;
    RECT 126.73 42.1 126.99 42.17 ;
    RECT 128.705 42.1 128.935 42.17 ;
    RECT 129.42 42.1 129.68 42.17 ;
    RECT 130.59 42.1 130.66 42.17 ;
    RECT 133.925 42.1 134.135 42.17 ;
    RECT 134.31 42.1 134.58 42.17 ;
    RECT 138.365 42.1 138.435 42.17 ;
    RECT 138.695 42.1 138.96 42.17 ;
    RECT 140.45 42.1 140.71 42.17 ;
    RECT 140.895 42.1 140.965 42.17 ;
    RECT 141.385 42.1 141.645 42.17 ;
    RECT 142.51 42.1 142.72 42.17 ;
    RECT 144.32 42.275 145.135 42.345 ;
    RECT 146.125 41.83 146.395 41.9 ;
    RECT 146.125 42.185 146.395 42.255 ;
    RECT 146.125 42.55 146.395 42.62 ;
    RECT 121.44 41.11 121.51 41.9 ;
    RECT 122.04 41.11 122.25 41.18 ;
    RECT 122.04 41.465 122.25 41.535 ;
    RECT 122.04 41.83 122.25 41.9 ;
    RECT 123.205 41.555 124.005 41.625 ;
    RECT 125.67 41.38 125.905 41.45 ;
    RECT 126.73 41.38 126.99 41.45 ;
    RECT 128.705 41.38 128.935 41.45 ;
    RECT 129.42 41.38 129.68 41.45 ;
    RECT 130.59 41.38 130.66 41.45 ;
    RECT 133.925 41.38 134.135 41.45 ;
    RECT 134.31 41.38 134.58 41.45 ;
    RECT 138.365 41.38 138.435 41.45 ;
    RECT 138.695 41.38 138.96 41.45 ;
    RECT 140.45 41.38 140.71 41.45 ;
    RECT 140.895 41.38 140.965 41.45 ;
    RECT 141.385 41.38 141.645 41.45 ;
    RECT 142.51 41.38 142.72 41.45 ;
    RECT 144.32 41.555 145.135 41.625 ;
    RECT 146.125 41.11 146.395 41.18 ;
    RECT 146.125 41.465 146.395 41.535 ;
    RECT 146.125 41.83 146.395 41.9 ;
    RECT 121.44 40.39 121.51 41.18 ;
    RECT 122.04 40.39 122.25 40.46 ;
    RECT 122.04 40.745 122.25 40.815 ;
    RECT 122.04 41.11 122.25 41.18 ;
    RECT 123.205 40.835 124.005 40.905 ;
    RECT 125.67 40.66 125.905 40.73 ;
    RECT 126.73 40.66 126.99 40.73 ;
    RECT 128.705 40.66 128.935 40.73 ;
    RECT 129.42 40.66 129.68 40.73 ;
    RECT 130.59 40.66 130.66 40.73 ;
    RECT 133.925 40.66 134.135 40.73 ;
    RECT 134.31 40.66 134.58 40.73 ;
    RECT 138.365 40.66 138.435 40.73 ;
    RECT 138.695 40.66 138.96 40.73 ;
    RECT 140.45 40.66 140.71 40.73 ;
    RECT 140.895 40.66 140.965 40.73 ;
    RECT 141.385 40.66 141.645 40.73 ;
    RECT 142.51 40.66 142.72 40.73 ;
    RECT 144.32 40.835 145.135 40.905 ;
    RECT 146.125 40.39 146.395 40.46 ;
    RECT 146.125 40.745 146.395 40.815 ;
    RECT 146.125 41.11 146.395 41.18 ;
    RECT 121.44 39.67 121.51 40.46 ;
    RECT 122.04 39.67 122.25 39.74 ;
    RECT 122.04 40.025 122.25 40.095 ;
    RECT 122.04 40.39 122.25 40.46 ;
    RECT 123.205 40.115 124.005 40.185 ;
    RECT 125.67 39.94 125.905 40.01 ;
    RECT 126.73 39.94 126.99 40.01 ;
    RECT 128.705 39.94 128.935 40.01 ;
    RECT 129.42 39.94 129.68 40.01 ;
    RECT 130.59 39.94 130.66 40.01 ;
    RECT 133.925 39.94 134.135 40.01 ;
    RECT 134.31 39.94 134.58 40.01 ;
    RECT 138.365 39.94 138.435 40.01 ;
    RECT 138.695 39.94 138.96 40.01 ;
    RECT 140.45 39.94 140.71 40.01 ;
    RECT 140.895 39.94 140.965 40.01 ;
    RECT 141.385 39.94 141.645 40.01 ;
    RECT 142.51 39.94 142.72 40.01 ;
    RECT 144.32 40.115 145.135 40.185 ;
    RECT 146.125 39.67 146.395 39.74 ;
    RECT 146.125 40.025 146.395 40.095 ;
    RECT 146.125 40.39 146.395 40.46 ;
    RECT 121.44 38.95 121.51 39.74 ;
    RECT 122.04 38.95 122.25 39.02 ;
    RECT 122.04 39.305 122.25 39.375 ;
    RECT 122.04 39.67 122.25 39.74 ;
    RECT 123.205 39.395 124.005 39.465 ;
    RECT 125.67 39.22 125.905 39.29 ;
    RECT 126.73 39.22 126.99 39.29 ;
    RECT 128.705 39.22 128.935 39.29 ;
    RECT 129.42 39.22 129.68 39.29 ;
    RECT 130.59 39.22 130.66 39.29 ;
    RECT 133.925 39.22 134.135 39.29 ;
    RECT 134.31 39.22 134.58 39.29 ;
    RECT 138.365 39.22 138.435 39.29 ;
    RECT 138.695 39.22 138.96 39.29 ;
    RECT 140.45 39.22 140.71 39.29 ;
    RECT 140.895 39.22 140.965 39.29 ;
    RECT 141.385 39.22 141.645 39.29 ;
    RECT 142.51 39.22 142.72 39.29 ;
    RECT 144.32 39.395 145.135 39.465 ;
    RECT 146.125 38.95 146.395 39.02 ;
    RECT 146.125 39.305 146.395 39.375 ;
    RECT 146.125 39.67 146.395 39.74 ;
    RECT 121.44 38.23 121.51 39.02 ;
    RECT 122.04 38.23 122.25 38.3 ;
    RECT 122.04 38.585 122.25 38.655 ;
    RECT 122.04 38.95 122.25 39.02 ;
    RECT 123.205 38.675 124.005 38.745 ;
    RECT 125.67 38.5 125.905 38.57 ;
    RECT 126.73 38.5 126.99 38.57 ;
    RECT 128.705 38.5 128.935 38.57 ;
    RECT 129.42 38.5 129.68 38.57 ;
    RECT 130.59 38.5 130.66 38.57 ;
    RECT 133.925 38.5 134.135 38.57 ;
    RECT 134.31 38.5 134.58 38.57 ;
    RECT 138.365 38.5 138.435 38.57 ;
    RECT 138.695 38.5 138.96 38.57 ;
    RECT 140.45 38.5 140.71 38.57 ;
    RECT 140.895 38.5 140.965 38.57 ;
    RECT 141.385 38.5 141.645 38.57 ;
    RECT 142.51 38.5 142.72 38.57 ;
    RECT 144.32 38.675 145.135 38.745 ;
    RECT 146.125 38.23 146.395 38.3 ;
    RECT 146.125 38.585 146.395 38.655 ;
    RECT 146.125 38.95 146.395 39.02 ;
    RECT 121.44 37.51 121.51 38.3 ;
    RECT 122.04 37.51 122.25 37.58 ;
    RECT 122.04 37.865 122.25 37.935 ;
    RECT 122.04 38.23 122.25 38.3 ;
    RECT 123.205 37.955 124.005 38.025 ;
    RECT 125.67 37.78 125.905 37.85 ;
    RECT 126.73 37.78 126.99 37.85 ;
    RECT 128.705 37.78 128.935 37.85 ;
    RECT 129.42 37.78 129.68 37.85 ;
    RECT 130.59 37.78 130.66 37.85 ;
    RECT 133.925 37.78 134.135 37.85 ;
    RECT 134.31 37.78 134.58 37.85 ;
    RECT 138.365 37.78 138.435 37.85 ;
    RECT 138.695 37.78 138.96 37.85 ;
    RECT 140.45 37.78 140.71 37.85 ;
    RECT 140.895 37.78 140.965 37.85 ;
    RECT 141.385 37.78 141.645 37.85 ;
    RECT 142.51 37.78 142.72 37.85 ;
    RECT 144.32 37.955 145.135 38.025 ;
    RECT 146.125 37.51 146.395 37.58 ;
    RECT 146.125 37.865 146.395 37.935 ;
    RECT 146.125 38.23 146.395 38.3 ;
    RECT 125.67 60.992 125.88 61.062 ;
    RECT 145.485 52.27 145.695 52.34 ;
    RECT 139.73 52.18 139.94 52.25 ;
    RECT 127.69 52.177 127.9 52.247 ;
    RECT 145.485 93.33 145.695 93.4 ;
    RECT 127.69 42.097 127.9 42.167 ;
    RECT 139.73 93.24 139.94 93.31 ;
    RECT 122.63 42.19 122.84 42.26 ;
    RECT 135.5 98.277 135.57 98.347 ;
    RECT 145.485 59.47 145.695 59.54 ;
    RECT 123.235 60.627 123.445 60.697 ;
    RECT 122.63 52.27 122.84 52.34 ;
    RECT 139.73 59.38 139.94 59.45 ;
    RECT 121.44 14.47 121.51 37.58 ;
    RECT 122.04 14.47 122.25 14.895 ;
    RECT 122.04 15.19 122.25 15.26 ;
    RECT 122.04 15.55 122.25 15.62 ;
    RECT 122.04 15.91 122.25 15.98 ;
    RECT 122.04 16.27 122.25 16.34 ;
    RECT 122.04 16.63 122.25 16.7 ;
    RECT 122.04 16.99 122.25 17.06 ;
    RECT 122.04 17.35 122.25 17.42 ;
    RECT 122.04 17.71 122.25 17.78 ;
    RECT 122.04 18.07 122.25 18.14 ;
    RECT 122.04 18.43 122.25 18.5 ;
    RECT 122.04 18.79 122.25 18.86 ;
    RECT 122.04 19.15 122.25 19.22 ;
    RECT 122.04 19.51 122.25 19.58 ;
    RECT 122.04 19.87 122.25 19.94 ;
    RECT 122.04 20.23 122.25 20.3 ;
    RECT 122.04 20.59 122.25 20.66 ;
    RECT 122.04 20.95 122.25 21.02 ;
    RECT 122.04 21.31 122.25 21.38 ;
    RECT 122.04 21.67 122.25 21.74 ;
    RECT 122.04 22.03 122.25 22.1 ;
    RECT 122.04 22.39 122.25 22.46 ;
    RECT 122.04 22.75 122.25 22.82 ;
    RECT 122.04 23.11 122.25 23.18 ;
    RECT 122.04 23.47 122.25 23.54 ;
    RECT 122.04 23.83 122.25 23.9 ;
    RECT 122.04 24.19 122.25 24.26 ;
    RECT 122.04 24.55 122.25 24.62 ;
    RECT 122.04 24.91 122.25 24.98 ;
    RECT 122.04 25.27 122.25 25.34 ;
    RECT 122.04 25.63 122.25 25.7 ;
    RECT 122.04 25.99 122.25 26.06 ;
    RECT 122.04 26.35 122.25 26.42 ;
    RECT 122.04 26.71 122.25 26.78 ;
    RECT 122.04 27.07 122.25 27.14 ;
    RECT 122.04 27.43 122.25 27.5 ;
    RECT 122.04 27.79 122.25 27.86 ;
    RECT 122.04 28.15 122.25 28.22 ;
    RECT 122.04 28.51 122.25 28.58 ;
    RECT 122.04 28.87 122.25 28.94 ;
    RECT 122.04 29.23 122.25 29.3 ;
    RECT 122.04 29.59 122.25 29.66 ;
    RECT 122.04 29.95 122.25 30.02 ;
    RECT 122.04 30.31 122.25 30.38 ;
    RECT 122.04 30.67 122.25 30.74 ;
    RECT 122.04 31.03 122.25 31.1 ;
    RECT 122.04 31.39 122.25 31.46 ;
    RECT 122.04 31.75 122.25 31.82 ;
    RECT 122.04 32.11 122.25 32.18 ;
    RECT 122.04 32.47 122.25 32.54 ;
    RECT 122.04 32.83 122.25 32.9 ;
    RECT 122.04 33.19 122.25 33.26 ;
    RECT 122.04 33.55 122.25 33.62 ;
    RECT 122.04 33.91 122.25 33.98 ;
    RECT 122.04 34.27 122.25 34.34 ;
    RECT 122.04 34.63 122.25 34.7 ;
    RECT 122.04 34.99 122.25 35.06 ;
    RECT 122.04 35.35 122.25 35.42 ;
    RECT 122.04 35.71 122.25 35.78 ;
    RECT 122.04 36.07 122.25 36.14 ;
    RECT 122.04 36.43 122.25 36.5 ;
    RECT 122.04 36.79 122.25 36.86 ;
    RECT 122.04 37.15 122.25 37.22 ;
    RECT 122.04 37.51 122.25 37.58 ;
    RECT 123.235 14.915 123.975 14.985 ;
    RECT 123.235 15.635 123.975 15.705 ;
    RECT 123.235 16.35 123.975 16.42 ;
    RECT 123.235 17.075 123.975 17.145 ;
    RECT 123.235 17.795 123.975 17.865 ;
    RECT 123.235 18.515 123.975 18.585 ;
    RECT 123.235 19.23 123.975 19.3 ;
    RECT 123.235 19.955 123.975 20.025 ;
    RECT 123.235 20.675 123.975 20.745 ;
    RECT 123.235 21.39 123.975 21.46 ;
    RECT 123.235 22.115 123.975 22.185 ;
    RECT 123.235 22.835 123.975 22.905 ;
    RECT 123.235 23.555 123.975 23.625 ;
    RECT 123.235 24.275 123.975 24.345 ;
    RECT 123.235 24.995 123.975 25.065 ;
    RECT 123.235 25.715 123.975 25.785 ;
    RECT 123.235 26.435 123.975 26.505 ;
    RECT 123.235 27.155 123.975 27.225 ;
    RECT 123.235 27.875 123.975 27.945 ;
    RECT 123.235 28.595 123.975 28.665 ;
    RECT 123.235 29.315 123.975 29.385 ;
    RECT 123.235 30.035 123.975 30.105 ;
    RECT 123.235 30.75 123.975 30.82 ;
    RECT 123.235 31.47 123.975 31.54 ;
    RECT 123.235 32.195 123.975 32.265 ;
    RECT 123.235 32.915 123.975 32.985 ;
    RECT 123.235 33.635 123.975 33.705 ;
    RECT 123.235 34.355 123.975 34.425 ;
    RECT 123.235 35.075 123.975 35.145 ;
    RECT 123.235 35.79 123.975 35.86 ;
    RECT 123.235 36.51 123.975 36.58 ;
    RECT 123.235 37.235 123.975 37.305 ;
    RECT 125.68 37.055 125.89 37.125 ;
    RECT 125.695 14.74 125.905 14.81 ;
    RECT 125.695 15.455 125.905 15.525 ;
    RECT 125.695 16.17 125.905 16.24 ;
    RECT 125.695 16.885 125.905 16.955 ;
    RECT 125.695 17.6 125.905 17.67 ;
    RECT 125.695 18.34 125.905 18.41 ;
    RECT 125.695 19.055 125.905 19.125 ;
    RECT 125.695 19.775 125.905 19.845 ;
    RECT 125.695 20.495 125.905 20.565 ;
    RECT 125.695 21.215 125.905 21.285 ;
    RECT 125.695 21.935 125.905 22.005 ;
    RECT 125.695 22.655 125.905 22.725 ;
    RECT 125.695 25.535 125.905 25.605 ;
    RECT 125.695 26.255 125.905 26.325 ;
    RECT 125.695 27.695 125.905 27.765 ;
    RECT 125.695 29.14 125.905 29.21 ;
    RECT 125.695 29.86 125.905 29.93 ;
    RECT 125.695 30.58 125.905 30.65 ;
    RECT 125.695 31.295 125.905 31.365 ;
    RECT 125.695 32.015 125.905 32.085 ;
    RECT 125.695 32.735 125.905 32.805 ;
    RECT 125.695 33.455 125.905 33.525 ;
    RECT 125.695 34.18 125.905 34.25 ;
    RECT 125.695 34.9 125.905 34.97 ;
    RECT 125.695 35.62 125.905 35.69 ;
    RECT 125.695 36.335 125.905 36.405 ;
    RECT 126.73 14.74 126.99 14.81 ;
    RECT 126.73 15.455 126.99 15.525 ;
    RECT 126.73 16.17 126.99 16.24 ;
    RECT 126.73 18.34 126.99 18.41 ;
    RECT 126.73 19.055 126.99 19.125 ;
    RECT 126.73 19.775 126.99 19.845 ;
    RECT 126.73 20.495 126.99 20.565 ;
    RECT 126.73 22.655 126.99 22.725 ;
    RECT 126.73 26.255 126.99 26.325 ;
    RECT 126.73 29.14 126.99 29.21 ;
    RECT 126.73 29.86 126.99 29.93 ;
    RECT 126.73 30.58 126.99 30.65 ;
    RECT 126.73 32.735 126.99 32.805 ;
    RECT 126.73 33.455 126.99 33.525 ;
    RECT 126.73 34.18 126.99 34.25 ;
    RECT 126.73 34.9 126.99 34.97 ;
    RECT 126.73 35.62 126.99 35.69 ;
    RECT 126.73 36.335 126.99 36.405 ;
    RECT 126.76 16.89 126.97 16.96 ;
    RECT 126.76 17.605 126.97 17.675 ;
    RECT 126.76 21.22 126.97 21.29 ;
    RECT 126.76 21.935 126.97 22.005 ;
    RECT 126.76 32.025 126.97 32.095 ;
    RECT 126.76 37.06 126.97 37.13 ;
    RECT 127.67 14.74 127.92 14.81 ;
    RECT 127.67 15.455 127.92 15.525 ;
    RECT 127.67 16.17 127.92 16.24 ;
    RECT 127.67 19.055 127.92 19.125 ;
    RECT 127.67 19.775 127.92 19.845 ;
    RECT 127.67 20.495 127.92 20.565 ;
    RECT 127.67 22.655 127.92 22.725 ;
    RECT 127.67 23.375 127.92 23.445 ;
    RECT 127.67 24.82 127.92 24.89 ;
    RECT 127.67 32.735 127.89 32.805 ;
    RECT 127.675 26.255 127.92 26.325 ;
    RECT 127.675 30.58 127.895 30.65 ;
    RECT 127.68 33.455 127.9 33.525 ;
    RECT 127.68 34.18 127.9 34.25 ;
    RECT 127.68 34.9 127.9 34.97 ;
    RECT 127.685 28.415 127.92 28.485 ;
    RECT 127.685 36.335 127.92 36.405 ;
    RECT 127.69 26.97 127.9 27.04 ;
    RECT 127.69 29.13 127.9 29.2 ;
    RECT 127.69 29.85 127.9 29.92 ;
    RECT 127.69 35.62 127.91 35.69 ;
    RECT 128.125 16.17 128.195 16.24 ;
    RECT 128.125 19.775 128.195 19.845 ;
    RECT 128.125 22.655 128.195 22.725 ;
    RECT 128.125 23.375 128.195 23.445 ;
    RECT 128.125 24.82 128.195 24.89 ;
    RECT 128.125 26.255 128.195 26.325 ;
    RECT 128.125 28.415 128.195 28.485 ;
    RECT 128.335 17.605 128.405 17.675 ;
    RECT 128.335 21.22 128.545 21.29 ;
    RECT 128.335 21.935 128.545 22.005 ;
    RECT 128.335 32.025 128.545 32.095 ;
    RECT 128.37 16.89 128.44 16.96 ;
    RECT 128.475 17.605 128.545 17.675 ;
    RECT 128.705 16.17 128.935 16.24 ;
    RECT 128.705 16.885 128.935 16.955 ;
    RECT 128.705 19.775 128.935 19.845 ;
    RECT 128.705 22.655 128.935 22.725 ;
    RECT 128.705 23.375 128.935 23.445 ;
    RECT 128.705 24.82 128.935 24.89 ;
    RECT 128.705 25.535 128.935 25.605 ;
    RECT 128.705 26.255 128.935 26.325 ;
    RECT 128.705 27.695 128.935 27.765 ;
    RECT 128.705 28.415 128.935 28.485 ;
    RECT 129.415 16.885 129.685 16.955 ;
    RECT 129.415 19.775 129.685 19.845 ;
    RECT 129.415 22.655 129.685 22.725 ;
    RECT 129.415 23.375 129.685 23.445 ;
    RECT 129.415 24.82 129.685 24.89 ;
    RECT 129.415 25.535 129.685 25.605 ;
    RECT 129.415 26.255 129.685 26.325 ;
    RECT 129.415 27.695 129.685 27.765 ;
    RECT 129.415 28.415 129.685 28.485 ;
    RECT 129.42 16.17 129.68 16.24 ;
    RECT 129.42 30.58 129.68 30.65 ;
    RECT 129.94 16.17 130.2 16.24 ;
    RECT 129.965 26.97 130.175 27.04 ;
    RECT 129.965 29.13 130.175 29.2 ;
    RECT 129.965 29.85 130.175 29.92 ;
    RECT 130.59 18.335 130.66 18.405 ;
    RECT 130.985 16.17 131.225 16.24 ;
    RECT 131.0 26.97 131.21 27.04 ;
    RECT 131.0 29.13 131.21 29.2 ;
    RECT 131.0 29.85 131.21 29.92 ;
    RECT 131.385 16.885 131.655 16.955 ;
    RECT 131.385 19.775 131.655 19.845 ;
    RECT 131.385 21.94 131.655 22.01 ;
    RECT 131.385 22.655 131.655 22.725 ;
    RECT 131.385 23.375 131.655 23.445 ;
    RECT 131.385 24.82 131.655 24.89 ;
    RECT 131.385 25.535 131.655 25.605 ;
    RECT 131.385 26.255 131.655 26.325 ;
    RECT 131.385 27.695 131.655 27.765 ;
    RECT 131.385 28.415 131.655 28.485 ;
    RECT 131.795 17.605 131.865 17.675 ;
    RECT 131.795 17.605 131.865 17.675 ;
    RECT 131.795 37.06 131.865 37.13 ;
    RECT 131.995 36.34 132.065 36.41 ;
    RECT 132.195 33.46 132.265 33.53 ;
    RECT 132.395 30.58 132.465 30.65 ;
    RECT 132.395 34.895 132.465 34.965 ;
    RECT 132.595 28.415 132.665 28.485 ;
    RECT 132.595 34.175 132.665 34.245 ;
    RECT 132.79 25.535 132.86 25.605 ;
    RECT 132.79 35.615 132.86 35.685 ;
    RECT 132.99 21.935 133.06 22.005 ;
    RECT 132.99 22.655 133.06 22.725 ;
    RECT 132.99 32.74 133.06 32.81 ;
    RECT 133.19 19.775 133.26 19.845 ;
    RECT 133.19 32.02 133.26 32.09 ;
    RECT 133.39 16.885 133.46 16.955 ;
    RECT 133.39 31.295 133.46 31.365 ;
    RECT 133.61 23.375 133.68 23.445 ;
    RECT 133.61 24.1 133.68 24.17 ;
    RECT 133.61 24.82 133.68 24.89 ;
    RECT 133.61 26.255 133.68 26.325 ;
    RECT 133.61 27.695 133.68 27.765 ;
    RECT 133.925 16.885 134.135 16.955 ;
    RECT 133.925 19.775 134.135 19.845 ;
    RECT 133.925 21.215 134.135 21.285 ;
    RECT 133.925 21.935 134.135 22.005 ;
    RECT 133.925 22.655 134.135 22.725 ;
    RECT 133.925 25.535 134.135 25.605 ;
    RECT 133.925 28.42 134.135 28.49 ;
    RECT 133.925 30.58 134.135 30.65 ;
    RECT 133.925 31.3 134.135 31.37 ;
    RECT 133.925 32.02 134.135 32.09 ;
    RECT 133.925 32.74 134.135 32.81 ;
    RECT 133.925 33.46 134.135 33.53 ;
    RECT 133.925 34.185 134.135 34.255 ;
    RECT 133.925 34.905 134.135 34.975 ;
    RECT 133.925 35.625 134.135 35.695 ;
    RECT 133.925 36.34 134.135 36.41 ;
    RECT 134.34 17.605 134.55 17.675 ;
    RECT 134.34 19.775 134.55 19.845 ;
    RECT 134.34 21.22 134.55 21.29 ;
    RECT 134.34 21.94 134.565 22.01 ;
    RECT 134.34 22.66 134.55 22.73 ;
    RECT 134.34 24.1 134.58 24.17 ;
    RECT 134.34 25.535 134.575 25.605 ;
    RECT 134.34 28.415 134.57 28.485 ;
    RECT 134.34 37.06 134.55 37.13 ;
    RECT 134.345 16.885 134.585 16.955 ;
    RECT 134.35 33.46 134.585 33.53 ;
    RECT 134.35 34.185 134.585 34.255 ;
    RECT 134.35 34.905 134.585 34.975 ;
    RECT 134.35 35.625 134.585 35.695 ;
    RECT 134.35 36.34 134.585 36.41 ;
    RECT 134.355 32.02 134.585 32.09 ;
    RECT 134.355 32.74 134.585 32.81 ;
    RECT 134.375 30.58 134.585 30.65 ;
    RECT 134.375 31.3 134.585 31.37 ;
    RECT 134.715 23.375 134.785 23.445 ;
    RECT 134.715 23.375 134.785 23.445 ;
    RECT 134.715 24.82 134.785 24.89 ;
    RECT 134.715 24.82 134.785 24.89 ;
    RECT 134.715 26.255 134.785 26.325 ;
    RECT 134.715 26.255 134.785 26.325 ;
    RECT 134.715 27.695 134.785 27.765 ;
    RECT 134.715 27.695 134.785 27.765 ;
    RECT 134.905 31.3 134.975 31.37 ;
    RECT 135.095 32.015 135.165 32.085 ;
    RECT 135.3 32.74 135.37 32.81 ;
    RECT 135.5 35.615 135.57 35.685 ;
    RECT 135.7 34.18 135.77 34.25 ;
    RECT 135.9 34.895 135.97 34.965 ;
    RECT 136.1 33.46 136.17 33.53 ;
    RECT 136.295 36.335 136.365 36.405 ;
    RECT 136.5 23.375 136.735 23.445 ;
    RECT 136.5 24.82 136.735 24.89 ;
    RECT 136.5 25.535 136.735 25.605 ;
    RECT 136.5 26.255 136.735 26.325 ;
    RECT 136.5 28.415 136.75 28.485 ;
    RECT 136.505 27.695 136.755 27.765 ;
    RECT 136.515 17.6 136.75 17.67 ;
    RECT 136.515 21.94 136.75 22.01 ;
    RECT 136.92 16.885 137.13 16.955 ;
    RECT 136.92 19.775 137.13 19.845 ;
    RECT 136.92 21.22 137.13 21.29 ;
    RECT 136.92 22.66 137.13 22.73 ;
    RECT 136.92 25.535 137.13 25.605 ;
    RECT 136.92 37.06 137.13 37.13 ;
    RECT 137.64 23.375 137.71 23.445 ;
    RECT 137.64 24.82 137.71 24.89 ;
    RECT 137.64 26.255 137.71 26.325 ;
    RECT 137.87 24.095 138.14 24.165 ;
    RECT 137.87 25.535 138.11 25.605 ;
    RECT 137.89 16.885 138.1 16.955 ;
    RECT 137.89 27.7 138.1 27.77 ;
    RECT 137.9 26.97 138.11 27.04 ;
    RECT 137.9 28.42 138.11 28.49 ;
    RECT 137.9 29.13 138.11 29.2 ;
    RECT 137.9 29.85 138.11 29.92 ;
    RECT 138.365 25.535 138.435 25.605 ;
    RECT 138.365 27.695 138.435 27.765 ;
    RECT 138.365 28.415 138.435 28.485 ;
    RECT 138.37 16.17 138.44 16.24 ;
    RECT 138.37 30.575 138.44 30.645 ;
    RECT 138.39 16.895 138.46 16.965 ;
    RECT 138.4 24.095 138.47 24.165 ;
    RECT 138.69 23.375 138.96 23.445 ;
    RECT 138.69 24.82 138.96 24.89 ;
    RECT 138.69 26.255 138.955 26.325 ;
    RECT 138.7 25.535 138.96 25.605 ;
    RECT 138.7 30.575 138.96 30.645 ;
    RECT 138.715 27.695 138.96 27.765 ;
    RECT 138.735 16.17 138.96 16.24 ;
    RECT 138.735 16.885 138.96 16.955 ;
    RECT 138.735 24.095 138.96 24.165 ;
    RECT 138.735 28.415 138.96 28.485 ;
    RECT 139.7 16.89 139.97 16.96 ;
    RECT 139.705 14.415 139.965 14.485 ;
    RECT 139.73 14.745 139.94 14.815 ;
    RECT 139.73 16.175 139.94 16.245 ;
    RECT 139.73 18.34 139.94 18.41 ;
    RECT 139.73 19.06 139.94 19.13 ;
    RECT 139.73 19.775 139.94 19.845 ;
    RECT 139.73 21.22 139.94 21.29 ;
    RECT 139.73 21.935 139.94 22.005 ;
    RECT 139.73 22.66 139.94 22.73 ;
    RECT 139.73 23.375 139.94 23.445 ;
    RECT 139.73 24.82 139.94 24.89 ;
    RECT 139.73 26.26 139.94 26.33 ;
    RECT 139.73 28.42 139.94 28.49 ;
    RECT 139.73 30.58 139.94 30.65 ;
    RECT 139.76 20.495 139.97 20.565 ;
    RECT 140.445 15.46 140.715 15.53 ;
    RECT 140.445 16.89 140.715 16.96 ;
    RECT 140.45 14.74 140.71 14.81 ;
    RECT 140.45 17.605 140.71 17.675 ;
    RECT 140.45 32.015 140.66 32.085 ;
    RECT 140.45 32.735 140.66 32.805 ;
    RECT 140.45 33.455 140.71 33.525 ;
    RECT 140.45 34.18 140.71 34.25 ;
    RECT 140.45 34.9 140.71 34.97 ;
    RECT 140.45 35.62 140.71 35.69 ;
    RECT 140.45 36.335 140.71 36.405 ;
    RECT 140.475 26.97 140.685 27.04 ;
    RECT 140.475 29.13 140.685 29.2 ;
    RECT 140.475 29.85 140.685 29.92 ;
    RECT 140.5 18.34 140.71 18.41 ;
    RECT 140.5 20.5 140.71 20.57 ;
    RECT 140.5 23.38 140.71 23.45 ;
    RECT 140.5 24.82 140.71 24.89 ;
    RECT 140.5 26.26 140.71 26.33 ;
    RECT 140.5 28.42 140.71 28.49 ;
    RECT 140.5 30.58 140.71 30.65 ;
    RECT 140.505 19.06 140.715 19.13 ;
    RECT 140.895 29.13 140.965 29.2 ;
    RECT 140.895 29.85 140.965 29.92 ;
    RECT 140.895 30.58 140.965 30.65 ;
    RECT 140.895 32.015 140.965 32.085 ;
    RECT 140.895 32.735 140.965 32.805 ;
    RECT 140.895 33.455 140.965 33.525 ;
    RECT 140.895 34.18 140.965 34.25 ;
    RECT 140.895 34.9 140.965 34.97 ;
    RECT 140.895 35.62 140.965 35.69 ;
    RECT 140.895 36.335 140.965 36.405 ;
    RECT 140.895 37.06 140.965 37.13 ;
    RECT 141.385 14.74 141.645 14.81 ;
    RECT 141.385 15.455 141.645 15.525 ;
    RECT 141.385 16.89 141.645 16.96 ;
    RECT 141.385 17.605 141.645 17.675 ;
    RECT 141.385 18.34 141.645 18.41 ;
    RECT 141.385 19.055 141.645 19.125 ;
    RECT 141.385 20.495 141.645 20.565 ;
    RECT 141.385 26.255 141.645 26.325 ;
    RECT 141.385 29.13 141.645 29.2 ;
    RECT 141.385 29.85 141.645 29.92 ;
    RECT 141.385 30.58 141.645 30.65 ;
    RECT 141.385 32.015 141.645 32.085 ;
    RECT 141.385 32.735 141.645 32.805 ;
    RECT 141.385 33.455 141.645 33.525 ;
    RECT 141.385 34.18 141.645 34.25 ;
    RECT 141.385 34.9 141.645 34.97 ;
    RECT 141.385 35.62 141.645 35.69 ;
    RECT 141.385 36.335 141.645 36.405 ;
    RECT 141.385 37.055 141.645 37.125 ;
    RECT 141.415 16.175 141.625 16.245 ;
    RECT 141.415 19.775 141.625 19.845 ;
    RECT 141.415 21.22 141.625 21.29 ;
    RECT 141.415 21.935 141.625 22.005 ;
    RECT 141.415 22.66 141.625 22.73 ;
    RECT 142.51 14.74 142.72 14.81 ;
    RECT 142.51 15.455 142.72 15.525 ;
    RECT 142.51 16.17 142.72 16.24 ;
    RECT 142.51 16.89 142.72 16.96 ;
    RECT 142.51 17.62 142.72 17.69 ;
    RECT 142.51 18.34 142.72 18.41 ;
    RECT 142.51 19.055 142.72 19.125 ;
    RECT 142.51 19.775 142.72 19.845 ;
    RECT 142.51 20.495 142.72 20.565 ;
    RECT 142.51 21.215 142.72 21.285 ;
    RECT 142.51 21.94 142.72 22.01 ;
    RECT 142.51 22.66 142.72 22.73 ;
    RECT 142.51 25.535 142.72 25.605 ;
    RECT 142.51 26.255 142.72 26.325 ;
    RECT 142.51 27.7 142.72 27.77 ;
    RECT 142.51 29.13 142.72 29.2 ;
    RECT 142.51 29.85 142.72 29.92 ;
    RECT 142.51 30.58 142.72 30.65 ;
    RECT 142.51 31.295 142.72 31.365 ;
    RECT 142.51 32.015 142.72 32.085 ;
    RECT 142.51 32.735 142.72 32.805 ;
    RECT 142.51 33.455 142.72 33.525 ;
    RECT 142.51 34.18 142.72 34.25 ;
    RECT 142.51 34.9 142.72 34.97 ;
    RECT 142.51 35.62 142.72 35.69 ;
    RECT 142.51 36.335 142.72 36.405 ;
    RECT 142.51 37.055 142.72 37.125 ;
    RECT 144.345 14.915 145.135 14.985 ;
    RECT 144.345 15.635 145.135 15.705 ;
    RECT 144.345 16.35 145.135 16.42 ;
    RECT 144.345 17.075 145.135 17.145 ;
    RECT 144.345 17.795 145.135 17.865 ;
    RECT 144.345 18.515 145.135 18.585 ;
    RECT 144.345 19.23 145.135 19.3 ;
    RECT 144.345 19.955 145.135 20.025 ;
    RECT 144.345 20.675 145.135 20.745 ;
    RECT 144.345 21.39 145.135 21.46 ;
    RECT 144.345 22.115 145.135 22.185 ;
    RECT 144.345 22.835 145.135 22.905 ;
    RECT 144.345 23.555 145.135 23.625 ;
    RECT 144.345 24.275 145.135 24.345 ;
    RECT 144.345 24.995 145.135 25.065 ;
    RECT 144.345 25.715 145.135 25.785 ;
    RECT 144.345 26.435 145.135 26.505 ;
    RECT 144.345 27.155 145.135 27.225 ;
    RECT 144.345 27.875 145.135 27.945 ;
    RECT 144.345 28.595 145.135 28.665 ;
    RECT 144.345 29.315 145.135 29.385 ;
    RECT 144.345 30.035 145.135 30.105 ;
    RECT 144.345 30.75 145.135 30.82 ;
    RECT 144.345 31.47 145.135 31.54 ;
    RECT 144.345 32.195 145.135 32.265 ;
    RECT 144.345 32.915 145.135 32.985 ;
    RECT 144.345 33.635 145.135 33.705 ;
    RECT 144.345 34.355 145.135 34.425 ;
    RECT 144.345 35.075 145.135 35.145 ;
    RECT 144.345 35.79 145.135 35.86 ;
    RECT 144.345 36.51 145.135 36.58 ;
    RECT 144.345 37.235 145.135 37.305 ;
    RECT 146.125 14.47 146.395 37.58 ;
    RECT 146.125 35.35 146.395 35.42 ;
    RECT 135.305 83.877 135.375 83.947 ;
    RECT 127.69 59.377 127.9 59.447 ;
    RECT 135.105 43.537 135.175 43.607 ;
    RECT 145.485 89.01 145.695 89.08 ;
    RECT 132.195 56.497 132.265 56.567 ;
    RECT 139.73 88.92 139.94 88.99 ;
    RECT 133.39 84.597 133.46 84.667 ;
    RECT 127.69 88.917 127.9 88.987 ;
    RECT 122.63 59.47 122.84 59.54 ;
    RECT 135.305 69.477 135.375 69.547 ;
    RECT 135.305 78.837 135.375 78.907 ;
    RECT 122.63 89.01 122.84 89.08 ;
    RECT 122.63 67.41 122.84 67.48 ;
    RECT 132.79 70.197 132.86 70.267 ;
    RECT 135.305 64.437 135.375 64.507 ;
    RECT 132.195 79.557 132.265 79.627 ;
    RECT 133.19 65.157 133.26 65.227 ;
    RECT 135.5 91.797 135.57 91.867 ;
    RECT 135.105 49.297 135.175 49.367 ;
    RECT 133.39 39.217 133.46 39.287 ;
    RECT 132.99 92.517 133.06 92.587 ;
    RECT 145.485 44.35 145.695 44.42 ;
    RECT 139.73 44.26 139.94 44.33 ;
    RECT 132.595 50.017 132.665 50.087 ;
    RECT 145.485 95.49 145.695 95.56 ;
    RECT 127.69 44.257 127.9 44.327 ;
    RECT 139.73 95.4 139.94 95.47 ;
    RECT 122.63 44.35 122.84 44.42 ;
    RECT 127.69 95.397 127.9 95.467 ;
    RECT 135.105 57.217 135.175 57.287 ;
    RECT 122.63 95.49 122.84 95.56 ;
    RECT 145.485 91.17 145.695 91.24 ;
    RECT 139.73 91.08 139.94 91.15 ;
    RECT 131.995 57.937 132.065 58.007 ;
    RECT 127.69 91.077 127.9 91.147 ;
    RECT 145.485 46.51 145.695 46.58 ;
    RECT 139.73 46.42 139.94 46.49 ;
    RECT 135.5 86.037 135.57 86.107 ;
    RECT 127.69 46.417 127.9 46.487 ;
    RECT 122.63 91.17 122.84 91.24 ;
    RECT 145.485 76.05 145.695 76.12 ;
    RECT 139.73 75.96 139.94 76.03 ;
    RECT 122.63 29.95 122.84 30.02 ;
    RECT 133.39 86.757 133.46 86.827 ;
    RECT 127.69 75.957 127.9 76.027 ;
    RECT 122.63 29.23 122.84 29.3 ;
    RECT 122.63 46.51 122.84 46.58 ;
    RECT 135.305 71.637 135.375 71.707 ;
    RECT 132.79 72.357 132.86 72.427 ;
    RECT 145.485 83.25 145.695 83.32 ;
    RECT 122.63 76.05 122.84 76.12 ;
    RECT 139.73 83.16 139.94 83.23 ;
    RECT 122.63 28.51 122.84 28.58 ;
    RECT 122.63 27.79 122.84 27.86 ;
    RECT 145.485 60.19 145.695 60.26 ;
    RECT 122.63 27.07 122.84 27.14 ;
    RECT 139.73 60.1 139.94 60.17 ;
    RECT 127.69 83.157 127.9 83.227 ;
    RECT 122.63 26.35 122.84 26.42 ;
    RECT 127.69 60.097 127.9 60.167 ;
    RECT 135.305 66.597 135.375 66.667 ;
    RECT 122.63 83.25 122.84 83.32 ;
    RECT 145.485 37.87 145.695 37.94 ;
    RECT 122.63 25.63 122.84 25.7 ;
    RECT 145.485 68.13 145.695 68.2 ;
    RECT 139.73 37.78 139.94 37.85 ;
    RECT 139.73 68.04 139.94 68.11 ;
    RECT 122.63 24.91 122.84 24.98 ;
    RECT 135.5 93.957 135.57 94.027 ;
    RECT 127.69 37.777 127.9 37.847 ;
    RECT 132.79 94.677 132.86 94.747 ;
    RECT 127.69 68.037 127.9 68.107 ;
    RECT 122.63 24.19 122.84 24.26 ;
    RECT 135.105 51.457 135.175 51.527 ;
    RECT 135.305 79.557 135.375 79.627 ;
    RECT 133.19 41.377 133.26 41.447 ;
    RECT 122.63 37.87 122.84 37.94 ;
    RECT 122.63 68.13 122.84 68.2 ;
    RECT 145.485 60.627 145.695 60.697 ;
    RECT 122.63 23.47 122.84 23.54 ;
    RECT 140.475 60.812 140.685 60.882 ;
    RECT 137.9 60.812 138.11 60.882 ;
    RECT 122.63 22.75 122.84 22.82 ;
    RECT 132.195 80.277 132.265 80.347 ;
    RECT 145.485 71.01 145.695 71.08 ;
    RECT 145.485 96.21 145.695 96.28 ;
    RECT 139.73 96.12 139.94 96.19 ;
    RECT 131.795 60.812 131.865 60.882 ;
    RECT 131.0 60.812 131.21 60.882 ;
    RECT 127.69 96.117 127.9 96.187 ;
    RECT 135.105 37.777 135.175 37.847 ;
    RECT 122.63 22.03 122.84 22.1 ;
    RECT 129.965 60.812 130.175 60.882 ;
    RECT 127.69 60.812 127.9 60.882 ;
    RECT 122.63 60.627 122.84 60.697 ;
    RECT 145.485 37.15 145.695 37.22 ;
    RECT 122.63 21.31 122.84 21.38 ;
    RECT 135.105 44.977 135.175 45.047 ;
    RECT 145.485 36.43 145.695 36.5 ;
    RECT 122.63 20.59 122.84 20.66 ;
    RECT 145.485 35.71 145.695 35.78 ;
    RECT 139.73 70.92 139.94 70.99 ;
    RECT 127.69 93.237 127.9 93.307 ;
    RECT 127.69 70.917 127.9 70.987 ;
    RECT 122.63 93.33 122.84 93.4 ;
    RECT 145.485 78.21 145.695 78.28 ;
    RECT 122.63 71.01 122.84 71.08 ;
    RECT 122.63 96.21 122.84 96.28 ;
    RECT 145.485 55.15 145.695 55.22 ;
    RECT 132.99 45.697 133.06 45.767 ;
    RECT 145.485 34.99 145.695 35.06 ;
    RECT 145.485 34.27 145.695 34.34 ;
    RECT 145.485 33.55 145.695 33.62 ;
    RECT 122.63 19.87 122.84 19.94 ;
    RECT 145.485 32.83 145.695 32.9 ;
    RECT 145.485 32.11 145.695 32.18 ;
    RECT 145.485 31.39 145.695 31.46 ;
    RECT 145.485 30.67 145.695 30.74 ;
    RECT 122.63 19.15 122.84 19.22 ;
    RECT 145.485 29.95 145.695 30.02 ;
    RECT 122.63 18.43 122.84 18.5 ;
    RECT 145.485 29.23 145.695 29.3 ;
    RECT 122.63 17.71 122.84 17.78 ;
    RECT 122.63 16.99 122.84 17.06 ;
    RECT 122.63 16.27 122.84 16.34 ;
    RECT 122.63 15.55 122.84 15.62 ;
    RECT 139.73 78.12 139.94 78.19 ;
    RECT 127.69 78.117 127.9 78.187 ;
    RECT 139.73 55.06 139.94 55.13 ;
    RECT 145.485 85.41 145.695 85.48 ;
    RECT 122.63 78.21 122.84 78.28 ;
    RECT 127.69 55.057 127.9 55.127 ;
    RECT 145.485 63.09 145.695 63.16 ;
    RECT 122.63 55.15 122.84 55.22 ;
    RECT 135.5 88.197 135.57 88.267 ;
    RECT 145.485 28.51 145.695 28.58 ;
    RECT 122.63 14.83 122.84 14.9 ;
    RECT 145.485 98.892 145.695 98.962 ;
    RECT 145.485 27.79 145.695 27.86 ;
    RECT 140.475 98.892 140.685 98.962 ;
    RECT 139.73 85.32 139.94 85.39 ;
    RECT 135.305 73.797 135.375 73.867 ;
    RECT 139.73 63.0 139.94 63.07 ;
    RECT 127.69 85.317 127.9 85.387 ;
    RECT 127.69 62.997 127.9 63.067 ;
    RECT 122.63 85.41 122.84 85.48 ;
    RECT 122.63 63.09 122.84 63.16 ;
    RECT 145.485 27.07 145.695 27.14 ;
    RECT 145.485 26.35 145.695 26.42 ;
    RECT 145.485 25.63 145.695 25.7 ;
    RECT 145.485 24.91 145.695 24.98 ;
    RECT 139.73 99.325 139.94 99.395 ;
    RECT 137.9 98.892 138.11 98.962 ;
    RECT 145.485 24.19 145.695 24.26 ;
    RECT 136.92 99.325 137.13 99.395 ;
    RECT 131.795 99.325 131.865 99.395 ;
    RECT 145.485 40.03 145.695 40.1 ;
    RECT 139.73 39.94 139.94 40.01 ;
    RECT 145.485 47.23 145.695 47.3 ;
    RECT 127.69 39.937 127.9 40.007 ;
    RECT 139.73 47.14 139.94 47.21 ;
    RECT 127.69 47.137 127.9 47.207 ;
    RECT 145.485 23.47 145.695 23.54 ;
    RECT 131.0 98.892 131.21 98.962 ;
    RECT 145.485 22.75 145.695 22.82 ;
    RECT 129.965 98.892 130.175 98.962 ;
    RECT 145.485 22.03 145.695 22.1 ;
    RECT 145.485 21.31 145.695 21.38 ;
    RECT 127.69 98.892 127.9 98.962 ;
    RECT 145.485 20.59 145.695 20.66 ;
    RECT 145.485 19.87 145.695 19.94 ;
    RECT 126.76 99.325 126.97 99.395 ;
    RECT 122.63 98.892 122.84 98.962 ;
    RECT 122.63 40.03 122.84 40.1 ;
    RECT 135.305 67.317 135.375 67.387 ;
    RECT 145.485 73.17 145.695 73.24 ;
    RECT 139.73 73.08 139.94 73.15 ;
    RECT 145.485 98.37 145.695 98.44 ;
    RECT 135.105 52.177 135.175 52.247 ;
    RECT 139.73 98.28 139.94 98.35 ;
    RECT 132.99 43.537 133.06 43.607 ;
    RECT 132.99 68.037 133.06 68.107 ;
    RECT 127.69 98.277 127.9 98.347 ;
    RECT 132.395 52.897 132.465 52.967 ;
    RECT 127.69 73.077 127.9 73.147 ;
    RECT 122.63 73.17 122.84 73.24 ;
    RECT 135.5 89.637 135.57 89.707 ;
    RECT 122.63 98.37 122.84 98.44 ;
    RECT 145.485 57.31 145.695 57.38 ;
    RECT 139.73 57.22 139.94 57.29 ;
    RECT 135.105 39.937 135.175 40.007 ;
    RECT 135.305 75.237 135.375 75.307 ;
    RECT 127.69 80.277 127.9 80.347 ;
    RECT 144.925 60.627 145.135 60.697 ;
    RECT 122.63 80.37 122.84 80.44 ;
    RECT 127.69 57.217 127.9 57.287 ;
    RECT 145.485 65.25 145.695 65.32 ;
    RECT 122.63 57.31 122.84 57.38 ;
    RECT 139.73 65.16 139.94 65.23 ;
    RECT 132.395 75.957 132.465 76.027 ;
    RECT 135.105 60.097 135.175 60.167 ;
    RECT 127.69 65.157 127.9 65.227 ;
    RECT 122.63 65.25 122.84 65.32 ;
    RECT 145.485 49.39 145.695 49.46 ;
    RECT 139.73 49.3 139.94 49.37 ;
    RECT 133.39 61.557 133.46 61.627 ;
    RECT 121.44 98.01 121.51 98.8 ;
    RECT 122.04 98.01 122.25 98.08 ;
    RECT 122.04 98.365 122.25 98.435 ;
    RECT 122.04 98.73 122.25 98.8 ;
    RECT 123.205 98.455 124.005 98.525 ;
    RECT 125.67 98.28 125.905 98.35 ;
    RECT 126.73 98.28 126.99 98.35 ;
    RECT 128.705 98.28 128.935 98.35 ;
    RECT 129.42 98.28 129.68 98.35 ;
    RECT 130.59 98.28 130.66 98.35 ;
    RECT 133.925 98.28 134.135 98.35 ;
    RECT 134.31 98.28 134.58 98.35 ;
    RECT 138.365 98.28 138.435 98.35 ;
    RECT 138.695 98.28 138.96 98.35 ;
    RECT 140.45 98.28 140.71 98.35 ;
    RECT 140.895 98.28 140.965 98.35 ;
    RECT 141.385 98.28 141.645 98.35 ;
    RECT 142.51 98.28 142.72 98.35 ;
    RECT 144.32 98.455 145.135 98.525 ;
    RECT 146.125 98.01 146.395 98.08 ;
    RECT 146.125 98.365 146.395 98.435 ;
    RECT 146.125 98.73 146.395 98.8 ;
    RECT 133.19 89.637 133.26 89.707 ;
    RECT 127.69 49.297 127.9 49.367 ;
    RECT 122.63 49.39 122.84 49.46 ;
    RECT 135.105 55.057 135.175 55.127 ;
    RECT 145.485 40.75 145.695 40.82 ;
    RECT 135.5 96.837 135.57 96.907 ;
    RECT 135.305 82.437 135.375 82.507 ;
    RECT 139.73 40.66 139.94 40.73 ;
    RECT 132.595 97.557 132.665 97.627 ;
    RECT 127.69 40.657 127.9 40.727 ;
    RECT 122.63 40.75 122.84 40.82 ;
    RECT 132.195 55.057 132.265 55.127 ;
    RECT 131.995 83.157 132.065 83.227 ;
    RECT 135.105 42.097 135.175 42.167 ;
    RECT 135.305 77.397 135.375 77.467 ;
    RECT 145.485 73.89 145.695 73.96 ;
    RECT 139.73 73.8 139.94 73.87 ;
    RECT 145.485 51.55 145.695 51.62 ;
    RECT 139.73 51.46 139.94 51.53 ;
    RECT 132.395 78.117 132.465 78.187 ;
    RECT 145.485 81.09 145.695 81.16 ;
    RECT 139.73 81.0 139.94 81.07 ;
    RECT 135.305 62.997 135.375 63.067 ;
    RECT 127.69 51.457 127.9 51.527 ;
    RECT 135.5 90.357 135.57 90.427 ;
    RECT 122.63 51.55 122.84 51.62 ;
    RECT 135.105 47.857 135.175 47.927 ;
    RECT 133.39 63.717 133.46 63.787 ;
    RECT 133.39 37.777 133.46 37.847 ;
    RECT 127.69 80.997 127.9 81.067 ;
    RECT 132.99 91.077 133.06 91.147 ;
    RECT 145.485 88.29 145.695 88.36 ;
    RECT 122.63 81.09 122.84 81.16 ;
    RECT 139.73 88.2 139.94 88.27 ;
    RECT 132.79 48.577 132.86 48.647 ;
    RECT 127.69 88.197 127.9 88.267 ;
    RECT 122.63 88.29 122.84 88.36 ;
    RECT 145.485 42.91 145.695 42.98 ;
    RECT 139.73 42.82 139.94 42.89 ;
    RECT 145.485 52.99 145.695 53.06 ;
    RECT 139.73 52.9 139.94 52.97 ;
    RECT 127.69 52.897 127.9 52.967 ;
    RECT 145.485 94.05 145.695 94.12 ;
    RECT 127.69 42.817 127.9 42.887 ;
    RECT 139.73 93.96 139.94 94.03 ;
    RECT 122.63 42.91 122.84 42.98 ;
    RECT 122.63 52.99 122.84 53.06 ;
    RECT 127.69 93.957 127.9 94.027 ;
    RECT 122.63 94.05 122.84 94.12 ;
    RECT 145.485 89.73 145.695 89.8 ;
    RECT 135.105 44.257 135.175 44.327 ;
    RECT 139.73 89.64 139.94 89.71 ;
    RECT 132.195 57.217 132.265 57.287 ;
    RECT 127.69 89.637 127.9 89.707 ;
    RECT 122.63 60.19 122.84 60.26 ;
    RECT 135.5 84.597 135.57 84.667 ;
    RECT 133.39 85.317 133.46 85.387 ;
    RECT 145.485 45.07 145.695 45.14 ;
    RECT 139.73 44.98 139.94 45.05 ;
    RECT 127.69 44.977 127.9 45.047 ;
    RECT 135.305 70.197 135.375 70.267 ;
    RECT 122.63 89.73 122.84 89.8 ;
    RECT 145.485 74.61 145.695 74.68 ;
    RECT 139.73 74.52 139.94 74.59 ;
    RECT 127.69 74.517 127.9 74.587 ;
    RECT 122.63 45.07 122.84 45.14 ;
    RECT 132.79 70.917 132.86 70.987 ;
    RECT 145.485 81.81 145.695 81.88 ;
    RECT 122.63 74.61 122.84 74.68 ;
    RECT 139.73 81.72 139.94 81.79 ;
    RECT 127.69 81.717 127.9 81.787 ;
    RECT 135.305 65.157 135.375 65.227 ;
    RECT 133.19 65.877 133.26 65.947 ;
    RECT 135.5 92.517 135.57 92.587 ;
    RECT 135.105 50.017 135.175 50.087 ;
    RECT 133.39 39.937 133.46 40.007 ;
    RECT 122.63 81.81 122.84 81.88 ;
    RECT 132.79 93.237 132.86 93.307 ;
    RECT 132.595 50.737 132.665 50.807 ;
    RECT 145.485 91.89 145.695 91.96 ;
    RECT 139.73 91.8 139.94 91.87 ;
    RECT 127.69 91.797 127.9 91.867 ;
    RECT 122.63 91.89 122.84 91.96 ;
    RECT 135.105 57.937 135.175 58.007 ;
    RECT 135.5 86.757 135.57 86.827 ;
    RECT 131.995 58.657 132.065 58.727 ;
    RECT 145.485 76.77 145.695 76.84 ;
    RECT 139.73 76.68 139.94 76.75 ;
    RECT 145.485 53.71 145.695 53.78 ;
    RECT 127.69 76.677 127.9 76.747 ;
    RECT 139.73 53.62 139.94 53.69 ;
    RECT 122.63 47.23 122.84 47.3 ;
    RECT 133.19 87.477 133.26 87.547 ;
    RECT 127.69 53.617 127.9 53.687 ;
    RECT 145.485 19.15 145.695 19.22 ;
    RECT 145.485 18.43 145.695 18.5 ;
    RECT 145.485 17.71 145.695 17.78 ;
    RECT 145.485 16.99 145.695 17.06 ;
    RECT 145.485 16.27 145.695 16.34 ;
    RECT 145.485 15.55 145.695 15.62 ;
    RECT 145.485 14.83 145.695 14.9 ;
    RECT 135.305 72.357 135.375 72.427 ;
    RECT 145.485 83.97 145.695 84.04 ;
    RECT 122.63 76.77 122.84 76.84 ;
    RECT 139.73 83.88 139.94 83.95 ;
    RECT 145.485 61.65 145.695 61.72 ;
    RECT 139.73 61.56 139.94 61.63 ;
    RECT 127.69 83.877 127.9 83.947 ;
    RECT 127.69 61.557 127.9 61.627 ;
    RECT 132.595 73.077 132.665 73.147 ;
    RECT 122.63 83.97 122.84 84.04 ;
    RECT 145.485 38.59 145.695 38.66 ;
    RECT 145.485 68.85 145.695 68.92 ;
    RECT 122.63 61.65 122.84 61.72 ;
    RECT 139.73 38.5 139.94 38.57 ;
    RECT 139.73 68.76 139.94 68.83 ;
    RECT 127.69 38.497 127.9 38.567 ;
    RECT 127.69 68.757 127.9 68.827 ;
    RECT 135.5 94.677 135.57 94.747 ;
    RECT 140.475 22.657 140.685 22.727 ;
    RECT 133.19 42.097 133.26 42.167 ;
    RECT 135.305 80.277 135.375 80.347 ;
    RECT 122.63 38.59 122.84 38.66 ;
    RECT 122.63 68.85 122.84 68.92 ;
    RECT 132.79 95.397 132.86 95.467 ;
    RECT 140.475 21.937 140.685 22.007 ;
    RECT 132.195 80.997 132.265 81.067 ;
    RECT 140.475 21.217 140.685 21.287 ;
    RECT 140.475 19.777 140.685 19.847 ;
    RECT 145.485 71.73 145.695 71.8 ;
    RECT 140.475 16.175 140.685 16.245 ;
    RECT 139.73 71.64 139.94 71.71 ;
    RECT 145.485 96.93 145.695 97.0 ;
    RECT 139.73 96.84 139.94 96.91 ;
    RECT 127.69 96.837 127.9 96.907 ;
    RECT 135.105 38.497 135.175 38.567 ;
    RECT 135.105 45.697 135.175 45.767 ;
    RECT 127.69 71.637 127.9 71.707 ;
    RECT 145.485 78.93 145.695 79.0 ;
    RECT 122.63 71.73 122.84 71.8 ;
    RECT 139.73 78.84 139.94 78.91 ;
    RECT 122.63 96.93 122.84 97.0 ;
    RECT 145.485 55.87 145.695 55.94 ;
    RECT 132.79 46.417 132.86 46.487 ;
    RECT 132.595 74.517 132.665 74.587 ;
    RECT 127.69 78.837 127.9 78.907 ;
    RECT 139.73 55.78 139.94 55.85 ;
    RECT 139.73 29.85 139.94 29.92 ;
    RECT 145.485 86.13 145.695 86.2 ;
    RECT 139.73 29.13 139.94 29.2 ;
    RECT 122.63 78.93 122.84 79.0 ;
    RECT 127.69 55.777 127.9 55.847 ;
    RECT 139.73 26.97 139.94 27.04 ;
    RECT 139.73 86.04 139.94 86.11 ;
    RECT 145.485 63.81 145.695 63.88 ;
    RECT 122.63 55.87 122.84 55.94 ;
    RECT 137.9 22.657 138.11 22.727 ;
    RECT 131.995 59.377 132.065 59.447 ;
    RECT 139.73 63.72 139.94 63.79 ;
    RECT 127.69 86.037 127.9 86.107 ;
    RECT 137.9 21.217 138.11 21.287 ;
    RECT 127.69 63.717 127.9 63.787 ;
    RECT 122.63 86.13 122.84 86.2 ;
    RECT 137.9 19.777 138.11 19.847 ;
    RECT 137.9 14.745 138.11 14.815 ;
    RECT 122.63 63.81 122.84 63.88 ;
    RECT 145.485 47.95 145.695 48.02 ;
    RECT 139.73 47.86 139.94 47.93 ;
    RECT 127.69 47.857 127.9 47.927 ;
    RECT 122.63 47.95 122.84 48.02 ;
    RECT 135.305 68.037 135.375 68.107 ;
    RECT 135.105 52.897 135.175 52.967 ;
    RECT 132.99 68.757 133.06 68.827 ;
    RECT 132.99 44.257 133.06 44.327 ;
    RECT 137.002 27.697 137.072 27.767 ;
    RECT 132.595 96.117 132.665 96.187 ;
    RECT 136.92 29.85 137.13 29.92 ;
    RECT 136.92 29.13 137.13 29.2 ;
    RECT 136.92 28.417 137.13 28.487 ;
    RECT 136.92 26.97 137.13 27.04 ;
    RECT 127.69 73.797 127.9 73.867 ;
    RECT 132.395 53.617 132.465 53.687 ;
    RECT 122.63 73.89 122.84 73.96 ;
    RECT 145.485 58.03 145.695 58.1 ;
    RECT 139.73 57.94 139.94 58.01 ;
    RECT 135.105 40.657 135.175 40.727 ;
    RECT 131.995 81.717 132.065 81.787 ;
    RECT 127.69 57.937 127.9 58.007 ;
    RECT 146.16 61.05 146.37 61.12 ;
    RECT 143.69 61.177 143.9 61.247 ;
    RECT 143.065 61.177 143.135 61.247 ;
    RECT 145.485 65.97 145.695 66.04 ;
    RECT 122.63 58.03 122.84 58.1 ;
    RECT 141.415 61.177 141.625 61.247 ;
    RECT 139.73 65.88 139.94 65.95 ;
    RECT 135.305 75.957 135.375 76.027 ;
    RECT 127.69 65.877 127.9 65.947 ;
    RECT 135.305 61.557 135.375 61.627 ;
    RECT 122.63 65.97 122.84 66.04 ;
    RECT 145.485 50.11 145.695 50.18 ;
    RECT 132.395 76.677 132.465 76.747 ;
    RECT 139.73 50.02 139.94 50.09 ;
    RECT 133.39 62.277 133.46 62.347 ;
    RECT 127.69 50.017 127.9 50.087 ;
    RECT 122.63 50.11 122.84 50.18 ;
    RECT 135.105 55.777 135.175 55.847 ;
    RECT 132.99 90.357 133.06 90.427 ;
    RECT 145.485 86.85 145.695 86.92 ;
    RECT 139.73 86.76 139.94 86.83 ;
    RECT 145.485 41.47 145.695 41.54 ;
    RECT 135.5 97.557 135.57 97.627 ;
    RECT 139.73 41.38 139.94 41.45 ;
    RECT 127.69 41.377 127.9 41.447 ;
    RECT 122.63 41.47 122.84 41.54 ;
    RECT 132.595 98.277 132.665 98.347 ;
    RECT 132.195 55.777 132.265 55.847 ;
    RECT 135.305 83.157 135.375 83.227 ;
    RECT 135.105 42.817 135.175 42.887 ;
    RECT 135.305 68.757 135.375 68.827 ;
    RECT 131.995 83.877 132.065 83.947 ;
    RECT 132.99 69.477 133.06 69.547 ;
    RECT 135.305 78.117 135.375 78.187 ;
    RECT 132.195 78.837 132.265 78.907 ;
    RECT 121.44 97.29 121.51 98.08 ;
    RECT 122.04 97.29 122.25 97.36 ;
    RECT 122.04 97.645 122.25 97.715 ;
    RECT 122.04 98.01 122.25 98.08 ;
    RECT 123.205 97.735 124.005 97.805 ;
    RECT 125.67 97.56 125.905 97.63 ;
    RECT 126.73 97.56 126.99 97.63 ;
    RECT 128.705 97.56 128.935 97.63 ;
    RECT 129.42 97.56 129.68 97.63 ;
    RECT 130.59 97.56 130.66 97.63 ;
    RECT 133.925 97.56 134.135 97.63 ;
    RECT 134.31 97.56 134.58 97.63 ;
    RECT 138.365 97.56 138.435 97.63 ;
    RECT 138.695 97.56 138.96 97.63 ;
    RECT 140.45 97.56 140.71 97.63 ;
    RECT 140.895 97.56 140.965 97.63 ;
    RECT 141.385 97.56 141.645 97.63 ;
    RECT 142.51 97.56 142.72 97.63 ;
    RECT 144.32 97.735 145.135 97.805 ;
    RECT 146.125 97.29 146.395 97.36 ;
    RECT 146.125 97.645 146.395 97.715 ;
    RECT 146.125 98.01 146.395 98.08 ;
    RECT 121.44 96.57 121.51 97.36 ;
    RECT 122.04 96.57 122.25 96.64 ;
    RECT 122.04 96.925 122.25 96.995 ;
    RECT 122.04 97.29 122.25 97.36 ;
    RECT 123.205 97.015 124.005 97.085 ;
    RECT 125.67 96.84 125.905 96.91 ;
    RECT 126.73 96.84 126.99 96.91 ;
    RECT 128.705 96.84 128.935 96.91 ;
    RECT 129.42 96.84 129.68 96.91 ;
    RECT 130.59 96.84 130.66 96.91 ;
    RECT 133.925 96.84 134.135 96.91 ;
    RECT 134.31 96.84 134.58 96.91 ;
    RECT 138.365 96.84 138.435 96.91 ;
    RECT 138.695 96.84 138.96 96.91 ;
    RECT 140.45 96.84 140.71 96.91 ;
    RECT 140.895 96.84 140.965 96.91 ;
    RECT 141.385 96.84 141.645 96.91 ;
    RECT 142.51 96.84 142.72 96.91 ;
    RECT 144.32 97.015 145.135 97.085 ;
    RECT 146.125 96.57 146.395 96.64 ;
    RECT 146.125 96.925 146.395 96.995 ;
    RECT 146.125 97.29 146.395 97.36 ;
    RECT 121.44 95.85 121.51 96.64 ;
    RECT 122.04 95.85 122.25 95.92 ;
    RECT 122.04 96.205 122.25 96.275 ;
    RECT 122.04 96.57 122.25 96.64 ;
    RECT 123.205 96.295 124.005 96.365 ;
    RECT 125.67 96.12 125.905 96.19 ;
    RECT 126.73 96.12 126.99 96.19 ;
    RECT 128.705 96.12 128.935 96.19 ;
    RECT 129.42 96.12 129.68 96.19 ;
    RECT 130.59 96.12 130.66 96.19 ;
    RECT 133.925 96.12 134.135 96.19 ;
    RECT 134.31 96.12 134.58 96.19 ;
    RECT 138.365 96.12 138.435 96.19 ;
    RECT 138.695 96.12 138.96 96.19 ;
    RECT 140.45 96.12 140.71 96.19 ;
    RECT 140.895 96.12 140.965 96.19 ;
    RECT 141.385 96.12 141.645 96.19 ;
    RECT 142.51 96.12 142.72 96.19 ;
    RECT 144.32 96.295 145.135 96.365 ;
    RECT 146.125 95.85 146.395 95.92 ;
    RECT 146.125 96.205 146.395 96.275 ;
    RECT 146.125 96.57 146.395 96.64 ;
    RECT 121.44 98.73 121.51 98.8 ;
    RECT 122.04 98.73 122.25 98.8 ;
    RECT 122.395 99.75 122.465 99.82 ;
    RECT 123.235 99.185 123.975 99.255 ;
    RECT 124.255 98.895 124.465 98.965 ;
    RECT 124.715 99.75 124.925 99.82 ;
    RECT 125.11 98.895 125.32 98.965 ;
    RECT 126.76 98.895 126.97 98.965 ;
    RECT 127.32 99.75 127.53 99.82 ;
    RECT 127.69 99.325 127.9 99.395 ;
    RECT 128.105 99.75 128.175 99.82 ;
    RECT 128.715 99.75 128.925 99.82 ;
    RECT 129.445 99.75 129.655 99.82 ;
    RECT 129.965 99.325 130.175 99.395 ;
    RECT 131.0 99.325 131.21 99.395 ;
    RECT 131.415 99.75 131.625 99.82 ;
    RECT 131.795 98.895 131.865 98.965 ;
    RECT 133.575 99.75 133.785 99.82 ;
    RECT 134.34 98.895 134.55 98.965 ;
    RECT 134.715 99.75 134.785 99.82 ;
    RECT 136.535 99.75 136.745 99.82 ;
    RECT 136.92 98.895 137.13 98.965 ;
    RECT 137.625 99.75 137.695 99.82 ;
    RECT 137.9 99.325 138.11 99.395 ;
    RECT 138.37 99.04 138.44 99.11 ;
    RECT 138.72 99.75 138.93 99.82 ;
    RECT 139.73 98.895 139.94 98.965 ;
    RECT 140.475 99.325 140.685 99.395 ;
    RECT 141.415 98.895 141.625 98.965 ;
    RECT 141.935 99.75 142.145 99.82 ;
    RECT 143.065 98.895 143.135 98.965 ;
    RECT 143.31 99.75 143.52 99.82 ;
    RECT 143.69 98.895 143.9 98.965 ;
    RECT 144.345 99.185 145.135 99.255 ;
    RECT 145.87 99.75 145.94 99.82 ;
    RECT 146.125 98.73 146.395 98.8 ;
    RECT 146.765 99.75 146.975 99.82 ;
    RECT 135.305 63.717 135.375 63.787 ;
    RECT 135.5 91.077 135.57 91.147 ;
    RECT 121.44 95.13 121.51 95.92 ;
    RECT 122.04 95.13 122.25 95.2 ;
    RECT 122.04 95.485 122.25 95.555 ;
    RECT 122.04 95.85 122.25 95.92 ;
    RECT 123.205 95.575 124.005 95.645 ;
    RECT 125.67 95.4 125.905 95.47 ;
    RECT 126.73 95.4 126.99 95.47 ;
    RECT 128.705 95.4 128.935 95.47 ;
    RECT 129.42 95.4 129.68 95.47 ;
    RECT 130.59 95.4 130.66 95.47 ;
    RECT 133.925 95.4 134.135 95.47 ;
    RECT 134.31 95.4 134.58 95.47 ;
    RECT 138.365 95.4 138.435 95.47 ;
    RECT 138.695 95.4 138.96 95.47 ;
    RECT 140.45 95.4 140.71 95.47 ;
    RECT 140.895 95.4 140.965 95.47 ;
    RECT 141.385 95.4 141.645 95.47 ;
    RECT 142.51 95.4 142.72 95.47 ;
    RECT 144.32 95.575 145.135 95.645 ;
    RECT 146.125 95.13 146.395 95.2 ;
    RECT 146.125 95.485 146.395 95.555 ;
    RECT 146.125 95.85 146.395 95.92 ;
    RECT 121.44 94.41 121.51 95.2 ;
    RECT 122.04 94.41 122.25 94.48 ;
    RECT 122.04 94.765 122.25 94.835 ;
    RECT 122.04 95.13 122.25 95.2 ;
    RECT 123.205 94.855 124.005 94.925 ;
    RECT 125.67 94.68 125.905 94.75 ;
    RECT 126.73 94.68 126.99 94.75 ;
    RECT 128.705 94.68 128.935 94.75 ;
    RECT 129.42 94.68 129.68 94.75 ;
    RECT 130.59 94.68 130.66 94.75 ;
    RECT 133.925 94.68 134.135 94.75 ;
    RECT 134.31 94.68 134.58 94.75 ;
    RECT 138.365 94.68 138.435 94.75 ;
    RECT 138.695 94.68 138.96 94.75 ;
    RECT 140.45 94.68 140.71 94.75 ;
    RECT 140.895 94.68 140.965 94.75 ;
    RECT 141.385 94.68 141.645 94.75 ;
    RECT 142.51 94.68 142.72 94.75 ;
    RECT 144.32 94.855 145.135 94.925 ;
    RECT 146.125 94.41 146.395 94.48 ;
    RECT 146.125 94.765 146.395 94.835 ;
    RECT 146.125 95.13 146.395 95.2 ;
    RECT 121.44 93.69 121.51 94.48 ;
    RECT 122.04 93.69 122.25 93.76 ;
    RECT 122.04 94.045 122.25 94.115 ;
    RECT 122.04 94.41 122.25 94.48 ;
    RECT 123.205 94.135 124.005 94.205 ;
    RECT 125.67 93.96 125.905 94.03 ;
    RECT 126.73 93.96 126.99 94.03 ;
    RECT 128.705 93.96 128.935 94.03 ;
    RECT 129.42 93.96 129.68 94.03 ;
    RECT 130.59 93.96 130.66 94.03 ;
    RECT 133.925 93.96 134.135 94.03 ;
    RECT 134.31 93.96 134.58 94.03 ;
    RECT 138.365 93.96 138.435 94.03 ;
    RECT 138.695 93.96 138.96 94.03 ;
    RECT 140.45 93.96 140.71 94.03 ;
    RECT 140.895 93.96 140.965 94.03 ;
    RECT 141.385 93.96 141.645 94.03 ;
    RECT 142.51 93.96 142.72 94.03 ;
    RECT 144.32 94.135 145.135 94.205 ;
    RECT 146.125 93.69 146.395 93.76 ;
    RECT 146.125 94.045 146.395 94.115 ;
    RECT 146.125 94.41 146.395 94.48 ;
    RECT 121.44 92.97 121.51 93.76 ;
    RECT 122.04 92.97 122.25 93.04 ;
    RECT 122.04 93.325 122.25 93.395 ;
    RECT 122.04 93.69 122.25 93.76 ;
    RECT 123.205 93.415 124.005 93.485 ;
    RECT 125.67 93.24 125.905 93.31 ;
    RECT 126.73 93.24 126.99 93.31 ;
    RECT 128.705 93.24 128.935 93.31 ;
    RECT 129.42 93.24 129.68 93.31 ;
    RECT 130.59 93.24 130.66 93.31 ;
    RECT 133.925 93.24 134.135 93.31 ;
    RECT 134.31 93.24 134.58 93.31 ;
    RECT 138.365 93.24 138.435 93.31 ;
    RECT 138.695 93.24 138.96 93.31 ;
    RECT 140.45 93.24 140.71 93.31 ;
    RECT 140.895 93.24 140.965 93.31 ;
    RECT 141.385 93.24 141.645 93.31 ;
    RECT 142.51 93.24 142.72 93.31 ;
    RECT 144.32 93.415 145.135 93.485 ;
    RECT 146.125 92.97 146.395 93.04 ;
    RECT 146.125 93.325 146.395 93.395 ;
    RECT 146.125 93.69 146.395 93.76 ;
    RECT 121.44 92.25 121.51 93.04 ;
    RECT 122.04 92.25 122.25 92.32 ;
    RECT 122.04 92.605 122.25 92.675 ;
    RECT 122.04 92.97 122.25 93.04 ;
    RECT 123.205 92.695 124.005 92.765 ;
    RECT 125.67 92.52 125.905 92.59 ;
    RECT 126.73 92.52 126.99 92.59 ;
    RECT 128.705 92.52 128.935 92.59 ;
    RECT 129.42 92.52 129.68 92.59 ;
    RECT 130.59 92.52 130.66 92.59 ;
    RECT 133.925 92.52 134.135 92.59 ;
    RECT 134.31 92.52 134.58 92.59 ;
    RECT 138.365 92.52 138.435 92.59 ;
    RECT 138.695 92.52 138.96 92.59 ;
    RECT 140.45 92.52 140.71 92.59 ;
    RECT 140.895 92.52 140.965 92.59 ;
    RECT 141.385 92.52 141.645 92.59 ;
    RECT 142.51 92.52 142.72 92.59 ;
    RECT 144.32 92.695 145.135 92.765 ;
    RECT 146.125 92.25 146.395 92.32 ;
    RECT 146.125 92.605 146.395 92.675 ;
    RECT 146.125 92.97 146.395 93.04 ;
    RECT 121.44 91.53 121.51 92.32 ;
    RECT 122.04 91.53 122.25 91.6 ;
    RECT 122.04 91.885 122.25 91.955 ;
    RECT 122.04 92.25 122.25 92.32 ;
    RECT 123.205 91.975 124.005 92.045 ;
    RECT 125.67 91.8 125.905 91.87 ;
    RECT 126.73 91.8 126.99 91.87 ;
    RECT 128.705 91.8 128.935 91.87 ;
    RECT 129.42 91.8 129.68 91.87 ;
    RECT 130.59 91.8 130.66 91.87 ;
    RECT 133.925 91.8 134.135 91.87 ;
    RECT 134.31 91.8 134.58 91.87 ;
    RECT 138.365 91.8 138.435 91.87 ;
    RECT 138.695 91.8 138.96 91.87 ;
    RECT 140.45 91.8 140.71 91.87 ;
    RECT 140.895 91.8 140.965 91.87 ;
    RECT 141.385 91.8 141.645 91.87 ;
    RECT 142.51 91.8 142.72 91.87 ;
    RECT 144.32 91.975 145.135 92.045 ;
    RECT 146.125 91.53 146.395 91.6 ;
    RECT 146.125 91.885 146.395 91.955 ;
    RECT 146.125 92.25 146.395 92.32 ;
    RECT 121.44 90.81 121.51 91.6 ;
    RECT 122.04 90.81 122.25 90.88 ;
    RECT 122.04 91.165 122.25 91.235 ;
    RECT 122.04 91.53 122.25 91.6 ;
    RECT 123.205 91.255 124.005 91.325 ;
    RECT 125.67 91.08 125.905 91.15 ;
    RECT 126.73 91.08 126.99 91.15 ;
    RECT 128.705 91.08 128.935 91.15 ;
    RECT 129.42 91.08 129.68 91.15 ;
    RECT 130.59 91.08 130.66 91.15 ;
    RECT 133.925 91.08 134.135 91.15 ;
    RECT 134.31 91.08 134.58 91.15 ;
    RECT 138.365 91.08 138.435 91.15 ;
    RECT 138.695 91.08 138.96 91.15 ;
    RECT 140.45 91.08 140.71 91.15 ;
    RECT 140.895 91.08 140.965 91.15 ;
    RECT 141.385 91.08 141.645 91.15 ;
    RECT 142.51 91.08 142.72 91.15 ;
    RECT 144.32 91.255 145.135 91.325 ;
    RECT 146.125 90.81 146.395 90.88 ;
    RECT 146.125 91.165 146.395 91.235 ;
    RECT 146.125 91.53 146.395 91.6 ;
    RECT 121.44 90.09 121.51 90.88 ;
    RECT 122.04 90.09 122.25 90.16 ;
    RECT 122.04 90.445 122.25 90.515 ;
    RECT 122.04 90.81 122.25 90.88 ;
    RECT 123.205 90.535 124.005 90.605 ;
    RECT 125.67 90.36 125.905 90.43 ;
    RECT 126.73 90.36 126.99 90.43 ;
    RECT 128.705 90.36 128.935 90.43 ;
    RECT 129.42 90.36 129.68 90.43 ;
    RECT 130.59 90.36 130.66 90.43 ;
    RECT 133.925 90.36 134.135 90.43 ;
    RECT 134.31 90.36 134.58 90.43 ;
    RECT 138.365 90.36 138.435 90.43 ;
    RECT 138.695 90.36 138.96 90.43 ;
    RECT 140.45 90.36 140.71 90.43 ;
    RECT 140.895 90.36 140.965 90.43 ;
    RECT 141.385 90.36 141.645 90.43 ;
    RECT 142.51 90.36 142.72 90.43 ;
    RECT 144.32 90.535 145.135 90.605 ;
    RECT 146.125 90.09 146.395 90.16 ;
    RECT 146.125 90.445 146.395 90.515 ;
    RECT 146.125 90.81 146.395 90.88 ;
    RECT 121.44 89.37 121.51 90.16 ;
    RECT 122.04 89.37 122.25 89.44 ;
    RECT 122.04 89.725 122.25 89.795 ;
    RECT 122.04 90.09 122.25 90.16 ;
    RECT 123.205 89.815 124.005 89.885 ;
    RECT 125.67 89.64 125.905 89.71 ;
    RECT 126.73 89.64 126.99 89.71 ;
    RECT 128.705 89.64 128.935 89.71 ;
    RECT 129.42 89.64 129.68 89.71 ;
    RECT 130.59 89.64 130.66 89.71 ;
    RECT 133.925 89.64 134.135 89.71 ;
    RECT 134.31 89.64 134.58 89.71 ;
    RECT 138.365 89.64 138.435 89.71 ;
    RECT 138.695 89.64 138.96 89.71 ;
    RECT 140.45 89.64 140.71 89.71 ;
    RECT 140.895 89.64 140.965 89.71 ;
    RECT 141.385 89.64 141.645 89.71 ;
    RECT 142.51 89.64 142.72 89.71 ;
    RECT 144.32 89.815 145.135 89.885 ;
    RECT 146.125 89.37 146.395 89.44 ;
    RECT 146.125 89.725 146.395 89.795 ;
    RECT 146.125 90.09 146.395 90.16 ;
    RECT 121.44 88.65 121.51 89.44 ;
    RECT 122.04 88.65 122.25 88.72 ;
    RECT 122.04 89.005 122.25 89.075 ;
    RECT 122.04 89.37 122.25 89.44 ;
    RECT 123.205 89.095 124.005 89.165 ;
    RECT 125.67 88.92 125.905 88.99 ;
    RECT 126.73 88.92 126.99 88.99 ;
    RECT 128.705 88.92 128.935 88.99 ;
    RECT 129.42 88.92 129.68 88.99 ;
    RECT 130.59 88.92 130.66 88.99 ;
    RECT 133.925 88.92 134.135 88.99 ;
    RECT 134.31 88.92 134.58 88.99 ;
    RECT 138.365 88.92 138.435 88.99 ;
    RECT 138.695 88.92 138.96 88.99 ;
    RECT 140.45 88.92 140.71 88.99 ;
    RECT 140.895 88.92 140.965 88.99 ;
    RECT 141.385 88.92 141.645 88.99 ;
    RECT 142.51 88.92 142.72 88.99 ;
    RECT 144.32 89.095 145.135 89.165 ;
    RECT 146.125 88.65 146.395 88.72 ;
    RECT 146.125 89.005 146.395 89.075 ;
    RECT 146.125 89.37 146.395 89.44 ;
    RECT 133.19 64.437 133.26 64.507 ;
    RECT 121.44 60.55 121.51 60.62 ;
    RECT 121.44 61.29 121.51 61.36 ;
    RECT 122.04 60.55 122.25 60.62 ;
    RECT 122.04 61.29 122.25 61.36 ;
    RECT 124.225 60.81 124.495 60.88 ;
    RECT 125.19 60.81 125.26 60.88 ;
    RECT 125.645 60.63 125.905 60.7 ;
    RECT 126.73 60.81 126.995 60.88 ;
    RECT 130.59 61.175 130.66 61.245 ;
    RECT 134.305 60.81 134.565 60.88 ;
    RECT 136.92 60.815 137.13 60.885 ;
    RECT 139.7 60.81 139.97 60.88 ;
    RECT 140.895 61.175 140.965 61.245 ;
    RECT 141.385 60.81 141.635 60.88 ;
    RECT 142.51 60.63 142.72 60.7 ;
    RECT 143.065 60.81 143.135 60.88 ;
    RECT 143.66 60.81 143.93 60.88 ;
    RECT 146.125 60.55 146.395 60.62 ;
    RECT 146.125 61.29 146.395 61.36 ;
    RECT 132.99 91.797 133.06 91.867 ;
    RECT 135.105 48.577 135.175 48.647 ;
    RECT 132.595 49.297 132.665 49.367 ;
    RECT 121.44 87.93 121.51 88.72 ;
    RECT 122.04 87.93 122.25 88.0 ;
    RECT 122.04 88.285 122.25 88.355 ;
    RECT 122.04 88.65 122.25 88.72 ;
    RECT 123.205 88.375 124.005 88.445 ;
    RECT 125.67 88.2 125.905 88.27 ;
    RECT 126.73 88.2 126.99 88.27 ;
    RECT 128.705 88.2 128.935 88.27 ;
    RECT 129.42 88.2 129.68 88.27 ;
    RECT 130.59 88.2 130.66 88.27 ;
    RECT 133.925 88.2 134.135 88.27 ;
    RECT 134.31 88.2 134.58 88.27 ;
    RECT 138.365 88.2 138.435 88.27 ;
    RECT 138.695 88.2 138.96 88.27 ;
    RECT 140.45 88.2 140.71 88.27 ;
    RECT 140.895 88.2 140.965 88.27 ;
    RECT 141.385 88.2 141.645 88.27 ;
    RECT 142.51 88.2 142.72 88.27 ;
    RECT 144.32 88.375 145.135 88.445 ;
    RECT 146.125 87.93 146.395 88.0 ;
    RECT 146.125 88.285 146.395 88.355 ;
    RECT 146.125 88.65 146.395 88.72 ;
    RECT 121.44 87.21 121.51 88.0 ;
    RECT 122.04 87.21 122.25 87.28 ;
    RECT 122.04 87.565 122.25 87.635 ;
    RECT 122.04 87.93 122.25 88.0 ;
    RECT 123.205 87.655 124.005 87.725 ;
    RECT 125.67 87.48 125.905 87.55 ;
    RECT 126.73 87.48 126.99 87.55 ;
    RECT 128.705 87.48 128.935 87.55 ;
    RECT 129.42 87.48 129.68 87.55 ;
    RECT 130.59 87.48 130.66 87.55 ;
    RECT 133.925 87.48 134.135 87.55 ;
    RECT 134.31 87.48 134.58 87.55 ;
    RECT 138.365 87.48 138.435 87.55 ;
    RECT 138.695 87.48 138.96 87.55 ;
    RECT 140.45 87.48 140.71 87.55 ;
    RECT 140.895 87.48 140.965 87.55 ;
    RECT 141.385 87.48 141.645 87.55 ;
    RECT 142.51 87.48 142.72 87.55 ;
    RECT 144.32 87.655 145.135 87.725 ;
    RECT 146.125 87.21 146.395 87.28 ;
    RECT 146.125 87.565 146.395 87.635 ;
    RECT 146.125 87.93 146.395 88.0 ;
    RECT 121.44 86.49 121.51 87.28 ;
    RECT 122.04 86.49 122.25 86.56 ;
    RECT 122.04 86.845 122.25 86.915 ;
    RECT 122.04 87.21 122.25 87.28 ;
    RECT 123.205 86.935 124.005 87.005 ;
    RECT 125.67 86.76 125.905 86.83 ;
    RECT 126.73 86.76 126.99 86.83 ;
    RECT 128.705 86.76 128.935 86.83 ;
    RECT 129.42 86.76 129.68 86.83 ;
    RECT 130.59 86.76 130.66 86.83 ;
    RECT 133.925 86.76 134.135 86.83 ;
    RECT 134.31 86.76 134.58 86.83 ;
    RECT 138.365 86.76 138.435 86.83 ;
    RECT 138.695 86.76 138.96 86.83 ;
    RECT 140.45 86.76 140.71 86.83 ;
    RECT 140.895 86.76 140.965 86.83 ;
    RECT 141.385 86.76 141.645 86.83 ;
    RECT 142.51 86.76 142.72 86.83 ;
    RECT 144.32 86.935 145.135 87.005 ;
    RECT 146.125 86.49 146.395 86.56 ;
    RECT 146.125 86.845 146.395 86.915 ;
    RECT 146.125 87.21 146.395 87.28 ;
    RECT 121.44 85.77 121.51 86.56 ;
    RECT 122.04 85.77 122.25 85.84 ;
    RECT 122.04 86.125 122.25 86.195 ;
    RECT 122.04 86.49 122.25 86.56 ;
    RECT 123.205 86.215 124.005 86.285 ;
    RECT 125.67 86.04 125.905 86.11 ;
    RECT 126.73 86.04 126.99 86.11 ;
    RECT 128.705 86.04 128.935 86.11 ;
    RECT 129.42 86.04 129.68 86.11 ;
    RECT 130.59 86.04 130.66 86.11 ;
    RECT 133.925 86.04 134.135 86.11 ;
    RECT 134.31 86.04 134.58 86.11 ;
    RECT 138.365 86.04 138.435 86.11 ;
    RECT 138.695 86.04 138.96 86.11 ;
    RECT 140.45 86.04 140.71 86.11 ;
    RECT 140.895 86.04 140.965 86.11 ;
    RECT 141.385 86.04 141.645 86.11 ;
    RECT 142.51 86.04 142.72 86.11 ;
    RECT 144.32 86.215 145.135 86.285 ;
    RECT 146.125 85.77 146.395 85.84 ;
    RECT 146.125 86.125 146.395 86.195 ;
    RECT 146.125 86.49 146.395 86.56 ;
    RECT 121.44 85.05 121.51 85.84 ;
    RECT 122.04 85.05 122.25 85.12 ;
    RECT 122.04 85.405 122.25 85.475 ;
    RECT 122.04 85.77 122.25 85.84 ;
    RECT 123.205 85.495 124.005 85.565 ;
    RECT 125.67 85.32 125.905 85.39 ;
    RECT 126.73 85.32 126.99 85.39 ;
    RECT 128.705 85.32 128.935 85.39 ;
    RECT 129.42 85.32 129.68 85.39 ;
    RECT 130.59 85.32 130.66 85.39 ;
    RECT 133.925 85.32 134.135 85.39 ;
    RECT 134.31 85.32 134.58 85.39 ;
    RECT 138.365 85.32 138.435 85.39 ;
    RECT 138.695 85.32 138.96 85.39 ;
    RECT 140.45 85.32 140.71 85.39 ;
    RECT 140.895 85.32 140.965 85.39 ;
    RECT 141.385 85.32 141.645 85.39 ;
    RECT 142.51 85.32 142.72 85.39 ;
    RECT 144.32 85.495 145.135 85.565 ;
    RECT 146.125 85.05 146.395 85.12 ;
    RECT 146.125 85.405 146.395 85.475 ;
    RECT 146.125 85.77 146.395 85.84 ;
    RECT 133.39 38.497 133.46 38.567 ;
    RECT 121.44 84.33 121.51 85.12 ;
    RECT 122.04 84.33 122.25 84.4 ;
    RECT 122.04 84.685 122.25 84.755 ;
    RECT 122.04 85.05 122.25 85.12 ;
    RECT 123.205 84.775 124.005 84.845 ;
    RECT 125.67 84.6 125.905 84.67 ;
    RECT 126.73 84.6 126.99 84.67 ;
    RECT 128.705 84.6 128.935 84.67 ;
    RECT 129.42 84.6 129.68 84.67 ;
    RECT 130.59 84.6 130.66 84.67 ;
    RECT 133.925 84.6 134.135 84.67 ;
    RECT 134.31 84.6 134.58 84.67 ;
    RECT 138.365 84.6 138.435 84.67 ;
    RECT 138.695 84.6 138.96 84.67 ;
    RECT 140.45 84.6 140.71 84.67 ;
    RECT 140.895 84.6 140.965 84.67 ;
    RECT 141.385 84.6 141.645 84.67 ;
    RECT 142.51 84.6 142.72 84.67 ;
    RECT 144.32 84.775 145.135 84.845 ;
    RECT 146.125 84.33 146.395 84.4 ;
    RECT 146.125 84.685 146.395 84.755 ;
    RECT 146.125 85.05 146.395 85.12 ;
    RECT 121.44 83.61 121.51 84.4 ;
    RECT 122.04 83.61 122.25 83.68 ;
    RECT 122.04 83.965 122.25 84.035 ;
    RECT 122.04 84.33 122.25 84.4 ;
    RECT 123.205 84.055 124.005 84.125 ;
    RECT 125.67 83.88 125.905 83.95 ;
    RECT 126.73 83.88 126.99 83.95 ;
    RECT 128.705 83.88 128.935 83.95 ;
    RECT 129.42 83.88 129.68 83.95 ;
    RECT 130.59 83.88 130.66 83.95 ;
    RECT 133.925 83.88 134.135 83.95 ;
    RECT 134.31 83.88 134.58 83.95 ;
    RECT 138.365 83.88 138.435 83.95 ;
    RECT 138.695 83.88 138.96 83.95 ;
    RECT 140.45 83.88 140.71 83.95 ;
    RECT 140.895 83.88 140.965 83.95 ;
    RECT 141.385 83.88 141.645 83.95 ;
    RECT 142.51 83.88 142.72 83.95 ;
    RECT 144.32 84.055 145.135 84.125 ;
    RECT 146.125 83.61 146.395 83.68 ;
    RECT 146.125 83.965 146.395 84.035 ;
    RECT 146.125 84.33 146.395 84.4 ;
    RECT 121.44 82.89 121.51 83.68 ;
    RECT 122.04 82.89 122.25 82.96 ;
    RECT 122.04 83.245 122.25 83.315 ;
    RECT 122.04 83.61 122.25 83.68 ;
    RECT 123.205 83.335 124.005 83.405 ;
    RECT 125.67 83.16 125.905 83.23 ;
    RECT 126.73 83.16 126.99 83.23 ;
    RECT 128.705 83.16 128.935 83.23 ;
    RECT 129.42 83.16 129.68 83.23 ;
    RECT 130.59 83.16 130.66 83.23 ;
    RECT 133.925 83.16 134.135 83.23 ;
    RECT 134.31 83.16 134.58 83.23 ;
    RECT 138.365 83.16 138.435 83.23 ;
    RECT 138.695 83.16 138.96 83.23 ;
    RECT 140.45 83.16 140.71 83.23 ;
    RECT 140.895 83.16 140.965 83.23 ;
    RECT 141.385 83.16 141.645 83.23 ;
    RECT 142.51 83.16 142.72 83.23 ;
    RECT 144.32 83.335 145.135 83.405 ;
    RECT 146.125 82.89 146.395 82.96 ;
    RECT 146.125 83.245 146.395 83.315 ;
    RECT 146.125 83.61 146.395 83.68 ;
    RECT 121.44 82.17 121.51 82.96 ;
    RECT 122.04 82.17 122.25 82.24 ;
    RECT 122.04 82.525 122.25 82.595 ;
    RECT 122.04 82.89 122.25 82.96 ;
    RECT 123.205 82.615 124.005 82.685 ;
    RECT 125.67 82.44 125.905 82.51 ;
    RECT 126.73 82.44 126.99 82.51 ;
    RECT 128.705 82.44 128.935 82.51 ;
    RECT 129.42 82.44 129.68 82.51 ;
    RECT 130.59 82.44 130.66 82.51 ;
    RECT 133.925 82.44 134.135 82.51 ;
    RECT 134.31 82.44 134.58 82.51 ;
    RECT 138.365 82.44 138.435 82.51 ;
    RECT 138.695 82.44 138.96 82.51 ;
    RECT 140.45 82.44 140.71 82.51 ;
    RECT 140.895 82.44 140.965 82.51 ;
    RECT 141.385 82.44 141.645 82.51 ;
    RECT 142.51 82.44 142.72 82.51 ;
    RECT 144.32 82.615 145.135 82.685 ;
    RECT 146.125 82.17 146.395 82.24 ;
    RECT 146.125 82.525 146.395 82.595 ;
    RECT 146.125 82.89 146.395 82.96 ;
    RECT 121.44 81.45 121.51 82.24 ;
    RECT 122.04 81.45 122.25 81.52 ;
    RECT 122.04 81.805 122.25 81.875 ;
    RECT 122.04 82.17 122.25 82.24 ;
    RECT 123.205 81.895 124.005 81.965 ;
    RECT 125.67 81.72 125.905 81.79 ;
    RECT 126.73 81.72 126.99 81.79 ;
    RECT 128.705 81.72 128.935 81.79 ;
    RECT 129.42 81.72 129.68 81.79 ;
    RECT 130.59 81.72 130.66 81.79 ;
    RECT 133.925 81.72 134.135 81.79 ;
    RECT 134.31 81.72 134.58 81.79 ;
    RECT 138.365 81.72 138.435 81.79 ;
    RECT 138.695 81.72 138.96 81.79 ;
    RECT 140.45 81.72 140.71 81.79 ;
    RECT 140.895 81.72 140.965 81.79 ;
    RECT 141.385 81.72 141.645 81.79 ;
    RECT 142.51 81.72 142.72 81.79 ;
    RECT 144.32 81.895 145.135 81.965 ;
    RECT 146.125 81.45 146.395 81.52 ;
    RECT 146.125 81.805 146.395 81.875 ;
    RECT 146.125 82.17 146.395 82.24 ;
    RECT 145.485 43.63 145.695 43.7 ;
    RECT 139.73 43.54 139.94 43.61 ;
    RECT 121.44 80.73 121.51 81.52 ;
    RECT 122.04 80.73 122.25 80.8 ;
    RECT 122.04 81.085 122.25 81.155 ;
    RECT 122.04 81.45 122.25 81.52 ;
    RECT 123.205 81.175 124.005 81.245 ;
    RECT 125.67 81.0 125.905 81.07 ;
    RECT 126.73 81.0 126.99 81.07 ;
    RECT 128.705 81.0 128.935 81.07 ;
    RECT 129.42 81.0 129.68 81.07 ;
    RECT 130.59 81.0 130.66 81.07 ;
    RECT 133.925 81.0 134.135 81.07 ;
    RECT 134.31 81.0 134.58 81.07 ;
    RECT 138.365 81.0 138.435 81.07 ;
    RECT 138.695 81.0 138.96 81.07 ;
    RECT 140.45 81.0 140.71 81.07 ;
    RECT 140.895 81.0 140.965 81.07 ;
    RECT 141.385 81.0 141.645 81.07 ;
    RECT 142.51 81.0 142.72 81.07 ;
    RECT 144.32 81.175 145.135 81.245 ;
    RECT 146.125 80.73 146.395 80.8 ;
    RECT 146.125 81.085 146.395 81.155 ;
    RECT 146.125 81.45 146.395 81.52 ;
    RECT 121.44 80.01 121.51 80.8 ;
    RECT 122.04 80.01 122.25 80.08 ;
    RECT 122.04 80.365 122.25 80.435 ;
    RECT 122.04 80.73 122.25 80.8 ;
    RECT 123.205 80.455 124.005 80.525 ;
    RECT 125.67 80.28 125.905 80.35 ;
    RECT 126.73 80.28 126.99 80.35 ;
    RECT 128.705 80.28 128.935 80.35 ;
    RECT 129.42 80.28 129.68 80.35 ;
    RECT 130.59 80.28 130.66 80.35 ;
    RECT 133.925 80.28 134.135 80.35 ;
    RECT 134.31 80.28 134.58 80.35 ;
    RECT 138.365 80.28 138.435 80.35 ;
    RECT 138.695 80.28 138.96 80.35 ;
    RECT 140.45 80.28 140.71 80.35 ;
    RECT 140.895 80.28 140.965 80.35 ;
    RECT 141.385 80.28 141.645 80.35 ;
    RECT 142.51 80.28 142.72 80.35 ;
    RECT 144.32 80.455 145.135 80.525 ;
    RECT 146.125 80.01 146.395 80.08 ;
    RECT 146.125 80.365 146.395 80.435 ;
    RECT 146.125 80.73 146.395 80.8 ;
    RECT 121.44 79.29 121.51 80.08 ;
    RECT 122.04 79.29 122.25 79.36 ;
    RECT 122.04 79.645 122.25 79.715 ;
    RECT 122.04 80.01 122.25 80.08 ;
    RECT 123.205 79.735 124.005 79.805 ;
    RECT 125.67 79.56 125.905 79.63 ;
    RECT 126.73 79.56 126.99 79.63 ;
    RECT 128.705 79.56 128.935 79.63 ;
    RECT 129.42 79.56 129.68 79.63 ;
    RECT 130.59 79.56 130.66 79.63 ;
    RECT 133.925 79.56 134.135 79.63 ;
    RECT 134.31 79.56 134.58 79.63 ;
    RECT 138.365 79.56 138.435 79.63 ;
    RECT 138.695 79.56 138.96 79.63 ;
    RECT 140.45 79.56 140.71 79.63 ;
    RECT 140.895 79.56 140.965 79.63 ;
    RECT 141.385 79.56 141.645 79.63 ;
    RECT 142.51 79.56 142.72 79.63 ;
    RECT 144.32 79.735 145.135 79.805 ;
    RECT 146.125 79.29 146.395 79.36 ;
    RECT 146.125 79.645 146.395 79.715 ;
    RECT 146.125 80.01 146.395 80.08 ;
    RECT 121.44 78.57 121.51 79.36 ;
    RECT 122.04 78.57 122.25 78.64 ;
    RECT 122.04 78.925 122.25 78.995 ;
    RECT 122.04 79.29 122.25 79.36 ;
    RECT 123.205 79.015 124.005 79.085 ;
    RECT 125.67 78.84 125.905 78.91 ;
    RECT 126.73 78.84 126.99 78.91 ;
    RECT 128.705 78.84 128.935 78.91 ;
    RECT 129.42 78.84 129.68 78.91 ;
    RECT 130.59 78.84 130.66 78.91 ;
    RECT 133.925 78.84 134.135 78.91 ;
    RECT 134.31 78.84 134.58 78.91 ;
    RECT 138.365 78.84 138.435 78.91 ;
    RECT 138.695 78.84 138.96 78.91 ;
    RECT 140.45 78.84 140.71 78.91 ;
    RECT 140.895 78.84 140.965 78.91 ;
    RECT 141.385 78.84 141.645 78.91 ;
    RECT 142.51 78.84 142.72 78.91 ;
    RECT 144.32 79.015 145.135 79.085 ;
    RECT 146.125 78.57 146.395 78.64 ;
    RECT 146.125 78.925 146.395 78.995 ;
    RECT 146.125 79.29 146.395 79.36 ;
    RECT 121.44 77.85 121.51 78.64 ;
    RECT 122.04 77.85 122.25 77.92 ;
    RECT 122.04 78.205 122.25 78.275 ;
    RECT 122.04 78.57 122.25 78.64 ;
    RECT 123.205 78.295 124.005 78.365 ;
    RECT 125.67 78.12 125.905 78.19 ;
    RECT 126.73 78.12 126.99 78.19 ;
    RECT 128.705 78.12 128.935 78.19 ;
    RECT 129.42 78.12 129.68 78.19 ;
    RECT 130.59 78.12 130.66 78.19 ;
    RECT 133.925 78.12 134.135 78.19 ;
    RECT 134.31 78.12 134.58 78.19 ;
    RECT 138.365 78.12 138.435 78.19 ;
    RECT 138.695 78.12 138.96 78.19 ;
    RECT 140.45 78.12 140.71 78.19 ;
    RECT 140.895 78.12 140.965 78.19 ;
    RECT 141.385 78.12 141.645 78.19 ;
    RECT 142.51 78.12 142.72 78.19 ;
    RECT 144.32 78.295 145.135 78.365 ;
    RECT 146.125 77.85 146.395 77.92 ;
    RECT 146.125 78.205 146.395 78.275 ;
    RECT 146.125 78.57 146.395 78.64 ;
    RECT 121.44 77.13 121.51 77.92 ;
    RECT 122.04 77.13 122.25 77.2 ;
    RECT 122.04 77.485 122.25 77.555 ;
    RECT 122.04 77.85 122.25 77.92 ;
    RECT 123.205 77.575 124.005 77.645 ;
    RECT 125.67 77.4 125.905 77.47 ;
    RECT 126.73 77.4 126.99 77.47 ;
    RECT 128.705 77.4 128.935 77.47 ;
    RECT 129.42 77.4 129.68 77.47 ;
    RECT 130.59 77.4 130.66 77.47 ;
    RECT 133.925 77.4 134.135 77.47 ;
    RECT 134.31 77.4 134.58 77.47 ;
    RECT 138.365 77.4 138.435 77.47 ;
    RECT 138.695 77.4 138.96 77.47 ;
    RECT 140.45 77.4 140.71 77.47 ;
    RECT 140.895 77.4 140.965 77.47 ;
    RECT 141.385 77.4 141.645 77.47 ;
    RECT 142.51 77.4 142.72 77.47 ;
    RECT 144.32 77.575 145.135 77.645 ;
    RECT 146.125 77.13 146.395 77.2 ;
    RECT 146.125 77.485 146.395 77.555 ;
    RECT 146.125 77.85 146.395 77.92 ;
    RECT 121.44 76.41 121.51 77.2 ;
    RECT 122.04 76.41 122.25 76.48 ;
    RECT 122.04 76.765 122.25 76.835 ;
    RECT 122.04 77.13 122.25 77.2 ;
    RECT 123.205 76.855 124.005 76.925 ;
    RECT 125.67 76.68 125.905 76.75 ;
    RECT 126.73 76.68 126.99 76.75 ;
    RECT 128.705 76.68 128.935 76.75 ;
    RECT 129.42 76.68 129.68 76.75 ;
    RECT 130.59 76.68 130.66 76.75 ;
    RECT 133.925 76.68 134.135 76.75 ;
    RECT 134.31 76.68 134.58 76.75 ;
    RECT 138.365 76.68 138.435 76.75 ;
    RECT 138.695 76.68 138.96 76.75 ;
    RECT 140.45 76.68 140.71 76.75 ;
    RECT 140.895 76.68 140.965 76.75 ;
    RECT 141.385 76.68 141.645 76.75 ;
    RECT 142.51 76.68 142.72 76.75 ;
    RECT 144.32 76.855 145.135 76.925 ;
    RECT 146.125 76.41 146.395 76.48 ;
    RECT 146.125 76.765 146.395 76.835 ;
    RECT 146.125 77.13 146.395 77.2 ;
    RECT 121.44 75.69 121.51 76.48 ;
    RECT 122.04 75.69 122.25 75.76 ;
    RECT 122.04 76.045 122.25 76.115 ;
    RECT 122.04 76.41 122.25 76.48 ;
    RECT 123.205 76.135 124.005 76.205 ;
    RECT 125.67 75.96 125.905 76.03 ;
    RECT 126.73 75.96 126.99 76.03 ;
    RECT 128.705 75.96 128.935 76.03 ;
    RECT 129.42 75.96 129.68 76.03 ;
    RECT 130.59 75.96 130.66 76.03 ;
    RECT 133.925 75.96 134.135 76.03 ;
    RECT 134.31 75.96 134.58 76.03 ;
    RECT 138.365 75.96 138.435 76.03 ;
    RECT 138.695 75.96 138.96 76.03 ;
    RECT 140.45 75.96 140.71 76.03 ;
    RECT 140.895 75.96 140.965 76.03 ;
    RECT 141.385 75.96 141.645 76.03 ;
    RECT 142.51 75.96 142.72 76.03 ;
    RECT 144.32 76.135 145.135 76.205 ;
    RECT 146.125 75.69 146.395 75.76 ;
    RECT 146.125 76.045 146.395 76.115 ;
    RECT 146.125 76.41 146.395 76.48 ;
    RECT 121.44 74.97 121.51 75.76 ;
    RECT 122.04 74.97 122.25 75.04 ;
    RECT 122.04 75.325 122.25 75.395 ;
    RECT 122.04 75.69 122.25 75.76 ;
    RECT 123.205 75.415 124.005 75.485 ;
    RECT 125.67 75.24 125.905 75.31 ;
    RECT 126.73 75.24 126.99 75.31 ;
    RECT 128.705 75.24 128.935 75.31 ;
    RECT 129.42 75.24 129.68 75.31 ;
    RECT 130.59 75.24 130.66 75.31 ;
    RECT 133.925 75.24 134.135 75.31 ;
    RECT 134.31 75.24 134.58 75.31 ;
    RECT 138.365 75.24 138.435 75.31 ;
    RECT 138.695 75.24 138.96 75.31 ;
    RECT 140.45 75.24 140.71 75.31 ;
    RECT 140.895 75.24 140.965 75.31 ;
    RECT 141.385 75.24 141.645 75.31 ;
    RECT 142.51 75.24 142.72 75.31 ;
    RECT 144.32 75.415 145.135 75.485 ;
    RECT 146.125 74.97 146.395 75.04 ;
    RECT 146.125 75.325 146.395 75.395 ;
    RECT 146.125 75.69 146.395 75.76 ;
    RECT 121.44 74.25 121.51 75.04 ;
    RECT 122.04 74.25 122.25 74.32 ;
    RECT 122.04 74.605 122.25 74.675 ;
    RECT 122.04 74.97 122.25 75.04 ;
    RECT 123.205 74.695 124.005 74.765 ;
    RECT 125.67 74.52 125.905 74.59 ;
    RECT 126.73 74.52 126.99 74.59 ;
    RECT 128.705 74.52 128.935 74.59 ;
    RECT 129.42 74.52 129.68 74.59 ;
    RECT 130.59 74.52 130.66 74.59 ;
    RECT 133.925 74.52 134.135 74.59 ;
    RECT 134.31 74.52 134.58 74.59 ;
    RECT 138.365 74.52 138.435 74.59 ;
    RECT 138.695 74.52 138.96 74.59 ;
    RECT 140.45 74.52 140.71 74.59 ;
    RECT 140.895 74.52 140.965 74.59 ;
    RECT 141.385 74.52 141.645 74.59 ;
    RECT 142.51 74.52 142.72 74.59 ;
    RECT 144.32 74.695 145.135 74.765 ;
    RECT 146.125 74.25 146.395 74.32 ;
    RECT 146.125 74.605 146.395 74.675 ;
    RECT 146.125 74.97 146.395 75.04 ;
    RECT 145.485 94.77 145.695 94.84 ;
    RECT 127.69 43.537 127.9 43.607 ;
    RECT 139.73 94.68 139.94 94.75 ;
    RECT 122.63 43.63 122.84 43.7 ;
    RECT 121.44 73.53 121.51 74.32 ;
    RECT 122.04 73.53 122.25 73.6 ;
    RECT 122.04 73.885 122.25 73.955 ;
    RECT 122.04 74.25 122.25 74.32 ;
    RECT 123.205 73.975 124.005 74.045 ;
    RECT 125.67 73.8 125.905 73.87 ;
    RECT 126.73 73.8 126.99 73.87 ;
    RECT 128.705 73.8 128.935 73.87 ;
    RECT 129.42 73.8 129.68 73.87 ;
    RECT 130.59 73.8 130.66 73.87 ;
    RECT 133.925 73.8 134.135 73.87 ;
    RECT 134.31 73.8 134.58 73.87 ;
    RECT 138.365 73.8 138.435 73.87 ;
    RECT 138.695 73.8 138.96 73.87 ;
    RECT 140.45 73.8 140.71 73.87 ;
    RECT 140.895 73.8 140.965 73.87 ;
    RECT 141.385 73.8 141.645 73.87 ;
    RECT 142.51 73.8 142.72 73.87 ;
    RECT 144.32 73.975 145.135 74.045 ;
    RECT 146.125 73.53 146.395 73.6 ;
    RECT 146.125 73.885 146.395 73.955 ;
    RECT 146.125 74.25 146.395 74.32 ;
    RECT 121.44 72.81 121.51 73.6 ;
    RECT 122.04 72.81 122.25 72.88 ;
    RECT 122.04 73.165 122.25 73.235 ;
    RECT 122.04 73.53 122.25 73.6 ;
    RECT 123.205 73.255 124.005 73.325 ;
    RECT 125.67 73.08 125.905 73.15 ;
    RECT 126.73 73.08 126.99 73.15 ;
    RECT 128.705 73.08 128.935 73.15 ;
    RECT 129.42 73.08 129.68 73.15 ;
    RECT 130.59 73.08 130.66 73.15 ;
    RECT 133.925 73.08 134.135 73.15 ;
    RECT 134.31 73.08 134.58 73.15 ;
    RECT 138.365 73.08 138.435 73.15 ;
    RECT 138.695 73.08 138.96 73.15 ;
    RECT 140.45 73.08 140.71 73.15 ;
    RECT 140.895 73.08 140.965 73.15 ;
    RECT 141.385 73.08 141.645 73.15 ;
    RECT 142.51 73.08 142.72 73.15 ;
    RECT 144.32 73.255 145.135 73.325 ;
    RECT 146.125 72.81 146.395 72.88 ;
    RECT 146.125 73.165 146.395 73.235 ;
    RECT 146.125 73.53 146.395 73.6 ;
    RECT 121.44 72.09 121.51 72.88 ;
    RECT 122.04 72.09 122.25 72.16 ;
    RECT 122.04 72.445 122.25 72.515 ;
    RECT 122.04 72.81 122.25 72.88 ;
    RECT 123.205 72.535 124.005 72.605 ;
    RECT 125.67 72.36 125.905 72.43 ;
    RECT 126.73 72.36 126.99 72.43 ;
    RECT 128.705 72.36 128.935 72.43 ;
    RECT 129.42 72.36 129.68 72.43 ;
    RECT 130.59 72.36 130.66 72.43 ;
    RECT 133.925 72.36 134.135 72.43 ;
    RECT 134.31 72.36 134.58 72.43 ;
    RECT 138.365 72.36 138.435 72.43 ;
    RECT 138.695 72.36 138.96 72.43 ;
    RECT 140.45 72.36 140.71 72.43 ;
    RECT 140.895 72.36 140.965 72.43 ;
    RECT 141.385 72.36 141.645 72.43 ;
    RECT 142.51 72.36 142.72 72.43 ;
    RECT 144.32 72.535 145.135 72.605 ;
    RECT 146.125 72.09 146.395 72.16 ;
    RECT 146.125 72.445 146.395 72.515 ;
    RECT 146.125 72.81 146.395 72.88 ;
    RECT 121.44 71.37 121.51 72.16 ;
    RECT 122.04 71.37 122.25 71.44 ;
    RECT 122.04 71.725 122.25 71.795 ;
    RECT 122.04 72.09 122.25 72.16 ;
    RECT 123.205 71.815 124.005 71.885 ;
    RECT 125.67 71.64 125.905 71.71 ;
    RECT 126.73 71.64 126.99 71.71 ;
    RECT 128.705 71.64 128.935 71.71 ;
    RECT 129.42 71.64 129.68 71.71 ;
    RECT 130.59 71.64 130.66 71.71 ;
    RECT 133.925 71.64 134.135 71.71 ;
    RECT 134.31 71.64 134.58 71.71 ;
    RECT 138.365 71.64 138.435 71.71 ;
    RECT 138.695 71.64 138.96 71.71 ;
    RECT 140.45 71.64 140.71 71.71 ;
    RECT 140.895 71.64 140.965 71.71 ;
    RECT 141.385 71.64 141.645 71.71 ;
    RECT 142.51 71.64 142.72 71.71 ;
    RECT 144.32 71.815 145.135 71.885 ;
    RECT 146.125 71.37 146.395 71.44 ;
    RECT 146.125 71.725 146.395 71.795 ;
    RECT 146.125 72.09 146.395 72.16 ;
    RECT 122.63 53.71 122.84 53.78 ;
    RECT 121.44 70.65 121.51 71.44 ;
    RECT 122.04 70.65 122.25 70.72 ;
    RECT 122.04 71.005 122.25 71.075 ;
    RECT 122.04 71.37 122.25 71.44 ;
    RECT 123.205 71.095 124.005 71.165 ;
    RECT 125.67 70.92 125.905 70.99 ;
    RECT 126.73 70.92 126.99 70.99 ;
    RECT 128.705 70.92 128.935 70.99 ;
    RECT 129.42 70.92 129.68 70.99 ;
    RECT 130.59 70.92 130.66 70.99 ;
    RECT 133.925 70.92 134.135 70.99 ;
    RECT 134.31 70.92 134.58 70.99 ;
    RECT 138.365 70.92 138.435 70.99 ;
    RECT 138.695 70.92 138.96 70.99 ;
    RECT 140.45 70.92 140.71 70.99 ;
    RECT 140.895 70.92 140.965 70.99 ;
    RECT 141.385 70.92 141.645 70.99 ;
    RECT 142.51 70.92 142.72 70.99 ;
    RECT 144.32 71.095 145.135 71.165 ;
    RECT 146.125 70.65 146.395 70.72 ;
    RECT 146.125 71.005 146.395 71.075 ;
    RECT 146.125 71.37 146.395 71.44 ;
    RECT 121.44 69.93 121.51 70.72 ;
    RECT 122.04 69.93 122.25 70.0 ;
    RECT 122.04 70.285 122.25 70.355 ;
    RECT 122.04 70.65 122.25 70.72 ;
    RECT 123.205 70.375 124.005 70.445 ;
    RECT 125.67 70.2 125.905 70.27 ;
    RECT 126.73 70.2 126.99 70.27 ;
    RECT 128.705 70.2 128.935 70.27 ;
    RECT 129.42 70.2 129.68 70.27 ;
    RECT 130.59 70.2 130.66 70.27 ;
    RECT 133.925 70.2 134.135 70.27 ;
    RECT 134.31 70.2 134.58 70.27 ;
    RECT 138.365 70.2 138.435 70.27 ;
    RECT 138.695 70.2 138.96 70.27 ;
    RECT 140.45 70.2 140.71 70.27 ;
    RECT 140.895 70.2 140.965 70.27 ;
    RECT 141.385 70.2 141.645 70.27 ;
    RECT 142.51 70.2 142.72 70.27 ;
    RECT 144.32 70.375 145.135 70.445 ;
    RECT 146.125 69.93 146.395 70.0 ;
    RECT 146.125 70.285 146.395 70.355 ;
    RECT 146.125 70.65 146.395 70.72 ;
    RECT 134.34 29.85 134.55 29.92 ;
    RECT 121.44 69.21 121.51 70.0 ;
    RECT 122.04 69.21 122.25 69.28 ;
    RECT 122.04 69.565 122.25 69.635 ;
    RECT 122.04 69.93 122.25 70.0 ;
    RECT 123.205 69.655 124.005 69.725 ;
    RECT 125.67 69.48 125.905 69.55 ;
    RECT 126.73 69.48 126.99 69.55 ;
    RECT 128.705 69.48 128.935 69.55 ;
    RECT 129.42 69.48 129.68 69.55 ;
    RECT 130.59 69.48 130.66 69.55 ;
    RECT 133.925 69.48 134.135 69.55 ;
    RECT 134.31 69.48 134.58 69.55 ;
    RECT 138.365 69.48 138.435 69.55 ;
    RECT 138.695 69.48 138.96 69.55 ;
    RECT 140.45 69.48 140.71 69.55 ;
    RECT 140.895 69.48 140.965 69.55 ;
    RECT 141.385 69.48 141.645 69.55 ;
    RECT 142.51 69.48 142.72 69.55 ;
    RECT 144.32 69.655 145.135 69.725 ;
    RECT 146.125 69.21 146.395 69.28 ;
    RECT 146.125 69.565 146.395 69.635 ;
    RECT 146.125 69.93 146.395 70.0 ;
    RECT 127.69 94.677 127.9 94.747 ;
    RECT 134.34 29.13 134.55 29.2 ;
    RECT 121.44 68.49 121.51 69.28 ;
    RECT 122.04 68.49 122.25 68.56 ;
    RECT 122.04 68.845 122.25 68.915 ;
    RECT 122.04 69.21 122.25 69.28 ;
    RECT 123.205 68.935 124.005 69.005 ;
    RECT 125.67 68.76 125.905 68.83 ;
    RECT 126.73 68.76 126.99 68.83 ;
    RECT 128.705 68.76 128.935 68.83 ;
    RECT 129.42 68.76 129.68 68.83 ;
    RECT 130.59 68.76 130.66 68.83 ;
    RECT 133.925 68.76 134.135 68.83 ;
    RECT 134.31 68.76 134.58 68.83 ;
    RECT 138.365 68.76 138.435 68.83 ;
    RECT 138.695 68.76 138.96 68.83 ;
    RECT 140.45 68.76 140.71 68.83 ;
    RECT 140.895 68.76 140.965 68.83 ;
    RECT 141.385 68.76 141.645 68.83 ;
    RECT 142.51 68.76 142.72 68.83 ;
    RECT 144.32 68.935 145.135 69.005 ;
    RECT 146.125 68.49 146.395 68.56 ;
    RECT 146.125 68.845 146.395 68.915 ;
    RECT 146.125 69.21 146.395 69.28 ;
    RECT 134.34 26.97 134.55 27.04 ;
    RECT 121.44 67.77 121.51 68.56 ;
    RECT 122.04 67.77 122.25 67.84 ;
    RECT 122.04 68.125 122.25 68.195 ;
    RECT 122.04 68.49 122.25 68.56 ;
    RECT 123.205 68.215 124.005 68.285 ;
    RECT 125.67 68.04 125.905 68.11 ;
    RECT 126.73 68.04 126.99 68.11 ;
    RECT 128.705 68.04 128.935 68.11 ;
    RECT 129.42 68.04 129.68 68.11 ;
    RECT 130.59 68.04 130.66 68.11 ;
    RECT 133.925 68.04 134.135 68.11 ;
    RECT 134.31 68.04 134.58 68.11 ;
    RECT 138.365 68.04 138.435 68.11 ;
    RECT 138.695 68.04 138.96 68.11 ;
    RECT 140.45 68.04 140.71 68.11 ;
    RECT 140.895 68.04 140.965 68.11 ;
    RECT 141.385 68.04 141.645 68.11 ;
    RECT 142.51 68.04 142.72 68.11 ;
    RECT 144.32 68.215 145.135 68.285 ;
    RECT 146.125 67.77 146.395 67.84 ;
    RECT 146.125 68.125 146.395 68.195 ;
    RECT 146.125 68.49 146.395 68.56 ;
    RECT 131.795 29.85 131.865 29.92 ;
    RECT 121.44 67.05 121.51 67.84 ;
    RECT 122.04 67.05 122.25 67.12 ;
    RECT 122.04 67.405 122.25 67.475 ;
    RECT 122.04 67.77 122.25 67.84 ;
    RECT 123.205 67.495 124.005 67.565 ;
    RECT 125.67 67.32 125.905 67.39 ;
    RECT 126.73 67.32 126.99 67.39 ;
    RECT 128.705 67.32 128.935 67.39 ;
    RECT 129.42 67.32 129.68 67.39 ;
    RECT 130.59 67.32 130.66 67.39 ;
    RECT 133.925 67.32 134.135 67.39 ;
    RECT 134.31 67.32 134.58 67.39 ;
    RECT 138.365 67.32 138.435 67.39 ;
    RECT 138.695 67.32 138.96 67.39 ;
    RECT 140.45 67.32 140.71 67.39 ;
    RECT 140.895 67.32 140.965 67.39 ;
    RECT 141.385 67.32 141.645 67.39 ;
    RECT 142.51 67.32 142.72 67.39 ;
    RECT 144.32 67.495 145.135 67.565 ;
    RECT 146.125 67.05 146.395 67.12 ;
    RECT 146.125 67.405 146.395 67.475 ;
    RECT 146.125 67.77 146.395 67.84 ;
    RECT 131.795 29.13 131.865 29.2 ;
    RECT 122.63 94.77 122.84 94.84 ;
    RECT 131.795 26.97 131.865 27.04 ;
    RECT 131.0 37.057 131.21 37.127 ;
    RECT 131.0 17.602 131.21 17.672 ;
    RECT 145.485 90.45 145.695 90.52 ;
    RECT 139.73 90.36 139.94 90.43 ;
    RECT 127.69 90.357 127.9 90.427 ;
    RECT 121.44 66.33 121.51 67.12 ;
    RECT 122.04 66.33 122.25 66.4 ;
    RECT 122.04 66.685 122.25 66.755 ;
    RECT 122.04 67.05 122.25 67.12 ;
    RECT 123.205 66.775 124.005 66.845 ;
    RECT 125.67 66.6 125.905 66.67 ;
    RECT 126.73 66.6 126.99 66.67 ;
    RECT 128.705 66.6 128.935 66.67 ;
    RECT 129.42 66.6 129.68 66.67 ;
    RECT 130.59 66.6 130.66 66.67 ;
    RECT 133.925 66.6 134.135 66.67 ;
    RECT 134.31 66.6 134.58 66.67 ;
    RECT 138.365 66.6 138.435 66.67 ;
    RECT 138.695 66.6 138.96 66.67 ;
    RECT 140.45 66.6 140.71 66.67 ;
    RECT 140.895 66.6 140.965 66.67 ;
    RECT 141.385 66.6 141.645 66.67 ;
    RECT 142.51 66.6 142.72 66.67 ;
    RECT 144.32 66.775 145.135 66.845 ;
    RECT 146.125 66.33 146.395 66.4 ;
    RECT 146.125 66.685 146.395 66.755 ;
    RECT 146.125 67.05 146.395 67.12 ;
    RECT 121.44 65.61 121.51 66.4 ;
    RECT 122.04 65.61 122.25 65.68 ;
    RECT 122.04 65.965 122.25 66.035 ;
    RECT 122.04 66.33 122.25 66.4 ;
    RECT 123.205 66.055 124.005 66.125 ;
    RECT 125.67 65.88 125.905 65.95 ;
    RECT 126.73 65.88 126.99 65.95 ;
    RECT 128.705 65.88 128.935 65.95 ;
    RECT 129.42 65.88 129.68 65.95 ;
    RECT 130.59 65.88 130.66 65.95 ;
    RECT 133.925 65.88 134.135 65.95 ;
    RECT 134.31 65.88 134.58 65.95 ;
    RECT 138.365 65.88 138.435 65.95 ;
    RECT 138.695 65.88 138.96 65.95 ;
    RECT 140.45 65.88 140.71 65.95 ;
    RECT 140.895 65.88 140.965 65.95 ;
    RECT 141.385 65.88 141.645 65.95 ;
    RECT 142.51 65.88 142.72 65.95 ;
    RECT 144.32 66.055 145.135 66.125 ;
    RECT 146.125 65.61 146.395 65.68 ;
    RECT 146.125 65.965 146.395 66.035 ;
    RECT 146.125 66.33 146.395 66.4 ;
    RECT 121.44 64.89 121.51 65.68 ;
    RECT 122.04 64.89 122.25 64.96 ;
    RECT 122.04 65.245 122.25 65.315 ;
    RECT 122.04 65.61 122.25 65.68 ;
    RECT 123.205 65.335 124.005 65.405 ;
    RECT 125.67 65.16 125.905 65.23 ;
    RECT 126.73 65.16 126.99 65.23 ;
    RECT 128.705 65.16 128.935 65.23 ;
    RECT 129.42 65.16 129.68 65.23 ;
    RECT 130.59 65.16 130.66 65.23 ;
    RECT 133.925 65.16 134.135 65.23 ;
    RECT 134.31 65.16 134.58 65.23 ;
    RECT 138.365 65.16 138.435 65.23 ;
    RECT 138.695 65.16 138.96 65.23 ;
    RECT 140.45 65.16 140.71 65.23 ;
    RECT 140.895 65.16 140.965 65.23 ;
    RECT 141.385 65.16 141.645 65.23 ;
    RECT 142.51 65.16 142.72 65.23 ;
    RECT 144.32 65.335 145.135 65.405 ;
    RECT 146.125 64.89 146.395 64.96 ;
    RECT 146.125 65.245 146.395 65.315 ;
    RECT 146.125 65.61 146.395 65.68 ;
    RECT 121.44 64.17 121.51 64.96 ;
    RECT 122.04 64.17 122.25 64.24 ;
    RECT 122.04 64.525 122.25 64.595 ;
    RECT 122.04 64.89 122.25 64.96 ;
    RECT 123.205 64.615 124.005 64.685 ;
    RECT 125.67 64.44 125.905 64.51 ;
    RECT 126.73 64.44 126.99 64.51 ;
    RECT 128.705 64.44 128.935 64.51 ;
    RECT 129.42 64.44 129.68 64.51 ;
    RECT 130.59 64.44 130.66 64.51 ;
    RECT 133.925 64.44 134.135 64.51 ;
    RECT 134.31 64.44 134.58 64.51 ;
    RECT 138.365 64.44 138.435 64.51 ;
    RECT 138.695 64.44 138.96 64.51 ;
    RECT 140.45 64.44 140.71 64.51 ;
    RECT 140.895 64.44 140.965 64.51 ;
    RECT 141.385 64.44 141.645 64.51 ;
    RECT 142.51 64.44 142.72 64.51 ;
    RECT 144.32 64.615 145.135 64.685 ;
    RECT 146.125 64.17 146.395 64.24 ;
    RECT 146.125 64.525 146.395 64.595 ;
    RECT 146.125 64.89 146.395 64.96 ;
    RECT 135.5 85.317 135.57 85.387 ;
    RECT 121.44 63.45 121.51 64.24 ;
    RECT 122.04 63.45 122.25 63.52 ;
    RECT 122.04 63.805 122.25 63.875 ;
    RECT 122.04 64.17 122.25 64.24 ;
    RECT 123.205 63.895 124.005 63.965 ;
    RECT 125.67 63.72 125.905 63.79 ;
    RECT 126.73 63.72 126.99 63.79 ;
    RECT 128.705 63.72 128.935 63.79 ;
    RECT 129.42 63.72 129.68 63.79 ;
    RECT 130.59 63.72 130.66 63.79 ;
    RECT 133.925 63.72 134.135 63.79 ;
    RECT 134.31 63.72 134.58 63.79 ;
    RECT 138.365 63.72 138.435 63.79 ;
    RECT 138.695 63.72 138.96 63.79 ;
    RECT 140.45 63.72 140.71 63.79 ;
    RECT 140.895 63.72 140.965 63.79 ;
    RECT 141.385 63.72 141.645 63.79 ;
    RECT 142.51 63.72 142.72 63.79 ;
    RECT 144.32 63.895 145.135 63.965 ;
    RECT 146.125 63.45 146.395 63.52 ;
    RECT 146.125 63.805 146.395 63.875 ;
    RECT 146.125 64.17 146.395 64.24 ;
    RECT 121.44 62.73 121.51 63.52 ;
    RECT 122.04 62.73 122.25 62.8 ;
    RECT 122.04 63.085 122.25 63.155 ;
    RECT 122.04 63.45 122.25 63.52 ;
    RECT 123.205 63.175 124.005 63.245 ;
    RECT 125.67 63.0 125.905 63.07 ;
    RECT 126.73 63.0 126.99 63.07 ;
    RECT 128.705 63.0 128.935 63.07 ;
    RECT 129.42 63.0 129.68 63.07 ;
    RECT 130.59 63.0 130.66 63.07 ;
    RECT 133.925 63.0 134.135 63.07 ;
    RECT 134.31 63.0 134.58 63.07 ;
    RECT 138.365 63.0 138.435 63.07 ;
    RECT 138.695 63.0 138.96 63.07 ;
    RECT 140.45 63.0 140.71 63.07 ;
    RECT 140.895 63.0 140.965 63.07 ;
    RECT 141.385 63.0 141.645 63.07 ;
    RECT 142.51 63.0 142.72 63.07 ;
    RECT 144.32 63.175 145.135 63.245 ;
    RECT 146.125 62.73 146.395 62.8 ;
    RECT 146.125 63.085 146.395 63.155 ;
    RECT 146.125 63.45 146.395 63.52 ;
    RECT 145.485 45.79 145.695 45.86 ;
    RECT 121.44 62.01 121.51 62.8 ;
    RECT 122.04 62.01 122.25 62.08 ;
    RECT 122.04 62.365 122.25 62.435 ;
    RECT 122.04 62.73 122.25 62.8 ;
    RECT 123.205 62.455 124.005 62.525 ;
    RECT 125.67 62.28 125.905 62.35 ;
    RECT 126.73 62.28 126.99 62.35 ;
    RECT 128.705 62.28 128.935 62.35 ;
    RECT 129.42 62.28 129.68 62.35 ;
    RECT 130.59 62.28 130.66 62.35 ;
    RECT 133.925 62.28 134.135 62.35 ;
    RECT 134.31 62.28 134.58 62.35 ;
    RECT 138.365 62.28 138.435 62.35 ;
    RECT 138.695 62.28 138.96 62.35 ;
    RECT 140.45 62.28 140.71 62.35 ;
    RECT 140.895 62.28 140.965 62.35 ;
    RECT 141.385 62.28 141.645 62.35 ;
    RECT 142.51 62.28 142.72 62.35 ;
    RECT 144.32 62.455 145.135 62.525 ;
    RECT 146.125 62.01 146.395 62.08 ;
    RECT 146.125 62.365 146.395 62.435 ;
    RECT 146.125 62.73 146.395 62.8 ;
    RECT 129.965 37.057 130.175 37.127 ;
    RECT 121.44 61.29 121.51 62.08 ;
    RECT 122.04 61.29 122.25 61.36 ;
    RECT 122.04 61.645 122.25 61.715 ;
    RECT 122.04 62.01 122.25 62.08 ;
    RECT 123.205 61.735 124.005 61.805 ;
    RECT 125.67 61.56 125.905 61.63 ;
    RECT 126.73 61.56 126.99 61.63 ;
    RECT 128.705 61.56 128.935 61.63 ;
    RECT 129.42 61.56 129.68 61.63 ;
    RECT 130.59 61.56 130.66 61.63 ;
    RECT 133.925 61.56 134.135 61.63 ;
    RECT 134.31 61.56 134.58 61.63 ;
    RECT 138.365 61.56 138.435 61.63 ;
    RECT 138.695 61.56 138.96 61.63 ;
    RECT 140.45 61.56 140.71 61.63 ;
    RECT 140.895 61.56 140.965 61.63 ;
    RECT 141.385 61.56 141.645 61.63 ;
    RECT 142.51 61.56 142.72 61.63 ;
    RECT 144.32 61.735 145.135 61.805 ;
    RECT 146.125 61.29 146.395 61.36 ;
    RECT 146.125 61.645 146.395 61.715 ;
    RECT 146.125 62.01 146.395 62.08 ;
    RECT 139.73 45.7 139.94 45.77 ;
    RECT 129.965 17.602 130.175 17.672 ;
    RECT 121.44 59.83 121.51 60.62 ;
    RECT 122.04 59.83 122.25 59.9 ;
    RECT 122.04 60.185 122.25 60.255 ;
    RECT 122.04 60.55 122.25 60.62 ;
    RECT 123.205 60.275 124.005 60.345 ;
    RECT 125.67 60.1 125.905 60.17 ;
    RECT 126.73 60.1 126.99 60.17 ;
    RECT 128.705 60.1 128.935 60.17 ;
    RECT 129.42 60.1 129.68 60.17 ;
    RECT 130.59 60.1 130.66 60.17 ;
    RECT 133.925 60.1 134.135 60.17 ;
    RECT 134.31 60.1 134.58 60.17 ;
    RECT 138.365 60.1 138.435 60.17 ;
    RECT 138.695 60.1 138.96 60.17 ;
    RECT 140.45 60.1 140.71 60.17 ;
    RECT 140.895 60.1 140.965 60.17 ;
    RECT 141.385 60.1 141.645 60.17 ;
    RECT 142.51 60.1 142.72 60.17 ;
    RECT 144.32 60.275 145.135 60.345 ;
    RECT 146.125 59.83 146.395 59.9 ;
    RECT 146.125 60.185 146.395 60.255 ;
    RECT 146.125 60.55 146.395 60.62 ;
    RECT 128.335 29.85 128.545 29.92 ;
    RECT 121.44 59.11 121.51 59.9 ;
    RECT 122.04 59.11 122.25 59.18 ;
    RECT 122.04 59.465 122.25 59.535 ;
    RECT 122.04 59.83 122.25 59.9 ;
    RECT 123.205 59.555 124.005 59.625 ;
    RECT 125.67 59.38 125.905 59.45 ;
    RECT 126.73 59.38 126.99 59.45 ;
    RECT 128.705 59.38 128.935 59.45 ;
    RECT 129.42 59.38 129.68 59.45 ;
    RECT 130.59 59.38 130.66 59.45 ;
    RECT 133.925 59.38 134.135 59.45 ;
    RECT 134.31 59.38 134.58 59.45 ;
    RECT 138.365 59.38 138.435 59.45 ;
    RECT 138.695 59.38 138.96 59.45 ;
    RECT 140.45 59.38 140.71 59.45 ;
    RECT 140.895 59.38 140.965 59.45 ;
    RECT 141.385 59.38 141.645 59.45 ;
    RECT 142.51 59.38 142.72 59.45 ;
    RECT 144.32 59.555 145.135 59.625 ;
    RECT 146.125 59.11 146.395 59.18 ;
    RECT 146.125 59.465 146.395 59.535 ;
    RECT 146.125 59.83 146.395 59.9 ;
    RECT 128.335 29.13 128.545 29.2 ;
    RECT 128.335 26.97 128.545 27.04 ;
    RECT 127.69 45.697 127.9 45.767 ;
    RECT 135.305 70.917 135.375 70.987 ;
    RECT 122.63 90.45 122.84 90.52 ;
    RECT 133.39 86.037 133.46 86.107 ;
    RECT 145.485 75.33 145.695 75.4 ;
    RECT 139.73 75.24 139.94 75.31 ;
    RECT 121.44 58.39 121.51 59.18 ;
    RECT 122.04 58.39 122.25 58.46 ;
    RECT 122.04 58.745 122.25 58.815 ;
    RECT 122.04 59.11 122.25 59.18 ;
    RECT 123.205 58.835 124.005 58.905 ;
    RECT 125.67 58.66 125.905 58.73 ;
    RECT 126.73 58.66 126.99 58.73 ;
    RECT 128.705 58.66 128.935 58.73 ;
    RECT 129.42 58.66 129.68 58.73 ;
    RECT 130.59 58.66 130.66 58.73 ;
    RECT 133.925 58.66 134.135 58.73 ;
    RECT 134.31 58.66 134.58 58.73 ;
    RECT 138.365 58.66 138.435 58.73 ;
    RECT 138.695 58.66 138.96 58.73 ;
    RECT 140.45 58.66 140.71 58.73 ;
    RECT 140.895 58.66 140.965 58.73 ;
    RECT 141.385 58.66 141.645 58.73 ;
    RECT 142.51 58.66 142.72 58.73 ;
    RECT 144.32 58.835 145.135 58.905 ;
    RECT 146.125 58.39 146.395 58.46 ;
    RECT 146.125 58.745 146.395 58.815 ;
    RECT 146.125 59.11 146.395 59.18 ;
    RECT 121.44 57.67 121.51 58.46 ;
    RECT 122.04 57.67 122.25 57.74 ;
    RECT 122.04 58.025 122.25 58.095 ;
    RECT 122.04 58.39 122.25 58.46 ;
    RECT 123.205 58.115 124.005 58.185 ;
    RECT 125.67 57.94 125.905 58.01 ;
    RECT 126.73 57.94 126.99 58.01 ;
    RECT 128.705 57.94 128.935 58.01 ;
    RECT 129.42 57.94 129.68 58.01 ;
    RECT 130.59 57.94 130.66 58.01 ;
    RECT 133.925 57.94 134.135 58.01 ;
    RECT 134.31 57.94 134.58 58.01 ;
    RECT 138.365 57.94 138.435 58.01 ;
    RECT 138.695 57.94 138.96 58.01 ;
    RECT 140.45 57.94 140.71 58.01 ;
    RECT 140.895 57.94 140.965 58.01 ;
    RECT 141.385 57.94 141.645 58.01 ;
    RECT 142.51 57.94 142.72 58.01 ;
    RECT 144.32 58.115 145.135 58.185 ;
    RECT 146.125 57.67 146.395 57.74 ;
    RECT 146.125 58.025 146.395 58.095 ;
    RECT 146.125 58.39 146.395 58.46 ;
    RECT 121.44 56.95 121.51 57.74 ;
    RECT 122.04 56.95 122.25 57.02 ;
    RECT 122.04 57.305 122.25 57.375 ;
    RECT 122.04 57.67 122.25 57.74 ;
    RECT 123.205 57.395 124.005 57.465 ;
    RECT 125.67 57.22 125.905 57.29 ;
    RECT 126.73 57.22 126.99 57.29 ;
    RECT 128.705 57.22 128.935 57.29 ;
    RECT 129.42 57.22 129.68 57.29 ;
    RECT 130.59 57.22 130.66 57.29 ;
    RECT 133.925 57.22 134.135 57.29 ;
    RECT 134.31 57.22 134.58 57.29 ;
    RECT 138.365 57.22 138.435 57.29 ;
    RECT 138.695 57.22 138.96 57.29 ;
    RECT 140.45 57.22 140.71 57.29 ;
    RECT 140.895 57.22 140.965 57.29 ;
    RECT 141.385 57.22 141.645 57.29 ;
    RECT 142.51 57.22 142.72 57.29 ;
    RECT 144.32 57.395 145.135 57.465 ;
    RECT 146.125 56.95 146.395 57.02 ;
    RECT 146.125 57.305 146.395 57.375 ;
    RECT 146.125 57.67 146.395 57.74 ;
    RECT 127.69 75.237 127.9 75.307 ;
    RECT 121.44 56.23 121.51 57.02 ;
    RECT 122.04 56.23 122.25 56.3 ;
    RECT 122.04 56.585 122.25 56.655 ;
    RECT 122.04 56.95 122.25 57.02 ;
    RECT 123.205 56.675 124.005 56.745 ;
    RECT 125.67 56.5 125.905 56.57 ;
    RECT 126.73 56.5 126.99 56.57 ;
    RECT 128.705 56.5 128.935 56.57 ;
    RECT 129.42 56.5 129.68 56.57 ;
    RECT 130.59 56.5 130.66 56.57 ;
    RECT 133.925 56.5 134.135 56.57 ;
    RECT 134.31 56.5 134.58 56.57 ;
    RECT 138.365 56.5 138.435 56.57 ;
    RECT 138.695 56.5 138.96 56.57 ;
    RECT 140.45 56.5 140.71 56.57 ;
    RECT 140.895 56.5 140.965 56.57 ;
    RECT 141.385 56.5 141.645 56.57 ;
    RECT 142.51 56.5 142.72 56.57 ;
    RECT 144.32 56.675 145.135 56.745 ;
    RECT 146.125 56.23 146.395 56.3 ;
    RECT 146.125 56.585 146.395 56.655 ;
    RECT 146.125 56.95 146.395 57.02 ;
    RECT 121.44 55.51 121.51 56.3 ;
    RECT 122.04 55.51 122.25 55.58 ;
    RECT 122.04 55.865 122.25 55.935 ;
    RECT 122.04 56.23 122.25 56.3 ;
    RECT 123.205 55.955 124.005 56.025 ;
    RECT 125.67 55.78 125.905 55.85 ;
    RECT 126.73 55.78 126.99 55.85 ;
    RECT 128.705 55.78 128.935 55.85 ;
    RECT 129.42 55.78 129.68 55.85 ;
    RECT 130.59 55.78 130.66 55.85 ;
    RECT 133.925 55.78 134.135 55.85 ;
    RECT 134.31 55.78 134.58 55.85 ;
    RECT 138.365 55.78 138.435 55.85 ;
    RECT 138.695 55.78 138.96 55.85 ;
    RECT 140.45 55.78 140.71 55.85 ;
    RECT 140.895 55.78 140.965 55.85 ;
    RECT 141.385 55.78 141.645 55.85 ;
    RECT 142.51 55.78 142.72 55.85 ;
    RECT 144.32 55.955 145.135 56.025 ;
    RECT 146.125 55.51 146.395 55.58 ;
    RECT 146.125 55.865 146.395 55.935 ;
    RECT 146.125 56.23 146.395 56.3 ;
    RECT 121.44 54.79 121.51 55.58 ;
    RECT 122.04 54.79 122.25 54.86 ;
    RECT 122.04 55.145 122.25 55.215 ;
    RECT 122.04 55.51 122.25 55.58 ;
    RECT 123.205 55.235 124.005 55.305 ;
    RECT 125.67 55.06 125.905 55.13 ;
    RECT 126.73 55.06 126.99 55.13 ;
    RECT 128.705 55.06 128.935 55.13 ;
    RECT 129.42 55.06 129.68 55.13 ;
    RECT 130.59 55.06 130.66 55.13 ;
    RECT 133.925 55.06 134.135 55.13 ;
    RECT 134.31 55.06 134.58 55.13 ;
    RECT 138.365 55.06 138.435 55.13 ;
    RECT 138.695 55.06 138.96 55.13 ;
    RECT 140.45 55.06 140.71 55.13 ;
    RECT 140.895 55.06 140.965 55.13 ;
    RECT 141.385 55.06 141.645 55.13 ;
    RECT 142.51 55.06 142.72 55.13 ;
    RECT 144.32 55.235 145.135 55.305 ;
    RECT 146.125 54.79 146.395 54.86 ;
    RECT 146.125 55.145 146.395 55.215 ;
    RECT 146.125 55.51 146.395 55.58 ;
    RECT 122.63 45.79 122.84 45.86 ;
    RECT 121.44 54.07 121.51 54.86 ;
    RECT 122.04 54.07 122.25 54.14 ;
    RECT 122.04 54.425 122.25 54.495 ;
    RECT 122.04 54.79 122.25 54.86 ;
    RECT 123.205 54.515 124.005 54.585 ;
    RECT 125.67 54.34 125.905 54.41 ;
    RECT 126.73 54.34 126.99 54.41 ;
    RECT 128.705 54.34 128.935 54.41 ;
    RECT 129.42 54.34 129.68 54.41 ;
    RECT 130.59 54.34 130.66 54.41 ;
    RECT 133.925 54.34 134.135 54.41 ;
    RECT 134.31 54.34 134.58 54.41 ;
    RECT 138.365 54.34 138.435 54.41 ;
    RECT 138.695 54.34 138.96 54.41 ;
    RECT 140.45 54.34 140.71 54.41 ;
    RECT 140.895 54.34 140.965 54.41 ;
    RECT 141.385 54.34 141.645 54.41 ;
    RECT 142.51 54.34 142.72 54.41 ;
    RECT 144.32 54.515 145.135 54.585 ;
    RECT 146.125 54.07 146.395 54.14 ;
    RECT 146.125 54.425 146.395 54.495 ;
    RECT 146.125 54.79 146.395 54.86 ;
    RECT 121.44 53.35 121.51 54.14 ;
    RECT 122.04 53.35 122.25 53.42 ;
    RECT 122.04 53.705 122.25 53.775 ;
    RECT 122.04 54.07 122.25 54.14 ;
    RECT 123.205 53.795 124.005 53.865 ;
    RECT 125.67 53.62 125.905 53.69 ;
    RECT 126.73 53.62 126.99 53.69 ;
    RECT 128.705 53.62 128.935 53.69 ;
    RECT 129.42 53.62 129.68 53.69 ;
    RECT 130.59 53.62 130.66 53.69 ;
    RECT 133.925 53.62 134.135 53.69 ;
    RECT 134.31 53.62 134.58 53.69 ;
    RECT 138.365 53.62 138.435 53.69 ;
    RECT 138.695 53.62 138.96 53.69 ;
    RECT 140.45 53.62 140.71 53.69 ;
    RECT 140.895 53.62 140.965 53.69 ;
    RECT 141.385 53.62 141.645 53.69 ;
    RECT 142.51 53.62 142.72 53.69 ;
    RECT 144.32 53.795 145.135 53.865 ;
    RECT 146.125 53.35 146.395 53.42 ;
    RECT 146.125 53.705 146.395 53.775 ;
    RECT 146.125 54.07 146.395 54.14 ;
    RECT 121.44 52.63 121.51 53.42 ;
    RECT 122.04 52.63 122.25 52.7 ;
    RECT 122.04 52.985 122.25 53.055 ;
    RECT 122.04 53.35 122.25 53.42 ;
    RECT 123.205 53.075 124.005 53.145 ;
    RECT 125.67 52.9 125.905 52.97 ;
    RECT 126.73 52.9 126.99 52.97 ;
    RECT 128.705 52.9 128.935 52.97 ;
    RECT 129.42 52.9 129.68 52.97 ;
    RECT 130.59 52.9 130.66 52.97 ;
    RECT 133.925 52.9 134.135 52.97 ;
    RECT 134.31 52.9 134.58 52.97 ;
    RECT 138.365 52.9 138.435 52.97 ;
    RECT 138.695 52.9 138.96 52.97 ;
    RECT 140.45 52.9 140.71 52.97 ;
    RECT 140.895 52.9 140.965 52.97 ;
    RECT 141.385 52.9 141.645 52.97 ;
    RECT 142.51 52.9 142.72 52.97 ;
    RECT 144.32 53.075 145.135 53.145 ;
    RECT 146.125 52.63 146.395 52.7 ;
    RECT 146.125 52.985 146.395 53.055 ;
    RECT 146.125 53.35 146.395 53.42 ;
    RECT 121.44 51.91 121.51 52.7 ;
    RECT 122.04 51.91 122.25 51.98 ;
    RECT 122.04 52.265 122.25 52.335 ;
    RECT 122.04 52.63 122.25 52.7 ;
    RECT 123.205 52.355 124.005 52.425 ;
    RECT 125.67 52.18 125.905 52.25 ;
    RECT 126.73 52.18 126.99 52.25 ;
    RECT 128.705 52.18 128.935 52.25 ;
    RECT 129.42 52.18 129.68 52.25 ;
    RECT 130.59 52.18 130.66 52.25 ;
    RECT 133.925 52.18 134.135 52.25 ;
    RECT 134.31 52.18 134.58 52.25 ;
    RECT 138.365 52.18 138.435 52.25 ;
    RECT 138.695 52.18 138.96 52.25 ;
    RECT 140.45 52.18 140.71 52.25 ;
    RECT 140.895 52.18 140.965 52.25 ;
    RECT 141.385 52.18 141.645 52.25 ;
    RECT 142.51 52.18 142.72 52.25 ;
    RECT 144.32 52.355 145.135 52.425 ;
    RECT 146.125 51.91 146.395 51.98 ;
    RECT 146.125 52.265 146.395 52.335 ;
    RECT 146.125 52.63 146.395 52.7 ;
    RECT 132.79 71.637 132.86 71.707 ;
    RECT 145.485 82.53 145.695 82.6 ;
    RECT 122.63 75.33 122.84 75.4 ;
    RECT 139.73 82.44 139.94 82.51 ;
    RECT 121.44 51.19 121.51 51.98 ;
    RECT 122.04 51.19 122.25 51.26 ;
    RECT 122.04 51.545 122.25 51.615 ;
    RECT 122.04 51.91 122.25 51.98 ;
    RECT 123.205 51.635 124.005 51.705 ;
    RECT 125.67 51.46 125.905 51.53 ;
    RECT 126.73 51.46 126.99 51.53 ;
    RECT 128.705 51.46 128.935 51.53 ;
    RECT 129.42 51.46 129.68 51.53 ;
    RECT 130.59 51.46 130.66 51.53 ;
    RECT 133.925 51.46 134.135 51.53 ;
    RECT 134.31 51.46 134.58 51.53 ;
    RECT 138.365 51.46 138.435 51.53 ;
    RECT 138.695 51.46 138.96 51.53 ;
    RECT 140.45 51.46 140.71 51.53 ;
    RECT 140.895 51.46 140.965 51.53 ;
    RECT 141.385 51.46 141.645 51.53 ;
    RECT 142.51 51.46 142.72 51.53 ;
    RECT 144.32 51.635 145.135 51.705 ;
    RECT 146.125 51.19 146.395 51.26 ;
    RECT 146.125 51.545 146.395 51.615 ;
    RECT 146.125 51.91 146.395 51.98 ;
    RECT 121.44 50.47 121.51 51.26 ;
    RECT 122.04 50.47 122.25 50.54 ;
    RECT 122.04 50.825 122.25 50.895 ;
    RECT 122.04 51.19 122.25 51.26 ;
    RECT 123.205 50.915 124.005 50.985 ;
    RECT 125.67 50.74 125.905 50.81 ;
    RECT 126.73 50.74 126.99 50.81 ;
    RECT 128.705 50.74 128.935 50.81 ;
    RECT 129.42 50.74 129.68 50.81 ;
    RECT 130.59 50.74 130.66 50.81 ;
    RECT 133.925 50.74 134.135 50.81 ;
    RECT 134.31 50.74 134.58 50.81 ;
    RECT 138.365 50.74 138.435 50.81 ;
    RECT 138.695 50.74 138.96 50.81 ;
    RECT 140.45 50.74 140.71 50.81 ;
    RECT 140.895 50.74 140.965 50.81 ;
    RECT 141.385 50.74 141.645 50.81 ;
    RECT 142.51 50.74 142.72 50.81 ;
    RECT 144.32 50.915 145.135 50.985 ;
    RECT 146.125 50.47 146.395 50.54 ;
    RECT 146.125 50.825 146.395 50.895 ;
    RECT 146.125 51.19 146.395 51.26 ;
    RECT 127.69 82.437 127.9 82.507 ;
    RECT 267.7 11.985 267.77 12.195 ;
    RECT 267.7 7.972 267.77 8.182 ;
    RECT 268.12 13.97 268.19 14.04 ;
    RECT 267.91 14.23 267.98 14.3 ;
    RECT 267.7 6.12 267.77 6.19 ;
    RECT 267.7 4.445 267.77 4.655 ;
    RECT 267.7 3.32 267.77 3.53 ;
    RECT 267.91 7.58 267.98 7.65 ;
    RECT 267.695 4.22 267.765 4.29 ;
    RECT 267.695 7.125 267.765 7.195 ;
    RECT 246.79 4.445 246.86 4.655 ;
    RECT 262.9 9.995 263.11 10.205 ;
    RECT 262.9 8.902 263.11 9.112 ;
    RECT 262.9 8.705 263.11 8.775 ;
    RECT 247.22 7.125 247.43 7.195 ;
    RECT 262.9 8.325 263.11 8.395 ;
    RECT 247.22 4.22 247.43 4.29 ;
    RECT 262.9 6.315 263.11 6.385 ;
    RECT 262.9 4.815 263.11 5.025 ;
    RECT 262.9 3.742 263.11 3.952 ;
    RECT 262.9 2.99 263.11 3.2 ;
    RECT 243.47 6.12 243.54 6.19 ;
    RECT 243.47 5.182 243.54 5.392 ;
    RECT 259.58 9.995 259.79 10.205 ;
    RECT 243.47 4.445 243.54 4.655 ;
    RECT 259.58 8.902 259.79 9.112 ;
    RECT 259.58 8.705 259.79 8.775 ;
    RECT 259.58 8.325 259.79 8.395 ;
    RECT 243.9 7.125 244.11 7.195 ;
    RECT 259.58 6.315 259.79 6.385 ;
    RECT 243.9 4.22 244.11 4.29 ;
    RECT 259.58 4.815 259.79 5.025 ;
    RECT 259.58 3.742 259.79 3.952 ;
    RECT 259.58 2.99 259.79 3.2 ;
    RECT 240.15 6.12 240.22 6.19 ;
    RECT 256.26 9.995 256.47 10.205 ;
    RECT 240.15 5.182 240.22 5.392 ;
    RECT 256.26 8.902 256.47 9.112 ;
    RECT 240.15 4.445 240.22 4.655 ;
    RECT 256.26 8.705 256.47 8.775 ;
    RECT 256.26 8.325 256.47 8.395 ;
    RECT 240.58 7.125 240.79 7.195 ;
    RECT 240.58 4.22 240.79 4.29 ;
    RECT 236.83 6.12 236.9 6.19 ;
    RECT 236.83 5.182 236.9 5.392 ;
    RECT 236.83 4.445 236.9 4.655 ;
    RECT 180.785 5.255 181.065 5.325 ;
    RECT 180.785 8.065 181.065 8.135 ;
    RECT 180.785 11.985 181.065 12.195 ;
    RECT 180.82 3.32 181.03 3.53 ;
    RECT 180.82 4.445 181.03 4.655 ;
    RECT 180.82 6.12 181.03 6.19 ;
    RECT 180.59 3.035 180.66 3.105 ;
    RECT 180.59 3.78 180.66 3.85 ;
    RECT 180.59 4.86 180.66 4.93 ;
    RECT 180.59 6.315 180.66 6.385 ;
    RECT 180.59 6.745 180.66 6.815 ;
    RECT 180.59 12.31 180.66 12.38 ;
    RECT 180.39 4.23 180.46 4.3 ;
    RECT 180.39 7.135 180.46 7.205 ;
    RECT 180.39 8.325 180.46 8.395 ;
    RECT 180.39 8.71 180.46 9.115 ;
    RECT 180.39 9.995 180.46 10.205 ;
    RECT 179.385 12.605 179.65 12.675 ;
    RECT 179.12 8.325 179.19 8.395 ;
    RECT 178.92 8.325 179.19 9.115 ;
    RECT 179.12 8.71 179.19 8.97 ;
    RECT 178.92 9.995 179.19 10.205 ;
    RECT 178.95 2.99 179.16 3.955 ;
    RECT 178.95 4.815 179.16 5.025 ;
    RECT 178.95 6.315 179.16 6.385 ;
    RECT 177.465 5.255 177.745 5.325 ;
    RECT 177.465 8.065 177.745 8.135 ;
    RECT 177.465 11.985 177.745 12.195 ;
    RECT 177.5 3.32 177.71 3.53 ;
    RECT 177.5 4.445 177.71 4.655 ;
    RECT 177.5 6.12 177.71 6.19 ;
    RECT 177.27 3.035 177.34 3.105 ;
    RECT 177.27 3.78 177.34 3.85 ;
    RECT 177.27 4.86 177.34 4.93 ;
    RECT 177.27 6.315 177.34 6.385 ;
    RECT 177.27 6.745 177.34 6.815 ;
    RECT 177.27 12.31 177.34 12.38 ;
    RECT 177.07 4.23 177.14 4.3 ;
    RECT 177.07 7.135 177.14 7.205 ;
    RECT 177.07 8.325 177.14 8.395 ;
    RECT 177.07 8.71 177.14 9.115 ;
    RECT 177.07 9.995 177.14 10.205 ;
    RECT 176.065 12.605 176.33 12.675 ;
    RECT 175.8 8.325 175.87 8.395 ;
    RECT 175.6 8.325 175.87 9.115 ;
    RECT 175.8 8.71 175.87 8.97 ;
    RECT 175.6 9.995 175.87 10.205 ;
    RECT 175.63 2.99 175.84 3.955 ;
    RECT 175.63 4.815 175.84 5.025 ;
    RECT 175.63 6.315 175.84 6.385 ;
    RECT 174.145 5.255 174.425 5.325 ;
    RECT 174.145 8.065 174.425 8.135 ;
    RECT 174.145 11.985 174.425 12.195 ;
    RECT 174.18 3.32 174.39 3.53 ;
    RECT 174.18 4.445 174.39 4.655 ;
    RECT 174.18 6.12 174.39 6.19 ;
    RECT 173.95 3.035 174.02 3.105 ;
    RECT 173.95 3.78 174.02 3.85 ;
    RECT 173.95 4.86 174.02 4.93 ;
    RECT 173.95 6.315 174.02 6.385 ;
    RECT 173.95 6.745 174.02 6.815 ;
    RECT 173.95 12.31 174.02 12.38 ;
    RECT 173.75 4.23 173.82 4.3 ;
    RECT 173.75 7.135 173.82 7.205 ;
    RECT 173.75 8.325 173.82 8.395 ;
    RECT 173.75 8.71 173.82 9.115 ;
    RECT 173.75 9.995 173.82 10.205 ;
    RECT 172.745 12.605 173.01 12.675 ;
    RECT 172.48 8.325 172.55 8.395 ;
    RECT 172.28 8.325 172.55 9.115 ;
    RECT 172.48 8.71 172.55 8.97 ;
    RECT 172.28 9.995 172.55 10.205 ;
    RECT 172.31 2.99 172.52 3.955 ;
    RECT 172.31 4.815 172.52 5.025 ;
    RECT 172.31 6.315 172.52 6.385 ;
    RECT 170.825 5.255 171.105 5.325 ;
    RECT 170.825 8.065 171.105 8.135 ;
    RECT 170.825 11.985 171.105 12.195 ;
    RECT 170.86 3.32 171.07 3.53 ;
    RECT 170.86 4.445 171.07 4.655 ;
    RECT 170.86 6.12 171.07 6.19 ;
    RECT 170.63 3.035 170.7 3.105 ;
    RECT 170.63 3.78 170.7 3.85 ;
    RECT 170.63 4.86 170.7 4.93 ;
    RECT 170.63 6.315 170.7 6.385 ;
    RECT 170.63 6.745 170.7 6.815 ;
    RECT 170.63 12.31 170.7 12.38 ;
    RECT 170.43 4.23 170.5 4.3 ;
    RECT 170.43 7.135 170.5 7.205 ;
    RECT 170.43 8.325 170.5 8.395 ;
    RECT 170.43 8.71 170.5 9.115 ;
    RECT 170.43 9.995 170.5 10.205 ;
    RECT 169.425 12.605 169.69 12.675 ;
    RECT 169.16 8.325 169.23 8.395 ;
    RECT 168.96 8.325 169.23 9.115 ;
    RECT 169.16 8.71 169.23 8.97 ;
    RECT 168.96 9.995 169.23 10.205 ;
    RECT 168.99 2.99 169.2 3.955 ;
    RECT 168.99 4.815 169.2 5.025 ;
    RECT 168.99 6.315 169.2 6.385 ;
    RECT 167.505 5.255 167.785 5.325 ;
    RECT 167.505 8.065 167.785 8.135 ;
    RECT 167.505 11.985 167.785 12.195 ;
    RECT 167.54 3.32 167.75 3.53 ;
    RECT 167.54 4.445 167.75 4.655 ;
    RECT 167.54 6.12 167.75 6.19 ;
    RECT 167.31 3.035 167.38 3.105 ;
    RECT 167.31 3.78 167.38 3.85 ;
    RECT 167.31 4.86 167.38 4.93 ;
    RECT 167.31 6.315 167.38 6.385 ;
    RECT 167.31 6.745 167.38 6.815 ;
    RECT 167.31 12.31 167.38 12.38 ;
    RECT 167.11 4.23 167.18 4.3 ;
    RECT 167.11 7.135 167.18 7.205 ;
    RECT 167.11 8.325 167.18 8.395 ;
    RECT 167.11 8.71 167.18 9.115 ;
    RECT 167.11 9.995 167.18 10.205 ;
    RECT 166.105 12.605 166.37 12.675 ;
    RECT 165.84 8.325 165.91 8.395 ;
    RECT 165.64 8.325 165.91 9.115 ;
    RECT 165.84 8.71 165.91 8.97 ;
    RECT 165.64 9.995 165.91 10.205 ;
    RECT 165.67 2.99 165.88 3.955 ;
    RECT 165.67 4.815 165.88 5.025 ;
    RECT 165.67 6.315 165.88 6.385 ;
    RECT 164.185 5.255 164.465 5.325 ;
    RECT 164.185 8.065 164.465 8.135 ;
    RECT 164.185 11.985 164.465 12.195 ;
    RECT 164.22 3.32 164.43 3.53 ;
    RECT 164.22 4.445 164.43 4.655 ;
    RECT 164.22 6.12 164.43 6.19 ;
    RECT 163.99 3.035 164.06 3.105 ;
    RECT 163.99 3.78 164.06 3.85 ;
    RECT 163.99 4.86 164.06 4.93 ;
    RECT 163.99 6.315 164.06 6.385 ;
    RECT 163.99 6.745 164.06 6.815 ;
    RECT 163.99 12.31 164.06 12.38 ;
    RECT 163.79 4.23 163.86 4.3 ;
    RECT 163.79 7.135 163.86 7.205 ;
    RECT 163.79 8.325 163.86 8.395 ;
    RECT 163.79 8.71 163.86 9.115 ;
    RECT 163.79 9.995 163.86 10.205 ;
    RECT 162.785 12.605 163.05 12.675 ;
    RECT 162.52 8.325 162.59 8.395 ;
    RECT 162.32 8.325 162.59 9.115 ;
    RECT 162.52 8.71 162.59 8.97 ;
    RECT 162.32 9.995 162.59 10.205 ;
    RECT 162.35 2.99 162.56 3.955 ;
    RECT 162.35 4.815 162.56 5.025 ;
    RECT 162.35 6.315 162.56 6.385 ;
    RECT 160.865 5.255 161.145 5.325 ;
    RECT 160.865 8.065 161.145 8.135 ;
    RECT 160.865 11.985 161.145 12.195 ;
    RECT 160.9 3.32 161.11 3.53 ;
    RECT 160.9 4.445 161.11 4.655 ;
    RECT 160.9 6.12 161.11 6.19 ;
    RECT 160.67 3.035 160.74 3.105 ;
    RECT 160.67 3.78 160.74 3.85 ;
    RECT 160.67 4.86 160.74 4.93 ;
    RECT 160.67 6.315 160.74 6.385 ;
    RECT 160.67 6.745 160.74 6.815 ;
    RECT 160.67 12.31 160.74 12.38 ;
    RECT 160.47 4.23 160.54 4.3 ;
    RECT 160.47 7.135 160.54 7.205 ;
    RECT 160.47 8.325 160.54 8.395 ;
    RECT 160.47 8.71 160.54 9.115 ;
    RECT 160.47 9.995 160.54 10.205 ;
    RECT 159.465 12.605 159.73 12.675 ;
    RECT 159.2 8.325 159.27 8.395 ;
    RECT 159.0 8.325 159.27 9.115 ;
    RECT 159.2 8.71 159.27 8.97 ;
    RECT 159.0 9.995 159.27 10.205 ;
    RECT 159.03 2.99 159.24 3.955 ;
    RECT 159.03 4.815 159.24 5.025 ;
    RECT 159.03 6.315 159.24 6.385 ;
    RECT 157.545 5.255 157.825 5.325 ;
    RECT 157.545 8.065 157.825 8.135 ;
    RECT 157.545 11.985 157.825 12.195 ;
    RECT 157.58 3.32 157.79 3.53 ;
    RECT 157.58 4.445 157.79 4.655 ;
    RECT 157.58 6.12 157.79 6.19 ;
    RECT 157.35 3.035 157.42 3.105 ;
    RECT 157.35 3.78 157.42 3.85 ;
    RECT 157.35 4.86 157.42 4.93 ;
    RECT 157.35 6.315 157.42 6.385 ;
    RECT 157.35 6.745 157.42 6.815 ;
    RECT 157.35 12.31 157.42 12.38 ;
    RECT 157.15 4.23 157.22 4.3 ;
    RECT 157.15 7.135 157.22 7.205 ;
    RECT 157.15 8.325 157.22 8.395 ;
    RECT 157.15 8.71 157.22 9.115 ;
    RECT 157.15 9.995 157.22 10.205 ;
    RECT 156.145 12.605 156.41 12.675 ;
    RECT 155.88 8.325 155.95 8.395 ;
    RECT 155.68 8.325 155.95 9.115 ;
    RECT 155.88 8.71 155.95 8.97 ;
    RECT 155.68 9.995 155.95 10.205 ;
    RECT 155.71 2.99 155.92 3.955 ;
    RECT 155.71 4.815 155.92 5.025 ;
    RECT 155.71 6.315 155.92 6.385 ;
    RECT 154.225 5.255 154.505 5.325 ;
    RECT 154.225 8.065 154.505 8.135 ;
    RECT 154.225 11.985 154.505 12.195 ;
    RECT 154.26 3.32 154.47 3.53 ;
    RECT 154.26 4.445 154.47 4.655 ;
    RECT 154.26 6.12 154.47 6.19 ;
    RECT 154.03 3.035 154.1 3.105 ;
    RECT 154.03 3.78 154.1 3.85 ;
    RECT 154.03 4.86 154.1 4.93 ;
    RECT 154.03 6.315 154.1 6.385 ;
    RECT 154.03 6.745 154.1 6.815 ;
    RECT 154.03 12.31 154.1 12.38 ;
    RECT 153.83 4.23 153.9 4.3 ;
    RECT 153.83 7.135 153.9 7.205 ;
    RECT 153.83 8.325 153.9 8.395 ;
    RECT 153.83 8.71 153.9 9.115 ;
    RECT 153.83 9.995 153.9 10.205 ;
    RECT 152.825 12.605 153.09 12.675 ;
    RECT 152.56 8.325 152.63 8.395 ;
    RECT 152.36 8.325 152.63 9.115 ;
    RECT 152.56 8.71 152.63 8.97 ;
    RECT 152.36 9.995 152.63 10.205 ;
    RECT 152.39 2.99 152.6 3.955 ;
    RECT 152.39 4.815 152.6 5.025 ;
    RECT 152.39 6.315 152.6 6.385 ;
    RECT 266.22 7.565 266.43 7.635 ;
    RECT 267.105 5.255 267.385 5.325 ;
    RECT 267.105 8.065 267.385 8.135 ;
    RECT 267.105 11.985 267.385 12.195 ;
    RECT 267.14 3.32 267.35 3.53 ;
    RECT 267.14 4.445 267.35 4.655 ;
    RECT 267.14 6.12 267.35 6.19 ;
    RECT 266.91 3.035 266.98 3.105 ;
    RECT 266.91 3.78 266.98 3.85 ;
    RECT 266.91 4.86 266.98 4.93 ;
    RECT 266.91 6.315 266.98 6.385 ;
    RECT 266.91 6.745 266.98 6.815 ;
    RECT 266.91 12.31 266.98 12.38 ;
    RECT 266.71 4.23 266.78 4.3 ;
    RECT 266.71 7.135 266.78 7.205 ;
    RECT 266.71 8.325 266.78 8.395 ;
    RECT 266.71 8.71 266.78 9.115 ;
    RECT 266.71 9.995 266.78 10.205 ;
    RECT 265.705 12.605 265.97 12.675 ;
    RECT 265.44 8.325 265.51 8.395 ;
    RECT 265.24 8.325 265.51 9.115 ;
    RECT 265.44 8.71 265.51 8.97 ;
    RECT 265.24 9.995 265.51 10.205 ;
    RECT 265.27 2.99 265.48 3.955 ;
    RECT 265.27 4.815 265.48 5.025 ;
    RECT 265.27 6.315 265.48 6.385 ;
    RECT 150.905 5.255 151.185 5.325 ;
    RECT 150.905 8.065 151.185 8.135 ;
    RECT 150.905 11.985 151.185 12.195 ;
    RECT 150.94 3.32 151.15 3.53 ;
    RECT 150.94 4.445 151.15 4.655 ;
    RECT 150.94 6.12 151.15 6.19 ;
    RECT 150.71 3.035 150.78 3.105 ;
    RECT 150.71 3.78 150.78 3.85 ;
    RECT 150.71 4.86 150.78 4.93 ;
    RECT 150.71 6.315 150.78 6.385 ;
    RECT 150.71 6.745 150.78 6.815 ;
    RECT 150.71 12.31 150.78 12.38 ;
    RECT 150.51 4.23 150.58 4.3 ;
    RECT 150.51 7.135 150.58 7.205 ;
    RECT 150.51 8.325 150.58 8.395 ;
    RECT 150.51 8.71 150.58 9.115 ;
    RECT 150.51 9.995 150.58 10.205 ;
    RECT 149.505 12.605 149.77 12.675 ;
    RECT 149.24 8.325 149.31 8.395 ;
    RECT 149.04 8.325 149.31 9.115 ;
    RECT 149.24 8.71 149.31 8.97 ;
    RECT 149.04 9.995 149.31 10.205 ;
    RECT 149.07 2.99 149.28 3.955 ;
    RECT 149.07 4.815 149.28 5.025 ;
    RECT 149.07 6.315 149.28 6.385 ;
    RECT 262.9 7.565 263.11 7.635 ;
    RECT 259.58 7.565 259.79 7.635 ;
    RECT 256.26 7.565 256.47 7.635 ;
    RECT 252.94 7.565 253.15 7.635 ;
    RECT 263.785 5.255 264.065 5.325 ;
    RECT 263.785 8.065 264.065 8.135 ;
    RECT 263.785 11.985 264.065 12.195 ;
    RECT 263.82 3.32 264.03 3.53 ;
    RECT 263.82 4.445 264.03 4.655 ;
    RECT 263.82 6.12 264.03 6.19 ;
    RECT 263.59 3.035 263.66 3.105 ;
    RECT 263.59 3.78 263.66 3.85 ;
    RECT 263.59 4.86 263.66 4.93 ;
    RECT 263.59 6.315 263.66 6.385 ;
    RECT 263.59 6.745 263.66 6.815 ;
    RECT 263.59 12.31 263.66 12.38 ;
    RECT 263.39 4.23 263.46 4.3 ;
    RECT 263.39 7.135 263.46 7.205 ;
    RECT 263.39 8.325 263.46 8.395 ;
    RECT 263.39 8.71 263.46 9.115 ;
    RECT 263.39 9.995 263.46 10.205 ;
    RECT 262.385 12.605 262.65 12.675 ;
    RECT 262.12 8.325 262.19 8.395 ;
    RECT 261.92 8.325 262.19 9.115 ;
    RECT 262.12 8.71 262.19 8.97 ;
    RECT 261.92 9.995 262.19 10.205 ;
    RECT 261.95 2.99 262.16 3.955 ;
    RECT 261.95 4.815 262.16 5.025 ;
    RECT 261.95 6.315 262.16 6.385 ;
    RECT 249.62 7.565 249.83 7.635 ;
    RECT 260.465 5.255 260.745 5.325 ;
    RECT 260.465 8.065 260.745 8.135 ;
    RECT 260.465 11.985 260.745 12.195 ;
    RECT 260.5 3.32 260.71 3.53 ;
    RECT 260.5 4.445 260.71 4.655 ;
    RECT 260.5 6.12 260.71 6.19 ;
    RECT 260.27 3.035 260.34 3.105 ;
    RECT 260.27 3.78 260.34 3.85 ;
    RECT 260.27 4.86 260.34 4.93 ;
    RECT 260.27 6.315 260.34 6.385 ;
    RECT 260.27 6.745 260.34 6.815 ;
    RECT 260.27 12.31 260.34 12.38 ;
    RECT 260.07 4.23 260.14 4.3 ;
    RECT 260.07 7.135 260.14 7.205 ;
    RECT 260.07 8.325 260.14 8.395 ;
    RECT 260.07 8.71 260.14 9.115 ;
    RECT 260.07 9.995 260.14 10.205 ;
    RECT 259.065 12.605 259.33 12.675 ;
    RECT 258.8 8.325 258.87 8.395 ;
    RECT 258.6 8.325 258.87 9.115 ;
    RECT 258.8 8.71 258.87 8.97 ;
    RECT 258.6 9.995 258.87 10.205 ;
    RECT 258.63 2.99 258.84 3.955 ;
    RECT 258.63 4.815 258.84 5.025 ;
    RECT 258.63 6.315 258.84 6.385 ;
    RECT 257.145 5.255 257.425 5.325 ;
    RECT 257.145 8.065 257.425 8.135 ;
    RECT 257.145 11.985 257.425 12.195 ;
    RECT 257.18 3.32 257.39 3.53 ;
    RECT 257.18 4.445 257.39 4.655 ;
    RECT 257.18 6.12 257.39 6.19 ;
    RECT 256.95 3.035 257.02 3.105 ;
    RECT 256.95 3.78 257.02 3.85 ;
    RECT 256.95 4.86 257.02 4.93 ;
    RECT 256.95 6.315 257.02 6.385 ;
    RECT 256.95 6.745 257.02 6.815 ;
    RECT 256.95 12.31 257.02 12.38 ;
    RECT 256.75 4.23 256.82 4.3 ;
    RECT 256.75 7.135 256.82 7.205 ;
    RECT 256.75 8.325 256.82 8.395 ;
    RECT 256.75 8.71 256.82 9.115 ;
    RECT 256.75 9.995 256.82 10.205 ;
    RECT 255.745 12.605 256.01 12.675 ;
    RECT 255.48 8.325 255.55 8.395 ;
    RECT 255.28 8.325 255.55 9.115 ;
    RECT 255.48 8.71 255.55 8.97 ;
    RECT 255.28 9.995 255.55 10.205 ;
    RECT 255.31 2.99 255.52 3.955 ;
    RECT 255.31 4.815 255.52 5.025 ;
    RECT 255.31 6.315 255.52 6.385 ;
    RECT 253.825 5.255 254.105 5.325 ;
    RECT 253.825 8.065 254.105 8.135 ;
    RECT 253.825 11.985 254.105 12.195 ;
    RECT 253.86 3.32 254.07 3.53 ;
    RECT 253.86 4.445 254.07 4.655 ;
    RECT 253.86 6.12 254.07 6.19 ;
    RECT 253.63 3.035 253.7 3.105 ;
    RECT 253.63 3.78 253.7 3.85 ;
    RECT 253.63 4.86 253.7 4.93 ;
    RECT 253.63 6.315 253.7 6.385 ;
    RECT 253.63 6.745 253.7 6.815 ;
    RECT 253.63 12.31 253.7 12.38 ;
    RECT 253.43 4.23 253.5 4.3 ;
    RECT 253.43 7.135 253.5 7.205 ;
    RECT 253.43 8.325 253.5 8.395 ;
    RECT 253.43 8.71 253.5 9.115 ;
    RECT 253.43 9.995 253.5 10.205 ;
    RECT 252.425 12.605 252.69 12.675 ;
    RECT 252.16 8.325 252.23 8.395 ;
    RECT 251.96 8.325 252.23 9.115 ;
    RECT 252.16 8.71 252.23 8.97 ;
    RECT 251.96 9.995 252.23 10.205 ;
    RECT 251.99 2.99 252.2 3.955 ;
    RECT 251.99 4.815 252.2 5.025 ;
    RECT 251.99 6.315 252.2 6.385 ;
    RECT 250.505 5.255 250.785 5.325 ;
    RECT 250.505 8.065 250.785 8.135 ;
    RECT 250.505 11.985 250.785 12.195 ;
    RECT 250.54 3.32 250.75 3.53 ;
    RECT 250.54 4.445 250.75 4.655 ;
    RECT 250.54 6.12 250.75 6.19 ;
    RECT 250.31 3.035 250.38 3.105 ;
    RECT 250.31 3.78 250.38 3.85 ;
    RECT 250.31 4.86 250.38 4.93 ;
    RECT 250.31 6.315 250.38 6.385 ;
    RECT 250.31 6.745 250.38 6.815 ;
    RECT 250.31 12.31 250.38 12.38 ;
    RECT 250.11 4.23 250.18 4.3 ;
    RECT 250.11 7.135 250.18 7.205 ;
    RECT 250.11 8.325 250.18 8.395 ;
    RECT 250.11 8.71 250.18 9.115 ;
    RECT 250.11 9.995 250.18 10.205 ;
    RECT 249.105 12.605 249.37 12.675 ;
    RECT 248.84 8.325 248.91 8.395 ;
    RECT 248.64 8.325 248.91 9.115 ;
    RECT 248.84 8.71 248.91 8.97 ;
    RECT 248.64 9.995 248.91 10.205 ;
    RECT 248.67 2.99 248.88 3.955 ;
    RECT 248.67 4.815 248.88 5.025 ;
    RECT 248.67 6.315 248.88 6.385 ;
    RECT 247.185 5.255 247.465 5.325 ;
    RECT 247.185 8.065 247.465 8.135 ;
    RECT 247.185 11.985 247.465 12.195 ;
    RECT 247.22 3.32 247.43 3.53 ;
    RECT 247.22 4.445 247.43 4.655 ;
    RECT 247.22 6.12 247.43 6.19 ;
    RECT 246.99 3.035 247.06 3.105 ;
    RECT 246.99 3.78 247.06 3.85 ;
    RECT 246.99 4.86 247.06 4.93 ;
    RECT 246.99 6.315 247.06 6.385 ;
    RECT 246.99 6.745 247.06 6.815 ;
    RECT 246.99 12.31 247.06 12.38 ;
    RECT 246.79 4.23 246.86 4.3 ;
    RECT 246.79 7.135 246.86 7.205 ;
    RECT 246.79 8.325 246.86 8.395 ;
    RECT 246.79 8.71 246.86 9.115 ;
    RECT 246.79 9.995 246.86 10.205 ;
    RECT 245.785 12.605 246.05 12.675 ;
    RECT 245.52 8.325 245.59 8.395 ;
    RECT 245.32 8.325 245.59 9.115 ;
    RECT 245.52 8.71 245.59 8.97 ;
    RECT 245.32 9.995 245.59 10.205 ;
    RECT 245.35 2.99 245.56 3.955 ;
    RECT 245.35 4.815 245.56 5.025 ;
    RECT 245.35 6.315 245.56 6.385 ;
    RECT 243.865 5.255 244.145 5.325 ;
    RECT 243.865 8.065 244.145 8.135 ;
    RECT 243.865 11.985 244.145 12.195 ;
    RECT 243.9 3.32 244.11 3.53 ;
    RECT 243.9 4.445 244.11 4.655 ;
    RECT 243.9 6.12 244.11 6.19 ;
    RECT 243.67 3.035 243.74 3.105 ;
    RECT 243.67 3.78 243.74 3.85 ;
    RECT 243.67 4.86 243.74 4.93 ;
    RECT 243.67 6.315 243.74 6.385 ;
    RECT 243.67 6.745 243.74 6.815 ;
    RECT 243.67 12.31 243.74 12.38 ;
    RECT 243.47 4.23 243.54 4.3 ;
    RECT 243.47 7.135 243.54 7.205 ;
    RECT 243.47 8.325 243.54 8.395 ;
    RECT 243.47 8.71 243.54 9.115 ;
    RECT 243.47 9.995 243.54 10.205 ;
    RECT 242.465 12.605 242.73 12.675 ;
    RECT 242.2 8.325 242.27 8.395 ;
    RECT 242.0 8.325 242.27 9.115 ;
    RECT 242.2 8.71 242.27 8.97 ;
    RECT 242.0 9.995 242.27 10.205 ;
    RECT 242.03 2.99 242.24 3.955 ;
    RECT 242.03 4.815 242.24 5.025 ;
    RECT 242.03 6.315 242.24 6.385 ;
    RECT 240.545 5.255 240.825 5.325 ;
    RECT 240.545 8.065 240.825 8.135 ;
    RECT 240.545 11.985 240.825 12.195 ;
    RECT 240.58 3.32 240.79 3.53 ;
    RECT 240.58 4.445 240.79 4.655 ;
    RECT 240.58 6.12 240.79 6.19 ;
    RECT 240.35 3.035 240.42 3.105 ;
    RECT 240.35 3.78 240.42 3.85 ;
    RECT 240.35 4.86 240.42 4.93 ;
    RECT 240.35 6.315 240.42 6.385 ;
    RECT 240.35 6.745 240.42 6.815 ;
    RECT 240.35 12.31 240.42 12.38 ;
    RECT 240.15 4.23 240.22 4.3 ;
    RECT 240.15 7.135 240.22 7.205 ;
    RECT 240.15 8.325 240.22 8.395 ;
    RECT 240.15 8.71 240.22 9.115 ;
    RECT 240.15 9.995 240.22 10.205 ;
    RECT 239.145 12.605 239.41 12.675 ;
    RECT 238.88 8.325 238.95 8.395 ;
    RECT 238.68 8.325 238.95 9.115 ;
    RECT 238.88 8.71 238.95 8.97 ;
    RECT 238.68 9.995 238.95 10.205 ;
    RECT 238.71 2.99 238.92 3.955 ;
    RECT 238.71 4.815 238.92 5.025 ;
    RECT 238.71 6.315 238.92 6.385 ;
    RECT 237.225 5.255 237.505 5.325 ;
    RECT 237.225 8.065 237.505 8.135 ;
    RECT 237.225 11.985 237.505 12.195 ;
    RECT 237.26 3.32 237.47 3.53 ;
    RECT 237.26 4.445 237.47 4.655 ;
    RECT 237.26 6.12 237.47 6.19 ;
    RECT 237.03 3.035 237.1 3.105 ;
    RECT 237.03 3.78 237.1 3.85 ;
    RECT 237.03 4.86 237.1 4.93 ;
    RECT 237.03 6.315 237.1 6.385 ;
    RECT 237.03 6.745 237.1 6.815 ;
    RECT 237.03 12.31 237.1 12.38 ;
    RECT 236.83 4.23 236.9 4.3 ;
    RECT 236.83 7.135 236.9 7.205 ;
    RECT 236.83 8.325 236.9 8.395 ;
    RECT 236.83 8.71 236.9 9.115 ;
    RECT 236.83 9.995 236.9 10.205 ;
    RECT 235.825 12.605 236.09 12.675 ;
    RECT 235.56 8.325 235.63 8.395 ;
    RECT 235.36 8.325 235.63 9.115 ;
    RECT 235.56 8.71 235.63 8.97 ;
    RECT 235.36 9.995 235.63 10.205 ;
    RECT 235.39 2.99 235.6 3.955 ;
    RECT 235.39 4.815 235.6 5.025 ;
    RECT 235.39 6.315 235.6 6.385 ;
    RECT 233.905 5.255 234.185 5.325 ;
    RECT 233.905 8.065 234.185 8.135 ;
    RECT 233.905 11.985 234.185 12.195 ;
    RECT 233.94 3.32 234.15 3.53 ;
    RECT 233.94 4.445 234.15 4.655 ;
    RECT 233.94 6.12 234.15 6.19 ;
    RECT 233.71 3.035 233.78 3.105 ;
    RECT 233.71 3.78 233.78 3.85 ;
    RECT 233.71 4.86 233.78 4.93 ;
    RECT 233.71 6.315 233.78 6.385 ;
    RECT 233.71 6.745 233.78 6.815 ;
    RECT 233.71 12.31 233.78 12.38 ;
    RECT 233.51 4.23 233.58 4.3 ;
    RECT 233.51 7.135 233.58 7.205 ;
    RECT 233.51 8.325 233.58 8.395 ;
    RECT 233.51 8.71 233.58 9.115 ;
    RECT 233.51 9.995 233.58 10.205 ;
    RECT 232.505 12.605 232.77 12.675 ;
    RECT 232.24 8.325 232.31 8.395 ;
    RECT 232.04 8.325 232.31 9.115 ;
    RECT 232.24 8.71 232.31 8.97 ;
    RECT 232.04 9.995 232.31 10.205 ;
    RECT 232.07 2.99 232.28 3.955 ;
    RECT 232.07 4.815 232.28 5.025 ;
    RECT 232.07 6.315 232.28 6.385 ;
    RECT 230.585 5.255 230.865 5.325 ;
    RECT 230.585 8.065 230.865 8.135 ;
    RECT 230.585 11.985 230.865 12.195 ;
    RECT 230.62 3.32 230.83 3.53 ;
    RECT 230.62 4.445 230.83 4.655 ;
    RECT 230.62 6.12 230.83 6.19 ;
    RECT 230.39 3.035 230.46 3.105 ;
    RECT 230.39 3.78 230.46 3.85 ;
    RECT 230.39 4.86 230.46 4.93 ;
    RECT 230.39 6.315 230.46 6.385 ;
    RECT 230.39 6.745 230.46 6.815 ;
    RECT 230.39 12.31 230.46 12.38 ;
    RECT 230.19 4.23 230.26 4.3 ;
    RECT 230.19 7.135 230.26 7.205 ;
    RECT 230.19 8.325 230.26 8.395 ;
    RECT 230.19 8.71 230.26 9.115 ;
    RECT 230.19 9.995 230.26 10.205 ;
    RECT 229.185 12.605 229.45 12.675 ;
    RECT 228.92 8.325 228.99 8.395 ;
    RECT 228.72 8.325 228.99 9.115 ;
    RECT 228.92 8.71 228.99 8.97 ;
    RECT 228.72 9.995 228.99 10.205 ;
    RECT 228.75 2.99 228.96 3.955 ;
    RECT 228.75 4.815 228.96 5.025 ;
    RECT 228.75 6.315 228.96 6.385 ;
    RECT 227.265 5.255 227.545 5.325 ;
    RECT 227.265 8.065 227.545 8.135 ;
    RECT 227.265 11.985 227.545 12.195 ;
    RECT 227.3 3.32 227.51 3.53 ;
    RECT 227.3 4.445 227.51 4.655 ;
    RECT 227.3 6.12 227.51 6.19 ;
    RECT 227.07 3.035 227.14 3.105 ;
    RECT 227.07 3.78 227.14 3.85 ;
    RECT 227.07 4.86 227.14 4.93 ;
    RECT 227.07 6.315 227.14 6.385 ;
    RECT 227.07 6.745 227.14 6.815 ;
    RECT 227.07 12.31 227.14 12.38 ;
    RECT 226.87 4.23 226.94 4.3 ;
    RECT 226.87 7.135 226.94 7.205 ;
    RECT 226.87 8.325 226.94 8.395 ;
    RECT 226.87 8.71 226.94 9.115 ;
    RECT 226.87 9.995 226.94 10.205 ;
    RECT 225.865 12.605 226.13 12.675 ;
    RECT 225.6 8.325 225.67 8.395 ;
    RECT 225.4 8.325 225.67 9.115 ;
    RECT 225.6 8.71 225.67 8.97 ;
    RECT 225.4 9.995 225.67 10.205 ;
    RECT 225.43 2.99 225.64 3.955 ;
    RECT 225.43 4.815 225.64 5.025 ;
    RECT 225.43 6.315 225.64 6.385 ;
    RECT 223.945 5.255 224.225 5.325 ;
    RECT 223.945 8.065 224.225 8.135 ;
    RECT 223.945 11.985 224.225 12.195 ;
    RECT 223.98 3.32 224.19 3.53 ;
    RECT 223.98 4.445 224.19 4.655 ;
    RECT 223.98 6.12 224.19 6.19 ;
    RECT 223.75 3.035 223.82 3.105 ;
    RECT 223.75 3.78 223.82 3.85 ;
    RECT 223.75 4.86 223.82 4.93 ;
    RECT 223.75 6.315 223.82 6.385 ;
    RECT 223.75 6.745 223.82 6.815 ;
    RECT 223.75 12.31 223.82 12.38 ;
    RECT 223.55 4.23 223.62 4.3 ;
    RECT 223.55 7.135 223.62 7.205 ;
    RECT 223.55 8.325 223.62 8.395 ;
    RECT 223.55 8.71 223.62 9.115 ;
    RECT 223.55 9.995 223.62 10.205 ;
    RECT 222.545 12.605 222.81 12.675 ;
    RECT 222.28 8.325 222.35 8.395 ;
    RECT 222.08 8.325 222.35 9.115 ;
    RECT 222.28 8.71 222.35 8.97 ;
    RECT 222.08 9.995 222.35 10.205 ;
    RECT 222.11 2.99 222.32 3.955 ;
    RECT 222.11 4.815 222.32 5.025 ;
    RECT 222.11 6.315 222.32 6.385 ;
    RECT 220.625 5.255 220.905 5.325 ;
    RECT 220.625 8.065 220.905 8.135 ;
    RECT 220.625 11.985 220.905 12.195 ;
    RECT 220.66 3.32 220.87 3.53 ;
    RECT 220.66 4.445 220.87 4.655 ;
    RECT 220.66 6.12 220.87 6.19 ;
    RECT 220.43 3.035 220.5 3.105 ;
    RECT 220.43 3.78 220.5 3.85 ;
    RECT 220.43 4.86 220.5 4.93 ;
    RECT 220.43 6.315 220.5 6.385 ;
    RECT 220.43 6.745 220.5 6.815 ;
    RECT 220.43 12.31 220.5 12.38 ;
    RECT 220.23 4.23 220.3 4.3 ;
    RECT 220.23 7.135 220.3 7.205 ;
    RECT 220.23 8.325 220.3 8.395 ;
    RECT 220.23 8.71 220.3 9.115 ;
    RECT 220.23 9.995 220.3 10.205 ;
    RECT 219.225 12.605 219.49 12.675 ;
    RECT 218.96 8.325 219.03 8.395 ;
    RECT 218.76 8.325 219.03 9.115 ;
    RECT 218.96 8.71 219.03 8.97 ;
    RECT 218.76 9.995 219.03 10.205 ;
    RECT 218.79 2.99 219.0 3.955 ;
    RECT 218.79 4.815 219.0 5.025 ;
    RECT 218.79 6.315 219.0 6.385 ;
    RECT 217.305 5.255 217.585 5.325 ;
    RECT 217.305 8.065 217.585 8.135 ;
    RECT 217.305 11.985 217.585 12.195 ;
    RECT 217.34 3.32 217.55 3.53 ;
    RECT 217.34 4.445 217.55 4.655 ;
    RECT 217.34 6.12 217.55 6.19 ;
    RECT 217.11 3.035 217.18 3.105 ;
    RECT 217.11 3.78 217.18 3.85 ;
    RECT 217.11 4.86 217.18 4.93 ;
    RECT 217.11 6.315 217.18 6.385 ;
    RECT 217.11 6.745 217.18 6.815 ;
    RECT 217.11 12.31 217.18 12.38 ;
    RECT 216.91 4.23 216.98 4.3 ;
    RECT 216.91 7.135 216.98 7.205 ;
    RECT 216.91 8.325 216.98 8.395 ;
    RECT 216.91 8.71 216.98 9.115 ;
    RECT 216.91 9.995 216.98 10.205 ;
    RECT 215.905 12.605 216.17 12.675 ;
    RECT 215.64 8.325 215.71 8.395 ;
    RECT 215.44 8.325 215.71 9.115 ;
    RECT 215.64 8.71 215.71 8.97 ;
    RECT 215.44 9.995 215.71 10.205 ;
    RECT 215.47 2.99 215.68 3.955 ;
    RECT 215.47 4.815 215.68 5.025 ;
    RECT 215.47 6.315 215.68 6.385 ;
    RECT 213.985 5.255 214.265 5.325 ;
    RECT 213.985 8.065 214.265 8.135 ;
    RECT 213.985 11.985 214.265 12.195 ;
    RECT 214.02 3.32 214.23 3.53 ;
    RECT 214.02 4.445 214.23 4.655 ;
    RECT 214.02 6.12 214.23 6.19 ;
    RECT 213.79 3.035 213.86 3.105 ;
    RECT 213.79 3.78 213.86 3.85 ;
    RECT 213.79 4.86 213.86 4.93 ;
    RECT 213.79 6.315 213.86 6.385 ;
    RECT 213.79 6.745 213.86 6.815 ;
    RECT 213.79 12.31 213.86 12.38 ;
    RECT 213.59 4.23 213.66 4.3 ;
    RECT 213.59 7.135 213.66 7.205 ;
    RECT 213.59 8.325 213.66 8.395 ;
    RECT 213.59 8.71 213.66 9.115 ;
    RECT 213.59 9.995 213.66 10.205 ;
    RECT 212.585 12.605 212.85 12.675 ;
    RECT 212.32 8.325 212.39 8.395 ;
    RECT 212.12 8.325 212.39 9.115 ;
    RECT 212.32 8.71 212.39 8.97 ;
    RECT 212.12 9.995 212.39 10.205 ;
    RECT 212.15 2.99 212.36 3.955 ;
    RECT 212.15 4.815 212.36 5.025 ;
    RECT 212.15 6.315 212.36 6.385 ;
    RECT 210.665 5.255 210.945 5.325 ;
    RECT 210.665 8.065 210.945 8.135 ;
    RECT 210.665 11.985 210.945 12.195 ;
    RECT 210.7 3.32 210.91 3.53 ;
    RECT 210.7 4.445 210.91 4.655 ;
    RECT 210.7 6.12 210.91 6.19 ;
    RECT 210.47 3.035 210.54 3.105 ;
    RECT 210.47 3.78 210.54 3.85 ;
    RECT 210.47 4.86 210.54 4.93 ;
    RECT 210.47 6.315 210.54 6.385 ;
    RECT 210.47 6.745 210.54 6.815 ;
    RECT 210.47 12.31 210.54 12.38 ;
    RECT 210.27 4.23 210.34 4.3 ;
    RECT 210.27 7.135 210.34 7.205 ;
    RECT 210.27 8.325 210.34 8.395 ;
    RECT 210.27 8.71 210.34 9.115 ;
    RECT 210.27 9.995 210.34 10.205 ;
    RECT 209.265 12.605 209.53 12.675 ;
    RECT 209.0 8.325 209.07 8.395 ;
    RECT 208.8 8.325 209.07 9.115 ;
    RECT 209.0 8.71 209.07 8.97 ;
    RECT 208.8 9.995 209.07 10.205 ;
    RECT 208.83 2.99 209.04 3.955 ;
    RECT 208.83 4.815 209.04 5.025 ;
    RECT 208.83 6.315 209.04 6.385 ;
    RECT 207.345 5.255 207.625 5.325 ;
    RECT 207.345 8.065 207.625 8.135 ;
    RECT 207.345 11.985 207.625 12.195 ;
    RECT 207.38 3.32 207.59 3.53 ;
    RECT 207.38 4.445 207.59 4.655 ;
    RECT 207.38 6.12 207.59 6.19 ;
    RECT 207.15 3.035 207.22 3.105 ;
    RECT 207.15 3.78 207.22 3.85 ;
    RECT 207.15 4.86 207.22 4.93 ;
    RECT 207.15 6.315 207.22 6.385 ;
    RECT 207.15 6.745 207.22 6.815 ;
    RECT 207.15 12.31 207.22 12.38 ;
    RECT 206.95 4.23 207.02 4.3 ;
    RECT 206.95 7.135 207.02 7.205 ;
    RECT 206.95 8.325 207.02 8.395 ;
    RECT 206.95 8.71 207.02 9.115 ;
    RECT 206.95 9.995 207.02 10.205 ;
    RECT 205.945 12.605 206.21 12.675 ;
    RECT 205.68 8.325 205.75 8.395 ;
    RECT 205.48 8.325 205.75 9.115 ;
    RECT 205.68 8.71 205.75 8.97 ;
    RECT 205.48 9.995 205.75 10.205 ;
    RECT 205.51 2.99 205.72 3.955 ;
    RECT 205.51 4.815 205.72 5.025 ;
    RECT 205.51 6.315 205.72 6.385 ;
    RECT 204.025 5.255 204.305 5.325 ;
    RECT 204.025 8.065 204.305 8.135 ;
    RECT 204.025 11.985 204.305 12.195 ;
    RECT 204.06 3.32 204.27 3.53 ;
    RECT 204.06 4.445 204.27 4.655 ;
    RECT 204.06 6.12 204.27 6.19 ;
    RECT 203.83 3.035 203.9 3.105 ;
    RECT 203.83 3.78 203.9 3.85 ;
    RECT 203.83 4.86 203.9 4.93 ;
    RECT 203.83 6.315 203.9 6.385 ;
    RECT 203.83 6.745 203.9 6.815 ;
    RECT 203.83 12.31 203.9 12.38 ;
    RECT 203.63 4.23 203.7 4.3 ;
    RECT 203.63 7.135 203.7 7.205 ;
    RECT 203.63 8.325 203.7 8.395 ;
    RECT 203.63 8.71 203.7 9.115 ;
    RECT 203.63 9.995 203.7 10.205 ;
    RECT 202.625 12.605 202.89 12.675 ;
    RECT 202.36 8.325 202.43 8.395 ;
    RECT 202.16 8.325 202.43 9.115 ;
    RECT 202.36 8.71 202.43 8.97 ;
    RECT 202.16 9.995 202.43 10.205 ;
    RECT 202.19 2.99 202.4 3.955 ;
    RECT 202.19 4.815 202.4 5.025 ;
    RECT 202.19 6.315 202.4 6.385 ;
    RECT 200.705 5.255 200.985 5.325 ;
    RECT 200.705 8.065 200.985 8.135 ;
    RECT 200.705 11.985 200.985 12.195 ;
    RECT 200.74 3.32 200.95 3.53 ;
    RECT 200.74 4.445 200.95 4.655 ;
    RECT 200.74 6.12 200.95 6.19 ;
    RECT 200.51 3.035 200.58 3.105 ;
    RECT 200.51 3.78 200.58 3.85 ;
    RECT 200.51 4.86 200.58 4.93 ;
    RECT 200.51 6.315 200.58 6.385 ;
    RECT 200.51 6.745 200.58 6.815 ;
    RECT 200.51 12.31 200.58 12.38 ;
    RECT 200.31 4.23 200.38 4.3 ;
    RECT 200.31 7.135 200.38 7.205 ;
    RECT 200.31 8.325 200.38 8.395 ;
    RECT 200.31 8.71 200.38 9.115 ;
    RECT 200.31 9.995 200.38 10.205 ;
    RECT 199.305 12.605 199.57 12.675 ;
    RECT 199.04 8.325 199.11 8.395 ;
    RECT 198.84 8.325 199.11 9.115 ;
    RECT 199.04 8.71 199.11 8.97 ;
    RECT 198.84 9.995 199.11 10.205 ;
    RECT 198.87 2.99 199.08 3.955 ;
    RECT 198.87 4.815 199.08 5.025 ;
    RECT 198.87 6.315 199.08 6.385 ;
    RECT 197.385 5.255 197.665 5.325 ;
    RECT 197.385 8.065 197.665 8.135 ;
    RECT 197.385 11.985 197.665 12.195 ;
    RECT 197.42 3.32 197.63 3.53 ;
    RECT 197.42 4.445 197.63 4.655 ;
    RECT 197.42 6.12 197.63 6.19 ;
    RECT 197.19 3.035 197.26 3.105 ;
    RECT 197.19 3.78 197.26 3.85 ;
    RECT 197.19 4.86 197.26 4.93 ;
    RECT 197.19 6.315 197.26 6.385 ;
    RECT 197.19 6.745 197.26 6.815 ;
    RECT 197.19 12.31 197.26 12.38 ;
    RECT 196.99 4.23 197.06 4.3 ;
    RECT 196.99 7.135 197.06 7.205 ;
    RECT 196.99 8.325 197.06 8.395 ;
    RECT 196.99 8.71 197.06 9.115 ;
    RECT 196.99 9.995 197.06 10.205 ;
    RECT 195.985 12.605 196.25 12.675 ;
    RECT 195.72 8.325 195.79 8.395 ;
    RECT 195.52 8.325 195.79 9.115 ;
    RECT 195.72 8.71 195.79 8.97 ;
    RECT 195.52 9.995 195.79 10.205 ;
    RECT 195.55 2.99 195.76 3.955 ;
    RECT 195.55 4.815 195.76 5.025 ;
    RECT 195.55 6.315 195.76 6.385 ;
    RECT 194.065 5.255 194.345 5.325 ;
    RECT 194.065 8.065 194.345 8.135 ;
    RECT 194.065 11.985 194.345 12.195 ;
    RECT 194.1 3.32 194.31 3.53 ;
    RECT 194.1 4.445 194.31 4.655 ;
    RECT 194.1 6.12 194.31 6.19 ;
    RECT 193.87 3.035 193.94 3.105 ;
    RECT 193.87 3.78 193.94 3.85 ;
    RECT 193.87 4.86 193.94 4.93 ;
    RECT 193.87 6.315 193.94 6.385 ;
    RECT 193.87 6.745 193.94 6.815 ;
    RECT 193.87 12.31 193.94 12.38 ;
    RECT 193.67 4.23 193.74 4.3 ;
    RECT 193.67 7.135 193.74 7.205 ;
    RECT 193.67 8.325 193.74 8.395 ;
    RECT 193.67 8.71 193.74 9.115 ;
    RECT 193.67 9.995 193.74 10.205 ;
    RECT 192.665 12.605 192.93 12.675 ;
    RECT 192.4 8.325 192.47 8.395 ;
    RECT 192.2 8.325 192.47 9.115 ;
    RECT 192.4 8.71 192.47 8.97 ;
    RECT 192.2 9.995 192.47 10.205 ;
    RECT 192.23 2.99 192.44 3.955 ;
    RECT 192.23 4.815 192.44 5.025 ;
    RECT 192.23 6.315 192.44 6.385 ;
    RECT 190.745 5.255 191.025 5.325 ;
    RECT 190.745 8.065 191.025 8.135 ;
    RECT 190.745 11.985 191.025 12.195 ;
    RECT 190.78 3.32 190.99 3.53 ;
    RECT 190.78 4.445 190.99 4.655 ;
    RECT 190.78 6.12 190.99 6.19 ;
    RECT 190.55 3.035 190.62 3.105 ;
    RECT 190.55 3.78 190.62 3.85 ;
    RECT 190.55 4.86 190.62 4.93 ;
    RECT 190.55 6.315 190.62 6.385 ;
    RECT 190.55 6.745 190.62 6.815 ;
    RECT 190.55 12.31 190.62 12.38 ;
    RECT 190.35 4.23 190.42 4.3 ;
    RECT 190.35 7.135 190.42 7.205 ;
    RECT 190.35 8.325 190.42 8.395 ;
    RECT 190.35 8.71 190.42 9.115 ;
    RECT 190.35 9.995 190.42 10.205 ;
    RECT 189.345 12.605 189.61 12.675 ;
    RECT 189.08 8.325 189.15 8.395 ;
    RECT 188.88 8.325 189.15 9.115 ;
    RECT 189.08 8.71 189.15 8.97 ;
    RECT 188.88 9.995 189.15 10.205 ;
    RECT 188.91 2.99 189.12 3.955 ;
    RECT 188.91 4.815 189.12 5.025 ;
    RECT 188.91 6.315 189.12 6.385 ;
    RECT 187.425 5.255 187.705 5.325 ;
    RECT 187.425 8.065 187.705 8.135 ;
    RECT 187.425 11.985 187.705 12.195 ;
    RECT 187.46 3.32 187.67 3.53 ;
    RECT 187.46 4.445 187.67 4.655 ;
    RECT 187.46 6.12 187.67 6.19 ;
    RECT 187.23 3.035 187.3 3.105 ;
    RECT 187.23 3.78 187.3 3.85 ;
    RECT 187.23 4.86 187.3 4.93 ;
    RECT 187.23 6.315 187.3 6.385 ;
    RECT 187.23 6.745 187.3 6.815 ;
    RECT 187.23 12.31 187.3 12.38 ;
    RECT 187.03 4.23 187.1 4.3 ;
    RECT 187.03 7.135 187.1 7.205 ;
    RECT 187.03 8.325 187.1 8.395 ;
    RECT 187.03 8.71 187.1 9.115 ;
    RECT 187.03 9.995 187.1 10.205 ;
    RECT 186.025 12.605 186.29 12.675 ;
    RECT 185.76 8.325 185.83 8.395 ;
    RECT 185.56 8.325 185.83 9.115 ;
    RECT 185.76 8.71 185.83 8.97 ;
    RECT 185.56 9.995 185.83 10.205 ;
    RECT 185.59 2.99 185.8 3.955 ;
    RECT 185.59 4.815 185.8 5.025 ;
    RECT 185.59 6.315 185.8 6.385 ;
    RECT 184.105 5.255 184.385 5.325 ;
    RECT 184.105 8.065 184.385 8.135 ;
    RECT 184.105 11.985 184.385 12.195 ;
    RECT 184.14 3.32 184.35 3.53 ;
    RECT 184.14 4.445 184.35 4.655 ;
    RECT 184.14 6.12 184.35 6.19 ;
    RECT 183.91 3.035 183.98 3.105 ;
    RECT 183.91 3.78 183.98 3.85 ;
    RECT 183.91 4.86 183.98 4.93 ;
    RECT 183.91 6.315 183.98 6.385 ;
    RECT 183.91 6.745 183.98 6.815 ;
    RECT 183.91 12.31 183.98 12.38 ;
    RECT 183.71 4.23 183.78 4.3 ;
    RECT 183.71 7.135 183.78 7.205 ;
    RECT 183.71 8.325 183.78 8.395 ;
    RECT 183.71 8.71 183.78 9.115 ;
    RECT 183.71 9.995 183.78 10.205 ;
    RECT 182.705 12.605 182.97 12.675 ;
    RECT 182.44 8.325 182.51 8.395 ;
    RECT 182.24 8.325 182.51 9.115 ;
    RECT 182.44 8.71 182.51 8.97 ;
    RECT 182.24 9.995 182.51 10.205 ;
    RECT 182.27 2.99 182.48 3.955 ;
    RECT 182.27 4.815 182.48 5.025 ;
    RECT 182.27 6.315 182.48 6.385 ;
    RECT 179.9 7.565 180.11 7.635 ;
    RECT 176.58 7.565 176.79 7.635 ;
    RECT 173.26 7.565 173.47 7.635 ;
    RECT 173.26 6.315 173.47 6.385 ;
    RECT 173.26 4.815 173.47 5.025 ;
    RECT 173.26 3.742 173.47 3.952 ;
    RECT 173.26 2.99 173.47 3.2 ;
    RECT 169.94 7.565 170.15 7.635 ;
    RECT 169.94 9.995 170.15 10.205 ;
    RECT 166.62 7.565 166.83 7.635 ;
    RECT 169.94 8.902 170.15 9.112 ;
    RECT 256.26 6.315 256.47 6.385 ;
    RECT 169.94 8.705 170.15 8.775 ;
    RECT 256.26 4.815 256.47 5.025 ;
    RECT 169.94 8.325 170.15 8.395 ;
    RECT 256.26 3.742 256.47 3.952 ;
    RECT 169.94 6.315 170.15 6.385 ;
    RECT 256.26 2.99 256.47 3.2 ;
    RECT 169.94 4.815 170.15 5.025 ;
    RECT 163.3 7.565 163.51 7.635 ;
    RECT 252.94 9.995 253.15 10.205 ;
    RECT 252.94 8.902 253.15 9.112 ;
    RECT 252.94 8.705 253.15 8.775 ;
    RECT 252.94 8.325 253.15 8.395 ;
    RECT 252.94 6.315 253.15 6.385 ;
    RECT 252.94 4.815 253.15 5.025 ;
    RECT 169.94 3.742 170.15 3.952 ;
    RECT 169.94 2.99 170.15 3.2 ;
    RECT 159.98 7.565 160.19 7.635 ;
    RECT 223.55 6.12 223.62 6.19 ;
    RECT 166.62 9.995 166.83 10.205 ;
    RECT 223.55 5.182 223.62 5.392 ;
    RECT 166.62 8.902 166.83 9.112 ;
    RECT 223.55 4.445 223.62 4.655 ;
    RECT 166.62 8.705 166.83 8.775 ;
    RECT 166.62 8.325 166.83 8.395 ;
    RECT 252.94 3.742 253.15 3.952 ;
    RECT 166.62 6.315 166.83 6.385 ;
    RECT 252.94 2.99 253.15 3.2 ;
    RECT 156.66 7.565 156.87 7.635 ;
    RECT 223.98 7.125 224.19 7.195 ;
    RECT 166.62 4.815 166.83 5.025 ;
    RECT 223.98 4.22 224.19 4.29 ;
    RECT 166.62 3.742 166.83 3.952 ;
    RECT 166.62 2.99 166.83 3.2 ;
    RECT 200.74 4.22 200.95 4.29 ;
    RECT 249.62 9.995 249.83 10.205 ;
    RECT 249.62 8.902 249.83 9.112 ;
    RECT 249.62 8.705 249.83 8.775 ;
    RECT 213.1 9.995 213.31 10.205 ;
    RECT 249.62 8.325 249.83 8.395 ;
    RECT 213.1 8.902 213.31 9.112 ;
    RECT 249.62 6.315 249.83 6.385 ;
    RECT 213.1 8.705 213.31 8.775 ;
    RECT 249.62 4.815 249.83 5.025 ;
    RECT 196.99 6.12 197.06 6.19 ;
    RECT 213.1 8.325 213.31 8.395 ;
    RECT 249.62 3.742 249.83 3.952 ;
    RECT 196.99 5.182 197.06 5.392 ;
    RECT 213.1 6.315 213.31 6.385 ;
    RECT 249.62 2.99 249.83 3.2 ;
    RECT 196.99 4.445 197.06 4.655 ;
    RECT 213.1 4.815 213.31 5.025 ;
    RECT 213.1 3.742 213.31 3.952 ;
    RECT 213.1 2.99 213.31 3.2 ;
    RECT 197.42 7.125 197.63 7.195 ;
    RECT 197.42 4.22 197.63 4.29 ;
    RECT 153.34 7.565 153.55 7.635 ;
    RECT 163.3 9.995 163.51 10.205 ;
    RECT 220.23 6.12 220.3 6.19 ;
    RECT 163.3 8.902 163.51 9.112 ;
    RECT 220.23 5.182 220.3 5.392 ;
    RECT 163.3 8.705 163.51 8.775 ;
    RECT 209.78 9.995 209.99 10.205 ;
    RECT 220.23 4.445 220.3 4.655 ;
    RECT 163.3 8.325 163.51 8.395 ;
    RECT 209.78 8.902 209.99 9.112 ;
    RECT 163.3 6.315 163.51 6.385 ;
    RECT 163.3 4.815 163.51 5.025 ;
    RECT 220.66 7.125 220.87 7.195 ;
    RECT 163.3 3.742 163.51 3.952 ;
    RECT 220.66 4.22 220.87 4.29 ;
    RECT 163.3 2.99 163.51 3.2 ;
    RECT 150.02 7.565 150.23 7.635 ;
    RECT 159.98 9.995 160.19 10.205 ;
    RECT 159.98 8.902 160.19 9.112 ;
    RECT 216.91 6.12 216.98 6.19 ;
    RECT 209.78 8.705 209.99 8.775 ;
    RECT 209.78 8.325 209.99 8.395 ;
    RECT 193.67 6.12 193.74 6.19 ;
    RECT 209.78 6.315 209.99 6.385 ;
    RECT 193.67 5.182 193.74 5.392 ;
    RECT 209.78 4.815 209.99 5.025 ;
    RECT 193.67 4.445 193.74 4.655 ;
    RECT 209.78 3.742 209.99 3.952 ;
    RECT 209.78 2.99 209.99 3.2 ;
    RECT 194.1 7.125 194.31 7.195 ;
    RECT 194.1 4.22 194.31 4.29 ;
    RECT 159.98 8.705 160.19 8.775 ;
    RECT 206.46 9.995 206.67 10.205 ;
    RECT 216.91 5.182 216.98 5.392 ;
    RECT 159.98 8.325 160.19 8.395 ;
    RECT 206.46 8.902 206.67 9.112 ;
    RECT 216.91 4.445 216.98 4.655 ;
    RECT 159.98 6.315 160.19 6.385 ;
    RECT 206.46 8.705 206.67 8.775 ;
    RECT 159.98 4.815 160.19 5.025 ;
    RECT 206.46 8.325 206.67 8.395 ;
    RECT 159.98 3.742 160.19 3.952 ;
    RECT 217.34 7.125 217.55 7.195 ;
    RECT 159.98 2.99 160.19 3.2 ;
    RECT 217.34 4.22 217.55 4.29 ;
    RECT 160.47 6.12 160.54 6.19 ;
    RECT 160.47 5.182 160.54 5.392 ;
    RECT 160.47 4.445 160.54 4.655 ;
    RECT 160.9 7.125 161.11 7.195 ;
    RECT 160.9 4.22 161.11 4.29 ;
    RECT 156.66 9.995 156.87 10.205 ;
    RECT 246.3 7.565 246.51 7.635 ;
    RECT 156.66 8.902 156.87 9.112 ;
    RECT 156.66 8.705 156.87 8.775 ;
    RECT 156.66 8.325 156.87 8.395 ;
    RECT 206.46 6.315 206.67 6.385 ;
    RECT 190.35 6.12 190.42 6.19 ;
    RECT 206.46 4.815 206.67 5.025 ;
    RECT 190.35 5.182 190.42 5.392 ;
    RECT 206.46 3.742 206.67 3.952 ;
    RECT 190.35 4.445 190.42 4.655 ;
    RECT 206.46 2.99 206.67 3.2 ;
    RECT 190.78 7.125 190.99 7.195 ;
    RECT 190.78 4.22 190.99 4.29 ;
    RECT 242.98 7.565 243.19 7.635 ;
    RECT 203.14 9.995 203.35 10.205 ;
    RECT 203.14 8.902 203.35 9.112 ;
    RECT 156.66 6.315 156.87 6.385 ;
    RECT 203.14 8.705 203.35 8.775 ;
    RECT 156.66 4.815 156.87 5.025 ;
    RECT 203.14 8.325 203.35 8.395 ;
    RECT 156.66 3.742 156.87 3.952 ;
    RECT 203.14 6.315 203.35 6.385 ;
    RECT 156.66 2.99 156.87 3.2 ;
    RECT 203.14 4.815 203.35 5.025 ;
    RECT 239.66 7.565 239.87 7.635 ;
    RECT 157.15 6.12 157.22 6.19 ;
    RECT 157.15 5.182 157.22 5.392 ;
    RECT 157.15 4.445 157.22 4.655 ;
    RECT 157.58 7.125 157.79 7.195 ;
    RECT 157.58 4.22 157.79 4.29 ;
    RECT 153.34 9.995 153.55 10.205 ;
    RECT 153.34 8.902 153.55 9.112 ;
    RECT 153.34 8.705 153.55 8.775 ;
    RECT 153.34 8.325 153.55 8.395 ;
    RECT 236.34 7.565 236.55 7.635 ;
    RECT 153.34 6.315 153.55 6.385 ;
    RECT 187.03 6.12 187.1 6.19 ;
    RECT 153.34 4.815 153.55 5.025 ;
    RECT 203.14 3.742 203.35 3.952 ;
    RECT 187.03 5.182 187.1 5.392 ;
    RECT 203.14 2.99 203.35 3.2 ;
    RECT 187.03 4.445 187.1 4.655 ;
    RECT 187.46 7.125 187.67 7.195 ;
    RECT 213.1 7.565 213.31 7.635 ;
    RECT 187.46 4.22 187.67 4.29 ;
    RECT 233.02 7.565 233.23 7.635 ;
    RECT 199.82 9.995 200.03 10.205 ;
    RECT 199.82 8.902 200.03 9.112 ;
    RECT 199.82 8.705 200.03 8.775 ;
    RECT 199.82 8.325 200.03 8.395 ;
    RECT 199.82 6.315 200.03 6.385 ;
    RECT 209.78 7.565 209.99 7.635 ;
    RECT 153.34 3.742 153.55 3.952 ;
    RECT 199.82 4.815 200.03 5.025 ;
    RECT 153.34 2.99 153.55 3.2 ;
    RECT 199.82 3.742 200.03 3.952 ;
    RECT 183.71 6.12 183.78 6.19 ;
    RECT 199.82 2.99 200.03 3.2 ;
    RECT 266.71 6.12 266.78 6.19 ;
    RECT 266.71 5.182 266.78 5.392 ;
    RECT 229.7 7.565 229.91 7.635 ;
    RECT 266.71 4.445 266.78 4.655 ;
    RECT 153.83 6.12 153.9 6.19 ;
    RECT 153.83 5.182 153.9 5.392 ;
    RECT 153.83 4.445 153.9 4.655 ;
    RECT 267.14 7.125 267.35 7.195 ;
    RECT 154.26 7.125 154.47 7.195 ;
    RECT 154.26 4.22 154.47 4.29 ;
    RECT 206.46 7.565 206.67 7.635 ;
    RECT 150.02 9.995 150.23 10.205 ;
    RECT 150.02 8.902 150.23 9.112 ;
    RECT 150.02 8.705 150.23 8.775 ;
    RECT 150.02 8.325 150.23 8.395 ;
    RECT 150.02 6.315 150.23 6.385 ;
    RECT 150.02 4.815 150.23 5.025 ;
    RECT 150.02 3.742 150.23 3.952 ;
    RECT 183.71 5.182 183.78 5.392 ;
    RECT 150.02 2.99 150.23 3.2 ;
    RECT 226.38 7.565 226.59 7.635 ;
    RECT 183.71 4.445 183.78 4.655 ;
    RECT 184.14 7.125 184.35 7.195 ;
    RECT 184.14 4.22 184.35 4.29 ;
    RECT 203.14 7.565 203.35 7.635 ;
    RECT 150.51 6.12 150.58 6.19 ;
    RECT 267.14 4.22 267.35 4.29 ;
    RECT 196.5 9.995 196.71 10.205 ;
    RECT 196.5 8.902 196.71 9.112 ;
    RECT 223.06 7.565 223.27 7.635 ;
    RECT 196.5 8.705 196.71 8.775 ;
    RECT 196.5 8.325 196.71 8.395 ;
    RECT 196.5 6.315 196.71 6.385 ;
    RECT 196.5 4.815 196.71 5.025 ;
    RECT 196.5 3.742 196.71 3.952 ;
    RECT 196.5 2.99 196.71 3.2 ;
    RECT 199.82 7.565 200.03 7.635 ;
    RECT 263.39 6.12 263.46 6.19 ;
    RECT 263.39 5.182 263.46 5.392 ;
    RECT 263.39 4.445 263.46 4.655 ;
    RECT 150.51 5.182 150.58 5.392 ;
    RECT 150.51 4.445 150.58 4.655 ;
    RECT 263.82 7.125 264.03 7.195 ;
    RECT 263.82 4.22 264.03 4.29 ;
    RECT 150.94 7.125 151.15 7.195 ;
    RECT 150.94 4.22 151.15 4.29 ;
    RECT 193.18 9.995 193.39 10.205 ;
    RECT 193.18 8.902 193.39 9.112 ;
    RECT 196.5 7.565 196.71 7.635 ;
    RECT 219.74 7.565 219.95 7.635 ;
    RECT 193.18 7.565 193.39 7.635 ;
    RECT 193.18 8.705 193.39 8.775 ;
    RECT 193.18 8.325 193.39 8.395 ;
    RECT 193.18 6.315 193.39 6.385 ;
    RECT 193.18 4.815 193.39 5.025 ;
    RECT 193.18 3.742 193.39 3.952 ;
    RECT 193.18 2.99 193.39 3.2 ;
    RECT 216.42 7.565 216.63 7.635 ;
    RECT 189.86 7.565 190.07 7.635 ;
    RECT 260.07 6.12 260.14 6.19 ;
    RECT 260.07 5.182 260.14 5.392 ;
    RECT 260.07 4.445 260.14 4.655 ;
    RECT 260.5 7.125 260.71 7.195 ;
    RECT 260.5 4.22 260.71 4.29 ;
    RECT 237.26 7.125 237.47 7.195 ;
    RECT 237.26 4.22 237.47 4.29 ;
    RECT 189.86 9.995 190.07 10.205 ;
    RECT 189.86 8.902 190.07 9.112 ;
    RECT 189.86 8.705 190.07 8.775 ;
    RECT 189.86 8.325 190.07 8.395 ;
    RECT 233.51 6.12 233.58 6.19 ;
    RECT 233.51 5.182 233.58 5.392 ;
    RECT 233.51 4.445 233.58 4.655 ;
    RECT 233.94 7.125 234.15 7.195 ;
    RECT 189.86 6.315 190.07 6.385 ;
    RECT 189.86 4.815 190.07 5.025 ;
    RECT 186.54 7.565 186.75 7.635 ;
    RECT 189.86 3.742 190.07 3.952 ;
    RECT 189.86 2.99 190.07 3.2 ;
    RECT 256.75 6.12 256.82 6.19 ;
    RECT 256.75 5.182 256.82 5.392 ;
    RECT 256.75 4.445 256.82 4.655 ;
    RECT 257.18 7.125 257.39 7.195 ;
    RECT 257.18 4.22 257.39 4.29 ;
    RECT 183.22 7.565 183.43 7.635 ;
    RECT 233.94 4.22 234.15 4.29 ;
    RECT 186.54 9.995 186.75 10.205 ;
    RECT 186.54 8.902 186.75 9.112 ;
    RECT 186.54 8.705 186.75 8.775 ;
    RECT 186.54 8.325 186.75 8.395 ;
    RECT 186.54 6.315 186.75 6.385 ;
    RECT 186.54 4.815 186.75 5.025 ;
    RECT 230.19 6.12 230.26 6.19 ;
    RECT 230.19 5.182 230.26 5.392 ;
    RECT 230.19 4.445 230.26 4.655 ;
    RECT 230.62 7.125 230.83 7.195 ;
    RECT 230.62 4.22 230.83 4.29 ;
    RECT 186.54 3.742 186.75 3.952 ;
    RECT 186.54 2.99 186.75 3.2 ;
    RECT 253.43 6.12 253.5 6.19 ;
    RECT 253.43 5.182 253.5 5.392 ;
    RECT 253.43 4.445 253.5 4.655 ;
    RECT 253.86 7.125 254.07 7.195 ;
    RECT 253.86 4.22 254.07 4.29 ;
    RECT 183.22 9.995 183.43 10.205 ;
    RECT 183.22 8.902 183.43 9.112 ;
    RECT 246.3 9.995 246.51 10.205 ;
    RECT 183.22 8.705 183.43 8.775 ;
    RECT 246.3 8.902 246.51 9.112 ;
    RECT 183.22 8.325 183.43 8.395 ;
    RECT 246.3 8.705 246.51 8.775 ;
    RECT 183.22 6.315 183.43 6.385 ;
    RECT 246.3 8.325 246.51 8.395 ;
    RECT 183.22 4.815 183.43 5.025 ;
    RECT 246.3 6.315 246.51 6.385 ;
    RECT 183.22 3.742 183.43 3.952 ;
    RECT 246.3 4.815 246.51 5.025 ;
    RECT 183.22 2.99 183.43 3.2 ;
    RECT 246.3 3.742 246.51 3.952 ;
    RECT 246.3 2.99 246.51 3.2 ;
    RECT 250.11 6.12 250.18 6.19 ;
    RECT 226.87 6.12 226.94 6.19 ;
    RECT 226.87 5.182 226.94 5.392 ;
    RECT 226.87 4.445 226.94 4.655 ;
    RECT 227.3 7.125 227.51 7.195 ;
    RECT 227.3 4.22 227.51 4.29 ;
    RECT 242.98 9.995 243.19 10.205 ;
    RECT 242.98 8.902 243.19 9.112 ;
    RECT 250.11 5.182 250.18 5.392 ;
    RECT 250.11 4.445 250.18 4.655 ;
    RECT 250.54 7.125 250.75 7.195 ;
    RECT 250.54 4.22 250.75 4.29 ;
    RECT 242.98 8.705 243.19 8.775 ;
    RECT 242.98 8.325 243.19 8.395 ;
    RECT 242.98 6.315 243.19 6.385 ;
    RECT 213.59 6.12 213.66 6.19 ;
    RECT 242.98 4.815 243.19 5.025 ;
    RECT 213.59 5.182 213.66 5.392 ;
    RECT 242.98 3.742 243.19 3.952 ;
    RECT 242.98 2.99 243.19 3.2 ;
    RECT 239.66 9.995 239.87 10.205 ;
    RECT 239.66 8.902 239.87 9.112 ;
    RECT 239.66 8.705 239.87 8.775 ;
    RECT 239.66 8.325 239.87 8.395 ;
    RECT 213.59 4.445 213.66 4.655 ;
    RECT 214.02 7.125 214.23 7.195 ;
    RECT 214.02 4.22 214.23 4.29 ;
    RECT 180.39 6.12 180.46 6.19 ;
    RECT 180.39 5.182 180.46 5.392 ;
    RECT 239.66 6.315 239.87 6.385 ;
    RECT 239.66 4.815 239.87 5.025 ;
    RECT 210.27 6.12 210.34 6.19 ;
    RECT 179.9 9.995 180.11 10.205 ;
    RECT 239.66 3.742 239.87 3.952 ;
    RECT 210.27 5.182 210.34 5.392 ;
    RECT 179.9 8.902 180.11 9.112 ;
    RECT 239.66 2.99 239.87 3.2 ;
    RECT 210.27 4.445 210.34 4.655 ;
    RECT 179.9 8.705 180.11 8.775 ;
    RECT 179.9 8.325 180.11 8.395 ;
    RECT 179.9 6.315 180.11 6.385 ;
    RECT 179.9 4.815 180.11 5.025 ;
    RECT 179.9 3.742 180.11 3.952 ;
    RECT 179.9 2.99 180.11 3.2 ;
    RECT 180.39 4.445 180.46 4.655 ;
    RECT 180.82 7.125 181.03 7.195 ;
    RECT 180.82 4.22 181.03 4.29 ;
    RECT 236.34 9.995 236.55 10.205 ;
    RECT 236.34 8.902 236.55 9.112 ;
    RECT 236.34 8.705 236.55 8.775 ;
    RECT 236.34 8.325 236.55 8.395 ;
    RECT 236.34 6.315 236.55 6.385 ;
    RECT 236.34 4.815 236.55 5.025 ;
    RECT 176.58 9.995 176.79 10.205 ;
    RECT 176.58 8.902 176.79 9.112 ;
    RECT 210.7 7.125 210.91 7.195 ;
    RECT 210.7 4.22 210.91 4.29 ;
    RECT 177.07 6.12 177.14 6.19 ;
    RECT 177.07 5.182 177.14 5.392 ;
    RECT 177.07 4.445 177.14 4.655 ;
    RECT 236.34 3.742 236.55 3.952 ;
    RECT 206.95 6.12 207.02 6.19 ;
    RECT 236.34 2.99 236.55 3.2 ;
    RECT 206.95 5.182 207.02 5.392 ;
    RECT 176.58 8.705 176.79 8.775 ;
    RECT 206.95 4.445 207.02 4.655 ;
    RECT 176.58 8.325 176.79 8.395 ;
    RECT 176.58 6.315 176.79 6.385 ;
    RECT 176.58 4.815 176.79 5.025 ;
    RECT 176.58 3.742 176.79 3.952 ;
    RECT 176.58 2.99 176.79 3.2 ;
    RECT 177.5 7.125 177.71 7.195 ;
    RECT 177.5 4.22 177.71 4.29 ;
    RECT 233.02 9.995 233.23 10.205 ;
    RECT 233.02 8.902 233.23 9.112 ;
    RECT 233.02 8.705 233.23 8.775 ;
    RECT 233.02 8.325 233.23 8.395 ;
    RECT 233.02 6.315 233.23 6.385 ;
    RECT 233.02 4.815 233.23 5.025 ;
    RECT 173.26 9.995 173.47 10.205 ;
    RECT 233.02 3.742 233.23 3.952 ;
    RECT 173.26 8.902 173.47 9.112 ;
    RECT 233.02 2.99 233.23 3.2 ;
    RECT 173.26 8.705 173.47 8.775 ;
    RECT 173.26 8.325 173.47 8.395 ;
    RECT 207.38 7.125 207.59 7.195 ;
    RECT 207.38 4.22 207.59 4.29 ;
    RECT 173.75 6.12 173.82 6.19 ;
    RECT 173.75 5.182 173.82 5.392 ;
    RECT 173.75 4.445 173.82 4.655 ;
    RECT 203.63 6.12 203.7 6.19 ;
    RECT 203.63 5.182 203.7 5.392 ;
    RECT 203.63 4.445 203.7 4.655 ;
    RECT 174.18 7.125 174.39 7.195 ;
    RECT 174.18 4.22 174.39 4.29 ;
    RECT 229.7 9.995 229.91 10.205 ;
    RECT 229.7 8.902 229.91 9.112 ;
    RECT 229.7 8.705 229.91 8.775 ;
    RECT 229.7 8.325 229.91 8.395 ;
    RECT 229.7 6.315 229.91 6.385 ;
    RECT 229.7 4.815 229.91 5.025 ;
    RECT 229.7 3.742 229.91 3.952 ;
    RECT 229.7 2.99 229.91 3.2 ;
    RECT 204.06 7.125 204.27 7.195 ;
    RECT 204.06 4.22 204.27 4.29 ;
    RECT 170.43 6.12 170.5 6.19 ;
    RECT 170.43 5.182 170.5 5.392 ;
    RECT 170.43 4.445 170.5 4.655 ;
    RECT 226.38 9.995 226.59 10.205 ;
    RECT 226.38 8.902 226.59 9.112 ;
    RECT 200.31 6.12 200.38 6.19 ;
    RECT 200.31 5.182 200.38 5.392 ;
    RECT 200.31 4.445 200.38 4.655 ;
    RECT 200.74 7.125 200.95 7.195 ;
    RECT 170.86 7.125 171.07 7.195 ;
    RECT 170.86 4.22 171.07 4.29 ;
    RECT 226.38 8.705 226.59 8.775 ;
    RECT 226.38 8.325 226.59 8.395 ;
    RECT 226.38 6.315 226.59 6.385 ;
    RECT 226.38 4.815 226.59 5.025 ;
    RECT 226.38 3.742 226.59 3.952 ;
    RECT 226.38 2.99 226.59 3.2 ;
    RECT 167.11 6.12 167.18 6.19 ;
    RECT 167.11 5.182 167.18 5.392 ;
    RECT 167.11 4.445 167.18 4.655 ;
    RECT 167.54 7.125 167.75 7.195 ;
    RECT 223.06 9.995 223.27 10.205 ;
    RECT 223.06 8.902 223.27 9.112 ;
    RECT 223.06 8.705 223.27 8.775 ;
    RECT 223.06 8.325 223.27 8.395 ;
    RECT 167.54 4.22 167.75 4.29 ;
    RECT 223.06 6.315 223.27 6.385 ;
    RECT 223.06 4.815 223.27 5.025 ;
    RECT 223.06 3.742 223.27 3.952 ;
    RECT 223.06 2.99 223.27 3.2 ;
    RECT 163.79 6.12 163.86 6.19 ;
    RECT 163.79 5.182 163.86 5.392 ;
    RECT 163.79 4.445 163.86 4.655 ;
    RECT 164.22 7.125 164.43 7.195 ;
    RECT 219.74 9.995 219.95 10.205 ;
    RECT 164.22 4.22 164.43 4.29 ;
    RECT 219.74 8.902 219.95 9.112 ;
    RECT 219.74 8.705 219.95 8.775 ;
    RECT 219.74 8.325 219.95 8.395 ;
    RECT 219.74 6.315 219.95 6.385 ;
    RECT 219.74 4.815 219.95 5.025 ;
    RECT 219.74 3.742 219.95 3.952 ;
    RECT 219.74 2.99 219.95 3.2 ;
    RECT 266.22 9.995 266.43 10.205 ;
    RECT 266.22 8.902 266.43 9.112 ;
    RECT 216.42 9.995 216.63 10.205 ;
    RECT 266.22 8.705 266.43 8.775 ;
    RECT 216.42 8.902 216.63 9.112 ;
    RECT 266.22 8.325 266.43 8.395 ;
    RECT 216.42 8.705 216.63 8.775 ;
    RECT 266.22 6.315 266.43 6.385 ;
    RECT 216.42 8.325 216.63 8.395 ;
    RECT 266.22 4.815 266.43 5.025 ;
    RECT 216.42 6.315 216.63 6.385 ;
    RECT 266.22 3.742 266.43 3.952 ;
    RECT 216.42 4.815 216.63 5.025 ;
    RECT 266.22 2.99 266.43 3.2 ;
    RECT 216.42 3.742 216.63 3.952 ;
    RECT 216.42 2.99 216.63 3.2 ;
    RECT 246.79 6.12 246.86 6.19 ;
    RECT 246.79 5.182 246.86 5.392 ;
    RECT 245.35 0.775 245.56 0.845 ;
    RECT 198.87 0.775 199.08 0.845 ;
    RECT 199.82 1.775 200.03 1.985 ;
    RECT 199.82 1.15 200.03 1.36 ;
    RECT 165.67 0.775 165.88 0.845 ;
    RECT 166.62 1.775 166.83 1.985 ;
    RECT 166.62 1.15 166.83 1.36 ;
    RECT 246.3 1.775 246.51 1.985 ;
    RECT 246.3 1.15 246.51 1.36 ;
    RECT 195.55 0.775 195.76 0.845 ;
    RECT 162.35 0.775 162.56 0.845 ;
    RECT 242.03 0.775 242.24 0.845 ;
    RECT 242.98 1.775 243.19 1.985 ;
    RECT 242.98 1.15 243.19 1.36 ;
    RECT 196.5 1.775 196.71 1.985 ;
    RECT 196.5 1.15 196.71 1.36 ;
    RECT 163.3 1.775 163.51 1.985 ;
    RECT 163.3 1.15 163.51 1.36 ;
    RECT 238.71 0.775 238.92 0.845 ;
    RECT 192.23 0.775 192.44 0.845 ;
    RECT 193.18 1.775 193.39 1.985 ;
    RECT 193.18 1.15 193.39 1.36 ;
    RECT 159.03 0.775 159.24 0.845 ;
    RECT 159.98 1.775 160.19 1.985 ;
    RECT 159.98 1.15 160.19 1.36 ;
    RECT 239.66 1.775 239.87 1.985 ;
    RECT 239.66 1.15 239.87 1.36 ;
    RECT 188.91 0.775 189.12 0.845 ;
    RECT 155.71 0.775 155.92 0.845 ;
    RECT 235.39 0.775 235.6 0.845 ;
    RECT 236.34 1.775 236.55 1.985 ;
    RECT 236.34 1.15 236.55 1.36 ;
    RECT 189.86 1.775 190.07 1.985 ;
    RECT 189.86 1.15 190.07 1.36 ;
    RECT 156.66 1.775 156.87 1.985 ;
    RECT 156.66 1.15 156.87 1.36 ;
    RECT 185.59 0.775 185.8 0.845 ;
    RECT 186.54 1.775 186.75 1.985 ;
    RECT 186.54 1.15 186.75 1.36 ;
    RECT 152.39 0.775 152.6 0.845 ;
    RECT 232.07 0.775 232.28 0.845 ;
    RECT 153.34 1.775 153.55 1.985 ;
    RECT 153.34 1.15 153.55 1.36 ;
    RECT 233.02 1.775 233.23 1.985 ;
    RECT 233.02 1.15 233.23 1.36 ;
    RECT 265.27 0.775 265.48 0.845 ;
    RECT 266.22 1.775 266.43 1.985 ;
    RECT 266.22 1.15 266.43 1.36 ;
    RECT 228.75 0.775 228.96 0.845 ;
    RECT 182.27 0.775 182.48 0.845 ;
    RECT 183.22 1.775 183.43 1.985 ;
    RECT 183.22 1.15 183.43 1.36 ;
    RECT 149.07 0.775 149.28 0.845 ;
    RECT 150.02 1.775 150.23 1.985 ;
    RECT 150.02 1.15 150.23 1.36 ;
    RECT 229.7 1.775 229.91 1.985 ;
    RECT 229.7 1.15 229.91 1.36 ;
    RECT 261.95 0.775 262.16 0.845 ;
    RECT 262.9 1.775 263.11 1.985 ;
    RECT 262.9 1.15 263.11 1.36 ;
    RECT 225.43 0.775 225.64 0.845 ;
    RECT 226.38 1.775 226.59 1.985 ;
    RECT 226.38 1.15 226.59 1.36 ;
    RECT 263.82 1.465 264.03 1.675 ;
    RECT 263.4 0.98 263.47 1.05 ;
    RECT 262.9 0.775 263.11 0.845 ;
    RECT 261.95 1.15 262.16 1.985 ;
    RECT 260.5 1.465 260.71 1.675 ;
    RECT 260.08 0.98 260.15 1.05 ;
    RECT 259.58 0.775 259.79 0.845 ;
    RECT 258.63 1.15 258.84 1.985 ;
    RECT 257.18 1.465 257.39 1.675 ;
    RECT 256.76 0.98 256.83 1.05 ;
    RECT 256.26 0.775 256.47 0.845 ;
    RECT 255.31 1.15 255.52 1.985 ;
    RECT 253.86 1.465 254.07 1.675 ;
    RECT 253.44 0.98 253.51 1.05 ;
    RECT 252.94 0.775 253.15 0.845 ;
    RECT 251.99 1.15 252.2 1.985 ;
    RECT 250.54 1.465 250.75 1.675 ;
    RECT 250.12 0.98 250.19 1.05 ;
    RECT 249.62 0.775 249.83 0.845 ;
    RECT 248.67 1.15 248.88 1.985 ;
    RECT 267.14 1.465 267.35 1.675 ;
    RECT 266.72 0.98 266.79 1.05 ;
    RECT 266.22 0.775 266.43 0.845 ;
    RECT 265.27 1.15 265.48 1.985 ;
    RECT 258.63 0.775 258.84 0.845 ;
    RECT 259.58 1.775 259.79 1.985 ;
    RECT 259.58 1.15 259.79 1.36 ;
    RECT 150.94 1.465 151.15 1.675 ;
    RECT 150.52 0.98 150.59 1.05 ;
    RECT 150.02 0.775 150.23 0.845 ;
    RECT 149.07 1.15 149.28 1.985 ;
    RECT 247.22 1.465 247.43 1.675 ;
    RECT 246.8 0.98 246.87 1.05 ;
    RECT 246.3 0.775 246.51 0.845 ;
    RECT 245.35 1.15 245.56 1.985 ;
    RECT 222.11 0.775 222.32 0.845 ;
    RECT 243.9 1.465 244.11 1.675 ;
    RECT 243.48 0.98 243.55 1.05 ;
    RECT 242.98 0.775 243.19 0.845 ;
    RECT 242.03 1.15 242.24 1.985 ;
    RECT 240.58 1.465 240.79 1.675 ;
    RECT 240.16 0.98 240.23 1.05 ;
    RECT 239.66 0.775 239.87 0.845 ;
    RECT 238.71 1.15 238.92 1.985 ;
    RECT 237.26 1.465 237.47 1.675 ;
    RECT 236.84 0.98 236.91 1.05 ;
    RECT 236.34 0.775 236.55 0.845 ;
    RECT 235.39 1.15 235.6 1.985 ;
    RECT 233.94 1.465 234.15 1.675 ;
    RECT 233.52 0.98 233.59 1.05 ;
    RECT 233.02 0.775 233.23 0.845 ;
    RECT 232.07 1.15 232.28 1.985 ;
    RECT 230.62 1.465 230.83 1.675 ;
    RECT 230.2 0.98 230.27 1.05 ;
    RECT 229.7 0.775 229.91 0.845 ;
    RECT 228.75 1.15 228.96 1.985 ;
    RECT 227.3 1.465 227.51 1.675 ;
    RECT 226.88 0.98 226.95 1.05 ;
    RECT 226.38 0.775 226.59 0.845 ;
    RECT 225.43 1.15 225.64 1.985 ;
    RECT 223.98 1.465 224.19 1.675 ;
    RECT 223.56 0.98 223.63 1.05 ;
    RECT 223.06 0.775 223.27 0.845 ;
    RECT 222.11 1.15 222.32 1.985 ;
    RECT 220.66 1.465 220.87 1.675 ;
    RECT 220.24 0.98 220.31 1.05 ;
    RECT 219.74 0.775 219.95 0.845 ;
    RECT 218.79 1.15 219.0 1.985 ;
    RECT 217.34 1.465 217.55 1.675 ;
    RECT 216.92 0.98 216.99 1.05 ;
    RECT 216.42 0.775 216.63 0.845 ;
    RECT 215.47 1.15 215.68 1.985 ;
    RECT 180.82 1.465 181.03 1.675 ;
    RECT 180.4 0.98 180.47 1.05 ;
    RECT 179.9 0.775 180.11 0.845 ;
    RECT 178.95 1.15 179.16 1.985 ;
    RECT 177.5 1.465 177.71 1.675 ;
    RECT 177.08 0.98 177.15 1.05 ;
    RECT 176.58 0.775 176.79 0.845 ;
    RECT 175.63 1.15 175.84 1.985 ;
    RECT 174.18 1.465 174.39 1.675 ;
    RECT 173.76 0.98 173.83 1.05 ;
    RECT 173.26 0.775 173.47 0.845 ;
    RECT 172.31 1.15 172.52 1.985 ;
    RECT 170.86 1.465 171.07 1.675 ;
    RECT 170.44 0.98 170.51 1.05 ;
    RECT 169.94 0.775 170.15 0.845 ;
    RECT 168.99 1.15 169.2 1.985 ;
    RECT 167.54 1.465 167.75 1.675 ;
    RECT 167.12 0.98 167.19 1.05 ;
    RECT 166.62 0.775 166.83 0.845 ;
    RECT 165.67 1.15 165.88 1.985 ;
    RECT 164.22 1.465 164.43 1.675 ;
    RECT 163.8 0.98 163.87 1.05 ;
    RECT 163.3 0.775 163.51 0.845 ;
    RECT 162.35 1.15 162.56 1.985 ;
    RECT 160.9 1.465 161.11 1.675 ;
    RECT 160.48 0.98 160.55 1.05 ;
    RECT 159.98 0.775 160.19 0.845 ;
    RECT 159.03 1.15 159.24 1.985 ;
    RECT 157.58 1.465 157.79 1.675 ;
    RECT 157.16 0.98 157.23 1.05 ;
    RECT 156.66 0.775 156.87 0.845 ;
    RECT 155.71 1.15 155.92 1.985 ;
    RECT 154.26 1.465 154.47 1.675 ;
    RECT 153.84 0.98 153.91 1.05 ;
    RECT 153.34 0.775 153.55 0.845 ;
    RECT 152.39 1.15 152.6 1.985 ;
    RECT 223.06 1.775 223.27 1.985 ;
    RECT 223.06 1.15 223.27 1.36 ;
    RECT 255.31 0.775 255.52 0.845 ;
    RECT 214.02 1.465 214.23 1.675 ;
    RECT 213.6 0.98 213.67 1.05 ;
    RECT 213.1 0.775 213.31 0.845 ;
    RECT 212.15 1.15 212.36 1.985 ;
    RECT 210.7 1.465 210.91 1.675 ;
    RECT 210.28 0.98 210.35 1.05 ;
    RECT 209.78 0.775 209.99 0.845 ;
    RECT 208.83 1.15 209.04 1.985 ;
    RECT 207.38 1.465 207.59 1.675 ;
    RECT 206.96 0.98 207.03 1.05 ;
    RECT 206.46 0.775 206.67 0.845 ;
    RECT 205.51 1.15 205.72 1.985 ;
    RECT 204.06 1.465 204.27 1.675 ;
    RECT 203.64 0.98 203.71 1.05 ;
    RECT 203.14 0.775 203.35 0.845 ;
    RECT 202.19 1.15 202.4 1.985 ;
    RECT 200.74 1.465 200.95 1.675 ;
    RECT 200.32 0.98 200.39 1.05 ;
    RECT 199.82 0.775 200.03 0.845 ;
    RECT 198.87 1.15 199.08 1.985 ;
    RECT 197.42 1.465 197.63 1.675 ;
    RECT 197.0 0.98 197.07 1.05 ;
    RECT 196.5 0.775 196.71 0.845 ;
    RECT 195.55 1.15 195.76 1.985 ;
    RECT 194.1 1.465 194.31 1.675 ;
    RECT 193.68 0.98 193.75 1.05 ;
    RECT 193.18 0.775 193.39 0.845 ;
    RECT 192.23 1.15 192.44 1.985 ;
    RECT 190.78 1.465 190.99 1.675 ;
    RECT 190.36 0.98 190.43 1.05 ;
    RECT 189.86 0.775 190.07 0.845 ;
    RECT 188.91 1.15 189.12 1.985 ;
    RECT 187.46 1.465 187.67 1.675 ;
    RECT 187.04 0.98 187.11 1.05 ;
    RECT 186.54 0.775 186.75 0.845 ;
    RECT 185.59 1.15 185.8 1.985 ;
    RECT 184.14 1.465 184.35 1.675 ;
    RECT 183.72 0.98 183.79 1.05 ;
    RECT 183.22 0.775 183.43 0.845 ;
    RECT 182.27 1.15 182.48 1.985 ;
    RECT 256.26 1.775 256.47 1.985 ;
    RECT 256.26 1.15 256.47 1.36 ;
    RECT 212.15 0.775 212.36 0.845 ;
    RECT 218.79 0.775 219.0 0.845 ;
    RECT 219.74 1.775 219.95 1.985 ;
    RECT 219.74 1.15 219.95 1.36 ;
    RECT 178.95 0.775 179.16 0.845 ;
    RECT 213.1 1.775 213.31 1.985 ;
    RECT 213.1 1.15 213.31 1.36 ;
    RECT 251.99 0.775 252.2 0.845 ;
    RECT 252.94 1.775 253.15 1.985 ;
    RECT 252.94 1.15 253.15 1.36 ;
    RECT 179.9 1.775 180.11 1.985 ;
    RECT 179.9 1.15 180.11 1.36 ;
    RECT 208.83 0.775 209.04 0.845 ;
    RECT 209.78 1.775 209.99 1.985 ;
    RECT 209.78 1.15 209.99 1.36 ;
    RECT 215.47 0.775 215.68 0.845 ;
    RECT 216.42 1.775 216.63 1.985 ;
    RECT 216.42 1.15 216.63 1.36 ;
    RECT 175.63 0.775 175.84 0.845 ;
    RECT 176.58 1.775 176.79 1.985 ;
    RECT 176.58 1.15 176.79 1.36 ;
    RECT 248.67 0.775 248.88 0.845 ;
    RECT 249.62 1.775 249.83 1.985 ;
    RECT 249.62 1.15 249.83 1.36 ;
    RECT 205.51 0.775 205.72 0.845 ;
    RECT 172.31 0.775 172.52 0.845 ;
    RECT 206.46 1.775 206.67 1.985 ;
    RECT 206.46 1.15 206.67 1.36 ;
    RECT 173.26 1.775 173.47 1.985 ;
    RECT 173.26 1.15 173.47 1.36 ;
    RECT 202.19 0.775 202.4 0.845 ;
    RECT 203.14 1.775 203.35 1.985 ;
    RECT 203.14 1.15 203.35 1.36 ;
    RECT 168.99 0.775 169.2 0.845 ;
    RECT 169.94 1.775 170.15 1.985 ;
    RECT 169.94 1.15 170.15 1.36 ;
    RECT 253.4 14.23 253.61 14.3 ;
    RECT 212.61 13.71 212.82 13.78 ;
    RECT 199.33 13.97 199.54 14.04 ;
    RECT 219.25 13.97 219.46 14.04 ;
    RECT 169.45 13.97 169.66 14.04 ;
    RECT 225.89 13.71 226.1 13.78 ;
    RECT 209.78 14.23 209.99 14.3 ;
    RECT 214.015 13.45 214.235 13.52 ;
    RECT 210.24 14.23 210.45 14.3 ;
    RECT 210.695 13.45 210.915 13.52 ;
    RECT 207.375 13.45 207.595 13.52 ;
    RECT 204.055 13.45 204.275 13.52 ;
    RECT 200.735 13.45 200.955 13.52 ;
    RECT 197.415 13.45 197.635 13.52 ;
    RECT 233.02 14.23 233.23 14.3 ;
    RECT 194.095 13.45 194.315 13.52 ;
    RECT 233.48 14.23 233.69 14.3 ;
    RECT 190.775 13.45 190.995 13.52 ;
    RECT 159.49 13.71 159.7 13.78 ;
    RECT 187.455 13.45 187.675 13.52 ;
    RECT 184.135 13.45 184.355 13.52 ;
    RECT 150.02 14.23 150.23 14.3 ;
    RECT 150.48 14.23 150.69 14.3 ;
    RECT 173.26 14.23 173.47 14.3 ;
    RECT 265.73 13.97 265.94 14.04 ;
    RECT 173.72 14.23 173.93 14.3 ;
    RECT 205.97 13.71 206.18 13.78 ;
    RECT 186.54 14.23 186.75 14.3 ;
    RECT 187.0 14.23 187.21 14.3 ;
    RECT 182.73 13.71 182.94 13.78 ;
    RECT 162.81 13.97 163.02 14.04 ;
    RECT 249.13 13.71 249.34 13.78 ;
    RECT 245.81 13.97 246.02 14.04 ;
    RECT 226.38 14.23 226.59 14.3 ;
    RECT 226.84 14.23 227.05 14.3 ;
    RECT 192.69 13.97 192.9 14.04 ;
    RECT 166.62 14.23 166.83 14.3 ;
    RECT 167.08 14.23 167.29 14.3 ;
    RECT 199.33 13.71 199.54 13.78 ;
    RECT 219.25 13.71 219.46 13.78 ;
    RECT 262.9 14.23 263.11 14.3 ;
    RECT 263.36 14.23 263.57 14.3 ;
    RECT 203.14 14.23 203.35 14.3 ;
    RECT 203.6 14.23 203.81 14.3 ;
    RECT 242.49 13.71 242.7 13.78 ;
    RECT 152.85 13.71 153.06 13.78 ;
    RECT 239.17 13.97 239.38 14.04 ;
    RECT 259.09 13.97 259.3 14.04 ;
    RECT 176.09 13.71 176.3 13.78 ;
    RECT 265.73 13.71 265.94 13.78 ;
    RECT 242.98 14.23 243.19 14.3 ;
    RECT 186.05 13.97 186.26 14.04 ;
    RECT 243.44 14.23 243.65 14.3 ;
    RECT 159.98 14.23 160.19 14.3 ;
    RECT 160.44 14.23 160.65 14.3 ;
    RECT 192.69 13.71 192.9 13.78 ;
    RECT 209.29 13.97 209.5 14.04 ;
    RECT 179.41 13.97 179.62 14.04 ;
    RECT 196.5 14.23 196.71 14.3 ;
    RECT 156.17 13.97 156.38 14.04 ;
    RECT 196.96 14.23 197.17 14.3 ;
    RECT 235.85 13.71 236.06 13.78 ;
    RECT 180.815 13.45 181.035 13.52 ;
    RECT 219.74 14.23 219.95 14.3 ;
    RECT 177.495 13.45 177.715 13.52 ;
    RECT 220.2 14.23 220.41 14.3 ;
    RECT 174.175 13.45 174.395 13.52 ;
    RECT 170.855 13.45 171.075 13.52 ;
    RECT 252.45 13.97 252.66 14.04 ;
    RECT 167.535 13.45 167.755 13.52 ;
    RECT 232.53 13.97 232.74 14.04 ;
    RECT 164.215 13.45 164.435 13.52 ;
    RECT 160.895 13.45 161.115 13.52 ;
    RECT 157.575 13.45 157.795 13.52 ;
    RECT 169.45 13.71 169.66 13.78 ;
    RECT 154.255 13.45 154.475 13.52 ;
    RECT 259.09 13.71 259.3 13.78 ;
    RECT 150.935 13.45 151.155 13.52 ;
    RECT 256.26 14.23 256.47 14.3 ;
    RECT 256.72 14.23 256.93 14.3 ;
    RECT 176.58 14.23 176.79 14.3 ;
    RECT 177.04 14.23 177.25 14.3 ;
    RECT 202.65 13.97 202.86 14.04 ;
    RECT 222.57 13.97 222.78 14.04 ;
    RECT 172.77 13.97 172.98 14.04 ;
    RECT 149.53 13.97 149.74 14.04 ;
    RECT 229.21 13.71 229.42 13.78 ;
    RECT 213.1 14.23 213.31 14.3 ;
    RECT 213.56 14.23 213.77 14.3 ;
    RECT 236.34 14.23 236.55 14.3 ;
    RECT 236.8 14.23 237.01 14.3 ;
    RECT 162.81 13.71 163.02 13.78 ;
    RECT 153.34 14.23 153.55 14.3 ;
    RECT 153.8 14.23 154.01 14.3 ;
    RECT 249.62 14.23 249.83 14.3 ;
    RECT 250.08 14.23 250.29 14.3 ;
    RECT 209.29 13.71 209.5 13.78 ;
    RECT 189.86 14.23 190.07 14.3 ;
    RECT 190.32 14.23 190.53 14.3 ;
    RECT 186.05 13.71 186.26 13.78 ;
    RECT 225.89 13.97 226.1 14.04 ;
    RECT 196.01 13.97 196.22 14.04 ;
    RECT 215.93 13.97 216.14 14.04 ;
    RECT 166.13 13.97 166.34 14.04 ;
    RECT 252.45 13.71 252.66 13.78 ;
    RECT 222.57 13.71 222.78 13.78 ;
    RECT 229.7 14.23 229.91 14.3 ;
    RECT 156.17 13.71 156.38 13.78 ;
    RECT 230.16 14.23 230.37 14.3 ;
    RECT 262.41 13.97 262.62 14.04 ;
    RECT 169.94 14.23 170.15 14.3 ;
    RECT 170.4 14.23 170.61 14.3 ;
    RECT 202.65 13.71 202.86 13.78 ;
    RECT 183.22 14.23 183.43 14.3 ;
    RECT 266.22 14.23 266.43 14.3 ;
    RECT 183.68 14.23 183.89 14.3 ;
    RECT 266.68 14.23 266.89 14.3 ;
    RECT 206.46 14.23 206.67 14.3 ;
    RECT 206.92 14.23 207.13 14.3 ;
    RECT 245.81 13.71 246.02 13.78 ;
    RECT 242.49 13.97 242.7 14.04 ;
    RECT 179.41 13.71 179.62 13.78 ;
    RECT 246.3 14.23 246.51 14.3 ;
    RECT 246.76 14.23 246.97 14.3 ;
    RECT 189.37 13.97 189.58 14.04 ;
    RECT 163.3 14.23 163.51 14.3 ;
    RECT 163.76 14.23 163.97 14.3 ;
    RECT 196.01 13.71 196.22 13.78 ;
    RECT 215.93 13.71 216.14 13.78 ;
    RECT 212.61 13.97 212.82 14.04 ;
    RECT 259.58 14.23 259.79 14.3 ;
    RECT 260.04 14.23 260.25 14.3 ;
    RECT 199.82 14.23 200.03 14.3 ;
    RECT 200.28 14.23 200.49 14.3 ;
    RECT 239.17 13.71 239.38 13.78 ;
    RECT 159.49 13.97 159.7 14.04 ;
    RECT 149.53 13.71 149.74 13.78 ;
    RECT 223.06 14.23 223.27 14.3 ;
    RECT 223.52 14.23 223.73 14.3 ;
    RECT 235.85 13.97 236.06 14.04 ;
    RECT 255.77 13.97 255.98 14.04 ;
    RECT 172.77 13.71 172.98 13.78 ;
    RECT 262.41 13.71 262.62 13.78 ;
    RECT 267.135 13.45 267.355 13.52 ;
    RECT 263.815 13.45 264.035 13.52 ;
    RECT 260.495 13.45 260.715 13.52 ;
    RECT 257.175 13.45 257.395 13.52 ;
    RECT 182.73 13.97 182.94 14.04 ;
    RECT 253.855 13.45 254.075 13.52 ;
    RECT 250.535 13.45 250.755 13.52 ;
    RECT 189.37 13.71 189.58 13.78 ;
    RECT 179.9 14.23 180.11 14.3 ;
    RECT 180.36 14.23 180.57 14.3 ;
    RECT 205.97 13.97 206.18 14.04 ;
    RECT 176.09 13.97 176.3 14.04 ;
    RECT 193.18 14.23 193.39 14.3 ;
    RECT 232.53 13.71 232.74 13.78 ;
    RECT 152.85 13.97 153.06 14.04 ;
    RECT 193.64 14.23 193.85 14.3 ;
    RECT 216.42 14.23 216.63 14.3 ;
    RECT 216.88 14.23 217.09 14.3 ;
    RECT 239.66 14.23 239.87 14.3 ;
    RECT 229.21 13.97 229.42 14.04 ;
    RECT 249.13 13.97 249.34 14.04 ;
    RECT 240.12 14.23 240.33 14.3 ;
    RECT 247.215 13.45 247.435 13.52 ;
    RECT 243.895 13.45 244.115 13.52 ;
    RECT 166.13 13.71 166.34 13.78 ;
    RECT 240.575 13.45 240.795 13.52 ;
    RECT 156.66 14.23 156.87 14.3 ;
    RECT 255.77 13.71 255.98 13.78 ;
    RECT 237.255 13.45 237.475 13.52 ;
    RECT 157.12 14.23 157.33 14.3 ;
    RECT 233.935 13.45 234.155 13.52 ;
    RECT 230.615 13.45 230.835 13.52 ;
    RECT 227.295 13.45 227.515 13.52 ;
    RECT 223.975 13.45 224.195 13.52 ;
    RECT 220.655 13.45 220.875 13.52 ;
    RECT 252.94 14.23 253.15 14.3 ;
    RECT 217.335 13.45 217.555 13.52 ;
    RECT 141.415 7.565 141.625 7.635 ;
    RECT 140.895 12.302 140.965 12.372 ;
    RECT 140.895 6.707 140.965 6.777 ;
    RECT 140.895 1.807 140.965 1.877 ;
    RECT 120.615 13.45 120.685 13.52 ;
    RECT 120.615 11.985 120.685 12.195 ;
    RECT 120.615 7.972 120.685 8.182 ;
    RECT 120.615 6.12 120.685 6.19 ;
    RECT 120.615 4.445 120.685 4.655 ;
    RECT 134.34 4.815 134.55 5.025 ;
    RECT 129.15 1.465 129.22 1.675 ;
    RECT 134.34 2.99 134.55 3.2 ;
    RECT 128.715 8.972 128.925 9.042 ;
    RECT 128.715 3.777 128.925 3.847 ;
    RECT 134.34 1.15 134.55 1.36 ;
    RECT 139.73 7.565 139.94 7.635 ;
    RECT 136.92 7.565 137.13 7.635 ;
    RECT 120.615 3.32 120.685 3.53 ;
    RECT 120.615 1.465 120.685 1.675 ;
    RECT 131.795 11.435 131.865 11.505 ;
    RECT 134.34 7.565 134.55 7.635 ;
    RECT 131.795 7.565 131.865 7.635 ;
    RECT 130.595 10.31 130.665 10.38 ;
    RECT 130.595 6.707 130.665 6.777 ;
    RECT 130.595 1.807 130.665 1.877 ;
    RECT 128.335 14.23 128.545 14.3 ;
    RECT 128.335 7.565 128.545 7.635 ;
    RECT 126.76 14.23 126.97 14.3 ;
    RECT 131.795 11.06 131.865 11.13 ;
    RECT 131.795 8.325 131.865 8.395 ;
    RECT 126.76 7.565 126.97 7.635 ;
    RECT 131.795 6.315 131.865 6.385 ;
    RECT 131.795 4.815 131.865 5.025 ;
    RECT 131.795 2.99 131.865 3.2 ;
    RECT 131.795 1.15 131.865 1.36 ;
    RECT 125.11 14.23 125.32 14.3 ;
    RECT 125.11 7.565 125.32 7.635 ;
    RECT 124.255 14.23 124.465 14.3 ;
    RECT 131.0 10.31 131.21 10.38 ;
    RECT 124.255 7.565 124.465 7.635 ;
    RECT 131.0 6.707 131.21 6.777 ;
    RECT 131.0 1.807 131.21 1.877 ;
    RECT 122.04 14.23 122.25 14.3 ;
    RECT 122.04 7.565 122.25 7.635 ;
    RECT 129.965 10.31 130.175 10.38 ;
    RECT 129.965 6.707 130.175 6.777 ;
    RECT 129.965 1.807 130.175 1.877 ;
    RECT 121.44 14.23 121.51 14.3 ;
    RECT 121.44 12.82 121.51 13.03 ;
    RECT 121.44 7.565 121.51 7.635 ;
    RECT 128.335 11.435 128.545 11.505 ;
    RECT 121.44 2.615 121.51 2.685 ;
    RECT 128.335 11.06 128.545 11.13 ;
    RECT 128.335 9.94 128.545 10.01 ;
    RECT 128.335 8.325 128.545 8.395 ;
    RECT 127.69 12.302 127.9 12.372 ;
    RECT 127.69 9.507 127.9 9.577 ;
    RECT 127.69 6.707 127.9 6.777 ;
    RECT 127.69 1.807 127.9 1.877 ;
    RECT 126.76 9.94 126.97 10.01 ;
    RECT 126.76 6.315 126.97 6.385 ;
    RECT 126.76 4.815 126.97 5.025 ;
    RECT 126.76 2.99 126.97 3.2 ;
    RECT 126.76 1.15 126.97 1.36 ;
    RECT 147.695 13.45 147.765 13.52 ;
    RECT 147.695 11.985 147.765 12.195 ;
    RECT 147.695 7.972 147.765 8.182 ;
    RECT 147.695 6.12 147.765 6.19 ;
    RECT 125.11 9.995 125.32 10.205 ;
    RECT 125.11 6.315 125.32 6.385 ;
    RECT 125.11 4.815 125.32 5.025 ;
    RECT 125.11 2.99 125.32 3.2 ;
    RECT 125.11 1.15 125.32 1.36 ;
    RECT 147.695 3.32 147.765 3.53 ;
    RECT 147.695 1.465 147.765 1.675 ;
    RECT 146.765 7.125 146.975 7.195 ;
    RECT 146.765 4.22 146.975 4.29 ;
    RECT 145.87 7.125 145.94 7.195 ;
    RECT 145.87 4.22 145.94 4.29 ;
    RECT 124.255 9.995 124.465 10.205 ;
    RECT 124.255 6.315 124.465 6.385 ;
    RECT 124.255 4.815 124.465 5.025 ;
    RECT 124.255 2.99 124.465 3.2 ;
    RECT 124.255 1.15 124.465 1.36 ;
    RECT 143.31 7.125 143.52 7.195 ;
    RECT 143.31 4.22 143.52 4.29 ;
    RECT 122.63 12.82 122.84 13.03 ;
    RECT 122.63 12.302 122.84 12.372 ;
    RECT 141.935 7.125 142.145 7.195 ;
    RECT 141.935 4.22 142.145 4.29 ;
    RECT 132.25 13.085 132.32 13.155 ;
    RECT 122.63 6.707 122.84 6.777 ;
    RECT 122.63 4.515 122.84 4.585 ;
    RECT 122.63 1.807 122.84 1.877 ;
    RECT 122.04 9.995 122.25 10.205 ;
    RECT 146.16 9.995 146.37 10.205 ;
    RECT 122.04 8.705 122.25 8.775 ;
    RECT 122.04 6.315 122.25 6.385 ;
    RECT 122.04 4.815 122.25 5.025 ;
    RECT 122.04 2.99 122.25 3.2 ;
    RECT 122.04 1.15 122.25 1.36 ;
    RECT 138.72 7.125 138.93 7.195 ;
    RECT 138.72 4.22 138.93 4.29 ;
    RECT 146.16 8.902 146.37 9.112 ;
    RECT 146.16 8.705 146.37 8.775 ;
    RECT 146.16 8.325 146.37 8.395 ;
    RECT 146.16 6.315 146.37 6.385 ;
    RECT 146.16 4.815 146.37 5.025 ;
    RECT 146.16 2.99 146.37 3.2 ;
    RECT 146.16 1.15 146.37 1.36 ;
    RECT 138.37 11.985 138.44 12.195 ;
    RECT 138.37 7.972 138.44 8.182 ;
    RECT 138.37 6.12 138.44 6.19 ;
    RECT 138.37 5.51 138.44 5.58 ;
    RECT 138.37 3.32 138.44 3.53 ;
    RECT 121.44 9.995 121.51 10.205 ;
    RECT 121.44 8.705 121.51 8.775 ;
    RECT 121.44 6.315 121.51 6.385 ;
    RECT 121.44 4.815 121.51 5.025 ;
    RECT 145.485 12.82 145.695 13.03 ;
    RECT 121.44 2.99 121.51 3.2 ;
    RECT 145.485 12.302 145.695 12.372 ;
    RECT 121.44 1.15 121.51 1.36 ;
    RECT 138.37 1.465 138.44 1.675 ;
    RECT 137.625 7.125 137.695 7.195 ;
    RECT 137.625 4.22 137.695 4.29 ;
    RECT 136.535 7.125 136.745 7.195 ;
    RECT 136.535 4.22 136.745 4.29 ;
    RECT 145.485 6.707 145.695 6.777 ;
    RECT 120.615 2.76 120.685 2.83 ;
    RECT 120.615 13.025 120.685 13.095 ;
    RECT 120.62 4.22 120.69 4.29 ;
    RECT 120.62 7.125 120.69 7.195 ;
    RECT 120.62 9.72 120.69 9.79 ;
    RECT 120.825 7.57 120.895 7.64 ;
    RECT 120.825 14.23 120.895 14.3 ;
    RECT 120.835 2.615 120.905 2.685 ;
    RECT 121.035 5.915 121.105 5.985 ;
    RECT 121.035 11.805 121.105 11.875 ;
    RECT 121.035 13.97 121.105 14.04 ;
    RECT 121.44 1.81 121.51 1.88 ;
    RECT 121.44 4.515 121.51 4.585 ;
    RECT 121.44 6.705 121.51 6.775 ;
    RECT 121.44 14.47 121.51 14.54 ;
    RECT 121.635 3.63 121.705 3.84 ;
    RECT 121.67 11.435 121.88 11.505 ;
    RECT 121.785 2.66 121.855 2.87 ;
    RECT 121.785 5.61 121.855 5.82 ;
    RECT 121.785 9.555 121.855 9.625 ;
    RECT 122.04 1.81 122.25 1.88 ;
    RECT 122.04 4.515 122.25 4.585 ;
    RECT 122.04 6.705 122.25 6.775 ;
    RECT 122.04 12.305 122.25 13.03 ;
    RECT 122.395 1.465 122.465 1.535 ;
    RECT 122.395 1.605 122.465 1.675 ;
    RECT 122.395 3.32 122.465 3.39 ;
    RECT 122.395 3.46 122.465 3.53 ;
    RECT 122.395 6.12 122.465 6.19 ;
    RECT 122.395 7.975 122.465 8.045 ;
    RECT 122.395 8.115 122.465 8.185 ;
    RECT 122.395 11.985 122.465 12.055 ;
    RECT 122.395 12.125 122.465 12.195 ;
    RECT 122.395 13.45 122.465 13.52 ;
    RECT 122.63 1.15 122.84 1.36 ;
    RECT 122.63 2.99 122.84 3.2 ;
    RECT 122.63 4.815 122.84 5.025 ;
    RECT 122.63 6.315 122.84 6.385 ;
    RECT 122.63 8.705 122.84 8.775 ;
    RECT 122.63 9.995 122.84 10.205 ;
    RECT 123.215 12.885 124.0 12.955 ;
    RECT 124.255 1.81 124.465 1.88 ;
    RECT 124.255 4.515 124.465 4.585 ;
    RECT 124.255 6.705 124.465 6.775 ;
    RECT 124.255 9.51 124.465 9.58 ;
    RECT 124.255 12.305 124.465 12.375 ;
    RECT 124.715 1.465 124.925 1.675 ;
    RECT 124.715 3.32 124.925 3.53 ;
    RECT 124.715 6.12 124.925 6.19 ;
    RECT 124.715 7.975 124.925 8.185 ;
    RECT 124.715 11.985 124.925 12.195 ;
    RECT 125.11 1.81 125.32 1.88 ;
    RECT 125.11 4.515 125.32 4.585 ;
    RECT 125.11 6.705 125.32 6.775 ;
    RECT 125.11 9.51 125.32 9.58 ;
    RECT 125.11 12.305 125.32 12.375 ;
    RECT 125.645 12.885 125.905 12.955 ;
    RECT 125.67 12.6 125.88 12.67 ;
    RECT 126.38 10.23 126.59 10.3 ;
    RECT 126.735 12.895 126.995 12.965 ;
    RECT 126.76 1.81 126.97 1.88 ;
    RECT 126.76 4.515 126.97 4.585 ;
    RECT 126.76 6.705 126.97 6.775 ;
    RECT 126.76 9.51 126.97 9.58 ;
    RECT 126.76 12.305 126.97 12.375 ;
    RECT 127.125 3.775 127.195 3.845 ;
    RECT 127.32 1.465 127.53 1.675 ;
    RECT 127.32 3.32 127.53 3.53 ;
    RECT 127.32 6.12 127.53 6.19 ;
    RECT 127.32 7.975 127.53 8.185 ;
    RECT 127.32 11.985 127.53 12.195 ;
    RECT 127.395 10.13 127.465 10.34 ;
    RECT 127.675 12.885 127.915 12.955 ;
    RECT 127.69 1.15 127.9 1.36 ;
    RECT 127.69 2.99 127.9 3.2 ;
    RECT 127.69 4.815 127.9 5.025 ;
    RECT 127.69 6.315 127.9 6.385 ;
    RECT 127.69 8.325 127.9 8.395 ;
    RECT 127.69 9.94 127.9 10.01 ;
    RECT 127.69 11.06 127.9 11.13 ;
    RECT 127.69 11.435 127.9 11.505 ;
    RECT 128.105 1.465 128.175 1.535 ;
    RECT 128.105 1.605 128.175 1.675 ;
    RECT 128.105 3.32 128.175 3.39 ;
    RECT 128.105 3.46 128.175 3.53 ;
    RECT 128.105 6.12 128.175 6.19 ;
    RECT 128.105 7.975 128.175 8.045 ;
    RECT 128.105 8.115 128.175 8.185 ;
    RECT 128.105 10.13 128.175 10.2 ;
    RECT 128.105 10.27 128.175 10.34 ;
    RECT 128.105 11.985 128.175 12.195 ;
    RECT 128.335 6.705 128.545 6.775 ;
    RECT 128.335 9.51 128.545 9.58 ;
    RECT 128.335 12.305 128.545 12.375 ;
    RECT 128.355 4.435 128.565 4.505 ;
    RECT 128.355 5.915 128.565 5.985 ;
    RECT 128.715 1.465 128.925 1.675 ;
    RECT 128.715 3.32 128.925 3.53 ;
    RECT 128.715 6.12 128.925 6.19 ;
    RECT 128.715 7.975 128.925 8.185 ;
    RECT 128.715 10.13 128.925 10.2 ;
    RECT 128.715 11.985 128.925 12.195 ;
    RECT 129.115 3.775 129.185 3.845 ;
    RECT 129.15 8.975 129.22 9.045 ;
    RECT 129.445 1.465 129.655 1.675 ;
    RECT 129.445 3.32 129.655 3.53 ;
    RECT 129.445 6.12 129.655 6.19 ;
    RECT 129.445 7.975 129.655 8.185 ;
    RECT 129.445 10.13 129.655 10.2 ;
    RECT 129.445 11.985 129.655 12.195 ;
    RECT 129.965 1.15 130.175 1.36 ;
    RECT 129.965 2.99 130.175 3.2 ;
    RECT 129.965 4.815 130.175 5.025 ;
    RECT 129.965 6.315 130.175 6.385 ;
    RECT 129.965 8.325 130.175 8.395 ;
    RECT 129.965 9.94 130.175 10.01 ;
    RECT 129.965 11.06 130.175 11.13 ;
    RECT 129.965 11.435 130.175 11.505 ;
    RECT 130.335 10.87 130.405 10.94 ;
    RECT 130.335 12.305 130.405 12.375 ;
    RECT 130.595 0.845 130.665 0.915 ;
    RECT 130.595 7.565 130.665 7.635 ;
    RECT 130.595 13.99 130.665 14.06 ;
    RECT 131.0 1.15 131.21 1.36 ;
    RECT 131.0 2.99 131.21 3.2 ;
    RECT 131.0 4.815 131.21 5.025 ;
    RECT 131.0 6.315 131.21 6.385 ;
    RECT 131.0 8.325 131.21 8.395 ;
    RECT 131.0 9.94 131.21 10.01 ;
    RECT 131.0 11.06 131.21 11.13 ;
    RECT 131.0 11.435 131.21 11.505 ;
    RECT 131.415 1.465 131.625 1.675 ;
    RECT 131.415 3.32 131.625 3.53 ;
    RECT 131.415 6.12 131.625 6.19 ;
    RECT 131.415 7.975 131.625 8.185 ;
    RECT 131.415 11.985 131.625 12.195 ;
    RECT 131.795 1.81 131.865 1.88 ;
    RECT 131.795 6.705 131.865 6.775 ;
    RECT 131.795 10.31 131.865 10.38 ;
    RECT 131.795 12.305 131.865 12.375 ;
    RECT 132.25 5.125 132.46 5.195 ;
    RECT 132.595 5.27 132.805 5.34 ;
    RECT 132.595 13.085 132.805 13.155 ;
    RECT 133.275 3.63 133.345 3.84 ;
    RECT 133.275 5.58 133.345 5.65 ;
    RECT 133.575 1.465 133.785 1.675 ;
    RECT 133.575 3.32 133.785 3.53 ;
    RECT 133.575 6.12 133.785 6.19 ;
    RECT 133.575 7.975 133.785 8.185 ;
    RECT 133.575 11.985 133.785 12.195 ;
    RECT 134.34 1.81 134.55 1.88 ;
    RECT 134.34 6.705 134.55 6.775 ;
    RECT 134.34 10.31 134.55 10.38 ;
    RECT 134.34 12.305 134.55 12.375 ;
    RECT 136.085 2.79 136.295 2.86 ;
    RECT 136.535 1.465 136.745 1.675 ;
    RECT 136.535 3.32 136.745 3.53 ;
    RECT 136.535 5.51 136.745 5.58 ;
    RECT 136.535 6.12 136.745 6.19 ;
    RECT 136.535 7.975 136.745 8.185 ;
    RECT 136.535 11.985 136.745 12.195 ;
    RECT 136.92 1.81 137.13 1.88 ;
    RECT 136.92 6.705 137.13 6.775 ;
    RECT 136.92 12.305 137.13 12.375 ;
    RECT 137.625 1.465 137.695 1.535 ;
    RECT 137.625 1.605 137.695 1.675 ;
    RECT 137.625 3.32 137.695 3.39 ;
    RECT 137.625 3.46 137.695 3.53 ;
    RECT 137.625 5.51 137.695 5.58 ;
    RECT 137.625 5.65 137.695 6.19 ;
    RECT 137.625 7.975 137.695 8.185 ;
    RECT 137.625 11.985 137.695 12.195 ;
    RECT 137.9 1.15 138.11 1.36 ;
    RECT 137.9 2.99 138.11 3.2 ;
    RECT 137.9 4.815 138.11 5.025 ;
    RECT 137.9 6.315 138.11 6.385 ;
    RECT 137.9 8.325 138.11 8.395 ;
    RECT 137.9 10.085 138.11 10.295 ;
    RECT 138.37 4.22 138.44 4.29 ;
    RECT 138.37 7.125 138.44 7.195 ;
    RECT 138.51 7.125 138.58 7.195 ;
    RECT 138.72 1.465 138.93 1.675 ;
    RECT 138.72 3.32 138.93 3.53 ;
    RECT 138.72 5.51 138.93 5.58 ;
    RECT 138.72 6.12 138.93 6.19 ;
    RECT 138.72 7.975 138.93 8.185 ;
    RECT 138.72 11.985 138.93 12.195 ;
    RECT 139.73 1.81 139.94 1.88 ;
    RECT 139.73 6.705 139.94 6.775 ;
    RECT 139.73 12.305 139.94 12.375 ;
    RECT 140.185 2.99 140.685 10.25 ;
    RECT 140.475 1.15 140.685 1.36 ;
    RECT 140.475 6.315 140.685 6.385 ;
    RECT 140.895 7.565 140.965 7.775 ;
    RECT 140.895 14.24 140.965 14.31 ;
    RECT 141.385 12.885 141.65 12.955 ;
    RECT 141.415 1.81 141.625 1.88 ;
    RECT 141.415 6.705 141.625 6.775 ;
    RECT 141.415 12.305 141.625 12.375 ;
    RECT 141.935 1.465 142.145 1.675 ;
    RECT 141.935 3.32 142.145 3.53 ;
    RECT 141.935 5.51 142.145 5.58 ;
    RECT 141.935 6.12 142.145 6.19 ;
    RECT 141.935 7.975 142.145 8.185 ;
    RECT 141.935 11.985 142.145 12.195 ;
    RECT 142.51 12.6 142.72 12.67 ;
    RECT 142.51 13.195 142.72 13.405 ;
    RECT 143.065 1.81 143.135 1.88 ;
    RECT 143.065 6.705 143.135 6.775 ;
    RECT 143.065 12.305 143.135 12.375 ;
    RECT 143.07 12.855 143.14 12.925 ;
    RECT 143.07 12.995 143.14 13.065 ;
    RECT 143.31 1.465 143.52 1.675 ;
    RECT 143.31 3.32 143.52 3.53 ;
    RECT 143.31 5.51 143.52 5.58 ;
    RECT 143.31 6.12 143.52 6.19 ;
    RECT 143.31 7.975 143.52 8.185 ;
    RECT 143.31 11.985 143.52 12.195 ;
    RECT 143.665 12.875 143.925 12.945 ;
    RECT 143.69 1.81 143.9 1.88 ;
    RECT 143.69 6.705 143.9 6.775 ;
    RECT 143.69 12.305 143.9 12.375 ;
    RECT 144.32 12.885 144.39 12.955 ;
    RECT 144.515 12.855 145.135 12.955 ;
    RECT 145.28 2.99 145.695 10.205 ;
    RECT 145.28 9.31 145.35 9.52 ;
    RECT 145.485 1.15 145.695 1.36 ;
    RECT 145.485 6.315 145.695 6.385 ;
    RECT 145.87 1.465 145.94 1.535 ;
    RECT 145.87 1.605 145.94 1.675 ;
    RECT 145.87 3.32 145.94 3.39 ;
    RECT 145.87 3.46 145.94 3.53 ;
    RECT 145.87 5.51 145.94 5.58 ;
    RECT 145.87 5.65 145.94 5.72 ;
    RECT 145.87 5.98 145.94 6.05 ;
    RECT 145.87 6.12 145.94 6.19 ;
    RECT 145.87 7.975 145.94 8.045 ;
    RECT 145.87 8.115 145.94 8.185 ;
    RECT 145.87 11.985 145.94 12.055 ;
    RECT 145.87 12.125 145.94 12.195 ;
    RECT 145.87 13.45 145.94 13.52 ;
    RECT 146.16 1.81 146.37 1.88 ;
    RECT 146.16 6.705 146.37 6.775 ;
    RECT 146.16 12.305 146.37 13.03 ;
    RECT 146.765 1.465 146.975 1.675 ;
    RECT 146.765 3.32 146.975 3.53 ;
    RECT 146.765 6.12 146.975 6.19 ;
    RECT 146.765 7.975 146.975 8.185 ;
    RECT 146.765 11.985 146.975 12.195 ;
    RECT 146.765 13.45 146.975 13.52 ;
    RECT 147.275 4.435 147.345 4.505 ;
    RECT 147.275 9.77 147.345 9.84 ;
    RECT 147.275 13.97 147.345 14.04 ;
    RECT 147.485 2.805 147.555 2.875 ;
    RECT 147.485 7.565 147.555 7.635 ;
    RECT 147.485 14.23 147.555 14.3 ;
    RECT 147.695 4.22 147.765 4.29 ;
    RECT 147.695 7.125 147.765 7.195 ;
    RECT 147.695 13.025 147.765 13.095 ;
    RECT 145.485 1.807 145.695 1.877 ;
    RECT 133.575 7.125 133.785 7.195 ;
    RECT 133.575 4.22 133.785 4.29 ;
    RECT 143.69 9.995 143.9 10.205 ;
    RECT 143.69 8.902 143.9 9.112 ;
    RECT 143.69 8.325 143.9 8.395 ;
    RECT 143.69 6.315 143.9 6.385 ;
    RECT 143.69 4.815 143.9 5.025 ;
    RECT 143.69 2.99 143.9 3.2 ;
    RECT 143.69 1.15 143.9 1.36 ;
    RECT 131.415 7.125 131.625 7.195 ;
    RECT 131.415 4.22 131.625 4.29 ;
    RECT 129.445 7.125 129.655 7.195 ;
    RECT 129.445 4.22 129.655 4.29 ;
    RECT 143.065 9.995 143.135 10.205 ;
    RECT 143.065 8.902 143.135 9.112 ;
    RECT 143.065 8.325 143.135 8.395 ;
    RECT 143.065 6.315 143.135 6.385 ;
    RECT 143.065 4.815 143.135 5.025 ;
    RECT 143.065 2.99 143.135 3.2 ;
    RECT 143.065 1.15 143.135 1.36 ;
    RECT 147.275 12.602 147.345 12.672 ;
    RECT 128.715 7.125 128.925 7.195 ;
    RECT 128.715 4.22 128.925 4.29 ;
    RECT 128.105 11.805 128.175 11.875 ;
    RECT 128.105 7.125 128.175 7.195 ;
    RECT 128.105 4.22 128.175 4.29 ;
    RECT 141.415 9.995 141.625 10.205 ;
    RECT 141.415 8.902 141.625 9.112 ;
    RECT 141.415 8.325 141.625 8.395 ;
    RECT 141.415 6.315 141.625 6.385 ;
    RECT 141.415 4.815 141.625 5.025 ;
    RECT 142.51 4.435 142.72 4.505 ;
    RECT 141.415 2.99 141.625 3.2 ;
    RECT 125.67 5.915 125.88 5.985 ;
    RECT 141.415 1.15 141.625 1.36 ;
    RECT 121.035 12.602 121.105 12.672 ;
    RECT 140.475 12.302 140.685 12.372 ;
    RECT 140.475 6.707 140.685 6.777 ;
    RECT 127.32 11.805 127.53 11.875 ;
    RECT 144.925 13.192 145.135 13.402 ;
    RECT 127.32 7.125 127.53 7.195 ;
    RECT 127.32 4.22 127.53 4.29 ;
    RECT 140.475 1.807 140.685 1.877 ;
    RECT 139.73 10.082 139.94 10.292 ;
    RECT 139.73 8.902 139.94 9.112 ;
    RECT 139.73 8.325 139.94 8.395 ;
    RECT 139.73 6.315 139.94 6.385 ;
    RECT 144.925 12.602 145.135 12.672 ;
    RECT 123.765 12.602 123.975 12.672 ;
    RECT 124.715 11.055 124.925 11.125 ;
    RECT 123.235 12.602 123.445 12.672 ;
    RECT 124.715 7.125 124.925 7.195 ;
    RECT 139.73 4.815 139.94 5.025 ;
    RECT 139.73 2.99 139.94 3.2 ;
    RECT 139.73 1.15 139.94 1.36 ;
    RECT 137.9 12.302 138.11 12.372 ;
    RECT 137.9 6.707 138.11 6.777 ;
    RECT 137.9 1.807 138.11 1.877 ;
    RECT 144.345 13.192 144.555 13.402 ;
    RECT 144.345 12.602 144.555 12.672 ;
    RECT 124.715 4.22 124.925 4.29 ;
    RECT 129.445 8.972 129.655 9.042 ;
    RECT 129.445 3.777 129.655 3.847 ;
    RECT 136.92 10.082 137.13 10.292 ;
    RECT 136.92 8.325 137.13 8.395 ;
    RECT 136.92 6.315 137.13 6.385 ;
    RECT 136.92 4.815 137.13 5.025 ;
    RECT 136.92 2.99 137.13 3.2 ;
    RECT 136.92 1.15 137.13 1.36 ;
    RECT 146.16 14.23 146.37 14.3 ;
    RECT 146.16 7.565 146.37 7.635 ;
    RECT 122.395 7.125 122.465 7.195 ;
    RECT 122.395 4.22 122.465 4.29 ;
    RECT 134.34 8.325 134.55 8.395 ;
    RECT 129.15 11.985 129.22 12.195 ;
    RECT 134.34 6.315 134.55 6.385 ;
    RECT 129.15 10.13 129.22 10.2 ;
    RECT 129.15 7.972 129.22 8.182 ;
    RECT 129.15 6.12 129.22 6.19 ;
    RECT 129.15 3.32 129.22 3.53 ;
    RECT 143.69 14.23 143.9 14.3 ;
    RECT 143.69 7.565 143.9 7.635 ;
    RECT 143.065 14.23 143.135 14.3 ;
    RECT 143.065 7.565 143.135 7.635 ;
    RECT 141.415 14.23 141.625 14.3 ;
    RECT 16.18 0.775 16.39 0.845 ;
    RECT 15.23 1.775 15.44 1.985 ;
    RECT 15.23 1.15 15.44 1.36 ;
    RECT 119.1 0.775 119.31 0.845 ;
    RECT 49.38 0.775 49.59 0.845 ;
    RECT 48.43 1.775 48.64 1.985 ;
    RECT 48.43 1.15 48.64 1.36 ;
    RECT 26.14 0.775 26.35 0.845 ;
    RECT 118.15 1.775 118.36 1.985 ;
    RECT 118.15 1.15 118.36 1.36 ;
    RECT 25.19 1.775 25.4 1.985 ;
    RECT 25.19 1.15 25.4 1.36 ;
    RECT 89.22 0.775 89.43 0.845 ;
    RECT 88.27 1.775 88.48 1.985 ;
    RECT 88.27 1.15 88.48 1.36 ;
    RECT 59.34 0.775 59.55 0.845 ;
    RECT 36.1 0.775 36.31 0.845 ;
    RECT 58.39 1.775 58.6 1.985 ;
    RECT 58.39 1.15 58.6 1.36 ;
    RECT 105.82 0.775 106.03 0.845 ;
    RECT 104.87 1.775 105.08 1.985 ;
    RECT 104.87 1.15 105.08 1.36 ;
    RECT 99.18 0.775 99.39 0.845 ;
    RECT 98.23 1.775 98.44 1.985 ;
    RECT 98.23 1.15 98.44 1.36 ;
    RECT 75.94 0.775 76.15 0.845 ;
    RECT 74.99 1.775 75.2 1.985 ;
    RECT 74.99 1.15 75.2 1.36 ;
    RECT 9.54 0.775 9.75 0.845 ;
    RECT 115.78 0.775 115.99 0.845 ;
    RECT 114.83 1.775 115.04 1.985 ;
    RECT 114.83 1.15 115.04 1.36 ;
    RECT 46.06 0.775 46.27 0.845 ;
    RECT 45.11 1.775 45.32 1.985 ;
    RECT 8.59 1.775 8.8 1.985 ;
    RECT 45.11 1.15 45.32 1.36 ;
    RECT 8.59 1.15 8.8 1.36 ;
    RECT 19.5 0.775 19.71 0.845 ;
    RECT 18.55 1.775 18.76 1.985 ;
    RECT 18.55 1.15 18.76 1.36 ;
    RECT 85.9 0.775 86.11 0.845 ;
    RECT 29.46 0.775 29.67 0.845 ;
    RECT 84.95 1.775 85.16 1.985 ;
    RECT 28.51 1.775 28.72 1.985 ;
    RECT 84.95 1.15 85.16 1.36 ;
    RECT 28.51 1.15 28.72 1.36 ;
    RECT 56.02 0.775 56.23 0.845 ;
    RECT 55.07 1.775 55.28 1.985 ;
    RECT 55.07 1.15 55.28 1.36 ;
    RECT 102.5 0.775 102.71 0.845 ;
    RECT 101.55 1.775 101.76 1.985 ;
    RECT 101.55 1.15 101.76 1.36 ;
    RECT 95.86 0.775 96.07 0.845 ;
    RECT 94.91 1.775 95.12 1.985 ;
    RECT 94.91 1.15 95.12 1.36 ;
    RECT 35.15 1.775 35.36 1.985 ;
    RECT 35.15 1.15 35.36 1.36 ;
    RECT 72.62 0.775 72.83 0.845 ;
    RECT 71.67 1.775 71.88 1.985 ;
    RECT 71.67 1.15 71.88 1.36 ;
    RECT 65.98 0.775 66.19 0.845 ;
    RECT 65.03 1.775 65.24 1.985 ;
    RECT 65.03 1.15 65.24 1.36 ;
    RECT 2.9 0.775 3.11 0.845 ;
    RECT 42.74 0.775 42.95 0.845 ;
    RECT 117.23 1.465 117.44 1.675 ;
    RECT 117.79 0.98 117.86 1.05 ;
    RECT 118.15 0.775 118.36 0.845 ;
    RECT 119.1 1.15 119.31 1.985 ;
    RECT 1.03 1.465 1.24 1.675 ;
    RECT 1.59 0.98 1.66 1.05 ;
    RECT 1.95 0.775 2.16 0.845 ;
    RECT 2.9 1.15 3.11 1.985 ;
    RECT 112.46 0.775 112.67 0.845 ;
    RECT 111.51 1.775 111.72 1.985 ;
    RECT 1.95 1.775 2.16 1.985 ;
    RECT 111.51 1.15 111.72 1.36 ;
    RECT 1.95 1.15 2.16 1.36 ;
    RECT 41.79 1.775 42.0 1.985 ;
    RECT 41.79 1.15 42.0 1.36 ;
    RECT 30.91 1.465 31.12 1.675 ;
    RECT 31.47 0.98 31.54 1.05 ;
    RECT 31.83 0.775 32.04 0.845 ;
    RECT 32.78 1.15 32.99 1.985 ;
    RECT 27.59 1.465 27.8 1.675 ;
    RECT 28.15 0.98 28.22 1.05 ;
    RECT 28.51 0.775 28.72 0.845 ;
    RECT 29.46 1.15 29.67 1.985 ;
    RECT 24.27 1.465 24.48 1.675 ;
    RECT 24.83 0.98 24.9 1.05 ;
    RECT 25.19 0.775 25.4 0.845 ;
    RECT 26.14 1.15 26.35 1.985 ;
    RECT 20.95 1.465 21.16 1.675 ;
    RECT 21.51 0.98 21.58 1.05 ;
    RECT 21.87 0.775 22.08 0.845 ;
    RECT 22.82 1.15 23.03 1.985 ;
    RECT 17.63 1.465 17.84 1.675 ;
    RECT 18.19 0.98 18.26 1.05 ;
    RECT 18.55 0.775 18.76 0.845 ;
    RECT 19.5 1.15 19.71 1.985 ;
    RECT 14.31 1.465 14.52 1.675 ;
    RECT 14.87 0.98 14.94 1.05 ;
    RECT 15.23 0.775 15.44 0.845 ;
    RECT 16.18 1.15 16.39 1.985 ;
    RECT 10.99 1.465 11.2 1.675 ;
    RECT 11.55 0.98 11.62 1.05 ;
    RECT 11.91 0.775 12.12 0.845 ;
    RECT 12.86 1.15 13.07 1.985 ;
    RECT 7.67 1.465 7.88 1.675 ;
    RECT 8.23 0.98 8.3 1.05 ;
    RECT 8.59 0.775 8.8 0.845 ;
    RECT 9.54 1.15 9.75 1.985 ;
    RECT 4.35 1.465 4.56 1.675 ;
    RECT 4.91 0.98 4.98 1.05 ;
    RECT 5.27 0.775 5.48 0.845 ;
    RECT 6.22 1.15 6.43 1.985 ;
    RECT 12.86 0.775 13.07 0.845 ;
    RECT 11.91 1.775 12.12 1.985 ;
    RECT 11.91 1.15 12.12 1.36 ;
    RECT 82.58 0.775 82.79 0.845 ;
    RECT 81.63 1.775 81.84 1.985 ;
    RECT 81.63 1.15 81.84 1.36 ;
    RECT 113.91 1.465 114.12 1.675 ;
    RECT 114.47 0.98 114.54 1.05 ;
    RECT 114.83 0.775 115.04 0.845 ;
    RECT 115.78 1.15 115.99 1.985 ;
    RECT 110.59 1.465 110.8 1.675 ;
    RECT 111.15 0.98 111.22 1.05 ;
    RECT 111.51 0.775 111.72 0.845 ;
    RECT 112.46 1.15 112.67 1.985 ;
    RECT 107.27 1.465 107.48 1.675 ;
    RECT 107.83 0.98 107.9 1.05 ;
    RECT 108.19 0.775 108.4 0.845 ;
    RECT 109.14 1.15 109.35 1.985 ;
    RECT 22.82 0.775 23.03 0.845 ;
    RECT 103.95 1.465 104.16 1.675 ;
    RECT 104.51 0.98 104.58 1.05 ;
    RECT 104.87 0.775 105.08 0.845 ;
    RECT 105.82 1.15 106.03 1.985 ;
    RECT 100.63 1.465 100.84 1.675 ;
    RECT 101.19 0.98 101.26 1.05 ;
    RECT 101.55 0.775 101.76 0.845 ;
    RECT 102.5 1.15 102.71 1.985 ;
    RECT 21.87 1.775 22.08 1.985 ;
    RECT 21.87 1.15 22.08 1.36 ;
    RECT 52.7 0.775 52.91 0.845 ;
    RECT 97.31 1.465 97.52 1.675 ;
    RECT 97.87 0.98 97.94 1.05 ;
    RECT 98.23 0.775 98.44 0.845 ;
    RECT 99.18 1.15 99.39 1.985 ;
    RECT 93.99 1.465 94.2 1.675 ;
    RECT 94.55 0.98 94.62 1.05 ;
    RECT 94.91 0.775 95.12 0.845 ;
    RECT 95.86 1.15 96.07 1.985 ;
    RECT 90.67 1.465 90.88 1.675 ;
    RECT 91.23 0.98 91.3 1.05 ;
    RECT 91.59 0.775 91.8 0.845 ;
    RECT 92.54 1.15 92.75 1.985 ;
    RECT 87.35 1.465 87.56 1.675 ;
    RECT 87.91 0.98 87.98 1.05 ;
    RECT 88.27 0.775 88.48 0.845 ;
    RECT 89.22 1.15 89.43 1.985 ;
    RECT 32.78 0.775 32.99 0.845 ;
    RECT 84.03 1.465 84.24 1.675 ;
    RECT 84.59 0.98 84.66 1.05 ;
    RECT 84.95 0.775 85.16 0.845 ;
    RECT 85.9 1.15 86.11 1.985 ;
    RECT 80.71 1.465 80.92 1.675 ;
    RECT 81.27 0.98 81.34 1.05 ;
    RECT 81.63 0.775 81.84 0.845 ;
    RECT 82.58 1.15 82.79 1.985 ;
    RECT 77.39 1.465 77.6 1.675 ;
    RECT 77.95 0.98 78.02 1.05 ;
    RECT 78.31 0.775 78.52 0.845 ;
    RECT 79.26 1.15 79.47 1.985 ;
    RECT 31.83 1.775 32.04 1.985 ;
    RECT 74.07 1.465 74.28 1.675 ;
    RECT 74.63 0.98 74.7 1.05 ;
    RECT 74.99 0.775 75.2 0.845 ;
    RECT 75.94 1.15 76.15 1.985 ;
    RECT 31.83 1.15 32.04 1.36 ;
    RECT 70.75 1.465 70.96 1.675 ;
    RECT 71.31 0.98 71.38 1.05 ;
    RECT 71.67 0.775 71.88 0.845 ;
    RECT 72.62 1.15 72.83 1.985 ;
    RECT 67.43 1.465 67.64 1.675 ;
    RECT 67.99 0.98 68.06 1.05 ;
    RECT 68.35 0.775 68.56 0.845 ;
    RECT 69.3 1.15 69.51 1.985 ;
    RECT 51.75 1.775 51.96 1.985 ;
    RECT 51.75 1.15 51.96 1.36 ;
    RECT 92.54 0.775 92.75 0.845 ;
    RECT 64.11 1.465 64.32 1.675 ;
    RECT 64.67 0.98 64.74 1.05 ;
    RECT 65.03 0.775 65.24 0.845 ;
    RECT 65.98 1.15 66.19 1.985 ;
    RECT 60.79 1.465 61.0 1.675 ;
    RECT 61.35 0.98 61.42 1.05 ;
    RECT 61.71 0.775 61.92 0.845 ;
    RECT 62.66 1.15 62.87 1.985 ;
    RECT 57.47 1.465 57.68 1.675 ;
    RECT 58.03 0.98 58.1 1.05 ;
    RECT 58.39 0.775 58.6 0.845 ;
    RECT 59.34 1.15 59.55 1.985 ;
    RECT 54.15 1.465 54.36 1.675 ;
    RECT 54.71 0.98 54.78 1.05 ;
    RECT 55.07 0.775 55.28 0.845 ;
    RECT 56.02 1.15 56.23 1.985 ;
    RECT 50.83 1.465 51.04 1.675 ;
    RECT 51.39 0.98 51.46 1.05 ;
    RECT 51.75 0.775 51.96 0.845 ;
    RECT 52.7 1.15 52.91 1.985 ;
    RECT 47.51 1.465 47.72 1.675 ;
    RECT 48.07 0.98 48.14 1.05 ;
    RECT 48.43 0.775 48.64 0.845 ;
    RECT 49.38 1.15 49.59 1.985 ;
    RECT 44.19 1.465 44.4 1.675 ;
    RECT 44.75 0.98 44.82 1.05 ;
    RECT 45.11 0.775 45.32 0.845 ;
    RECT 46.06 1.15 46.27 1.985 ;
    RECT 40.87 1.465 41.08 1.675 ;
    RECT 41.43 0.98 41.5 1.05 ;
    RECT 41.79 0.775 42.0 0.845 ;
    RECT 42.74 1.15 42.95 1.985 ;
    RECT 37.55 1.465 37.76 1.675 ;
    RECT 38.11 0.98 38.18 1.05 ;
    RECT 38.47 0.775 38.68 0.845 ;
    RECT 39.42 1.15 39.63 1.985 ;
    RECT 34.23 1.465 34.44 1.675 ;
    RECT 34.79 0.98 34.86 1.05 ;
    RECT 35.15 0.775 35.36 0.845 ;
    RECT 36.1 1.15 36.31 1.985 ;
    RECT 69.3 0.775 69.51 0.845 ;
    RECT 91.59 1.775 91.8 1.985 ;
    RECT 91.59 1.15 91.8 1.36 ;
    RECT 68.35 1.775 68.56 1.985 ;
    RECT 68.35 1.15 68.56 1.36 ;
    RECT 62.66 0.775 62.87 0.845 ;
    RECT 61.71 1.775 61.92 1.985 ;
    RECT 109.14 0.775 109.35 0.845 ;
    RECT 61.71 1.15 61.92 1.36 ;
    RECT 39.42 0.775 39.63 0.845 ;
    RECT 38.47 1.775 38.68 1.985 ;
    RECT 38.47 1.15 38.68 1.36 ;
    RECT 108.19 1.775 108.4 1.985 ;
    RECT 108.19 1.15 108.4 1.36 ;
    RECT 6.22 0.775 6.43 0.845 ;
    RECT 5.27 1.775 5.48 1.985 ;
    RECT 5.27 1.15 5.48 1.36 ;
    RECT 79.26 0.775 79.47 0.845 ;
    RECT 78.31 1.775 78.52 1.985 ;
    RECT 78.31 1.15 78.52 1.36 ;
    RECT 81.63 14.23 81.84 14.3 ;
    RECT 81.17 14.23 81.38 14.3 ;
    RECT 75.48 13.71 75.69 13.78 ;
    RECT 115.32 13.97 115.53 14.04 ;
    RECT 35.15 14.23 35.36 14.3 ;
    RECT 34.69 14.23 34.9 14.3 ;
    RECT 42.28 13.97 42.49 14.04 ;
    RECT 78.31 14.23 78.52 14.3 ;
    RECT 72.16 13.71 72.37 13.78 ;
    RECT 12.4 13.97 12.61 14.04 ;
    RECT 64.105 13.45 64.325 13.52 ;
    RECT 77.85 14.23 78.06 14.3 ;
    RECT 60.785 13.45 61.005 13.52 ;
    RECT 57.465 13.45 57.685 13.52 ;
    RECT 54.145 13.45 54.365 13.52 ;
    RECT 95.4 13.97 95.61 14.04 ;
    RECT 50.825 13.45 51.045 13.52 ;
    RECT 47.505 13.45 47.725 13.52 ;
    RECT 44.185 13.45 44.405 13.52 ;
    RECT 40.865 13.45 41.085 13.52 ;
    RECT 37.545 13.45 37.765 13.52 ;
    RECT 34.225 13.45 34.445 13.52 ;
    RECT 68.84 13.71 69.05 13.78 ;
    RECT 111.51 14.23 111.72 14.3 ;
    RECT 74.99 14.23 75.2 14.3 ;
    RECT 111.05 14.23 111.26 14.3 ;
    RECT 74.53 14.23 74.74 14.3 ;
    RECT 108.68 13.97 108.89 14.04 ;
    RECT 31.83 14.23 32.04 14.3 ;
    RECT 31.37 14.23 31.58 14.3 ;
    RECT 32.32 13.71 32.53 13.78 ;
    RECT 65.52 13.97 65.73 14.04 ;
    RECT 88.76 13.97 88.97 14.04 ;
    RECT 28.51 14.23 28.72 14.3 ;
    RECT 118.64 13.71 118.85 13.78 ;
    RECT 28.05 14.23 28.26 14.3 ;
    RECT 29.0 13.71 29.21 13.78 ;
    RECT 71.67 14.23 71.88 14.3 ;
    RECT 35.64 13.97 35.85 14.04 ;
    RECT 71.21 14.23 71.42 14.3 ;
    RECT 5.76 13.97 5.97 14.04 ;
    RECT 115.32 13.71 115.53 13.78 ;
    RECT 25.19 14.23 25.4 14.3 ;
    RECT 24.73 14.23 24.94 14.3 ;
    RECT 25.68 13.71 25.89 13.78 ;
    RECT 58.88 13.97 59.09 14.04 ;
    RECT 29.0 13.97 29.21 14.04 ;
    RECT 65.52 13.71 65.73 13.78 ;
    RECT 68.35 14.23 68.56 14.3 ;
    RECT 67.89 14.23 68.1 14.3 ;
    RECT 112.0 13.71 112.21 13.78 ;
    RECT 82.12 13.97 82.33 14.04 ;
    RECT 102.04 13.97 102.25 14.04 ;
    RECT 22.36 13.71 22.57 13.78 ;
    RECT 62.2 13.71 62.41 13.78 ;
    RECT 108.68 13.71 108.89 13.78 ;
    RECT 19.04 13.71 19.25 13.78 ;
    RECT 21.87 14.23 22.08 14.3 ;
    RECT 21.41 14.23 21.62 14.3 ;
    RECT 52.24 13.97 52.45 14.04 ;
    RECT 72.16 13.97 72.37 14.04 ;
    RECT 22.36 13.97 22.57 14.04 ;
    RECT 30.905 13.45 31.125 13.52 ;
    RECT 27.585 13.45 27.805 13.52 ;
    RECT 58.88 13.71 59.09 13.78 ;
    RECT 24.265 13.45 24.485 13.52 ;
    RECT 20.945 13.45 21.165 13.52 ;
    RECT 17.625 13.45 17.845 13.52 ;
    RECT 14.305 13.45 14.525 13.52 ;
    RECT 65.03 14.23 65.24 14.3 ;
    RECT 10.985 13.45 11.205 13.52 ;
    RECT 64.57 14.23 64.78 14.3 ;
    RECT 105.36 13.71 105.57 13.78 ;
    RECT 7.665 13.45 7.885 13.52 ;
    RECT 15.72 13.71 15.93 13.78 ;
    RECT 4.345 13.45 4.565 13.52 ;
    RECT 1.025 13.45 1.245 13.52 ;
    RECT 18.55 14.23 18.76 14.3 ;
    RECT 18.09 14.23 18.3 14.3 ;
    RECT 55.56 13.71 55.77 13.78 ;
    RECT 118.64 13.97 118.85 14.04 ;
    RECT 61.71 14.23 61.92 14.3 ;
    RECT 102.04 13.71 102.25 13.78 ;
    RECT 61.25 14.23 61.46 14.3 ;
    RECT 12.4 13.71 12.61 13.78 ;
    RECT 15.23 14.23 15.44 14.3 ;
    RECT 14.77 14.23 14.98 14.3 ;
    RECT 104.87 14.23 105.08 14.3 ;
    RECT 104.41 14.23 104.62 14.3 ;
    RECT 52.24 13.71 52.45 13.78 ;
    RECT 45.6 13.97 45.81 14.04 ;
    RECT 15.72 13.97 15.93 14.04 ;
    RECT 98.72 13.97 98.93 14.04 ;
    RECT 9.08 13.71 9.29 13.78 ;
    RECT 58.39 14.23 58.6 14.3 ;
    RECT 57.93 14.23 58.14 14.3 ;
    RECT 11.91 14.23 12.12 14.3 ;
    RECT 11.45 14.23 11.66 14.3 ;
    RECT 101.55 14.23 101.76 14.3 ;
    RECT 101.09 14.23 101.3 14.3 ;
    RECT 48.92 13.71 49.13 13.78 ;
    RECT 114.83 14.23 115.04 14.3 ;
    RECT 114.37 14.23 114.58 14.3 ;
    RECT 112.0 13.97 112.21 14.04 ;
    RECT 5.76 13.71 5.97 13.78 ;
    RECT 8.59 14.23 8.8 14.3 ;
    RECT 8.13 14.23 8.34 14.3 ;
    RECT 45.6 13.71 45.81 13.78 ;
    RECT 9.08 13.97 9.29 14.04 ;
    RECT 2.44 13.71 2.65 13.78 ;
    RECT 92.08 13.97 92.29 14.04 ;
    RECT 98.72 13.71 98.93 13.78 ;
    RECT 55.07 14.23 55.28 14.3 ;
    RECT 54.61 14.23 54.82 14.3 ;
    RECT 98.23 14.23 98.44 14.3 ;
    RECT 97.77 14.23 97.98 14.3 ;
    RECT 42.28 13.71 42.49 13.78 ;
    RECT 108.19 14.23 108.4 14.3 ;
    RECT 107.73 14.23 107.94 14.3 ;
    RECT 38.96 13.97 39.17 14.04 ;
    RECT 95.4 13.71 95.61 13.78 ;
    RECT 51.75 14.23 51.96 14.3 ;
    RECT 51.29 14.23 51.5 14.3 ;
    RECT 62.2 13.97 62.41 14.04 ;
    RECT 32.32 13.97 32.53 14.04 ;
    RECT 94.91 14.23 95.12 14.3 ;
    RECT 38.96 13.71 39.17 13.78 ;
    RECT 94.45 14.23 94.66 14.3 ;
    RECT 5.27 14.23 5.48 14.3 ;
    RECT 4.81 14.23 5.02 14.3 ;
    RECT 92.08 13.71 92.29 13.78 ;
    RECT 85.44 13.97 85.65 14.04 ;
    RECT 105.36 13.97 105.57 14.04 ;
    RECT 48.43 14.23 48.64 14.3 ;
    RECT 47.97 14.23 48.18 14.3 ;
    RECT 75.48 13.97 75.69 14.04 ;
    RECT 35.64 13.71 35.85 13.78 ;
    RECT 91.59 14.23 91.8 14.3 ;
    RECT 91.13 14.23 91.34 14.3 ;
    RECT 1.95 14.23 2.16 14.3 ;
    RECT 1.49 14.23 1.7 14.3 ;
    RECT 88.76 13.71 88.97 13.78 ;
    RECT 2.44 13.97 2.65 14.04 ;
    RECT 45.11 14.23 45.32 14.3 ;
    RECT 44.65 14.23 44.86 14.3 ;
    RECT 55.56 13.97 55.77 14.04 ;
    RECT 25.68 13.97 25.89 14.04 ;
    RECT 85.44 13.71 85.65 13.78 ;
    RECT 78.8 13.97 79.01 14.04 ;
    RECT 41.79 14.23 42.0 14.3 ;
    RECT 41.33 14.23 41.54 14.3 ;
    RECT 117.225 13.45 117.445 13.52 ;
    RECT 113.905 13.45 114.125 13.52 ;
    RECT 110.585 13.45 110.805 13.52 ;
    RECT 107.265 13.45 107.485 13.52 ;
    RECT 88.27 14.23 88.48 14.3 ;
    RECT 103.945 13.45 104.165 13.52 ;
    RECT 87.81 14.23 88.02 14.3 ;
    RECT 100.625 13.45 100.845 13.52 ;
    RECT 82.12 13.71 82.33 13.78 ;
    RECT 48.92 13.97 49.13 14.04 ;
    RECT 68.84 13.97 69.05 14.04 ;
    RECT 19.04 13.97 19.25 14.04 ;
    RECT 84.95 14.23 85.16 14.3 ;
    RECT 84.49 14.23 84.7 14.3 ;
    RECT 78.8 13.71 79.01 13.78 ;
    RECT 97.305 13.45 97.525 13.52 ;
    RECT 93.985 13.45 94.205 13.52 ;
    RECT 90.665 13.45 90.885 13.52 ;
    RECT 87.345 13.45 87.565 13.52 ;
    RECT 84.025 13.45 84.245 13.52 ;
    RECT 80.705 13.45 80.925 13.52 ;
    RECT 77.385 13.45 77.605 13.52 ;
    RECT 74.065 13.45 74.285 13.52 ;
    RECT 38.47 14.23 38.68 14.3 ;
    RECT 118.15 14.23 118.36 14.3 ;
    RECT 70.745 13.45 70.965 13.52 ;
    RECT 38.01 14.23 38.22 14.3 ;
    RECT 117.69 14.23 117.9 14.3 ;
    RECT 67.425 13.45 67.645 13.52 ;
    RECT 0.61 11.985 0.68 12.195 ;
    RECT 0.61 7.972 0.68 8.182 ;
    RECT 0.19 13.97 0.26 14.04 ;
    RECT 0.4 14.23 0.47 14.3 ;
    RECT 0.61 6.12 0.68 6.19 ;
    RECT 0.61 4.445 0.68 4.655 ;
    RECT 0.61 3.32 0.68 3.53 ;
    RECT 0.4 7.58 0.47 7.65 ;
    RECT 0.615 4.22 0.685 4.29 ;
    RECT 0.615 7.125 0.685 7.195 ;
    RECT 25.19 6.315 25.4 6.385 ;
    RECT 25.19 4.815 25.4 5.025 ;
    RECT 50.83 7.125 51.04 7.195 ;
    RECT 50.83 4.22 51.04 4.29 ;
    RECT 25.19 7.565 25.4 7.635 ;
    RECT 41.79 3.742 42.0 3.952 ;
    RECT 41.79 2.99 42.0 3.2 ;
    RECT 93.99 7.125 94.2 7.195 ;
    RECT 93.99 4.22 94.2 4.29 ;
    RECT 5.27 9.995 5.48 10.205 ;
    RECT 5.27 8.902 5.48 9.112 ;
    RECT 74.64 6.12 74.71 6.19 ;
    RECT 5.27 8.705 5.48 8.775 ;
    RECT 5.27 8.325 5.48 8.395 ;
    RECT 5.27 6.315 5.48 6.385 ;
    RECT 25.19 3.742 25.4 3.952 ;
    RECT 5.27 4.815 5.48 5.025 ;
    RECT 25.19 2.99 25.4 3.2 ;
    RECT 5.27 3.742 5.48 3.952 ;
    RECT 5.27 2.99 5.48 3.2 ;
    RECT 117.8 6.12 117.87 6.19 ;
    RECT 84.95 9.995 85.16 10.205 ;
    RECT 117.8 5.182 117.87 5.392 ;
    RECT 84.95 8.902 85.16 9.112 ;
    RECT 117.8 4.445 117.87 4.655 ;
    RECT 84.95 8.705 85.16 8.775 ;
    RECT 84.95 8.325 85.16 8.395 ;
    RECT 84.95 6.315 85.16 6.385 ;
    RECT 117.23 7.125 117.44 7.195 ;
    RECT 84.95 4.815 85.16 5.025 ;
    RECT 74.64 5.182 74.71 5.392 ;
    RECT 117.23 4.22 117.44 4.29 ;
    RECT 84.95 3.742 85.16 3.952 ;
    RECT 74.64 4.445 74.71 4.655 ;
    RECT 84.95 2.99 85.16 3.2 ;
    RECT 58.39 7.565 58.6 7.635 ;
    RECT 14.88 6.12 14.95 6.19 ;
    RECT 14.88 5.182 14.95 5.392 ;
    RECT 74.07 7.125 74.28 7.195 ;
    RECT 14.88 4.445 14.95 4.655 ;
    RECT 74.07 4.22 74.28 4.29 ;
    RECT 14.31 7.125 14.52 7.195 ;
    RECT 14.31 4.22 14.52 4.29 ;
    RECT 88.27 7.565 88.48 7.635 ;
    RECT 21.87 7.565 22.08 7.635 ;
    RECT 38.47 9.995 38.68 10.205 ;
    RECT 38.47 8.902 38.68 9.112 ;
    RECT 38.47 8.705 38.68 8.775 ;
    RECT 38.47 8.325 38.68 8.395 ;
    RECT 38.47 6.315 38.68 6.385 ;
    RECT 38.47 4.815 38.68 5.025 ;
    RECT 91.24 6.12 91.31 6.19 ;
    RECT 38.47 3.742 38.68 3.952 ;
    RECT 91.24 5.182 91.31 5.392 ;
    RECT 38.47 2.99 38.68 3.2 ;
    RECT 91.24 4.445 91.31 4.655 ;
    RECT 21.87 9.995 22.08 10.205 ;
    RECT 21.87 8.902 22.08 9.112 ;
    RECT 48.08 6.12 48.15 6.19 ;
    RECT 90.67 7.125 90.88 7.195 ;
    RECT 21.87 8.705 22.08 8.775 ;
    RECT 48.08 5.182 48.15 5.392 ;
    RECT 21.87 8.325 22.08 8.395 ;
    RECT 48.08 4.445 48.15 4.655 ;
    RECT 21.87 6.315 22.08 6.385 ;
    RECT 21.87 4.815 22.08 5.025 ;
    RECT 21.87 3.742 22.08 3.952 ;
    RECT 47.51 7.125 47.72 7.195 ;
    RECT 21.87 2.99 22.08 3.2 ;
    RECT 47.51 4.22 47.72 4.29 ;
    RECT 118.15 7.565 118.36 7.635 ;
    RECT 81.63 9.995 81.84 10.205 ;
    RECT 81.63 8.902 81.84 9.112 ;
    RECT 55.07 7.565 55.28 7.635 ;
    RECT 1.95 9.995 2.16 10.205 ;
    RECT 90.67 4.22 90.88 4.29 ;
    RECT 1.95 8.902 2.16 9.112 ;
    RECT 1.95 8.705 2.16 8.775 ;
    RECT 71.32 6.12 71.39 6.19 ;
    RECT 1.95 8.325 2.16 8.395 ;
    RECT 71.32 5.182 71.39 5.392 ;
    RECT 1.95 6.315 2.16 6.385 ;
    RECT 1.95 4.815 2.16 5.025 ;
    RECT 1.95 3.742 2.16 3.952 ;
    RECT 1.95 2.99 2.16 3.2 ;
    RECT 114.48 6.12 114.55 6.19 ;
    RECT 114.48 5.182 114.55 5.392 ;
    RECT 81.63 8.705 81.84 8.775 ;
    RECT 114.48 4.445 114.55 4.655 ;
    RECT 81.63 8.325 81.84 8.395 ;
    RECT 81.63 6.315 81.84 6.385 ;
    RECT 81.63 4.815 81.84 5.025 ;
    RECT 113.91 7.125 114.12 7.195 ;
    RECT 81.63 3.742 81.84 3.952 ;
    RECT 113.91 4.22 114.12 4.29 ;
    RECT 81.63 2.99 81.84 3.2 ;
    RECT 71.32 4.445 71.39 4.655 ;
    RECT 11.56 6.12 11.63 6.19 ;
    RECT 11.56 5.182 11.63 5.392 ;
    RECT 70.75 7.125 70.96 7.195 ;
    RECT 11.56 4.445 11.63 4.655 ;
    RECT 70.75 4.22 70.96 4.29 ;
    RECT 10.99 7.125 11.2 7.195 ;
    RECT 10.99 4.22 11.2 4.29 ;
    RECT 84.95 7.565 85.16 7.635 ;
    RECT 18.55 7.565 18.76 7.635 ;
    RECT 114.83 7.565 115.04 7.635 ;
    RECT 35.15 9.995 35.36 10.205 ;
    RECT 35.15 8.902 35.36 9.112 ;
    RECT 35.15 8.705 35.36 8.775 ;
    RECT 51.75 7.565 51.96 7.635 ;
    RECT 35.15 8.325 35.36 8.395 ;
    RECT 35.15 6.315 35.36 6.385 ;
    RECT 35.15 4.815 35.36 5.025 ;
    RECT 35.15 3.742 35.36 3.952 ;
    RECT 87.92 6.12 87.99 6.19 ;
    RECT 35.15 2.99 35.36 3.2 ;
    RECT 87.92 5.182 87.99 5.392 ;
    RECT 87.92 4.445 87.99 4.655 ;
    RECT 87.35 7.125 87.56 7.195 ;
    RECT 87.35 4.22 87.56 4.29 ;
    RECT 78.31 9.995 78.52 10.205 ;
    RECT 78.31 8.902 78.52 9.112 ;
    RECT 78.31 8.705 78.52 8.775 ;
    RECT 78.31 8.325 78.52 8.395 ;
    RECT 68.0 6.12 68.07 6.19 ;
    RECT 68.0 5.182 68.07 5.392 ;
    RECT 68.0 4.445 68.07 4.655 ;
    RECT 8.24 6.12 8.31 6.19 ;
    RECT 81.63 7.565 81.84 7.635 ;
    RECT 15.23 7.565 15.44 7.635 ;
    RECT 111.16 6.12 111.23 6.19 ;
    RECT 111.16 5.182 111.23 5.392 ;
    RECT 111.16 4.445 111.23 4.655 ;
    RECT 78.31 6.315 78.52 6.385 ;
    RECT 78.31 4.815 78.52 5.025 ;
    RECT 78.31 3.742 78.52 3.952 ;
    RECT 110.59 7.125 110.8 7.195 ;
    RECT 78.31 2.99 78.52 3.2 ;
    RECT 110.59 4.22 110.8 4.29 ;
    RECT 67.43 7.125 67.64 7.195 ;
    RECT 67.43 4.22 67.64 4.29 ;
    RECT 117.195 5.255 117.475 5.325 ;
    RECT 117.195 8.065 117.475 8.135 ;
    RECT 117.195 11.985 117.475 12.195 ;
    RECT 117.23 3.32 117.44 3.53 ;
    RECT 117.23 4.445 117.44 4.655 ;
    RECT 117.23 6.12 117.44 6.19 ;
    RECT 117.6 3.035 117.67 3.105 ;
    RECT 117.6 3.78 117.67 3.85 ;
    RECT 117.6 4.86 117.67 4.93 ;
    RECT 117.6 6.315 117.67 6.385 ;
    RECT 117.6 6.745 117.67 6.815 ;
    RECT 117.6 12.31 117.67 12.38 ;
    RECT 117.8 4.23 117.87 4.3 ;
    RECT 117.8 7.135 117.87 7.205 ;
    RECT 117.8 8.325 117.87 8.395 ;
    RECT 117.8 8.71 117.87 9.115 ;
    RECT 117.8 9.995 117.87 10.205 ;
    RECT 118.61 12.605 118.875 12.675 ;
    RECT 119.07 8.325 119.14 8.395 ;
    RECT 119.07 8.325 119.34 9.115 ;
    RECT 119.07 8.71 119.14 8.97 ;
    RECT 119.07 9.995 119.34 10.205 ;
    RECT 119.1 2.99 119.31 3.955 ;
    RECT 119.1 4.815 119.31 5.025 ;
    RECT 119.1 6.315 119.31 6.385 ;
    RECT 0.995 5.255 1.275 5.325 ;
    RECT 0.995 8.065 1.275 8.135 ;
    RECT 0.995 11.985 1.275 12.195 ;
    RECT 1.03 3.32 1.24 3.53 ;
    RECT 1.03 4.445 1.24 4.655 ;
    RECT 1.03 6.12 1.24 6.19 ;
    RECT 1.4 3.035 1.47 3.105 ;
    RECT 1.4 3.78 1.47 3.85 ;
    RECT 1.4 4.86 1.47 4.93 ;
    RECT 1.4 6.315 1.47 6.385 ;
    RECT 1.4 6.745 1.47 6.815 ;
    RECT 1.4 12.31 1.47 12.38 ;
    RECT 1.6 4.23 1.67 4.3 ;
    RECT 1.6 7.135 1.67 7.205 ;
    RECT 1.6 8.325 1.67 8.395 ;
    RECT 1.6 8.71 1.67 9.115 ;
    RECT 1.6 9.995 1.67 10.205 ;
    RECT 2.41 12.605 2.675 12.675 ;
    RECT 2.87 8.325 2.94 8.395 ;
    RECT 2.87 8.325 3.14 9.115 ;
    RECT 2.87 8.71 2.94 8.97 ;
    RECT 2.87 9.995 3.14 10.205 ;
    RECT 2.9 2.99 3.11 3.955 ;
    RECT 2.9 4.815 3.11 5.025 ;
    RECT 2.9 6.315 3.11 6.385 ;
    RECT 111.51 7.565 111.72 7.635 ;
    RECT 48.43 7.565 48.64 7.635 ;
    RECT 101.55 9.995 101.76 10.205 ;
    RECT 101.55 8.902 101.76 9.112 ;
    RECT 101.55 8.705 101.76 8.775 ;
    RECT 101.55 8.325 101.76 8.395 ;
    RECT 101.55 6.315 101.76 6.385 ;
    RECT 101.55 4.815 101.76 5.025 ;
    RECT 101.55 3.742 101.76 3.952 ;
    RECT 101.55 2.99 101.76 3.2 ;
    RECT 30.875 5.255 31.155 5.325 ;
    RECT 30.875 8.065 31.155 8.135 ;
    RECT 30.875 11.985 31.155 12.195 ;
    RECT 30.91 3.32 31.12 3.53 ;
    RECT 30.91 4.445 31.12 4.655 ;
    RECT 30.91 6.12 31.12 6.19 ;
    RECT 31.28 3.035 31.35 3.105 ;
    RECT 31.28 3.78 31.35 3.85 ;
    RECT 31.28 4.86 31.35 4.93 ;
    RECT 31.28 6.315 31.35 6.385 ;
    RECT 31.28 6.745 31.35 6.815 ;
    RECT 31.28 12.31 31.35 12.38 ;
    RECT 31.48 4.23 31.55 4.3 ;
    RECT 31.48 7.135 31.55 7.205 ;
    RECT 31.48 8.325 31.55 8.395 ;
    RECT 31.48 8.71 31.55 9.115 ;
    RECT 31.48 9.995 31.55 10.205 ;
    RECT 32.29 12.605 32.555 12.675 ;
    RECT 32.75 8.325 32.82 8.395 ;
    RECT 32.75 8.325 33.02 9.115 ;
    RECT 32.75 8.71 32.82 8.97 ;
    RECT 32.75 9.995 33.02 10.205 ;
    RECT 32.78 2.99 32.99 3.955 ;
    RECT 32.78 4.815 32.99 5.025 ;
    RECT 32.78 6.315 32.99 6.385 ;
    RECT 27.555 5.255 27.835 5.325 ;
    RECT 27.555 8.065 27.835 8.135 ;
    RECT 27.555 11.985 27.835 12.195 ;
    RECT 27.59 3.32 27.8 3.53 ;
    RECT 27.59 4.445 27.8 4.655 ;
    RECT 27.59 6.12 27.8 6.19 ;
    RECT 27.96 3.035 28.03 3.105 ;
    RECT 27.96 3.78 28.03 3.85 ;
    RECT 27.96 4.86 28.03 4.93 ;
    RECT 27.96 6.315 28.03 6.385 ;
    RECT 27.96 6.745 28.03 6.815 ;
    RECT 27.96 12.31 28.03 12.38 ;
    RECT 28.16 4.23 28.23 4.3 ;
    RECT 28.16 7.135 28.23 7.205 ;
    RECT 28.16 8.325 28.23 8.395 ;
    RECT 28.16 8.71 28.23 9.115 ;
    RECT 28.16 9.995 28.23 10.205 ;
    RECT 28.97 12.605 29.235 12.675 ;
    RECT 29.43 8.325 29.5 8.395 ;
    RECT 29.43 8.325 29.7 9.115 ;
    RECT 29.43 8.71 29.5 8.97 ;
    RECT 29.43 9.995 29.7 10.205 ;
    RECT 29.46 2.99 29.67 3.955 ;
    RECT 29.46 4.815 29.67 5.025 ;
    RECT 29.46 6.315 29.67 6.385 ;
    RECT 24.235 5.255 24.515 5.325 ;
    RECT 24.235 8.065 24.515 8.135 ;
    RECT 24.235 11.985 24.515 12.195 ;
    RECT 24.27 3.32 24.48 3.53 ;
    RECT 24.27 4.445 24.48 4.655 ;
    RECT 24.27 6.12 24.48 6.19 ;
    RECT 24.64 3.035 24.71 3.105 ;
    RECT 24.64 3.78 24.71 3.85 ;
    RECT 24.64 4.86 24.71 4.93 ;
    RECT 24.64 6.315 24.71 6.385 ;
    RECT 24.64 6.745 24.71 6.815 ;
    RECT 24.64 12.31 24.71 12.38 ;
    RECT 24.84 4.23 24.91 4.3 ;
    RECT 24.84 7.135 24.91 7.205 ;
    RECT 24.84 8.325 24.91 8.395 ;
    RECT 24.84 8.71 24.91 9.115 ;
    RECT 24.84 9.995 24.91 10.205 ;
    RECT 25.65 12.605 25.915 12.675 ;
    RECT 26.11 8.325 26.18 8.395 ;
    RECT 26.11 8.325 26.38 9.115 ;
    RECT 26.11 8.71 26.18 8.97 ;
    RECT 26.11 9.995 26.38 10.205 ;
    RECT 26.14 2.99 26.35 3.955 ;
    RECT 26.14 4.815 26.35 5.025 ;
    RECT 26.14 6.315 26.35 6.385 ;
    RECT 20.915 5.255 21.195 5.325 ;
    RECT 20.915 8.065 21.195 8.135 ;
    RECT 20.915 11.985 21.195 12.195 ;
    RECT 20.95 3.32 21.16 3.53 ;
    RECT 20.95 4.445 21.16 4.655 ;
    RECT 20.95 6.12 21.16 6.19 ;
    RECT 21.32 3.035 21.39 3.105 ;
    RECT 21.32 3.78 21.39 3.85 ;
    RECT 21.32 4.86 21.39 4.93 ;
    RECT 21.32 6.315 21.39 6.385 ;
    RECT 21.32 6.745 21.39 6.815 ;
    RECT 21.32 12.31 21.39 12.38 ;
    RECT 21.52 4.23 21.59 4.3 ;
    RECT 21.52 7.135 21.59 7.205 ;
    RECT 21.52 8.325 21.59 8.395 ;
    RECT 21.52 8.71 21.59 9.115 ;
    RECT 21.52 9.995 21.59 10.205 ;
    RECT 22.33 12.605 22.595 12.675 ;
    RECT 22.79 8.325 22.86 8.395 ;
    RECT 22.79 8.325 23.06 9.115 ;
    RECT 22.79 8.71 22.86 8.97 ;
    RECT 22.79 9.995 23.06 10.205 ;
    RECT 22.82 2.99 23.03 3.955 ;
    RECT 22.82 4.815 23.03 5.025 ;
    RECT 22.82 6.315 23.03 6.385 ;
    RECT 84.6 6.12 84.67 6.19 ;
    RECT 17.595 5.255 17.875 5.325 ;
    RECT 17.595 8.065 17.875 8.135 ;
    RECT 17.595 11.985 17.875 12.195 ;
    RECT 17.63 3.32 17.84 3.53 ;
    RECT 17.63 4.445 17.84 4.655 ;
    RECT 17.63 6.12 17.84 6.19 ;
    RECT 18.0 3.035 18.07 3.105 ;
    RECT 18.0 3.78 18.07 3.85 ;
    RECT 18.0 4.86 18.07 4.93 ;
    RECT 18.0 6.315 18.07 6.385 ;
    RECT 18.0 6.745 18.07 6.815 ;
    RECT 18.0 12.31 18.07 12.38 ;
    RECT 18.2 4.23 18.27 4.3 ;
    RECT 18.2 7.135 18.27 7.205 ;
    RECT 18.2 8.325 18.27 8.395 ;
    RECT 18.2 8.71 18.27 9.115 ;
    RECT 18.2 9.995 18.27 10.205 ;
    RECT 19.01 12.605 19.275 12.675 ;
    RECT 19.47 8.325 19.54 8.395 ;
    RECT 19.47 8.325 19.74 9.115 ;
    RECT 19.47 8.71 19.54 8.97 ;
    RECT 19.47 9.995 19.74 10.205 ;
    RECT 19.5 2.99 19.71 3.955 ;
    RECT 19.5 4.815 19.71 5.025 ;
    RECT 19.5 6.315 19.71 6.385 ;
    RECT 84.6 5.182 84.67 5.392 ;
    RECT 14.275 5.255 14.555 5.325 ;
    RECT 14.275 8.065 14.555 8.135 ;
    RECT 14.275 11.985 14.555 12.195 ;
    RECT 14.31 3.32 14.52 3.53 ;
    RECT 14.31 4.445 14.52 4.655 ;
    RECT 14.31 6.12 14.52 6.19 ;
    RECT 14.68 3.035 14.75 3.105 ;
    RECT 14.68 3.78 14.75 3.85 ;
    RECT 14.68 4.86 14.75 4.93 ;
    RECT 14.68 6.315 14.75 6.385 ;
    RECT 14.68 6.745 14.75 6.815 ;
    RECT 14.68 12.31 14.75 12.38 ;
    RECT 14.88 4.23 14.95 4.3 ;
    RECT 14.88 7.135 14.95 7.205 ;
    RECT 14.88 8.325 14.95 8.395 ;
    RECT 14.88 8.71 14.95 9.115 ;
    RECT 14.88 9.995 14.95 10.205 ;
    RECT 15.69 12.605 15.955 12.675 ;
    RECT 16.15 8.325 16.22 8.395 ;
    RECT 16.15 8.325 16.42 9.115 ;
    RECT 16.15 8.71 16.22 8.97 ;
    RECT 16.15 9.995 16.42 10.205 ;
    RECT 16.18 2.99 16.39 3.955 ;
    RECT 16.18 4.815 16.39 5.025 ;
    RECT 16.18 6.315 16.39 6.385 ;
    RECT 84.6 4.445 84.67 4.655 ;
    RECT 10.955 5.255 11.235 5.325 ;
    RECT 10.955 8.065 11.235 8.135 ;
    RECT 10.955 11.985 11.235 12.195 ;
    RECT 10.99 3.32 11.2 3.53 ;
    RECT 10.99 4.445 11.2 4.655 ;
    RECT 10.99 6.12 11.2 6.19 ;
    RECT 11.36 3.035 11.43 3.105 ;
    RECT 11.36 3.78 11.43 3.85 ;
    RECT 11.36 4.86 11.43 4.93 ;
    RECT 11.36 6.315 11.43 6.385 ;
    RECT 11.36 6.745 11.43 6.815 ;
    RECT 11.36 12.31 11.43 12.38 ;
    RECT 11.56 4.23 11.63 4.3 ;
    RECT 11.56 7.135 11.63 7.205 ;
    RECT 11.56 8.325 11.63 8.395 ;
    RECT 11.56 8.71 11.63 9.115 ;
    RECT 11.56 9.995 11.63 10.205 ;
    RECT 12.37 12.605 12.635 12.675 ;
    RECT 12.83 8.325 12.9 8.395 ;
    RECT 12.83 8.325 13.1 9.115 ;
    RECT 12.83 8.71 12.9 8.97 ;
    RECT 12.83 9.995 13.1 10.205 ;
    RECT 12.86 2.99 13.07 3.955 ;
    RECT 12.86 4.815 13.07 5.025 ;
    RECT 12.86 6.315 13.07 6.385 ;
    RECT 7.635 5.255 7.915 5.325 ;
    RECT 7.635 8.065 7.915 8.135 ;
    RECT 7.635 11.985 7.915 12.195 ;
    RECT 7.67 3.32 7.88 3.53 ;
    RECT 7.67 4.445 7.88 4.655 ;
    RECT 7.67 6.12 7.88 6.19 ;
    RECT 8.04 3.035 8.11 3.105 ;
    RECT 8.04 3.78 8.11 3.85 ;
    RECT 8.04 4.86 8.11 4.93 ;
    RECT 8.04 6.315 8.11 6.385 ;
    RECT 8.04 6.745 8.11 6.815 ;
    RECT 8.04 12.31 8.11 12.38 ;
    RECT 8.24 4.23 8.31 4.3 ;
    RECT 8.24 7.135 8.31 7.205 ;
    RECT 8.24 8.325 8.31 8.395 ;
    RECT 8.24 8.71 8.31 9.115 ;
    RECT 8.24 9.995 8.31 10.205 ;
    RECT 9.05 12.605 9.315 12.675 ;
    RECT 9.51 8.325 9.58 8.395 ;
    RECT 9.51 8.325 9.78 9.115 ;
    RECT 9.51 8.71 9.58 8.97 ;
    RECT 9.51 9.995 9.78 10.205 ;
    RECT 9.54 2.99 9.75 3.955 ;
    RECT 9.54 4.815 9.75 5.025 ;
    RECT 9.54 6.315 9.75 6.385 ;
    RECT 78.31 7.565 78.52 7.635 ;
    RECT 4.315 5.255 4.595 5.325 ;
    RECT 4.315 8.065 4.595 8.135 ;
    RECT 4.315 11.985 4.595 12.195 ;
    RECT 4.35 3.32 4.56 3.53 ;
    RECT 4.35 4.445 4.56 4.655 ;
    RECT 4.35 6.12 4.56 6.19 ;
    RECT 4.72 3.035 4.79 3.105 ;
    RECT 4.72 3.78 4.79 3.85 ;
    RECT 4.72 4.86 4.79 4.93 ;
    RECT 4.72 6.315 4.79 6.385 ;
    RECT 4.72 6.745 4.79 6.815 ;
    RECT 4.72 12.31 4.79 12.38 ;
    RECT 4.92 4.23 4.99 4.3 ;
    RECT 4.92 7.135 4.99 7.205 ;
    RECT 4.92 8.325 4.99 8.395 ;
    RECT 4.92 8.71 4.99 9.115 ;
    RECT 4.92 9.995 4.99 10.205 ;
    RECT 5.73 12.605 5.995 12.675 ;
    RECT 6.19 8.325 6.26 8.395 ;
    RECT 6.19 8.325 6.46 9.115 ;
    RECT 6.19 8.71 6.26 8.97 ;
    RECT 6.19 9.995 6.46 10.205 ;
    RECT 6.22 2.99 6.43 3.955 ;
    RECT 6.22 4.815 6.43 5.025 ;
    RECT 6.22 6.315 6.43 6.385 ;
    RECT 84.03 7.125 84.24 7.195 ;
    RECT 84.03 4.22 84.24 4.29 ;
    RECT 11.91 7.565 12.12 7.635 ;
    RECT 74.99 9.995 75.2 10.205 ;
    RECT 74.99 8.902 75.2 9.112 ;
    RECT 74.99 8.705 75.2 8.775 ;
    RECT 107.84 6.12 107.91 6.19 ;
    RECT 74.99 8.325 75.2 8.395 ;
    RECT 74.99 6.315 75.2 6.385 ;
    RECT 74.99 4.815 75.2 5.025 ;
    RECT 108.19 7.565 108.4 7.635 ;
    RECT 107.84 5.182 107.91 5.392 ;
    RECT 113.875 5.255 114.155 5.325 ;
    RECT 113.875 8.065 114.155 8.135 ;
    RECT 113.875 11.985 114.155 12.195 ;
    RECT 113.91 3.32 114.12 3.53 ;
    RECT 113.91 4.445 114.12 4.655 ;
    RECT 113.91 6.12 114.12 6.19 ;
    RECT 114.28 3.035 114.35 3.105 ;
    RECT 114.28 3.78 114.35 3.85 ;
    RECT 114.28 4.86 114.35 4.93 ;
    RECT 114.28 6.315 114.35 6.385 ;
    RECT 114.28 6.745 114.35 6.815 ;
    RECT 114.28 12.31 114.35 12.38 ;
    RECT 114.48 4.23 114.55 4.3 ;
    RECT 114.48 7.135 114.55 7.205 ;
    RECT 114.48 8.325 114.55 8.395 ;
    RECT 114.48 8.71 114.55 9.115 ;
    RECT 114.48 9.995 114.55 10.205 ;
    RECT 115.29 12.605 115.555 12.675 ;
    RECT 115.75 8.325 115.82 8.395 ;
    RECT 115.75 8.325 116.02 9.115 ;
    RECT 115.75 8.71 115.82 8.97 ;
    RECT 115.75 9.995 116.02 10.205 ;
    RECT 115.78 2.99 115.99 3.955 ;
    RECT 115.78 4.815 115.99 5.025 ;
    RECT 115.78 6.315 115.99 6.385 ;
    RECT 107.84 4.445 107.91 4.655 ;
    RECT 110.555 5.255 110.835 5.325 ;
    RECT 110.555 8.065 110.835 8.135 ;
    RECT 110.555 11.985 110.835 12.195 ;
    RECT 110.59 3.32 110.8 3.53 ;
    RECT 110.59 4.445 110.8 4.655 ;
    RECT 110.59 6.12 110.8 6.19 ;
    RECT 110.96 3.035 111.03 3.105 ;
    RECT 110.96 3.78 111.03 3.85 ;
    RECT 110.96 4.86 111.03 4.93 ;
    RECT 110.96 6.315 111.03 6.385 ;
    RECT 110.96 6.745 111.03 6.815 ;
    RECT 110.96 12.31 111.03 12.38 ;
    RECT 111.16 4.23 111.23 4.3 ;
    RECT 111.16 7.135 111.23 7.205 ;
    RECT 111.16 8.325 111.23 8.395 ;
    RECT 111.16 8.71 111.23 9.115 ;
    RECT 111.16 9.995 111.23 10.205 ;
    RECT 111.97 12.605 112.235 12.675 ;
    RECT 112.43 8.325 112.5 8.395 ;
    RECT 112.43 8.325 112.7 9.115 ;
    RECT 112.43 8.71 112.5 8.97 ;
    RECT 112.43 9.995 112.7 10.205 ;
    RECT 112.46 2.99 112.67 3.955 ;
    RECT 112.46 4.815 112.67 5.025 ;
    RECT 112.46 6.315 112.67 6.385 ;
    RECT 74.99 3.742 75.2 3.952 ;
    RECT 107.235 5.255 107.515 5.325 ;
    RECT 107.235 8.065 107.515 8.135 ;
    RECT 107.235 11.985 107.515 12.195 ;
    RECT 107.27 3.32 107.48 3.53 ;
    RECT 107.27 4.445 107.48 4.655 ;
    RECT 107.27 6.12 107.48 6.19 ;
    RECT 107.64 3.035 107.71 3.105 ;
    RECT 107.64 3.78 107.71 3.85 ;
    RECT 107.64 4.86 107.71 4.93 ;
    RECT 107.64 6.315 107.71 6.385 ;
    RECT 107.64 6.745 107.71 6.815 ;
    RECT 107.64 12.31 107.71 12.38 ;
    RECT 107.84 4.23 107.91 4.3 ;
    RECT 107.84 7.135 107.91 7.205 ;
    RECT 107.84 8.325 107.91 8.395 ;
    RECT 107.84 8.71 107.91 9.115 ;
    RECT 107.84 9.995 107.91 10.205 ;
    RECT 108.65 12.605 108.915 12.675 ;
    RECT 109.11 8.325 109.18 8.395 ;
    RECT 109.11 8.325 109.38 9.115 ;
    RECT 109.11 8.71 109.18 8.97 ;
    RECT 109.11 9.995 109.38 10.205 ;
    RECT 109.14 2.99 109.35 3.955 ;
    RECT 109.14 4.815 109.35 5.025 ;
    RECT 109.14 6.315 109.35 6.385 ;
    RECT 74.99 2.99 75.2 3.2 ;
    RECT 103.915 5.255 104.195 5.325 ;
    RECT 103.915 8.065 104.195 8.135 ;
    RECT 103.915 11.985 104.195 12.195 ;
    RECT 103.95 3.32 104.16 3.53 ;
    RECT 103.95 4.445 104.16 4.655 ;
    RECT 103.95 6.12 104.16 6.19 ;
    RECT 104.32 3.035 104.39 3.105 ;
    RECT 104.32 3.78 104.39 3.85 ;
    RECT 104.32 4.86 104.39 4.93 ;
    RECT 104.32 6.315 104.39 6.385 ;
    RECT 104.32 6.745 104.39 6.815 ;
    RECT 104.32 12.31 104.39 12.38 ;
    RECT 104.52 4.23 104.59 4.3 ;
    RECT 104.52 7.135 104.59 7.205 ;
    RECT 104.52 8.325 104.59 8.395 ;
    RECT 104.52 8.71 104.59 9.115 ;
    RECT 104.52 9.995 104.59 10.205 ;
    RECT 105.33 12.605 105.595 12.675 ;
    RECT 105.79 8.325 105.86 8.395 ;
    RECT 105.79 8.325 106.06 9.115 ;
    RECT 105.79 8.71 105.86 8.97 ;
    RECT 105.79 9.995 106.06 10.205 ;
    RECT 105.82 2.99 106.03 3.955 ;
    RECT 105.82 4.815 106.03 5.025 ;
    RECT 105.82 6.315 106.03 6.385 ;
    RECT 107.27 7.125 107.48 7.195 ;
    RECT 45.11 7.565 45.32 7.635 ;
    RECT 100.595 5.255 100.875 5.325 ;
    RECT 100.595 8.065 100.875 8.135 ;
    RECT 100.595 11.985 100.875 12.195 ;
    RECT 100.63 3.32 100.84 3.53 ;
    RECT 100.63 4.445 100.84 4.655 ;
    RECT 100.63 6.12 100.84 6.19 ;
    RECT 101.0 3.035 101.07 3.105 ;
    RECT 101.0 3.78 101.07 3.85 ;
    RECT 101.0 4.86 101.07 4.93 ;
    RECT 101.0 6.315 101.07 6.385 ;
    RECT 101.0 6.745 101.07 6.815 ;
    RECT 101.0 12.31 101.07 12.38 ;
    RECT 101.2 4.23 101.27 4.3 ;
    RECT 101.2 7.135 101.27 7.205 ;
    RECT 101.2 8.325 101.27 8.395 ;
    RECT 101.2 8.71 101.27 9.115 ;
    RECT 101.2 9.995 101.27 10.205 ;
    RECT 102.01 12.605 102.275 12.675 ;
    RECT 102.47 8.325 102.54 8.395 ;
    RECT 102.47 8.325 102.74 9.115 ;
    RECT 102.47 8.71 102.54 8.97 ;
    RECT 102.47 9.995 102.74 10.205 ;
    RECT 102.5 2.99 102.71 3.955 ;
    RECT 102.5 4.815 102.71 5.025 ;
    RECT 102.5 6.315 102.71 6.385 ;
    RECT 107.27 4.22 107.48 4.29 ;
    RECT 118.15 9.995 118.36 10.205 ;
    RECT 118.15 8.902 118.36 9.112 ;
    RECT 97.275 5.255 97.555 5.325 ;
    RECT 97.275 8.065 97.555 8.135 ;
    RECT 97.275 11.985 97.555 12.195 ;
    RECT 97.31 3.32 97.52 3.53 ;
    RECT 97.31 4.445 97.52 4.655 ;
    RECT 97.31 6.12 97.52 6.19 ;
    RECT 97.68 3.035 97.75 3.105 ;
    RECT 97.68 3.78 97.75 3.85 ;
    RECT 97.68 4.86 97.75 4.93 ;
    RECT 97.68 6.315 97.75 6.385 ;
    RECT 97.68 6.745 97.75 6.815 ;
    RECT 97.68 12.31 97.75 12.38 ;
    RECT 97.88 4.23 97.95 4.3 ;
    RECT 97.88 7.135 97.95 7.205 ;
    RECT 97.88 8.325 97.95 8.395 ;
    RECT 97.88 8.71 97.95 9.115 ;
    RECT 97.88 9.995 97.95 10.205 ;
    RECT 98.69 12.605 98.955 12.675 ;
    RECT 99.15 8.325 99.22 8.395 ;
    RECT 99.15 8.325 99.42 9.115 ;
    RECT 99.15 8.71 99.22 8.97 ;
    RECT 99.15 9.995 99.42 10.205 ;
    RECT 99.18 2.99 99.39 3.955 ;
    RECT 99.18 4.815 99.39 5.025 ;
    RECT 99.18 6.315 99.39 6.385 ;
    RECT 118.15 8.705 118.36 8.775 ;
    RECT 93.955 5.255 94.235 5.325 ;
    RECT 93.955 8.065 94.235 8.135 ;
    RECT 93.955 11.985 94.235 12.195 ;
    RECT 93.99 3.32 94.2 3.53 ;
    RECT 93.99 4.445 94.2 4.655 ;
    RECT 93.99 6.12 94.2 6.19 ;
    RECT 94.36 3.035 94.43 3.105 ;
    RECT 94.36 3.78 94.43 3.85 ;
    RECT 94.36 4.86 94.43 4.93 ;
    RECT 94.36 6.315 94.43 6.385 ;
    RECT 94.36 6.745 94.43 6.815 ;
    RECT 94.36 12.31 94.43 12.38 ;
    RECT 94.56 4.23 94.63 4.3 ;
    RECT 94.56 7.135 94.63 7.205 ;
    RECT 94.56 8.325 94.63 8.395 ;
    RECT 94.56 8.71 94.63 9.115 ;
    RECT 94.56 9.995 94.63 10.205 ;
    RECT 95.37 12.605 95.635 12.675 ;
    RECT 95.83 8.325 95.9 8.395 ;
    RECT 95.83 8.325 96.1 9.115 ;
    RECT 95.83 8.71 95.9 8.97 ;
    RECT 95.83 9.995 96.1 10.205 ;
    RECT 95.86 2.99 96.07 3.955 ;
    RECT 95.86 4.815 96.07 5.025 ;
    RECT 95.86 6.315 96.07 6.385 ;
    RECT 118.15 8.325 118.36 8.395 ;
    RECT 90.635 5.255 90.915 5.325 ;
    RECT 90.635 8.065 90.915 8.135 ;
    RECT 90.635 11.985 90.915 12.195 ;
    RECT 90.67 3.32 90.88 3.53 ;
    RECT 90.67 4.445 90.88 4.655 ;
    RECT 90.67 6.12 90.88 6.19 ;
    RECT 91.04 3.035 91.11 3.105 ;
    RECT 91.04 3.78 91.11 3.85 ;
    RECT 91.04 4.86 91.11 4.93 ;
    RECT 91.04 6.315 91.11 6.385 ;
    RECT 91.04 6.745 91.11 6.815 ;
    RECT 91.04 12.31 91.11 12.38 ;
    RECT 91.24 4.23 91.31 4.3 ;
    RECT 91.24 7.135 91.31 7.205 ;
    RECT 91.24 8.325 91.31 8.395 ;
    RECT 91.24 8.71 91.31 9.115 ;
    RECT 91.24 9.995 91.31 10.205 ;
    RECT 92.05 12.605 92.315 12.675 ;
    RECT 92.51 8.325 92.58 8.395 ;
    RECT 92.51 8.325 92.78 9.115 ;
    RECT 92.51 8.71 92.58 8.97 ;
    RECT 92.51 9.995 92.78 10.205 ;
    RECT 92.54 2.99 92.75 3.955 ;
    RECT 92.54 4.815 92.75 5.025 ;
    RECT 92.54 6.315 92.75 6.385 ;
    RECT 118.15 6.315 118.36 6.385 ;
    RECT 87.315 5.255 87.595 5.325 ;
    RECT 87.315 8.065 87.595 8.135 ;
    RECT 87.315 11.985 87.595 12.195 ;
    RECT 87.35 3.32 87.56 3.53 ;
    RECT 87.35 4.445 87.56 4.655 ;
    RECT 87.35 6.12 87.56 6.19 ;
    RECT 87.72 3.035 87.79 3.105 ;
    RECT 87.72 3.78 87.79 3.85 ;
    RECT 87.72 4.86 87.79 4.93 ;
    RECT 87.72 6.315 87.79 6.385 ;
    RECT 87.72 6.745 87.79 6.815 ;
    RECT 87.72 12.31 87.79 12.38 ;
    RECT 87.92 4.23 87.99 4.3 ;
    RECT 87.92 7.135 87.99 7.205 ;
    RECT 87.92 8.325 87.99 8.395 ;
    RECT 87.92 8.71 87.99 9.115 ;
    RECT 87.92 9.995 87.99 10.205 ;
    RECT 88.73 12.605 88.995 12.675 ;
    RECT 89.19 8.325 89.26 8.395 ;
    RECT 89.19 8.325 89.46 9.115 ;
    RECT 89.19 8.71 89.26 8.97 ;
    RECT 89.19 9.995 89.46 10.205 ;
    RECT 89.22 2.99 89.43 3.955 ;
    RECT 89.22 4.815 89.43 5.025 ;
    RECT 89.22 6.315 89.43 6.385 ;
    RECT 118.15 4.815 118.36 5.025 ;
    RECT 83.995 5.255 84.275 5.325 ;
    RECT 83.995 8.065 84.275 8.135 ;
    RECT 83.995 11.985 84.275 12.195 ;
    RECT 84.03 3.32 84.24 3.53 ;
    RECT 84.03 4.445 84.24 4.655 ;
    RECT 84.03 6.12 84.24 6.19 ;
    RECT 84.4 3.035 84.47 3.105 ;
    RECT 84.4 3.78 84.47 3.85 ;
    RECT 84.4 4.86 84.47 4.93 ;
    RECT 84.4 6.315 84.47 6.385 ;
    RECT 84.4 6.745 84.47 6.815 ;
    RECT 84.4 12.31 84.47 12.38 ;
    RECT 84.6 4.23 84.67 4.3 ;
    RECT 84.6 7.135 84.67 7.205 ;
    RECT 84.6 8.325 84.67 8.395 ;
    RECT 84.6 8.71 84.67 9.115 ;
    RECT 84.6 9.995 84.67 10.205 ;
    RECT 85.41 12.605 85.675 12.675 ;
    RECT 85.87 8.325 85.94 8.395 ;
    RECT 85.87 8.325 86.14 9.115 ;
    RECT 85.87 8.71 85.94 8.97 ;
    RECT 85.87 9.995 86.14 10.205 ;
    RECT 85.9 2.99 86.11 3.955 ;
    RECT 85.9 4.815 86.11 5.025 ;
    RECT 85.9 6.315 86.11 6.385 ;
    RECT 118.15 3.742 118.36 3.952 ;
    RECT 80.675 5.255 80.955 5.325 ;
    RECT 80.675 8.065 80.955 8.135 ;
    RECT 80.675 11.985 80.955 12.195 ;
    RECT 80.71 3.32 80.92 3.53 ;
    RECT 80.71 4.445 80.92 4.655 ;
    RECT 80.71 6.12 80.92 6.19 ;
    RECT 81.08 3.035 81.15 3.105 ;
    RECT 81.08 3.78 81.15 3.85 ;
    RECT 81.08 4.86 81.15 4.93 ;
    RECT 81.08 6.315 81.15 6.385 ;
    RECT 81.08 6.745 81.15 6.815 ;
    RECT 81.08 12.31 81.15 12.38 ;
    RECT 81.28 4.23 81.35 4.3 ;
    RECT 81.28 7.135 81.35 7.205 ;
    RECT 81.28 8.325 81.35 8.395 ;
    RECT 81.28 8.71 81.35 9.115 ;
    RECT 81.28 9.995 81.35 10.205 ;
    RECT 82.09 12.605 82.355 12.675 ;
    RECT 82.55 8.325 82.62 8.395 ;
    RECT 82.55 8.325 82.82 9.115 ;
    RECT 82.55 8.71 82.62 8.97 ;
    RECT 82.55 9.995 82.82 10.205 ;
    RECT 82.58 2.99 82.79 3.955 ;
    RECT 82.58 4.815 82.79 5.025 ;
    RECT 82.58 6.315 82.79 6.385 ;
    RECT 118.15 2.99 118.36 3.2 ;
    RECT 77.355 5.255 77.635 5.325 ;
    RECT 77.355 8.065 77.635 8.135 ;
    RECT 77.355 11.985 77.635 12.195 ;
    RECT 77.39 3.32 77.6 3.53 ;
    RECT 77.39 4.445 77.6 4.655 ;
    RECT 77.39 6.12 77.6 6.19 ;
    RECT 77.76 3.035 77.83 3.105 ;
    RECT 77.76 3.78 77.83 3.85 ;
    RECT 77.76 4.86 77.83 4.93 ;
    RECT 77.76 6.315 77.83 6.385 ;
    RECT 77.76 6.745 77.83 6.815 ;
    RECT 77.76 12.31 77.83 12.38 ;
    RECT 77.96 4.23 78.03 4.3 ;
    RECT 77.96 7.135 78.03 7.205 ;
    RECT 77.96 8.325 78.03 8.395 ;
    RECT 77.96 8.71 78.03 9.115 ;
    RECT 77.96 9.995 78.03 10.205 ;
    RECT 78.77 12.605 79.035 12.675 ;
    RECT 79.23 8.325 79.3 8.395 ;
    RECT 79.23 8.325 79.5 9.115 ;
    RECT 79.23 8.71 79.3 8.97 ;
    RECT 79.23 9.995 79.5 10.205 ;
    RECT 79.26 2.99 79.47 3.955 ;
    RECT 79.26 4.815 79.47 5.025 ;
    RECT 79.26 6.315 79.47 6.385 ;
    RECT 74.035 5.255 74.315 5.325 ;
    RECT 74.035 8.065 74.315 8.135 ;
    RECT 74.035 11.985 74.315 12.195 ;
    RECT 74.07 3.32 74.28 3.53 ;
    RECT 74.07 4.445 74.28 4.655 ;
    RECT 74.07 6.12 74.28 6.19 ;
    RECT 74.44 3.035 74.51 3.105 ;
    RECT 74.44 3.78 74.51 3.85 ;
    RECT 74.44 4.86 74.51 4.93 ;
    RECT 74.44 6.315 74.51 6.385 ;
    RECT 74.44 6.745 74.51 6.815 ;
    RECT 74.44 12.31 74.51 12.38 ;
    RECT 74.64 4.23 74.71 4.3 ;
    RECT 74.64 7.135 74.71 7.205 ;
    RECT 74.64 8.325 74.71 8.395 ;
    RECT 74.64 8.71 74.71 9.115 ;
    RECT 74.64 9.995 74.71 10.205 ;
    RECT 75.45 12.605 75.715 12.675 ;
    RECT 75.91 8.325 75.98 8.395 ;
    RECT 75.91 8.325 76.18 9.115 ;
    RECT 75.91 8.71 75.98 8.97 ;
    RECT 75.91 9.995 76.18 10.205 ;
    RECT 75.94 2.99 76.15 3.955 ;
    RECT 75.94 4.815 76.15 5.025 ;
    RECT 75.94 6.315 76.15 6.385 ;
    RECT 70.715 5.255 70.995 5.325 ;
    RECT 70.715 8.065 70.995 8.135 ;
    RECT 70.715 11.985 70.995 12.195 ;
    RECT 70.75 3.32 70.96 3.53 ;
    RECT 70.75 4.445 70.96 4.655 ;
    RECT 70.75 6.12 70.96 6.19 ;
    RECT 71.12 3.035 71.19 3.105 ;
    RECT 71.12 3.78 71.19 3.85 ;
    RECT 71.12 4.86 71.19 4.93 ;
    RECT 71.12 6.315 71.19 6.385 ;
    RECT 71.12 6.745 71.19 6.815 ;
    RECT 71.12 12.31 71.19 12.38 ;
    RECT 71.32 4.23 71.39 4.3 ;
    RECT 71.32 7.135 71.39 7.205 ;
    RECT 71.32 8.325 71.39 8.395 ;
    RECT 71.32 8.71 71.39 9.115 ;
    RECT 71.32 9.995 71.39 10.205 ;
    RECT 72.13 12.605 72.395 12.675 ;
    RECT 72.59 8.325 72.66 8.395 ;
    RECT 72.59 8.325 72.86 9.115 ;
    RECT 72.59 8.71 72.66 8.97 ;
    RECT 72.59 9.995 72.86 10.205 ;
    RECT 72.62 2.99 72.83 3.955 ;
    RECT 72.62 4.815 72.83 5.025 ;
    RECT 72.62 6.315 72.83 6.385 ;
    RECT 67.395 5.255 67.675 5.325 ;
    RECT 67.395 8.065 67.675 8.135 ;
    RECT 67.395 11.985 67.675 12.195 ;
    RECT 67.43 3.32 67.64 3.53 ;
    RECT 67.43 4.445 67.64 4.655 ;
    RECT 67.43 6.12 67.64 6.19 ;
    RECT 67.8 3.035 67.87 3.105 ;
    RECT 67.8 3.78 67.87 3.85 ;
    RECT 67.8 4.86 67.87 4.93 ;
    RECT 67.8 6.315 67.87 6.385 ;
    RECT 67.8 6.745 67.87 6.815 ;
    RECT 67.8 12.31 67.87 12.38 ;
    RECT 68.0 4.23 68.07 4.3 ;
    RECT 68.0 7.135 68.07 7.205 ;
    RECT 68.0 8.325 68.07 8.395 ;
    RECT 68.0 8.71 68.07 9.115 ;
    RECT 68.0 9.995 68.07 10.205 ;
    RECT 68.81 12.605 69.075 12.675 ;
    RECT 69.27 8.325 69.34 8.395 ;
    RECT 69.27 8.325 69.54 9.115 ;
    RECT 69.27 8.71 69.34 8.97 ;
    RECT 69.27 9.995 69.54 10.205 ;
    RECT 69.3 2.99 69.51 3.955 ;
    RECT 69.3 4.815 69.51 5.025 ;
    RECT 69.3 6.315 69.51 6.385 ;
    RECT 74.99 7.565 75.2 7.635 ;
    RECT 8.59 7.565 8.8 7.635 ;
    RECT 64.075 5.255 64.355 5.325 ;
    RECT 64.075 8.065 64.355 8.135 ;
    RECT 64.075 11.985 64.355 12.195 ;
    RECT 64.11 3.32 64.32 3.53 ;
    RECT 64.11 4.445 64.32 4.655 ;
    RECT 64.11 6.12 64.32 6.19 ;
    RECT 64.48 3.035 64.55 3.105 ;
    RECT 64.48 3.78 64.55 3.85 ;
    RECT 64.48 4.86 64.55 4.93 ;
    RECT 64.48 6.315 64.55 6.385 ;
    RECT 64.48 6.745 64.55 6.815 ;
    RECT 64.48 12.31 64.55 12.38 ;
    RECT 64.68 4.23 64.75 4.3 ;
    RECT 64.68 7.135 64.75 7.205 ;
    RECT 64.68 8.325 64.75 8.395 ;
    RECT 64.68 8.71 64.75 9.115 ;
    RECT 64.68 9.995 64.75 10.205 ;
    RECT 65.49 12.605 65.755 12.675 ;
    RECT 65.95 8.325 66.02 8.395 ;
    RECT 65.95 8.325 66.22 9.115 ;
    RECT 65.95 8.71 66.02 8.97 ;
    RECT 65.95 9.995 66.22 10.205 ;
    RECT 65.98 2.99 66.19 3.955 ;
    RECT 65.98 4.815 66.19 5.025 ;
    RECT 65.98 6.315 66.19 6.385 ;
    RECT 60.755 5.255 61.035 5.325 ;
    RECT 60.755 8.065 61.035 8.135 ;
    RECT 60.755 11.985 61.035 12.195 ;
    RECT 60.79 3.32 61.0 3.53 ;
    RECT 60.79 4.445 61.0 4.655 ;
    RECT 60.79 6.12 61.0 6.19 ;
    RECT 61.16 3.035 61.23 3.105 ;
    RECT 61.16 3.78 61.23 3.85 ;
    RECT 61.16 4.86 61.23 4.93 ;
    RECT 61.16 6.315 61.23 6.385 ;
    RECT 61.16 6.745 61.23 6.815 ;
    RECT 61.16 12.31 61.23 12.38 ;
    RECT 61.36 4.23 61.43 4.3 ;
    RECT 61.36 7.135 61.43 7.205 ;
    RECT 61.36 8.325 61.43 8.395 ;
    RECT 61.36 8.71 61.43 9.115 ;
    RECT 61.36 9.995 61.43 10.205 ;
    RECT 62.17 12.605 62.435 12.675 ;
    RECT 62.63 8.325 62.7 8.395 ;
    RECT 62.63 8.325 62.9 9.115 ;
    RECT 62.63 8.71 62.7 8.97 ;
    RECT 62.63 9.995 62.9 10.205 ;
    RECT 62.66 2.99 62.87 3.955 ;
    RECT 62.66 4.815 62.87 5.025 ;
    RECT 62.66 6.315 62.87 6.385 ;
    RECT 57.435 5.255 57.715 5.325 ;
    RECT 57.435 8.065 57.715 8.135 ;
    RECT 57.435 11.985 57.715 12.195 ;
    RECT 57.47 3.32 57.68 3.53 ;
    RECT 57.47 4.445 57.68 4.655 ;
    RECT 57.47 6.12 57.68 6.19 ;
    RECT 57.84 3.035 57.91 3.105 ;
    RECT 57.84 3.78 57.91 3.85 ;
    RECT 57.84 4.86 57.91 4.93 ;
    RECT 57.84 6.315 57.91 6.385 ;
    RECT 57.84 6.745 57.91 6.815 ;
    RECT 57.84 12.31 57.91 12.38 ;
    RECT 58.04 4.23 58.11 4.3 ;
    RECT 58.04 7.135 58.11 7.205 ;
    RECT 58.04 8.325 58.11 8.395 ;
    RECT 58.04 8.71 58.11 9.115 ;
    RECT 58.04 9.995 58.11 10.205 ;
    RECT 58.85 12.605 59.115 12.675 ;
    RECT 59.31 8.325 59.38 8.395 ;
    RECT 59.31 8.325 59.58 9.115 ;
    RECT 59.31 8.71 59.38 8.97 ;
    RECT 59.31 9.995 59.58 10.205 ;
    RECT 59.34 2.99 59.55 3.955 ;
    RECT 59.34 4.815 59.55 5.025 ;
    RECT 59.34 6.315 59.55 6.385 ;
    RECT 54.115 5.255 54.395 5.325 ;
    RECT 54.115 8.065 54.395 8.135 ;
    RECT 54.115 11.985 54.395 12.195 ;
    RECT 54.15 3.32 54.36 3.53 ;
    RECT 54.15 4.445 54.36 4.655 ;
    RECT 54.15 6.12 54.36 6.19 ;
    RECT 54.52 3.035 54.59 3.105 ;
    RECT 54.52 3.78 54.59 3.85 ;
    RECT 54.52 4.86 54.59 4.93 ;
    RECT 54.52 6.315 54.59 6.385 ;
    RECT 54.52 6.745 54.59 6.815 ;
    RECT 54.52 12.31 54.59 12.38 ;
    RECT 54.72 4.23 54.79 4.3 ;
    RECT 54.72 7.135 54.79 7.205 ;
    RECT 54.72 8.325 54.79 8.395 ;
    RECT 54.72 8.71 54.79 9.115 ;
    RECT 54.72 9.995 54.79 10.205 ;
    RECT 55.53 12.605 55.795 12.675 ;
    RECT 55.99 8.325 56.06 8.395 ;
    RECT 55.99 8.325 56.26 9.115 ;
    RECT 55.99 8.71 56.06 8.97 ;
    RECT 55.99 9.995 56.26 10.205 ;
    RECT 56.02 2.99 56.23 3.955 ;
    RECT 56.02 4.815 56.23 5.025 ;
    RECT 56.02 6.315 56.23 6.385 ;
    RECT 50.795 5.255 51.075 5.325 ;
    RECT 50.795 8.065 51.075 8.135 ;
    RECT 50.795 11.985 51.075 12.195 ;
    RECT 50.83 3.32 51.04 3.53 ;
    RECT 50.83 4.445 51.04 4.655 ;
    RECT 50.83 6.12 51.04 6.19 ;
    RECT 51.2 3.035 51.27 3.105 ;
    RECT 51.2 3.78 51.27 3.85 ;
    RECT 51.2 4.86 51.27 4.93 ;
    RECT 51.2 6.315 51.27 6.385 ;
    RECT 51.2 6.745 51.27 6.815 ;
    RECT 51.2 12.31 51.27 12.38 ;
    RECT 51.4 4.23 51.47 4.3 ;
    RECT 51.4 7.135 51.47 7.205 ;
    RECT 51.4 8.325 51.47 8.395 ;
    RECT 51.4 8.71 51.47 9.115 ;
    RECT 51.4 9.995 51.47 10.205 ;
    RECT 52.21 12.605 52.475 12.675 ;
    RECT 52.67 8.325 52.74 8.395 ;
    RECT 52.67 8.325 52.94 9.115 ;
    RECT 52.67 8.71 52.74 8.97 ;
    RECT 52.67 9.995 52.94 10.205 ;
    RECT 52.7 2.99 52.91 3.955 ;
    RECT 52.7 4.815 52.91 5.025 ;
    RECT 52.7 6.315 52.91 6.385 ;
    RECT 47.475 5.255 47.755 5.325 ;
    RECT 47.475 8.065 47.755 8.135 ;
    RECT 47.475 11.985 47.755 12.195 ;
    RECT 47.51 3.32 47.72 3.53 ;
    RECT 47.51 4.445 47.72 4.655 ;
    RECT 47.51 6.12 47.72 6.19 ;
    RECT 47.88 3.035 47.95 3.105 ;
    RECT 47.88 3.78 47.95 3.85 ;
    RECT 47.88 4.86 47.95 4.93 ;
    RECT 47.88 6.315 47.95 6.385 ;
    RECT 47.88 6.745 47.95 6.815 ;
    RECT 47.88 12.31 47.95 12.38 ;
    RECT 48.08 4.23 48.15 4.3 ;
    RECT 48.08 7.135 48.15 7.205 ;
    RECT 48.08 8.325 48.15 8.395 ;
    RECT 48.08 8.71 48.15 9.115 ;
    RECT 48.08 9.995 48.15 10.205 ;
    RECT 48.89 12.605 49.155 12.675 ;
    RECT 49.35 8.325 49.42 8.395 ;
    RECT 49.35 8.325 49.62 9.115 ;
    RECT 49.35 8.71 49.42 8.97 ;
    RECT 49.35 9.995 49.62 10.205 ;
    RECT 49.38 2.99 49.59 3.955 ;
    RECT 49.38 4.815 49.59 5.025 ;
    RECT 49.38 6.315 49.59 6.385 ;
    RECT 44.155 5.255 44.435 5.325 ;
    RECT 44.155 8.065 44.435 8.135 ;
    RECT 44.155 11.985 44.435 12.195 ;
    RECT 44.19 3.32 44.4 3.53 ;
    RECT 44.19 4.445 44.4 4.655 ;
    RECT 44.19 6.12 44.4 6.19 ;
    RECT 44.56 3.035 44.63 3.105 ;
    RECT 44.56 3.78 44.63 3.85 ;
    RECT 44.56 4.86 44.63 4.93 ;
    RECT 44.56 6.315 44.63 6.385 ;
    RECT 44.56 6.745 44.63 6.815 ;
    RECT 44.56 12.31 44.63 12.38 ;
    RECT 44.76 4.23 44.83 4.3 ;
    RECT 44.76 7.135 44.83 7.205 ;
    RECT 44.76 8.325 44.83 8.395 ;
    RECT 44.76 8.71 44.83 9.115 ;
    RECT 44.76 9.995 44.83 10.205 ;
    RECT 45.57 12.605 45.835 12.675 ;
    RECT 46.03 8.325 46.1 8.395 ;
    RECT 46.03 8.325 46.3 9.115 ;
    RECT 46.03 8.71 46.1 8.97 ;
    RECT 46.03 9.995 46.3 10.205 ;
    RECT 46.06 2.99 46.27 3.955 ;
    RECT 46.06 4.815 46.27 5.025 ;
    RECT 46.06 6.315 46.27 6.385 ;
    RECT 40.835 5.255 41.115 5.325 ;
    RECT 40.835 8.065 41.115 8.135 ;
    RECT 40.835 11.985 41.115 12.195 ;
    RECT 40.87 3.32 41.08 3.53 ;
    RECT 40.87 4.445 41.08 4.655 ;
    RECT 40.87 6.12 41.08 6.19 ;
    RECT 41.24 3.035 41.31 3.105 ;
    RECT 41.24 3.78 41.31 3.85 ;
    RECT 41.24 4.86 41.31 4.93 ;
    RECT 41.24 6.315 41.31 6.385 ;
    RECT 41.24 6.745 41.31 6.815 ;
    RECT 41.24 12.31 41.31 12.38 ;
    RECT 41.44 4.23 41.51 4.3 ;
    RECT 41.44 7.135 41.51 7.205 ;
    RECT 41.44 8.325 41.51 8.395 ;
    RECT 41.44 8.71 41.51 9.115 ;
    RECT 41.44 9.995 41.51 10.205 ;
    RECT 42.25 12.605 42.515 12.675 ;
    RECT 42.71 8.325 42.78 8.395 ;
    RECT 42.71 8.325 42.98 9.115 ;
    RECT 42.71 8.71 42.78 8.97 ;
    RECT 42.71 9.995 42.98 10.205 ;
    RECT 42.74 2.99 42.95 3.955 ;
    RECT 42.74 4.815 42.95 5.025 ;
    RECT 42.74 6.315 42.95 6.385 ;
    RECT 37.515 5.255 37.795 5.325 ;
    RECT 37.515 8.065 37.795 8.135 ;
    RECT 37.515 11.985 37.795 12.195 ;
    RECT 37.55 3.32 37.76 3.53 ;
    RECT 37.55 4.445 37.76 4.655 ;
    RECT 37.55 6.12 37.76 6.19 ;
    RECT 37.92 3.035 37.99 3.105 ;
    RECT 37.92 3.78 37.99 3.85 ;
    RECT 37.92 4.86 37.99 4.93 ;
    RECT 37.92 6.315 37.99 6.385 ;
    RECT 37.92 6.745 37.99 6.815 ;
    RECT 37.92 12.31 37.99 12.38 ;
    RECT 38.12 4.23 38.19 4.3 ;
    RECT 38.12 7.135 38.19 7.205 ;
    RECT 38.12 8.325 38.19 8.395 ;
    RECT 38.12 8.71 38.19 9.115 ;
    RECT 38.12 9.995 38.19 10.205 ;
    RECT 38.93 12.605 39.195 12.675 ;
    RECT 39.39 8.325 39.46 8.395 ;
    RECT 39.39 8.325 39.66 9.115 ;
    RECT 39.39 8.71 39.46 8.97 ;
    RECT 39.39 9.995 39.66 10.205 ;
    RECT 39.42 2.99 39.63 3.955 ;
    RECT 39.42 4.815 39.63 5.025 ;
    RECT 39.42 6.315 39.63 6.385 ;
    RECT 34.195 5.255 34.475 5.325 ;
    RECT 34.195 8.065 34.475 8.135 ;
    RECT 34.195 11.985 34.475 12.195 ;
    RECT 34.23 3.32 34.44 3.53 ;
    RECT 34.23 4.445 34.44 4.655 ;
    RECT 34.23 6.12 34.44 6.19 ;
    RECT 34.6 3.035 34.67 3.105 ;
    RECT 34.6 3.78 34.67 3.85 ;
    RECT 34.6 4.86 34.67 4.93 ;
    RECT 34.6 6.315 34.67 6.385 ;
    RECT 34.6 6.745 34.67 6.815 ;
    RECT 34.6 12.31 34.67 12.38 ;
    RECT 34.8 4.23 34.87 4.3 ;
    RECT 34.8 7.135 34.87 7.205 ;
    RECT 34.8 8.325 34.87 8.395 ;
    RECT 34.8 8.71 34.87 9.115 ;
    RECT 34.8 9.995 34.87 10.205 ;
    RECT 35.61 12.605 35.875 12.675 ;
    RECT 36.07 8.325 36.14 8.395 ;
    RECT 36.07 8.325 36.34 9.115 ;
    RECT 36.07 8.71 36.14 8.97 ;
    RECT 36.07 9.995 36.34 10.205 ;
    RECT 36.1 2.99 36.31 3.955 ;
    RECT 36.1 4.815 36.31 5.025 ;
    RECT 36.1 6.315 36.31 6.385 ;
    RECT 104.87 7.565 105.08 7.635 ;
    RECT 71.67 9.995 71.88 10.205 ;
    RECT 71.67 8.902 71.88 9.112 ;
    RECT 41.79 7.565 42.0 7.635 ;
    RECT 71.67 8.705 71.88 8.775 ;
    RECT 71.67 8.325 71.88 8.395 ;
    RECT 104.52 6.12 104.59 6.19 ;
    RECT 71.67 6.315 71.88 6.385 ;
    RECT 104.52 5.182 104.59 5.392 ;
    RECT 71.67 4.815 71.88 5.025 ;
    RECT 71.67 3.742 71.88 3.952 ;
    RECT 71.67 2.99 71.88 3.2 ;
    RECT 104.52 4.445 104.59 4.655 ;
    RECT 114.83 9.995 115.04 10.205 ;
    RECT 103.95 7.125 104.16 7.195 ;
    RECT 114.83 8.902 115.04 9.112 ;
    RECT 103.95 4.22 104.16 4.29 ;
    RECT 71.67 7.565 71.88 7.635 ;
    RECT 5.27 7.565 5.48 7.635 ;
    RECT 114.83 8.705 115.04 8.775 ;
    RECT 114.83 8.325 115.04 8.395 ;
    RECT 114.83 6.315 115.04 6.385 ;
    RECT 114.83 4.815 115.04 5.025 ;
    RECT 114.83 3.742 115.04 3.952 ;
    RECT 114.83 2.99 115.04 3.2 ;
    RECT 101.55 7.565 101.76 7.635 ;
    RECT 38.47 7.565 38.68 7.635 ;
    RECT 68.35 9.995 68.56 10.205 ;
    RECT 68.35 8.902 68.56 9.112 ;
    RECT 68.35 8.705 68.56 8.775 ;
    RECT 68.35 8.325 68.56 8.395 ;
    RECT 68.35 6.315 68.56 6.385 ;
    RECT 68.35 4.815 68.56 5.025 ;
    RECT 101.2 6.12 101.27 6.19 ;
    RECT 68.35 3.742 68.56 3.952 ;
    RECT 101.2 5.182 101.27 5.392 ;
    RECT 68.35 2.99 68.56 3.2 ;
    RECT 101.2 4.445 101.27 4.655 ;
    RECT 68.35 7.565 68.56 7.635 ;
    RECT 1.95 7.565 2.16 7.635 ;
    RECT 111.51 9.995 111.72 10.205 ;
    RECT 111.51 8.902 111.72 9.112 ;
    RECT 111.51 8.705 111.72 8.775 ;
    RECT 100.63 7.125 100.84 7.195 ;
    RECT 111.51 8.325 111.72 8.395 ;
    RECT 100.63 4.22 100.84 4.29 ;
    RECT 111.51 6.315 111.72 6.385 ;
    RECT 111.51 4.815 111.72 5.025 ;
    RECT 111.51 3.742 111.72 3.952 ;
    RECT 111.51 2.99 111.72 3.2 ;
    RECT 35.15 7.565 35.36 7.635 ;
    RECT 61.71 6.315 61.92 6.385 ;
    RECT 61.71 4.815 61.92 5.025 ;
    RECT 61.71 3.742 61.92 3.952 ;
    RECT 61.71 2.99 61.92 3.2 ;
    RECT 108.19 9.995 108.4 10.205 ;
    RECT 108.19 8.902 108.4 9.112 ;
    RECT 108.19 8.705 108.4 8.775 ;
    RECT 108.19 8.325 108.4 8.395 ;
    RECT 108.19 6.315 108.4 6.385 ;
    RECT 108.19 4.815 108.4 5.025 ;
    RECT 58.39 9.995 58.6 10.205 ;
    RECT 58.39 8.902 58.6 9.112 ;
    RECT 58.39 8.705 58.6 8.775 ;
    RECT 58.39 8.325 58.6 8.395 ;
    RECT 58.39 6.315 58.6 6.385 ;
    RECT 58.39 4.815 58.6 5.025 ;
    RECT 108.19 3.742 108.4 3.952 ;
    RECT 108.19 2.99 108.4 3.2 ;
    RECT 58.39 3.742 58.6 3.952 ;
    RECT 58.39 2.99 58.6 3.2 ;
    RECT 31.48 6.12 31.55 6.19 ;
    RECT 31.48 5.182 31.55 5.392 ;
    RECT 31.48 4.445 31.55 4.655 ;
    RECT 30.91 7.125 31.12 7.195 ;
    RECT 30.91 4.22 31.12 4.29 ;
    RECT 64.68 6.12 64.75 6.19 ;
    RECT 64.68 5.182 64.75 5.392 ;
    RECT 64.68 4.445 64.75 4.655 ;
    RECT 104.87 9.995 105.08 10.205 ;
    RECT 104.87 8.902 105.08 9.112 ;
    RECT 104.87 8.705 105.08 8.775 ;
    RECT 104.87 8.325 105.08 8.395 ;
    RECT 104.87 6.315 105.08 6.385 ;
    RECT 104.87 4.815 105.08 5.025 ;
    RECT 104.87 3.742 105.08 3.952 ;
    RECT 104.87 2.99 105.08 3.2 ;
    RECT 55.07 9.995 55.28 10.205 ;
    RECT 55.07 8.902 55.28 9.112 ;
    RECT 55.07 8.705 55.28 8.775 ;
    RECT 55.07 8.325 55.28 8.395 ;
    RECT 55.07 6.315 55.28 6.385 ;
    RECT 55.07 4.815 55.28 5.025 ;
    RECT 55.07 3.742 55.28 3.952 ;
    RECT 55.07 2.99 55.28 3.2 ;
    RECT 64.11 7.125 64.32 7.195 ;
    RECT 64.11 4.22 64.32 4.29 ;
    RECT 98.23 9.995 98.44 10.205 ;
    RECT 98.23 8.902 98.44 9.112 ;
    RECT 28.16 6.12 28.23 6.19 ;
    RECT 18.55 9.995 18.76 10.205 ;
    RECT 28.16 5.182 28.23 5.392 ;
    RECT 18.55 8.902 18.76 9.112 ;
    RECT 28.16 4.445 28.23 4.655 ;
    RECT 18.55 8.705 18.76 8.775 ;
    RECT 44.76 6.12 44.83 6.19 ;
    RECT 18.55 8.325 18.76 8.395 ;
    RECT 44.76 5.182 44.83 5.392 ;
    RECT 18.55 6.315 18.76 6.385 ;
    RECT 44.76 4.445 44.83 4.655 ;
    RECT 18.55 4.815 18.76 5.025 ;
    RECT 18.55 3.742 18.76 3.952 ;
    RECT 18.55 2.99 18.76 3.2 ;
    RECT 44.19 7.125 44.4 7.195 ;
    RECT 44.19 4.22 44.4 4.29 ;
    RECT 98.23 8.705 98.44 8.775 ;
    RECT 98.23 8.325 98.44 8.395 ;
    RECT 98.23 6.315 98.44 6.385 ;
    RECT 98.23 4.815 98.44 5.025 ;
    RECT 98.23 3.742 98.44 3.952 ;
    RECT 98.23 2.99 98.44 3.2 ;
    RECT 27.59 7.125 27.8 7.195 ;
    RECT 27.59 4.22 27.8 4.29 ;
    RECT 8.24 5.182 8.31 5.392 ;
    RECT 8.24 4.445 8.31 4.655 ;
    RECT 7.67 7.125 7.88 7.195 ;
    RECT 7.67 4.22 7.88 4.29 ;
    RECT 61.36 6.12 61.43 6.19 ;
    RECT 61.36 5.182 61.43 5.392 ;
    RECT 61.36 4.445 61.43 4.655 ;
    RECT 51.75 9.995 51.96 10.205 ;
    RECT 51.75 8.902 51.96 9.112 ;
    RECT 51.75 8.705 51.96 8.775 ;
    RECT 51.75 8.325 51.96 8.395 ;
    RECT 51.75 6.315 51.96 6.385 ;
    RECT 51.75 4.815 51.96 5.025 ;
    RECT 51.75 3.742 51.96 3.952 ;
    RECT 51.75 2.99 51.96 3.2 ;
    RECT 15.23 9.995 15.44 10.205 ;
    RECT 60.79 7.125 61.0 7.195 ;
    RECT 15.23 8.902 15.44 9.112 ;
    RECT 60.79 4.22 61.0 4.29 ;
    RECT 41.44 6.12 41.51 6.19 ;
    RECT 94.91 9.995 95.12 10.205 ;
    RECT 94.91 8.902 95.12 9.112 ;
    RECT 94.91 8.705 95.12 8.775 ;
    RECT 94.91 8.325 95.12 8.395 ;
    RECT 24.84 6.12 24.91 6.19 ;
    RECT 24.84 5.182 24.91 5.392 ;
    RECT 15.23 8.705 15.44 8.775 ;
    RECT 24.84 4.445 24.91 4.655 ;
    RECT 15.23 8.325 15.44 8.395 ;
    RECT 15.23 6.315 15.44 6.385 ;
    RECT 41.44 5.182 41.51 5.392 ;
    RECT 15.23 4.815 15.44 5.025 ;
    RECT 41.44 4.445 41.51 4.655 ;
    RECT 24.27 7.125 24.48 7.195 ;
    RECT 15.23 3.742 15.44 3.952 ;
    RECT 15.23 2.99 15.44 3.2 ;
    RECT 40.87 7.125 41.08 7.195 ;
    RECT 40.87 4.22 41.08 4.29 ;
    RECT 94.91 6.315 95.12 6.385 ;
    RECT 94.91 4.815 95.12 5.025 ;
    RECT 94.91 3.742 95.12 3.952 ;
    RECT 94.91 2.99 95.12 3.2 ;
    RECT 24.27 4.22 24.48 4.29 ;
    RECT 4.92 6.12 4.99 6.19 ;
    RECT 4.92 5.182 4.99 5.392 ;
    RECT 4.92 4.445 4.99 4.655 ;
    RECT 4.35 7.125 4.56 7.195 ;
    RECT 4.35 4.22 4.56 4.29 ;
    RECT 48.43 9.995 48.64 10.205 ;
    RECT 48.43 8.902 48.64 9.112 ;
    RECT 58.04 6.12 58.11 6.19 ;
    RECT 58.04 5.182 58.11 5.392 ;
    RECT 31.83 9.995 32.04 10.205 ;
    RECT 58.04 4.445 58.11 4.655 ;
    RECT 31.83 8.902 32.04 9.112 ;
    RECT 57.47 7.125 57.68 7.195 ;
    RECT 48.43 8.705 48.64 8.775 ;
    RECT 48.43 8.325 48.64 8.395 ;
    RECT 48.43 6.315 48.64 6.385 ;
    RECT 48.43 4.815 48.64 5.025 ;
    RECT 48.43 3.742 48.64 3.952 ;
    RECT 48.43 2.99 48.64 3.2 ;
    RECT 11.91 9.995 12.12 10.205 ;
    RECT 31.83 8.705 32.04 8.775 ;
    RECT 11.91 8.902 12.12 9.112 ;
    RECT 31.83 8.325 32.04 8.395 ;
    RECT 11.91 8.705 12.12 8.775 ;
    RECT 31.83 6.315 32.04 6.385 ;
    RECT 57.47 4.22 57.68 4.29 ;
    RECT 11.91 8.325 12.12 8.395 ;
    RECT 31.83 4.815 32.04 5.025 ;
    RECT 31.83 3.742 32.04 3.952 ;
    RECT 38.12 6.12 38.19 6.19 ;
    RECT 31.83 2.99 32.04 3.2 ;
    RECT 38.12 5.182 38.19 5.392 ;
    RECT 91.59 9.995 91.8 10.205 ;
    RECT 91.59 8.902 91.8 9.112 ;
    RECT 91.59 8.705 91.8 8.775 ;
    RECT 81.28 6.12 81.35 6.19 ;
    RECT 91.59 8.325 91.8 8.395 ;
    RECT 81.28 5.182 81.35 5.392 ;
    RECT 91.59 6.315 91.8 6.385 ;
    RECT 81.28 4.445 81.35 4.655 ;
    RECT 91.59 4.815 91.8 5.025 ;
    RECT 21.52 6.12 21.59 6.19 ;
    RECT 21.52 5.182 21.59 5.392 ;
    RECT 21.52 4.445 21.59 4.655 ;
    RECT 11.91 6.315 12.12 6.385 ;
    RECT 80.71 7.125 80.92 7.195 ;
    RECT 11.91 4.815 12.12 5.025 ;
    RECT 80.71 4.22 80.92 4.29 ;
    RECT 11.91 3.742 12.12 3.952 ;
    RECT 38.12 4.445 38.19 4.655 ;
    RECT 20.95 7.125 21.16 7.195 ;
    RECT 11.91 2.99 12.12 3.2 ;
    RECT 20.95 4.22 21.16 4.29 ;
    RECT 37.55 7.125 37.76 7.195 ;
    RECT 37.55 4.22 37.76 4.29 ;
    RECT 98.23 7.565 98.44 7.635 ;
    RECT 31.83 7.565 32.04 7.635 ;
    RECT 91.59 3.742 91.8 3.952 ;
    RECT 91.59 2.99 91.8 3.2 ;
    RECT 1.6 6.12 1.67 6.19 ;
    RECT 1.6 5.182 1.67 5.392 ;
    RECT 1.6 4.445 1.67 4.655 ;
    RECT 65.03 9.995 65.24 10.205 ;
    RECT 65.03 8.902 65.24 9.112 ;
    RECT 1.03 7.125 1.24 7.195 ;
    RECT 45.11 9.995 45.32 10.205 ;
    RECT 65.03 8.705 65.24 8.775 ;
    RECT 1.03 4.22 1.24 4.29 ;
    RECT 45.11 8.902 45.32 9.112 ;
    RECT 65.03 8.325 65.24 8.395 ;
    RECT 45.11 8.705 45.32 8.775 ;
    RECT 65.03 6.315 65.24 6.385 ;
    RECT 65.03 7.565 65.24 7.635 ;
    RECT 45.11 8.325 45.32 8.395 ;
    RECT 65.03 4.815 65.24 5.025 ;
    RECT 97.88 6.12 97.95 6.19 ;
    RECT 65.03 3.742 65.24 3.952 ;
    RECT 97.88 5.182 97.95 5.392 ;
    RECT 65.03 2.99 65.24 3.2 ;
    RECT 97.88 4.445 97.95 4.655 ;
    RECT 54.72 6.12 54.79 6.19 ;
    RECT 28.51 9.995 28.72 10.205 ;
    RECT 54.72 5.182 54.79 5.392 ;
    RECT 28.51 8.902 28.72 9.112 ;
    RECT 54.72 4.445 54.79 4.655 ;
    RECT 28.51 8.705 28.72 8.775 ;
    RECT 28.51 8.325 28.72 8.395 ;
    RECT 54.15 7.125 54.36 7.195 ;
    RECT 54.15 4.22 54.36 4.29 ;
    RECT 45.11 6.315 45.32 6.385 ;
    RECT 45.11 4.815 45.32 5.025 ;
    RECT 45.11 3.742 45.32 3.952 ;
    RECT 45.11 2.99 45.32 3.2 ;
    RECT 97.31 7.125 97.52 7.195 ;
    RECT 97.31 4.22 97.52 4.29 ;
    RECT 8.59 9.995 8.8 10.205 ;
    RECT 8.59 8.902 8.8 9.112 ;
    RECT 28.51 6.315 28.72 6.385 ;
    RECT 8.59 8.705 8.8 8.775 ;
    RECT 28.51 4.815 28.72 5.025 ;
    RECT 8.59 8.325 8.8 8.395 ;
    RECT 28.51 3.742 28.72 3.952 ;
    RECT 8.59 6.315 8.8 6.385 ;
    RECT 28.51 2.99 28.72 3.2 ;
    RECT 8.59 4.815 8.8 5.025 ;
    RECT 34.8 6.12 34.87 6.19 ;
    RECT 34.8 5.182 34.87 5.392 ;
    RECT 34.8 4.445 34.87 4.655 ;
    RECT 94.91 7.565 95.12 7.635 ;
    RECT 28.51 7.565 28.72 7.635 ;
    RECT 88.27 9.995 88.48 10.205 ;
    RECT 88.27 8.902 88.48 9.112 ;
    RECT 88.27 8.705 88.48 8.775 ;
    RECT 88.27 8.325 88.48 8.395 ;
    RECT 77.96 6.12 78.03 6.19 ;
    RECT 88.27 6.315 88.48 6.385 ;
    RECT 77.96 5.182 78.03 5.392 ;
    RECT 88.27 4.815 88.48 5.025 ;
    RECT 77.96 4.445 78.03 4.655 ;
    RECT 88.27 3.742 88.48 3.952 ;
    RECT 88.27 2.99 88.48 3.2 ;
    RECT 18.2 6.12 18.27 6.19 ;
    RECT 18.2 5.182 18.27 5.392 ;
    RECT 77.39 7.125 77.6 7.195 ;
    RECT 18.2 4.445 18.27 4.655 ;
    RECT 8.59 3.742 8.8 3.952 ;
    RECT 77.39 4.22 77.6 4.29 ;
    RECT 8.59 2.99 8.8 3.2 ;
    RECT 17.63 7.125 17.84 7.195 ;
    RECT 17.63 4.22 17.84 4.29 ;
    RECT 34.23 7.125 34.44 7.195 ;
    RECT 34.23 4.22 34.44 4.29 ;
    RECT 61.71 7.565 61.92 7.635 ;
    RECT 61.71 9.995 61.92 10.205 ;
    RECT 61.71 8.902 61.92 9.112 ;
    RECT 61.71 8.705 61.92 8.775 ;
    RECT 61.71 8.325 61.92 8.395 ;
    RECT 41.79 9.995 42.0 10.205 ;
    RECT 41.79 8.902 42.0 9.112 ;
    RECT 41.79 8.705 42.0 8.775 ;
    RECT 41.79 8.325 42.0 8.395 ;
    RECT 41.79 6.315 42.0 6.385 ;
    RECT 94.56 6.12 94.63 6.19 ;
    RECT 41.79 4.815 42.0 5.025 ;
    RECT 94.56 5.182 94.63 5.392 ;
    RECT 94.56 4.445 94.63 4.655 ;
    RECT 25.19 9.995 25.4 10.205 ;
    RECT 51.4 6.12 51.47 6.19 ;
    RECT 25.19 8.902 25.4 9.112 ;
    RECT 51.4 5.182 51.47 5.392 ;
    RECT 25.19 8.705 25.4 8.775 ;
    RECT 51.4 4.445 51.47 4.655 ;
    RECT 91.59 7.565 91.8 7.635 ;
    RECT 25.19 8.325 25.4 8.395 ;
    RECT 57.925 100.675 58.135 100.745 ;
    RECT 58.4 100.675 58.61 100.745 ;
    RECT 58.885 100.395 59.095 100.465 ;
    RECT 54.605 100.675 54.815 100.745 ;
    RECT 55.08 100.675 55.29 100.745 ;
    RECT 55.565 100.395 55.775 100.465 ;
    RECT 51.285 100.675 51.495 100.745 ;
    RECT 51.76 100.675 51.97 100.745 ;
    RECT 52.245 100.395 52.455 100.465 ;
    RECT 47.965 100.675 48.175 100.745 ;
    RECT 48.44 100.675 48.65 100.745 ;
    RECT 48.925 100.395 49.135 100.465 ;
    RECT 44.645 100.675 44.855 100.745 ;
    RECT 45.12 100.675 45.33 100.745 ;
    RECT 45.605 100.395 45.815 100.465 ;
    RECT 41.325 100.675 41.535 100.745 ;
    RECT 41.8 100.675 42.01 100.745 ;
    RECT 42.285 100.395 42.495 100.465 ;
    RECT 38.005 100.675 38.215 100.745 ;
    RECT 38.48 100.675 38.69 100.745 ;
    RECT 38.965 100.395 39.175 100.465 ;
    RECT 34.685 100.675 34.895 100.745 ;
    RECT 35.16 100.675 35.37 100.745 ;
    RECT 35.645 100.395 35.855 100.465 ;
    RECT 266.685 100.675 266.895 100.745 ;
    RECT 266.21 100.675 266.42 100.745 ;
    RECT 265.725 100.395 265.935 100.465 ;
    RECT 263.365 100.675 263.575 100.745 ;
    RECT 262.89 100.675 263.1 100.745 ;
    RECT 262.405 100.395 262.615 100.465 ;
    RECT 260.045 100.675 260.255 100.745 ;
    RECT 259.57 100.675 259.78 100.745 ;
    RECT 259.085 100.395 259.295 100.465 ;
    RECT 256.725 100.675 256.935 100.745 ;
    RECT 256.25 100.675 256.46 100.745 ;
    RECT 255.765 100.395 255.975 100.465 ;
    RECT 253.405 100.675 253.615 100.745 ;
    RECT 252.93 100.675 253.14 100.745 ;
    RECT 252.445 100.395 252.655 100.465 ;
    RECT 121.44 100.695 121.51 100.765 ;
    RECT 121.73 100.415 121.8 100.485 ;
    RECT 122.04 100.695 122.25 100.765 ;
    RECT 124.255 100.695 124.465 100.765 ;
    RECT 125.11 100.695 125.32 100.765 ;
    RECT 125.67 100.415 125.88 100.485 ;
    RECT 126.76 100.695 126.97 100.765 ;
    RECT 131.8 100.695 131.87 100.765 ;
    RECT 134.34 100.695 134.55 100.765 ;
    RECT 136.92 100.695 137.13 100.765 ;
    RECT 139.73 100.69 139.94 100.76 ;
    RECT 141.415 100.695 141.625 100.765 ;
    RECT 142.51 100.415 142.72 100.485 ;
    RECT 143.07 100.695 143.14 100.765 ;
    RECT 143.69 100.695 143.9 100.765 ;
    RECT 146.16 100.695 146.37 100.765 ;
    RECT 250.085 100.675 250.295 100.745 ;
    RECT 249.61 100.675 249.82 100.745 ;
    RECT 249.125 100.395 249.335 100.465 ;
    RECT 267.91 100.695 267.98 100.765 ;
    RECT 180.365 100.675 180.575 100.745 ;
    RECT 179.89 100.675 180.1 100.745 ;
    RECT 179.405 100.395 179.615 100.465 ;
    RECT 177.045 100.675 177.255 100.745 ;
    RECT 176.57 100.675 176.78 100.745 ;
    RECT 176.085 100.395 176.295 100.465 ;
    RECT 246.765 100.675 246.975 100.745 ;
    RECT 246.29 100.675 246.5 100.745 ;
    RECT 245.805 100.395 246.015 100.465 ;
    RECT 173.725 100.675 173.935 100.745 ;
    RECT 173.25 100.675 173.46 100.745 ;
    RECT 172.765 100.395 172.975 100.465 ;
    RECT 243.445 100.675 243.655 100.745 ;
    RECT 242.97 100.675 243.18 100.745 ;
    RECT 242.485 100.395 242.695 100.465 ;
    RECT 170.405 100.675 170.615 100.745 ;
    RECT 169.93 100.675 170.14 100.745 ;
    RECT 169.445 100.395 169.655 100.465 ;
    RECT 240.125 100.675 240.335 100.745 ;
    RECT 239.65 100.675 239.86 100.745 ;
    RECT 239.165 100.395 239.375 100.465 ;
    RECT 167.085 100.675 167.295 100.745 ;
    RECT 166.61 100.675 166.82 100.745 ;
    RECT 166.125 100.395 166.335 100.465 ;
    RECT 236.805 100.675 237.015 100.745 ;
    RECT 236.33 100.675 236.54 100.745 ;
    RECT 235.845 100.395 236.055 100.465 ;
    RECT 163.765 100.675 163.975 100.745 ;
    RECT 163.29 100.675 163.5 100.745 ;
    RECT 162.805 100.395 163.015 100.465 ;
    RECT 233.485 100.675 233.695 100.745 ;
    RECT 233.01 100.675 233.22 100.745 ;
    RECT 232.525 100.395 232.735 100.465 ;
    RECT 160.445 100.675 160.655 100.745 ;
    RECT 159.97 100.675 160.18 100.745 ;
    RECT 159.485 100.395 159.695 100.465 ;
    RECT 230.165 100.675 230.375 100.745 ;
    RECT 229.69 100.675 229.9 100.745 ;
    RECT 229.205 100.395 229.415 100.465 ;
    RECT 157.125 100.675 157.335 100.745 ;
    RECT 156.65 100.675 156.86 100.745 ;
    RECT 156.165 100.395 156.375 100.465 ;
    RECT 226.845 100.675 227.055 100.745 ;
    RECT 226.37 100.675 226.58 100.745 ;
    RECT 225.885 100.395 226.095 100.465 ;
    RECT 153.805 100.675 154.015 100.745 ;
    RECT 153.33 100.675 153.54 100.745 ;
    RECT 152.845 100.395 153.055 100.465 ;
    RECT 223.525 100.675 223.735 100.745 ;
    RECT 223.05 100.675 223.26 100.745 ;
    RECT 222.565 100.395 222.775 100.465 ;
    RECT 150.485 100.675 150.695 100.745 ;
    RECT 150.01 100.675 150.22 100.745 ;
    RECT 149.525 100.395 149.735 100.465 ;
    RECT 220.205 100.675 220.415 100.745 ;
    RECT 219.73 100.675 219.94 100.745 ;
    RECT 219.245 100.395 219.455 100.465 ;
    RECT 216.885 100.675 217.095 100.745 ;
    RECT 216.41 100.675 216.62 100.745 ;
    RECT 215.925 100.395 216.135 100.465 ;
    RECT 0.19 100.415 0.26 100.485 ;
    RECT 145.485 100.687 145.695 100.757 ;
    RECT 123.765 100.415 123.975 100.485 ;
    RECT 123.235 100.415 123.445 100.485 ;
    RECT 140.475 100.687 140.685 100.757 ;
    RECT 131.0 100.687 131.21 100.757 ;
    RECT 213.565 100.675 213.775 100.745 ;
    RECT 213.09 100.675 213.3 100.745 ;
    RECT 212.605 100.395 212.815 100.465 ;
    RECT 210.245 100.675 210.455 100.745 ;
    RECT 209.77 100.675 209.98 100.745 ;
    RECT 209.285 100.395 209.495 100.465 ;
    RECT 206.925 100.675 207.135 100.745 ;
    RECT 206.45 100.675 206.66 100.745 ;
    RECT 205.965 100.395 206.175 100.465 ;
    RECT 203.605 100.675 203.815 100.745 ;
    RECT 203.13 100.675 203.34 100.745 ;
    RECT 202.645 100.395 202.855 100.465 ;
    RECT 200.285 100.675 200.495 100.745 ;
    RECT 199.81 100.675 200.02 100.745 ;
    RECT 199.325 100.395 199.535 100.465 ;
    RECT 196.965 100.675 197.175 100.745 ;
    RECT 196.49 100.675 196.7 100.745 ;
    RECT 196.005 100.395 196.215 100.465 ;
    RECT 193.645 100.675 193.855 100.745 ;
    RECT 193.17 100.675 193.38 100.745 ;
    RECT 192.685 100.395 192.895 100.465 ;
    RECT 190.325 100.675 190.535 100.745 ;
    RECT 189.85 100.675 190.06 100.745 ;
    RECT 189.365 100.395 189.575 100.465 ;
    RECT 187.005 100.675 187.215 100.745 ;
    RECT 186.53 100.675 186.74 100.745 ;
    RECT 186.045 100.395 186.255 100.465 ;
    RECT 31.365 100.675 31.575 100.745 ;
    RECT 31.84 100.675 32.05 100.745 ;
    RECT 32.325 100.395 32.535 100.465 ;
    RECT 183.685 100.675 183.895 100.745 ;
    RECT 183.21 100.675 183.42 100.745 ;
    RECT 182.725 100.395 182.935 100.465 ;
    RECT 28.045 100.675 28.255 100.745 ;
    RECT 28.52 100.675 28.73 100.745 ;
    RECT 29.005 100.395 29.215 100.465 ;
    RECT 24.725 100.675 24.935 100.745 ;
    RECT 25.2 100.675 25.41 100.745 ;
    RECT 25.685 100.395 25.895 100.465 ;
    RECT 129.965 100.687 130.175 100.757 ;
    RECT 21.405 100.675 21.615 100.745 ;
    RECT 21.88 100.675 22.09 100.745 ;
    RECT 22.365 100.395 22.575 100.465 ;
    RECT 122.63 100.687 122.84 100.757 ;
    RECT 18.085 100.675 18.295 100.745 ;
    RECT 18.56 100.675 18.77 100.745 ;
    RECT 19.045 100.395 19.255 100.465 ;
    RECT 14.765 100.675 14.975 100.745 ;
    RECT 15.24 100.675 15.45 100.745 ;
    RECT 15.725 100.395 15.935 100.465 ;
    RECT 11.445 100.675 11.655 100.745 ;
    RECT 11.92 100.675 12.13 100.745 ;
    RECT 12.405 100.395 12.615 100.465 ;
    RECT 8.125 100.675 8.335 100.745 ;
    RECT 8.6 100.675 8.81 100.745 ;
    RECT 9.085 100.395 9.295 100.465 ;
    RECT 4.805 100.675 5.015 100.745 ;
    RECT 5.28 100.675 5.49 100.745 ;
    RECT 5.765 100.395 5.975 100.465 ;
    RECT 1.485 100.675 1.695 100.745 ;
    RECT 1.96 100.675 2.17 100.745 ;
    RECT 2.445 100.395 2.655 100.465 ;
    RECT 117.685 100.675 117.895 100.745 ;
    RECT 118.16 100.675 118.37 100.745 ;
    RECT 118.645 100.395 118.855 100.465 ;
    RECT 114.365 100.675 114.575 100.745 ;
    RECT 114.84 100.675 115.05 100.745 ;
    RECT 115.325 100.395 115.535 100.465 ;
    RECT 111.045 100.675 111.255 100.745 ;
    RECT 111.52 100.675 111.73 100.745 ;
    RECT 112.005 100.395 112.215 100.465 ;
    RECT 107.725 100.675 107.935 100.745 ;
    RECT 108.2 100.675 108.41 100.745 ;
    RECT 108.685 100.395 108.895 100.465 ;
    RECT 104.405 100.675 104.615 100.745 ;
    RECT 104.88 100.675 105.09 100.745 ;
    RECT 105.365 100.395 105.575 100.465 ;
    RECT 101.085 100.675 101.295 100.745 ;
    RECT 101.56 100.675 101.77 100.745 ;
    RECT 102.045 100.395 102.255 100.465 ;
    RECT 0.4 100.695 0.47 100.765 ;
    RECT 268.12 100.415 268.19 100.485 ;
    RECT 97.765 100.675 97.975 100.745 ;
    RECT 98.24 100.675 98.45 100.745 ;
    RECT 98.725 100.395 98.935 100.465 ;
    RECT 94.445 100.675 94.655 100.745 ;
    RECT 94.92 100.675 95.13 100.745 ;
    RECT 95.405 100.395 95.615 100.465 ;
    RECT 91.125 100.675 91.335 100.745 ;
    RECT 91.6 100.675 91.81 100.745 ;
    RECT 92.085 100.395 92.295 100.465 ;
    RECT 87.805 100.675 88.015 100.745 ;
    RECT 88.28 100.675 88.49 100.745 ;
    RECT 88.765 100.395 88.975 100.465 ;
    RECT 84.485 100.675 84.695 100.745 ;
    RECT 84.96 100.675 85.17 100.745 ;
    RECT 85.445 100.395 85.655 100.465 ;
    RECT 81.165 100.675 81.375 100.745 ;
    RECT 81.64 100.675 81.85 100.745 ;
    RECT 82.125 100.395 82.335 100.465 ;
    RECT 77.845 100.675 78.055 100.745 ;
    RECT 78.32 100.675 78.53 100.745 ;
    RECT 78.805 100.395 79.015 100.465 ;
    RECT 74.525 100.675 74.735 100.745 ;
    RECT 75.0 100.675 75.21 100.745 ;
    RECT 75.485 100.395 75.695 100.465 ;
    RECT 144.925 100.415 145.135 100.485 ;
    RECT 71.205 100.675 71.415 100.745 ;
    RECT 71.68 100.675 71.89 100.745 ;
    RECT 72.165 100.395 72.375 100.465 ;
    RECT 144.345 100.415 144.555 100.485 ;
    RECT 67.885 100.675 68.095 100.745 ;
    RECT 68.36 100.675 68.57 100.745 ;
    RECT 68.845 100.395 69.055 100.465 ;
    RECT 64.565 100.675 64.775 100.745 ;
    RECT 65.04 100.675 65.25 100.745 ;
    RECT 65.525 100.395 65.735 100.465 ;
    RECT 61.245 100.675 61.455 100.745 ;
    RECT 61.72 100.675 61.93 100.745 ;
    RECT 62.205 100.395 62.415 100.465 ;
    LAYER M4 DESIGNRULEWIDTH 0.165 ;
    RECT 57.96 0.0 58.03 0.33 ;
    RECT 58.03 0.0 58.1 0.695 ;
    RECT 59.305 0.385 59.585 0.695 ;
    RECT 54.64 0.0 54.71 0.33 ;
    RECT 54.71 0.0 54.78 0.695 ;
    RECT 55.985 0.385 56.265 0.695 ;
    RECT 51.32 0.0 51.39 0.33 ;
    RECT 51.39 0.0 51.46 0.695 ;
    RECT 52.665 0.385 52.945 0.695 ;
    RECT 48.0 0.0 48.07 0.33 ;
    RECT 48.07 0.0 48.14 0.695 ;
    RECT 49.345 0.385 49.625 0.695 ;
    RECT 44.68 0.0 44.75 0.33 ;
    RECT 44.75 0.0 44.82 0.695 ;
    RECT 46.025 0.385 46.305 0.695 ;
    RECT 41.36 0.0 41.43 0.33 ;
    RECT 41.43 0.0 41.5 0.695 ;
    RECT 42.705 0.385 42.985 0.695 ;
    RECT 38.04 0.0 38.11 0.33 ;
    RECT 38.11 0.0 38.18 0.695 ;
    RECT 39.385 0.385 39.665 0.695 ;
    RECT 34.72 0.0 34.79 0.33 ;
    RECT 34.79 0.0 34.86 0.695 ;
    RECT 36.065 0.385 36.345 0.695 ;
    RECT 266.79 0.0 266.86 0.33 ;
    RECT 266.72 0.0 266.79 0.695 ;
    RECT 265.235 0.385 265.515 0.695 ;
    RECT 263.47 0.0 263.54 0.33 ;
    RECT 263.4 0.0 263.47 0.695 ;
    RECT 261.915 0.385 262.195 0.695 ;
    RECT 260.15 0.0 260.22 0.33 ;
    RECT 260.08 0.0 260.15 0.695 ;
    RECT 258.595 0.385 258.875 0.695 ;
    RECT 256.83 0.0 256.9 0.33 ;
    RECT 256.76 0.0 256.83 0.695 ;
    RECT 255.275 0.385 255.555 0.695 ;
    RECT 253.51 0.0 253.58 0.33 ;
    RECT 253.44 0.0 253.51 0.695 ;
    RECT 251.955 0.385 252.235 0.695 ;
    RECT 120.445 0.0 120.525 0.695 ;
    RECT 121.195 0.0 121.33 0.695 ;
    RECT 121.62 0.0 121.97 0.695 ;
    RECT 122.555 0.0 124.12 0.695 ;
    RECT 125.39 0.0 125.545 0.695 ;
    RECT 126.005 0.32 126.63 0.695 ;
    RECT 126.005 0.0 126.24 0.32 ;
    RECT 127.1 0.0 127.25 0.695 ;
    RECT 127.6 0.0 127.995 0.695 ;
    RECT 128.285 0.0 128.605 0.695 ;
    RECT 129.035 0.0 129.315 0.695 ;
    RECT 129.785 0.0 130.485 0.695 ;
    RECT 130.775 0.0 131.285 0.695 ;
    RECT 131.955 0.0 133.505 0.695 ;
    RECT 133.855 0.0 134.205 0.695 ;
    RECT 134.685 0.0 136.4 0.695 ;
    RECT 137.2 0.0 137.52 0.695 ;
    RECT 137.8 0.0 138.26 0.695 ;
    RECT 139.06 0.0 140.785 0.695 ;
    RECT 141.075 0.0 141.28 0.695 ;
    RECT 142.28 0.0 142.44 0.695 ;
    RECT 142.79 0.0 142.96 0.695 ;
    RECT 144.03 0.0 145.765 0.695 ;
    RECT 146.505 0.0 146.695 0.695 ;
    RECT 147.045 0.0 147.185 0.695 ;
    RECT 147.855 0.0 147.935 0.695 ;
    RECT 250.19 0.0 250.26 0.33 ;
    RECT 250.12 0.0 250.19 0.695 ;
    RECT 248.635 0.385 248.915 0.695 ;
    RECT 180.47 0.0 180.54 0.33 ;
    RECT 180.4 0.0 180.47 0.695 ;
    RECT 178.915 0.385 179.195 0.695 ;
    RECT 177.15 0.0 177.22 0.33 ;
    RECT 177.08 0.0 177.15 0.695 ;
    RECT 175.595 0.385 175.875 0.695 ;
    RECT 246.87 0.0 246.94 0.33 ;
    RECT 246.8 0.0 246.87 0.695 ;
    RECT 245.315 0.385 245.595 0.695 ;
    RECT 173.83 0.0 173.9 0.33 ;
    RECT 173.76 0.0 173.83 0.695 ;
    RECT 172.275 0.385 172.555 0.695 ;
    RECT 243.55 0.0 243.62 0.33 ;
    RECT 243.48 0.0 243.55 0.695 ;
    RECT 241.995 0.385 242.275 0.695 ;
    RECT 170.51 0.0 170.58 0.33 ;
    RECT 170.44 0.0 170.51 0.695 ;
    RECT 168.955 0.385 169.235 0.695 ;
    RECT 240.23 0.0 240.3 0.33 ;
    RECT 240.16 0.0 240.23 0.695 ;
    RECT 238.675 0.385 238.955 0.695 ;
    RECT 167.19 0.0 167.26 0.33 ;
    RECT 167.12 0.0 167.19 0.695 ;
    RECT 165.635 0.385 165.915 0.695 ;
    RECT 236.91 0.0 236.98 0.33 ;
    RECT 236.84 0.0 236.91 0.695 ;
    RECT 235.355 0.385 235.635 0.695 ;
    RECT 163.87 0.0 163.94 0.33 ;
    RECT 163.8 0.0 163.87 0.695 ;
    RECT 162.315 0.385 162.595 0.695 ;
    RECT 233.59 0.0 233.66 0.33 ;
    RECT 233.52 0.0 233.59 0.695 ;
    RECT 232.035 0.385 232.315 0.695 ;
    RECT 160.55 0.0 160.62 0.33 ;
    RECT 160.48 0.0 160.55 0.695 ;
    RECT 158.995 0.385 159.275 0.695 ;
    RECT 230.27 0.0 230.34 0.33 ;
    RECT 230.2 0.0 230.27 0.695 ;
    RECT 228.715 0.385 228.995 0.695 ;
    RECT 157.23 0.0 157.3 0.33 ;
    RECT 157.16 0.0 157.23 0.695 ;
    RECT 155.675 0.385 155.955 0.695 ;
    RECT 226.95 0.0 227.02 0.33 ;
    RECT 226.88 0.0 226.95 0.695 ;
    RECT 225.395 0.385 225.675 0.695 ;
    RECT 153.91 0.0 153.98 0.33 ;
    RECT 153.84 0.0 153.91 0.695 ;
    RECT 152.355 0.385 152.635 0.695 ;
    RECT 223.63 0.0 223.7 0.33 ;
    RECT 223.56 0.0 223.63 0.695 ;
    RECT 222.075 0.385 222.355 0.695 ;
    RECT 150.59 0.0 150.66 0.33 ;
    RECT 150.52 0.0 150.59 0.695 ;
    RECT 149.035 0.385 149.315 0.695 ;
    RECT 220.31 0.0 220.38 0.33 ;
    RECT 220.24 0.0 220.31 0.695 ;
    RECT 218.755 0.385 219.035 0.695 ;
    RECT 216.99 0.0 217.06 0.33 ;
    RECT 216.92 0.0 216.99 0.695 ;
    RECT 215.435 0.385 215.715 0.695 ;
    RECT 213.67 0.0 213.74 0.33 ;
    RECT 213.6 0.0 213.67 0.695 ;
    RECT 212.115 0.385 212.395 0.695 ;
    RECT 210.35 0.0 210.42 0.33 ;
    RECT 210.28 0.0 210.35 0.695 ;
    RECT 208.795 0.385 209.075 0.695 ;
    RECT 207.03 0.0 207.1 0.33 ;
    RECT 206.96 0.0 207.03 0.695 ;
    RECT 205.475 0.385 205.755 0.695 ;
    RECT 203.71 0.0 203.78 0.33 ;
    RECT 203.64 0.0 203.71 0.695 ;
    RECT 202.155 0.385 202.435 0.695 ;
    RECT 200.39 0.0 200.46 0.33 ;
    RECT 200.32 0.0 200.39 0.695 ;
    RECT 198.835 0.385 199.115 0.695 ;
    RECT 197.07 0.0 197.14 0.33 ;
    RECT 197.0 0.0 197.07 0.695 ;
    RECT 195.515 0.385 195.795 0.695 ;
    RECT 193.75 0.0 193.82 0.33 ;
    RECT 193.68 0.0 193.75 0.695 ;
    RECT 192.195 0.385 192.475 0.695 ;
    RECT 190.43 0.0 190.5 0.33 ;
    RECT 190.36 0.0 190.43 0.695 ;
    RECT 188.875 0.385 189.155 0.695 ;
    RECT 187.11 0.0 187.18 0.33 ;
    RECT 187.04 0.0 187.11 0.695 ;
    RECT 185.555 0.385 185.835 0.695 ;
    RECT 31.4 0.0 31.47 0.33 ;
    RECT 31.47 0.0 31.54 0.695 ;
    RECT 32.745 0.385 33.025 0.695 ;
    RECT 183.79 0.0 183.86 0.33 ;
    RECT 183.72 0.0 183.79 0.695 ;
    RECT 182.235 0.385 182.515 0.695 ;
    RECT 28.08 0.0 28.15 0.33 ;
    RECT 28.15 0.0 28.22 0.695 ;
    RECT 29.425 0.385 29.705 0.695 ;
    RECT 24.76 0.0 24.83 0.33 ;
    RECT 24.83 0.0 24.9 0.695 ;
    RECT 26.105 0.385 26.385 0.695 ;
    RECT 21.44 0.0 21.51 0.33 ;
    RECT 21.51 0.0 21.58 0.695 ;
    RECT 22.785 0.385 23.065 0.695 ;
    RECT 18.12 0.0 18.19 0.33 ;
    RECT 18.19 0.0 18.26 0.695 ;
    RECT 19.465 0.385 19.745 0.695 ;
    RECT 14.8 0.0 14.87 0.33 ;
    RECT 14.87 0.0 14.94 0.695 ;
    RECT 16.145 0.385 16.425 0.695 ;
    RECT 11.48 0.0 11.55 0.33 ;
    RECT 11.55 0.0 11.62 0.695 ;
    RECT 12.825 0.385 13.105 0.695 ;
    RECT 8.16 0.0 8.23 0.33 ;
    RECT 8.23 0.0 8.3 0.695 ;
    RECT 9.505 0.385 9.785 0.695 ;
    RECT 4.84 0.0 4.91 0.33 ;
    RECT 4.91 0.0 4.98 0.695 ;
    RECT 6.185 0.385 6.465 0.695 ;
    RECT 1.52 0.0 1.59 0.33 ;
    RECT 1.59 0.0 1.66 0.695 ;
    RECT 2.865 0.385 3.145 0.695 ;
    RECT 117.72 0.0 117.79 0.33 ;
    RECT 117.79 0.0 117.86 0.695 ;
    RECT 119.065 0.385 119.345 0.695 ;
    RECT 114.4 0.0 114.47 0.33 ;
    RECT 114.47 0.0 114.54 0.695 ;
    RECT 115.745 0.385 116.025 0.695 ;
    RECT 111.08 0.0 111.15 0.33 ;
    RECT 111.15 0.0 111.22 0.695 ;
    RECT 112.425 0.385 112.705 0.695 ;
    RECT 107.76 0.0 107.83 0.33 ;
    RECT 107.83 0.0 107.9 0.695 ;
    RECT 109.105 0.385 109.385 0.695 ;
    RECT 104.44 0.0 104.51 0.33 ;
    RECT 104.51 0.0 104.58 0.695 ;
    RECT 105.785 0.385 106.065 0.695 ;
    RECT 101.12 0.0 101.19 0.33 ;
    RECT 101.19 0.0 101.26 0.695 ;
    RECT 102.465 0.385 102.745 0.695 ;
    RECT 97.8 0.0 97.87 0.33 ;
    RECT 97.87 0.0 97.94 0.695 ;
    RECT 99.145 0.385 99.425 0.695 ;
    RECT 94.48 0.0 94.55 0.33 ;
    RECT 94.55 0.0 94.62 0.695 ;
    RECT 95.825 0.385 96.105 0.695 ;
    RECT 91.16 0.0 91.23 0.33 ;
    RECT 91.23 0.0 91.3 0.695 ;
    RECT 92.505 0.385 92.785 0.695 ;
    RECT 87.84 0.0 87.91 0.33 ;
    RECT 87.91 0.0 87.98 0.695 ;
    RECT 89.185 0.385 89.465 0.695 ;
    RECT 84.52 0.0 84.59 0.33 ;
    RECT 84.59 0.0 84.66 0.695 ;
    RECT 85.865 0.385 86.145 0.695 ;
    RECT 81.2 0.0 81.27 0.33 ;
    RECT 81.27 0.0 81.34 0.695 ;
    RECT 82.545 0.385 82.825 0.695 ;
    RECT 77.88 0.0 77.95 0.33 ;
    RECT 77.95 0.0 78.02 0.695 ;
    RECT 79.225 0.385 79.505 0.695 ;
    RECT 74.56 0.0 74.63 0.33 ;
    RECT 74.63 0.0 74.7 0.695 ;
    RECT 75.905 0.385 76.185 0.695 ;
    RECT 71.24 0.0 71.31 0.33 ;
    RECT 71.31 0.0 71.38 0.695 ;
    RECT 72.585 0.385 72.865 0.695 ;
    RECT 67.92 0.0 67.99 0.33 ;
    RECT 67.99 0.0 68.06 0.695 ;
    RECT 69.265 0.385 69.545 0.695 ;
    RECT 64.6 0.0 64.67 0.33 ;
    RECT 64.67 0.0 64.74 0.695 ;
    RECT 65.945 0.385 66.225 0.695 ;
    RECT 61.28 0.0 61.35 0.33 ;
    RECT 61.35 0.0 61.42 0.695 ;
    RECT 62.625 0.385 62.905 0.695 ;
    RECT 121.21 49.785 121.33 50.505 ;
    RECT 121.62 49.785 121.97 50.505 ;
    RECT 122.555 49.785 124.12 50.505 ;
    RECT 125.39 49.785 125.545 50.505 ;
    RECT 126.005 49.785 126.63 50.505 ;
    RECT 127.1 49.785 127.25 50.505 ;
    RECT 127.6 49.785 127.995 50.505 ;
    RECT 128.285 49.785 128.605 50.505 ;
    RECT 129.035 49.785 129.315 50.505 ;
    RECT 129.785 49.785 130.485 50.505 ;
    RECT 130.775 49.785 131.285 50.505 ;
    RECT 131.955 49.785 133.505 50.505 ;
    RECT 133.855 49.785 134.205 50.505 ;
    RECT 134.86 49.785 136.4 50.505 ;
    RECT 137.2 49.785 137.52 50.505 ;
    RECT 137.8 49.785 138.26 50.505 ;
    RECT 139.06 49.785 139.6 50.505 ;
    RECT 140.07 49.785 140.785 50.505 ;
    RECT 141.075 49.785 141.28 50.505 ;
    RECT 142.28 49.785 142.44 50.505 ;
    RECT 142.79 49.785 142.96 50.505 ;
    RECT 144.03 49.785 145.765 50.505 ;
    RECT 146.505 49.785 146.695 50.505 ;
    RECT 147.045 49.785 147.17 50.505 ;
    RECT 121.21 49.065 121.33 49.785 ;
    RECT 121.62 49.065 121.97 49.785 ;
    RECT 122.555 49.065 124.12 49.785 ;
    RECT 125.39 49.065 125.545 49.785 ;
    RECT 126.005 49.065 126.63 49.785 ;
    RECT 127.1 49.065 127.25 49.785 ;
    RECT 127.6 49.065 127.995 49.785 ;
    RECT 128.285 49.065 128.605 49.785 ;
    RECT 129.035 49.065 129.315 49.785 ;
    RECT 129.785 49.065 130.485 49.785 ;
    RECT 130.775 49.065 131.285 49.785 ;
    RECT 131.955 49.065 133.505 49.785 ;
    RECT 133.855 49.065 134.205 49.785 ;
    RECT 134.86 49.065 136.4 49.785 ;
    RECT 137.2 49.065 137.52 49.785 ;
    RECT 137.8 49.065 138.26 49.785 ;
    RECT 139.06 49.065 139.6 49.785 ;
    RECT 140.07 49.065 140.785 49.785 ;
    RECT 141.075 49.065 141.28 49.785 ;
    RECT 142.28 49.065 142.44 49.785 ;
    RECT 142.79 49.065 142.96 49.785 ;
    RECT 144.03 49.065 145.765 49.785 ;
    RECT 146.505 49.065 146.695 49.785 ;
    RECT 147.045 49.065 147.17 49.785 ;
    RECT 121.21 48.345 121.33 49.065 ;
    RECT 121.62 48.345 121.97 49.065 ;
    RECT 122.555 48.345 124.12 49.065 ;
    RECT 125.39 48.345 125.545 49.065 ;
    RECT 126.005 48.345 126.63 49.065 ;
    RECT 127.1 48.345 127.25 49.065 ;
    RECT 127.6 48.345 127.995 49.065 ;
    RECT 128.285 48.345 128.605 49.065 ;
    RECT 129.035 48.345 129.315 49.065 ;
    RECT 129.785 48.345 130.485 49.065 ;
    RECT 130.775 48.345 131.285 49.065 ;
    RECT 131.955 48.345 133.505 49.065 ;
    RECT 133.855 48.345 134.205 49.065 ;
    RECT 134.86 48.345 136.4 49.065 ;
    RECT 137.2 48.345 137.52 49.065 ;
    RECT 137.8 48.345 138.26 49.065 ;
    RECT 139.06 48.345 139.6 49.065 ;
    RECT 140.07 48.345 140.785 49.065 ;
    RECT 141.075 48.345 141.28 49.065 ;
    RECT 142.28 48.345 142.44 49.065 ;
    RECT 142.79 48.345 142.96 49.065 ;
    RECT 144.03 48.345 145.765 49.065 ;
    RECT 146.505 48.345 146.695 49.065 ;
    RECT 147.045 48.345 147.17 49.065 ;
    RECT 121.21 47.625 121.33 48.345 ;
    RECT 121.62 47.625 121.97 48.345 ;
    RECT 122.555 47.625 124.12 48.345 ;
    RECT 125.39 47.625 125.545 48.345 ;
    RECT 126.005 47.625 126.63 48.345 ;
    RECT 127.1 47.625 127.25 48.345 ;
    RECT 127.6 47.625 127.995 48.345 ;
    RECT 128.285 47.625 128.605 48.345 ;
    RECT 129.035 47.625 129.315 48.345 ;
    RECT 129.785 47.625 130.485 48.345 ;
    RECT 130.775 47.625 131.285 48.345 ;
    RECT 131.955 47.625 133.505 48.345 ;
    RECT 133.855 47.625 134.205 48.345 ;
    RECT 134.86 47.625 136.4 48.345 ;
    RECT 137.2 47.625 137.52 48.345 ;
    RECT 137.8 47.625 138.26 48.345 ;
    RECT 139.06 47.625 139.6 48.345 ;
    RECT 140.07 47.625 140.785 48.345 ;
    RECT 141.075 47.625 141.28 48.345 ;
    RECT 142.28 47.625 142.44 48.345 ;
    RECT 142.79 47.625 142.96 48.345 ;
    RECT 144.03 47.625 145.765 48.345 ;
    RECT 146.505 47.625 146.695 48.345 ;
    RECT 147.045 47.625 147.17 48.345 ;
    RECT 121.21 46.905 121.33 47.625 ;
    RECT 121.62 46.905 121.97 47.625 ;
    RECT 122.555 46.905 124.12 47.625 ;
    RECT 125.39 46.905 125.545 47.625 ;
    RECT 126.005 46.905 126.63 47.625 ;
    RECT 127.1 46.905 127.25 47.625 ;
    RECT 127.6 46.905 127.995 47.625 ;
    RECT 128.285 46.905 128.605 47.625 ;
    RECT 129.035 46.905 129.315 47.625 ;
    RECT 129.785 46.905 130.485 47.625 ;
    RECT 130.775 46.905 131.285 47.625 ;
    RECT 131.955 46.905 133.505 47.625 ;
    RECT 133.855 46.905 134.205 47.625 ;
    RECT 134.86 46.905 136.4 47.625 ;
    RECT 137.2 46.905 137.52 47.625 ;
    RECT 137.8 46.905 138.26 47.625 ;
    RECT 139.06 46.905 139.6 47.625 ;
    RECT 140.07 46.905 140.785 47.625 ;
    RECT 141.075 46.905 141.28 47.625 ;
    RECT 142.28 46.905 142.44 47.625 ;
    RECT 142.79 46.905 142.96 47.625 ;
    RECT 144.03 46.905 145.765 47.625 ;
    RECT 146.505 46.905 146.695 47.625 ;
    RECT 147.045 46.905 147.17 47.625 ;
    RECT 121.21 46.185 121.33 46.905 ;
    RECT 121.62 46.185 121.97 46.905 ;
    RECT 122.555 46.185 124.12 46.905 ;
    RECT 125.39 46.185 125.545 46.905 ;
    RECT 126.005 46.185 126.63 46.905 ;
    RECT 127.1 46.185 127.25 46.905 ;
    RECT 127.6 46.185 127.995 46.905 ;
    RECT 128.285 46.185 128.605 46.905 ;
    RECT 129.035 46.185 129.315 46.905 ;
    RECT 129.785 46.185 130.485 46.905 ;
    RECT 130.775 46.185 131.285 46.905 ;
    RECT 131.955 46.185 133.505 46.905 ;
    RECT 133.855 46.185 134.205 46.905 ;
    RECT 134.86 46.185 136.4 46.905 ;
    RECT 137.2 46.185 137.52 46.905 ;
    RECT 137.8 46.185 138.26 46.905 ;
    RECT 139.06 46.185 139.6 46.905 ;
    RECT 140.07 46.185 140.785 46.905 ;
    RECT 141.075 46.185 141.28 46.905 ;
    RECT 142.28 46.185 142.44 46.905 ;
    RECT 142.79 46.185 142.96 46.905 ;
    RECT 144.03 46.185 145.765 46.905 ;
    RECT 146.505 46.185 146.695 46.905 ;
    RECT 147.045 46.185 147.17 46.905 ;
    RECT 121.21 45.465 121.33 46.185 ;
    RECT 121.62 45.465 121.97 46.185 ;
    RECT 122.555 45.465 124.12 46.185 ;
    RECT 125.39 45.465 125.545 46.185 ;
    RECT 126.005 45.465 126.63 46.185 ;
    RECT 127.1 45.465 127.25 46.185 ;
    RECT 127.6 45.465 127.995 46.185 ;
    RECT 128.285 45.465 128.605 46.185 ;
    RECT 129.035 45.465 129.315 46.185 ;
    RECT 129.785 45.465 130.485 46.185 ;
    RECT 130.775 45.465 131.285 46.185 ;
    RECT 131.955 45.465 133.505 46.185 ;
    RECT 133.855 45.465 134.205 46.185 ;
    RECT 134.86 45.465 136.4 46.185 ;
    RECT 137.2 45.465 137.52 46.185 ;
    RECT 137.8 45.465 138.26 46.185 ;
    RECT 139.06 45.465 139.6 46.185 ;
    RECT 140.07 45.465 140.785 46.185 ;
    RECT 141.075 45.465 141.28 46.185 ;
    RECT 142.28 45.465 142.44 46.185 ;
    RECT 142.79 45.465 142.96 46.185 ;
    RECT 144.03 45.465 145.765 46.185 ;
    RECT 146.505 45.465 146.695 46.185 ;
    RECT 147.045 45.465 147.17 46.185 ;
    RECT 121.21 44.745 121.33 45.465 ;
    RECT 121.62 44.745 121.97 45.465 ;
    RECT 122.555 44.745 124.12 45.465 ;
    RECT 125.39 44.745 125.545 45.465 ;
    RECT 126.005 44.745 126.63 45.465 ;
    RECT 127.1 44.745 127.25 45.465 ;
    RECT 127.6 44.745 127.995 45.465 ;
    RECT 128.285 44.745 128.605 45.465 ;
    RECT 129.035 44.745 129.315 45.465 ;
    RECT 129.785 44.745 130.485 45.465 ;
    RECT 130.775 44.745 131.285 45.465 ;
    RECT 131.955 44.745 133.505 45.465 ;
    RECT 133.855 44.745 134.205 45.465 ;
    RECT 134.86 44.745 136.4 45.465 ;
    RECT 137.2 44.745 137.52 45.465 ;
    RECT 137.8 44.745 138.26 45.465 ;
    RECT 139.06 44.745 139.6 45.465 ;
    RECT 140.07 44.745 140.785 45.465 ;
    RECT 141.075 44.745 141.28 45.465 ;
    RECT 142.28 44.745 142.44 45.465 ;
    RECT 142.79 44.745 142.96 45.465 ;
    RECT 144.03 44.745 145.765 45.465 ;
    RECT 146.505 44.745 146.695 45.465 ;
    RECT 147.045 44.745 147.17 45.465 ;
    RECT 121.21 44.025 121.33 44.745 ;
    RECT 121.62 44.025 121.97 44.745 ;
    RECT 122.555 44.025 124.12 44.745 ;
    RECT 125.39 44.025 125.545 44.745 ;
    RECT 126.005 44.025 126.63 44.745 ;
    RECT 127.1 44.025 127.25 44.745 ;
    RECT 127.6 44.025 127.995 44.745 ;
    RECT 128.285 44.025 128.605 44.745 ;
    RECT 129.035 44.025 129.315 44.745 ;
    RECT 129.785 44.025 130.485 44.745 ;
    RECT 130.775 44.025 131.285 44.745 ;
    RECT 131.955 44.025 133.505 44.745 ;
    RECT 133.855 44.025 134.205 44.745 ;
    RECT 134.86 44.025 136.4 44.745 ;
    RECT 137.2 44.025 137.52 44.745 ;
    RECT 137.8 44.025 138.26 44.745 ;
    RECT 139.06 44.025 139.6 44.745 ;
    RECT 140.07 44.025 140.785 44.745 ;
    RECT 141.075 44.025 141.28 44.745 ;
    RECT 142.28 44.025 142.44 44.745 ;
    RECT 142.79 44.025 142.96 44.745 ;
    RECT 144.03 44.025 145.765 44.745 ;
    RECT 146.505 44.025 146.695 44.745 ;
    RECT 147.045 44.025 147.17 44.745 ;
    RECT 121.21 43.305 121.33 44.025 ;
    RECT 121.62 43.305 121.97 44.025 ;
    RECT 122.555 43.305 124.12 44.025 ;
    RECT 125.39 43.305 125.545 44.025 ;
    RECT 126.005 43.305 126.63 44.025 ;
    RECT 127.1 43.305 127.25 44.025 ;
    RECT 127.6 43.305 127.995 44.025 ;
    RECT 128.285 43.305 128.605 44.025 ;
    RECT 129.035 43.305 129.315 44.025 ;
    RECT 129.785 43.305 130.485 44.025 ;
    RECT 130.775 43.305 131.285 44.025 ;
    RECT 131.955 43.305 133.505 44.025 ;
    RECT 133.855 43.305 134.205 44.025 ;
    RECT 134.86 43.305 136.4 44.025 ;
    RECT 137.2 43.305 137.52 44.025 ;
    RECT 137.8 43.305 138.26 44.025 ;
    RECT 139.06 43.305 139.6 44.025 ;
    RECT 140.07 43.305 140.785 44.025 ;
    RECT 141.075 43.305 141.28 44.025 ;
    RECT 142.28 43.305 142.44 44.025 ;
    RECT 142.79 43.305 142.96 44.025 ;
    RECT 144.03 43.305 145.765 44.025 ;
    RECT 146.505 43.305 146.695 44.025 ;
    RECT 147.045 43.305 147.17 44.025 ;
    RECT 121.21 42.585 121.33 43.305 ;
    RECT 121.62 42.585 121.97 43.305 ;
    RECT 122.555 42.585 124.12 43.305 ;
    RECT 125.39 42.585 125.545 43.305 ;
    RECT 126.005 42.585 126.63 43.305 ;
    RECT 127.1 42.585 127.25 43.305 ;
    RECT 127.6 42.585 127.995 43.305 ;
    RECT 128.285 42.585 128.605 43.305 ;
    RECT 129.035 42.585 129.315 43.305 ;
    RECT 129.785 42.585 130.485 43.305 ;
    RECT 130.775 42.585 131.285 43.305 ;
    RECT 131.955 42.585 133.505 43.305 ;
    RECT 133.855 42.585 134.205 43.305 ;
    RECT 134.86 42.585 136.4 43.305 ;
    RECT 137.2 42.585 137.52 43.305 ;
    RECT 137.8 42.585 138.26 43.305 ;
    RECT 139.06 42.585 139.6 43.305 ;
    RECT 140.07 42.585 140.785 43.305 ;
    RECT 141.075 42.585 141.28 43.305 ;
    RECT 142.28 42.585 142.44 43.305 ;
    RECT 142.79 42.585 142.96 43.305 ;
    RECT 144.03 42.585 145.765 43.305 ;
    RECT 146.505 42.585 146.695 43.305 ;
    RECT 147.045 42.585 147.17 43.305 ;
    RECT 121.21 41.865 121.33 42.585 ;
    RECT 121.62 41.865 121.97 42.585 ;
    RECT 122.555 41.865 124.12 42.585 ;
    RECT 125.39 41.865 125.545 42.585 ;
    RECT 126.005 41.865 126.63 42.585 ;
    RECT 127.1 41.865 127.25 42.585 ;
    RECT 127.6 41.865 127.995 42.585 ;
    RECT 128.285 41.865 128.605 42.585 ;
    RECT 129.035 41.865 129.315 42.585 ;
    RECT 129.785 41.865 130.485 42.585 ;
    RECT 130.775 41.865 131.285 42.585 ;
    RECT 131.955 41.865 133.505 42.585 ;
    RECT 133.855 41.865 134.205 42.585 ;
    RECT 134.86 41.865 136.4 42.585 ;
    RECT 137.2 41.865 137.52 42.585 ;
    RECT 137.8 41.865 138.26 42.585 ;
    RECT 139.06 41.865 139.6 42.585 ;
    RECT 140.07 41.865 140.785 42.585 ;
    RECT 141.075 41.865 141.28 42.585 ;
    RECT 142.28 41.865 142.44 42.585 ;
    RECT 142.79 41.865 142.96 42.585 ;
    RECT 144.03 41.865 145.765 42.585 ;
    RECT 146.505 41.865 146.695 42.585 ;
    RECT 147.045 41.865 147.17 42.585 ;
    RECT 121.21 41.145 121.33 41.865 ;
    RECT 121.62 41.145 121.97 41.865 ;
    RECT 122.555 41.145 124.12 41.865 ;
    RECT 125.39 41.145 125.545 41.865 ;
    RECT 126.005 41.145 126.63 41.865 ;
    RECT 127.1 41.145 127.25 41.865 ;
    RECT 127.6 41.145 127.995 41.865 ;
    RECT 128.285 41.145 128.605 41.865 ;
    RECT 129.035 41.145 129.315 41.865 ;
    RECT 129.785 41.145 130.485 41.865 ;
    RECT 130.775 41.145 131.285 41.865 ;
    RECT 131.955 41.145 133.505 41.865 ;
    RECT 133.855 41.145 134.205 41.865 ;
    RECT 134.86 41.145 136.4 41.865 ;
    RECT 137.2 41.145 137.52 41.865 ;
    RECT 137.8 41.145 138.26 41.865 ;
    RECT 139.06 41.145 139.6 41.865 ;
    RECT 140.07 41.145 140.785 41.865 ;
    RECT 141.075 41.145 141.28 41.865 ;
    RECT 142.28 41.145 142.44 41.865 ;
    RECT 142.79 41.145 142.96 41.865 ;
    RECT 144.03 41.145 145.765 41.865 ;
    RECT 146.505 41.145 146.695 41.865 ;
    RECT 147.045 41.145 147.17 41.865 ;
    RECT 121.21 40.425 121.33 41.145 ;
    RECT 121.62 40.425 121.97 41.145 ;
    RECT 122.555 40.425 124.12 41.145 ;
    RECT 125.39 40.425 125.545 41.145 ;
    RECT 126.005 40.425 126.63 41.145 ;
    RECT 127.1 40.425 127.25 41.145 ;
    RECT 127.6 40.425 127.995 41.145 ;
    RECT 128.285 40.425 128.605 41.145 ;
    RECT 129.035 40.425 129.315 41.145 ;
    RECT 129.785 40.425 130.485 41.145 ;
    RECT 130.775 40.425 131.285 41.145 ;
    RECT 131.955 40.425 133.505 41.145 ;
    RECT 133.855 40.425 134.205 41.145 ;
    RECT 134.86 40.425 136.4 41.145 ;
    RECT 137.2 40.425 137.52 41.145 ;
    RECT 137.8 40.425 138.26 41.145 ;
    RECT 139.06 40.425 139.6 41.145 ;
    RECT 140.07 40.425 140.785 41.145 ;
    RECT 141.075 40.425 141.28 41.145 ;
    RECT 142.28 40.425 142.44 41.145 ;
    RECT 142.79 40.425 142.96 41.145 ;
    RECT 144.03 40.425 145.765 41.145 ;
    RECT 146.505 40.425 146.695 41.145 ;
    RECT 147.045 40.425 147.17 41.145 ;
    RECT 121.21 39.705 121.33 40.425 ;
    RECT 121.62 39.705 121.97 40.425 ;
    RECT 122.555 39.705 124.12 40.425 ;
    RECT 125.39 39.705 125.545 40.425 ;
    RECT 126.005 39.705 126.63 40.425 ;
    RECT 127.1 39.705 127.25 40.425 ;
    RECT 127.6 39.705 127.995 40.425 ;
    RECT 128.285 39.705 128.605 40.425 ;
    RECT 129.035 39.705 129.315 40.425 ;
    RECT 129.785 39.705 130.485 40.425 ;
    RECT 130.775 39.705 131.285 40.425 ;
    RECT 131.955 39.705 133.505 40.425 ;
    RECT 133.855 39.705 134.205 40.425 ;
    RECT 134.86 39.705 136.4 40.425 ;
    RECT 137.2 39.705 137.52 40.425 ;
    RECT 137.8 39.705 138.26 40.425 ;
    RECT 139.06 39.705 139.6 40.425 ;
    RECT 140.07 39.705 140.785 40.425 ;
    RECT 141.075 39.705 141.28 40.425 ;
    RECT 142.28 39.705 142.44 40.425 ;
    RECT 142.79 39.705 142.96 40.425 ;
    RECT 144.03 39.705 145.765 40.425 ;
    RECT 146.505 39.705 146.695 40.425 ;
    RECT 147.045 39.705 147.17 40.425 ;
    RECT 121.21 38.985 121.33 39.705 ;
    RECT 121.62 38.985 121.97 39.705 ;
    RECT 122.555 38.985 124.12 39.705 ;
    RECT 125.39 38.985 125.545 39.705 ;
    RECT 126.005 38.985 126.63 39.705 ;
    RECT 127.1 38.985 127.25 39.705 ;
    RECT 127.6 38.985 127.995 39.705 ;
    RECT 128.285 38.985 128.605 39.705 ;
    RECT 129.035 38.985 129.315 39.705 ;
    RECT 129.785 38.985 130.485 39.705 ;
    RECT 130.775 38.985 131.285 39.705 ;
    RECT 131.955 38.985 133.505 39.705 ;
    RECT 133.855 38.985 134.205 39.705 ;
    RECT 134.86 38.985 136.4 39.705 ;
    RECT 137.2 38.985 137.52 39.705 ;
    RECT 137.8 38.985 138.26 39.705 ;
    RECT 139.06 38.985 139.6 39.705 ;
    RECT 140.07 38.985 140.785 39.705 ;
    RECT 141.075 38.985 141.28 39.705 ;
    RECT 142.28 38.985 142.44 39.705 ;
    RECT 142.79 38.985 142.96 39.705 ;
    RECT 144.03 38.985 145.765 39.705 ;
    RECT 146.505 38.985 146.695 39.705 ;
    RECT 147.045 38.985 147.17 39.705 ;
    RECT 121.21 38.265 121.33 38.985 ;
    RECT 121.62 38.265 121.97 38.985 ;
    RECT 122.555 38.265 124.12 38.985 ;
    RECT 125.39 38.265 125.545 38.985 ;
    RECT 126.005 38.265 126.63 38.985 ;
    RECT 127.1 38.265 127.25 38.985 ;
    RECT 127.6 38.265 127.995 38.985 ;
    RECT 128.285 38.265 128.605 38.985 ;
    RECT 129.035 38.265 129.315 38.985 ;
    RECT 129.785 38.265 130.485 38.985 ;
    RECT 130.775 38.265 131.285 38.985 ;
    RECT 131.955 38.265 133.505 38.985 ;
    RECT 133.855 38.265 134.205 38.985 ;
    RECT 134.86 38.265 136.4 38.985 ;
    RECT 137.2 38.265 137.52 38.985 ;
    RECT 137.8 38.265 138.26 38.985 ;
    RECT 139.06 38.265 139.6 38.985 ;
    RECT 140.07 38.265 140.785 38.985 ;
    RECT 141.075 38.265 141.28 38.985 ;
    RECT 142.28 38.265 142.44 38.985 ;
    RECT 142.79 38.265 142.96 38.985 ;
    RECT 144.03 38.265 145.765 38.985 ;
    RECT 146.505 38.265 146.695 38.985 ;
    RECT 147.045 38.265 147.17 38.985 ;
    RECT 121.21 37.545 121.33 38.265 ;
    RECT 121.62 37.545 121.97 38.265 ;
    RECT 122.555 37.545 124.12 38.265 ;
    RECT 125.39 37.545 125.545 38.265 ;
    RECT 126.005 37.545 126.63 38.265 ;
    RECT 127.1 37.545 127.25 38.265 ;
    RECT 127.6 37.545 127.995 38.265 ;
    RECT 128.285 37.545 128.605 38.265 ;
    RECT 129.035 37.545 129.315 38.265 ;
    RECT 129.785 37.545 130.485 38.265 ;
    RECT 130.775 37.545 131.285 38.265 ;
    RECT 131.955 37.545 133.505 38.265 ;
    RECT 133.855 37.545 134.205 38.265 ;
    RECT 134.86 37.545 136.4 38.265 ;
    RECT 137.2 37.545 137.52 38.265 ;
    RECT 137.8 37.545 138.26 38.265 ;
    RECT 139.06 37.545 139.6 38.265 ;
    RECT 140.07 37.545 140.785 38.265 ;
    RECT 141.075 37.545 141.28 38.265 ;
    RECT 142.28 37.545 142.44 38.265 ;
    RECT 142.79 37.545 142.96 38.265 ;
    RECT 144.03 37.545 145.765 38.265 ;
    RECT 146.505 37.545 146.695 38.265 ;
    RECT 147.045 37.545 147.17 38.265 ;
    RECT 121.21 14.505 121.33 37.545 ;
    RECT 121.62 14.505 121.97 37.545 ;
    RECT 122.555 14.505 124.12 37.545 ;
    RECT 125.39 14.505 125.545 37.545 ;
    RECT 126.005 14.505 126.63 37.545 ;
    RECT 127.1 14.505 127.25 37.545 ;
    RECT 127.6 14.505 127.995 37.545 ;
    RECT 128.285 32.215 128.605 37.545 ;
    RECT 129.035 14.505 129.315 37.545 ;
    RECT 129.785 14.505 130.485 37.545 ;
    RECT 130.775 14.505 131.285 37.545 ;
    RECT 131.755 15.295 131.955 26.405 ;
    RECT 131.755 27.68 131.955 28.565 ;
    RECT 131.755 30.56 131.955 36.485 ;
    RECT 131.955 14.505 131.98 37.545 ;
    RECT 131.98 14.505 132.08 37.69 ;
    RECT 132.08 14.505 132.18 37.545 ;
    RECT 132.18 14.505 132.28 37.69 ;
    RECT 132.28 14.505 132.38 37.545 ;
    RECT 132.38 14.505 132.48 37.69 ;
    RECT 132.48 14.505 132.58 37.545 ;
    RECT 132.58 14.505 132.68 37.69 ;
    RECT 132.68 14.505 132.775 37.545 ;
    RECT 132.775 14.505 132.875 37.69 ;
    RECT 132.875 14.505 132.975 37.545 ;
    RECT 132.975 14.505 133.075 37.69 ;
    RECT 133.075 14.505 133.175 37.545 ;
    RECT 133.175 14.505 133.275 37.69 ;
    RECT 133.275 14.505 133.375 37.545 ;
    RECT 133.375 14.505 133.475 37.69 ;
    RECT 133.475 14.505 133.505 37.545 ;
    RECT 133.855 14.505 134.205 37.545 ;
    RECT 134.685 14.505 134.86 36.485 ;
    RECT 134.86 14.505 134.89 37.545 ;
    RECT 134.89 14.505 134.99 37.69 ;
    RECT 134.99 14.505 135.09 37.545 ;
    RECT 135.09 14.505 135.19 37.69 ;
    RECT 135.19 14.505 135.29 37.545 ;
    RECT 135.29 14.505 135.39 37.69 ;
    RECT 135.39 14.505 135.485 37.545 ;
    RECT 135.485 14.505 135.585 37.69 ;
    RECT 135.585 14.505 135.685 37.545 ;
    RECT 135.685 14.505 135.785 37.69 ;
    RECT 135.785 14.505 135.885 37.545 ;
    RECT 135.885 14.505 135.985 37.69 ;
    RECT 135.985 14.505 136.085 37.545 ;
    RECT 136.085 14.505 136.185 37.69 ;
    RECT 136.185 14.505 136.28 37.545 ;
    RECT 136.28 14.505 136.38 37.69 ;
    RECT 136.38 14.505 136.4 37.545 ;
    RECT 137.2 14.505 137.52 37.545 ;
    RECT 137.8 14.505 138.26 37.545 ;
    RECT 139.06 14.505 139.6 37.545 ;
    RECT 140.07 14.505 140.785 37.545 ;
    RECT 141.075 14.505 141.28 37.545 ;
    RECT 142.28 14.505 142.44 37.545 ;
    RECT 142.79 14.505 142.96 37.545 ;
    RECT 144.03 14.505 145.765 37.545 ;
    RECT 146.505 14.505 146.695 37.545 ;
    RECT 147.045 14.505 147.17 37.545 ;
    RECT 121.21 98.045 121.33 98.765 ;
    RECT 121.62 98.045 121.97 98.765 ;
    RECT 122.555 98.045 124.12 98.765 ;
    RECT 125.39 98.045 125.545 98.765 ;
    RECT 126.005 98.045 126.63 98.765 ;
    RECT 127.1 98.045 127.25 98.765 ;
    RECT 127.6 98.045 127.995 98.765 ;
    RECT 128.285 98.045 128.605 98.765 ;
    RECT 129.035 98.045 129.315 98.765 ;
    RECT 129.785 98.045 130.485 98.765 ;
    RECT 130.775 98.045 131.285 98.765 ;
    RECT 131.955 98.045 133.505 98.765 ;
    RECT 133.855 98.045 134.205 98.765 ;
    RECT 134.86 98.045 136.4 98.765 ;
    RECT 137.2 98.045 137.52 98.765 ;
    RECT 137.8 98.045 138.26 98.765 ;
    RECT 139.06 98.045 139.6 98.765 ;
    RECT 140.07 98.045 140.785 98.765 ;
    RECT 141.075 98.045 141.28 98.765 ;
    RECT 142.28 98.045 142.44 98.765 ;
    RECT 142.79 98.045 142.96 98.765 ;
    RECT 144.03 98.045 145.765 98.765 ;
    RECT 146.505 98.045 146.695 98.765 ;
    RECT 147.045 98.045 147.17 98.765 ;
    RECT 121.21 97.325 121.33 98.045 ;
    RECT 121.62 97.325 121.97 98.045 ;
    RECT 122.555 97.325 124.12 98.045 ;
    RECT 125.39 97.325 125.545 98.045 ;
    RECT 126.005 97.325 126.63 98.045 ;
    RECT 127.1 97.325 127.25 98.045 ;
    RECT 127.6 97.325 127.995 98.045 ;
    RECT 128.285 97.325 128.605 98.045 ;
    RECT 129.035 97.325 129.315 98.045 ;
    RECT 129.785 97.325 130.485 98.045 ;
    RECT 130.775 97.325 131.285 98.045 ;
    RECT 131.955 97.325 133.505 98.045 ;
    RECT 133.855 97.325 134.205 98.045 ;
    RECT 134.86 97.325 136.4 98.045 ;
    RECT 137.2 97.325 137.52 98.045 ;
    RECT 137.8 97.325 138.26 98.045 ;
    RECT 139.06 97.325 139.6 98.045 ;
    RECT 140.07 97.325 140.785 98.045 ;
    RECT 141.075 97.325 141.28 98.045 ;
    RECT 142.28 97.325 142.44 98.045 ;
    RECT 142.79 97.325 142.96 98.045 ;
    RECT 144.03 97.325 145.765 98.045 ;
    RECT 146.505 97.325 146.695 98.045 ;
    RECT 147.045 97.325 147.17 98.045 ;
    RECT 121.21 96.605 121.33 97.325 ;
    RECT 121.62 96.605 121.97 97.325 ;
    RECT 122.555 96.605 124.12 97.325 ;
    RECT 125.39 96.605 125.545 97.325 ;
    RECT 126.005 96.605 126.63 97.325 ;
    RECT 127.1 96.605 127.25 97.325 ;
    RECT 127.6 96.605 127.995 97.325 ;
    RECT 128.285 96.605 128.605 97.325 ;
    RECT 129.035 96.605 129.315 97.325 ;
    RECT 129.785 96.605 130.485 97.325 ;
    RECT 130.775 96.605 131.285 97.325 ;
    RECT 131.955 96.605 133.505 97.325 ;
    RECT 133.855 96.605 134.205 97.325 ;
    RECT 134.86 96.605 136.4 97.325 ;
    RECT 137.2 96.605 137.52 97.325 ;
    RECT 137.8 96.605 138.26 97.325 ;
    RECT 139.06 96.605 139.6 97.325 ;
    RECT 140.07 96.605 140.785 97.325 ;
    RECT 141.075 96.605 141.28 97.325 ;
    RECT 142.28 96.605 142.44 97.325 ;
    RECT 142.79 96.605 142.96 97.325 ;
    RECT 144.03 96.605 145.765 97.325 ;
    RECT 146.505 96.605 146.695 97.325 ;
    RECT 147.045 96.605 147.17 97.325 ;
    RECT 121.21 95.885 121.33 96.605 ;
    RECT 121.62 95.885 121.97 96.605 ;
    RECT 122.555 95.885 124.12 96.605 ;
    RECT 125.39 95.885 125.545 96.605 ;
    RECT 126.005 95.885 126.63 96.605 ;
    RECT 127.1 95.885 127.25 96.605 ;
    RECT 127.6 95.885 127.995 96.605 ;
    RECT 128.285 95.885 128.605 96.605 ;
    RECT 129.035 95.885 129.315 96.605 ;
    RECT 129.785 95.885 130.485 96.605 ;
    RECT 130.775 95.885 131.285 96.605 ;
    RECT 131.955 95.885 133.505 96.605 ;
    RECT 133.855 95.885 134.205 96.605 ;
    RECT 134.86 95.885 136.4 96.605 ;
    RECT 137.2 95.885 137.52 96.605 ;
    RECT 137.8 95.885 138.26 96.605 ;
    RECT 139.06 95.885 139.6 96.605 ;
    RECT 140.07 95.885 140.785 96.605 ;
    RECT 141.075 95.885 141.28 96.605 ;
    RECT 142.28 95.885 142.44 96.605 ;
    RECT 142.79 95.885 142.96 96.605 ;
    RECT 144.03 95.885 145.765 96.605 ;
    RECT 146.505 95.885 146.695 96.605 ;
    RECT 147.045 95.885 147.17 96.605 ;
    RECT 121.21 98.765 121.33 100.295 ;
    RECT 121.62 98.765 121.97 99.73 ;
    RECT 122.555 98.765 124.12 100.295 ;
    RECT 125.39 98.765 125.545 100.295 ;
    RECT 126.005 98.765 126.63 100.295 ;
    RECT 127.1 98.765 127.25 100.295 ;
    RECT 127.6 98.765 127.995 100.295 ;
    RECT 128.285 98.765 128.605 100.295 ;
    RECT 129.035 98.765 129.315 100.295 ;
    RECT 129.785 98.765 130.485 100.295 ;
    RECT 130.775 98.765 131.285 100.295 ;
    RECT 131.955 98.765 131.98 100.295 ;
    RECT 131.98 98.74 132.08 100.295 ;
    RECT 132.08 98.765 133.505 100.295 ;
    RECT 133.855 98.765 134.205 100.295 ;
    RECT 134.86 98.765 136.4 100.295 ;
    RECT 137.2 98.765 137.52 100.295 ;
    RECT 137.8 98.765 138.26 100.295 ;
    RECT 139.06 98.765 139.6 100.295 ;
    RECT 140.07 98.765 140.785 100.295 ;
    RECT 141.075 98.765 141.28 100.295 ;
    RECT 142.28 98.765 142.44 100.295 ;
    RECT 142.79 98.765 142.96 100.295 ;
    RECT 144.03 98.765 145.765 100.295 ;
    RECT 146.505 98.765 146.695 100.295 ;
    RECT 147.045 98.765 147.17 100.295 ;
    RECT 121.21 95.165 121.33 95.885 ;
    RECT 121.62 95.165 121.97 95.885 ;
    RECT 122.555 95.165 124.12 95.885 ;
    RECT 125.39 95.165 125.545 95.885 ;
    RECT 126.005 95.165 126.63 95.885 ;
    RECT 127.1 95.165 127.25 95.885 ;
    RECT 127.6 95.165 127.995 95.885 ;
    RECT 128.285 95.165 128.605 95.885 ;
    RECT 129.035 95.165 129.315 95.885 ;
    RECT 129.785 95.165 130.485 95.885 ;
    RECT 130.775 95.165 131.285 95.885 ;
    RECT 131.955 95.165 133.505 95.885 ;
    RECT 133.855 95.165 134.205 95.885 ;
    RECT 134.86 95.165 136.4 95.885 ;
    RECT 137.2 95.165 137.52 95.885 ;
    RECT 137.8 95.165 138.26 95.885 ;
    RECT 139.06 95.165 139.6 95.885 ;
    RECT 140.07 95.165 140.785 95.885 ;
    RECT 141.075 95.165 141.28 95.885 ;
    RECT 142.28 95.165 142.44 95.885 ;
    RECT 142.79 95.165 142.96 95.885 ;
    RECT 144.03 95.165 145.765 95.885 ;
    RECT 146.505 95.165 146.695 95.885 ;
    RECT 147.045 95.165 147.17 95.885 ;
    RECT 121.21 94.445 121.33 95.165 ;
    RECT 121.62 94.445 121.97 95.165 ;
    RECT 122.555 94.445 124.12 95.165 ;
    RECT 125.39 94.445 125.545 95.165 ;
    RECT 126.005 94.445 126.63 95.165 ;
    RECT 127.1 94.445 127.25 95.165 ;
    RECT 127.6 94.445 127.995 95.165 ;
    RECT 128.285 94.445 128.605 95.165 ;
    RECT 129.035 94.445 129.315 95.165 ;
    RECT 129.785 94.445 130.485 95.165 ;
    RECT 130.775 94.445 131.285 95.165 ;
    RECT 131.955 94.445 133.505 95.165 ;
    RECT 133.855 94.445 134.205 95.165 ;
    RECT 134.86 94.445 136.4 95.165 ;
    RECT 137.2 94.445 137.52 95.165 ;
    RECT 137.8 94.445 138.26 95.165 ;
    RECT 139.06 94.445 139.6 95.165 ;
    RECT 140.07 94.445 140.785 95.165 ;
    RECT 141.075 94.445 141.28 95.165 ;
    RECT 142.28 94.445 142.44 95.165 ;
    RECT 142.79 94.445 142.96 95.165 ;
    RECT 144.03 94.445 145.765 95.165 ;
    RECT 146.505 94.445 146.695 95.165 ;
    RECT 147.045 94.445 147.17 95.165 ;
    RECT 121.21 93.725 121.33 94.445 ;
    RECT 121.62 93.725 121.97 94.445 ;
    RECT 122.555 93.725 124.12 94.445 ;
    RECT 125.39 93.725 125.545 94.445 ;
    RECT 126.005 93.725 126.63 94.445 ;
    RECT 127.1 93.725 127.25 94.445 ;
    RECT 127.6 93.725 127.995 94.445 ;
    RECT 128.285 93.725 128.605 94.445 ;
    RECT 129.035 93.725 129.315 94.445 ;
    RECT 129.785 93.725 130.485 94.445 ;
    RECT 130.775 93.725 131.285 94.445 ;
    RECT 131.955 93.725 133.505 94.445 ;
    RECT 133.855 93.725 134.205 94.445 ;
    RECT 134.86 93.725 136.4 94.445 ;
    RECT 137.2 93.725 137.52 94.445 ;
    RECT 137.8 93.725 138.26 94.445 ;
    RECT 139.06 93.725 139.6 94.445 ;
    RECT 140.07 93.725 140.785 94.445 ;
    RECT 141.075 93.725 141.28 94.445 ;
    RECT 142.28 93.725 142.44 94.445 ;
    RECT 142.79 93.725 142.96 94.445 ;
    RECT 144.03 93.725 145.765 94.445 ;
    RECT 146.505 93.725 146.695 94.445 ;
    RECT 147.045 93.725 147.17 94.445 ;
    RECT 121.21 93.005 121.33 93.725 ;
    RECT 121.62 93.005 121.97 93.725 ;
    RECT 122.555 93.005 124.12 93.725 ;
    RECT 125.39 93.005 125.545 93.725 ;
    RECT 126.005 93.005 126.63 93.725 ;
    RECT 127.1 93.005 127.25 93.725 ;
    RECT 127.6 93.005 127.995 93.725 ;
    RECT 128.285 93.005 128.605 93.725 ;
    RECT 129.035 93.005 129.315 93.725 ;
    RECT 129.785 93.005 130.485 93.725 ;
    RECT 130.775 93.005 131.285 93.725 ;
    RECT 131.955 93.005 133.505 93.725 ;
    RECT 133.855 93.005 134.205 93.725 ;
    RECT 134.86 93.005 136.4 93.725 ;
    RECT 137.2 93.005 137.52 93.725 ;
    RECT 137.8 93.005 138.26 93.725 ;
    RECT 139.06 93.005 139.6 93.725 ;
    RECT 140.07 93.005 140.785 93.725 ;
    RECT 141.075 93.005 141.28 93.725 ;
    RECT 142.28 93.005 142.44 93.725 ;
    RECT 142.79 93.005 142.96 93.725 ;
    RECT 144.03 93.005 145.765 93.725 ;
    RECT 146.505 93.005 146.695 93.725 ;
    RECT 147.045 93.005 147.17 93.725 ;
    RECT 121.21 92.285 121.33 93.005 ;
    RECT 121.62 92.285 121.97 93.005 ;
    RECT 122.555 92.285 124.12 93.005 ;
    RECT 125.39 92.285 125.545 93.005 ;
    RECT 126.005 92.285 126.63 93.005 ;
    RECT 127.1 92.285 127.25 93.005 ;
    RECT 127.6 92.285 127.995 93.005 ;
    RECT 128.285 92.285 128.605 93.005 ;
    RECT 129.035 92.285 129.315 93.005 ;
    RECT 129.785 92.285 130.485 93.005 ;
    RECT 130.775 92.285 131.285 93.005 ;
    RECT 131.955 92.285 133.505 93.005 ;
    RECT 133.855 92.285 134.205 93.005 ;
    RECT 134.86 92.285 136.4 93.005 ;
    RECT 137.2 92.285 137.52 93.005 ;
    RECT 137.8 92.285 138.26 93.005 ;
    RECT 139.06 92.285 139.6 93.005 ;
    RECT 140.07 92.285 140.785 93.005 ;
    RECT 141.075 92.285 141.28 93.005 ;
    RECT 142.28 92.285 142.44 93.005 ;
    RECT 142.79 92.285 142.96 93.005 ;
    RECT 144.03 92.285 145.765 93.005 ;
    RECT 146.505 92.285 146.695 93.005 ;
    RECT 147.045 92.285 147.17 93.005 ;
    RECT 121.21 91.565 121.33 92.285 ;
    RECT 121.62 91.565 121.97 92.285 ;
    RECT 122.555 91.565 124.12 92.285 ;
    RECT 125.39 91.565 125.545 92.285 ;
    RECT 126.005 91.565 126.63 92.285 ;
    RECT 127.1 91.565 127.25 92.285 ;
    RECT 127.6 91.565 127.995 92.285 ;
    RECT 128.285 91.565 128.605 92.285 ;
    RECT 129.035 91.565 129.315 92.285 ;
    RECT 129.785 91.565 130.485 92.285 ;
    RECT 130.775 91.565 131.285 92.285 ;
    RECT 131.955 91.565 133.505 92.285 ;
    RECT 133.855 91.565 134.205 92.285 ;
    RECT 134.86 91.565 136.4 92.285 ;
    RECT 137.2 91.565 137.52 92.285 ;
    RECT 137.8 91.565 138.26 92.285 ;
    RECT 139.06 91.565 139.6 92.285 ;
    RECT 140.07 91.565 140.785 92.285 ;
    RECT 141.075 91.565 141.28 92.285 ;
    RECT 142.28 91.565 142.44 92.285 ;
    RECT 142.79 91.565 142.96 92.285 ;
    RECT 144.03 91.565 145.765 92.285 ;
    RECT 146.505 91.565 146.695 92.285 ;
    RECT 147.045 91.565 147.17 92.285 ;
    RECT 121.21 90.845 121.33 91.565 ;
    RECT 121.62 90.845 121.97 91.565 ;
    RECT 122.555 90.845 124.12 91.565 ;
    RECT 125.39 90.845 125.545 91.565 ;
    RECT 126.005 90.845 126.63 91.565 ;
    RECT 127.1 90.845 127.25 91.565 ;
    RECT 127.6 90.845 127.995 91.565 ;
    RECT 128.285 90.845 128.605 91.565 ;
    RECT 129.035 90.845 129.315 91.565 ;
    RECT 129.785 90.845 130.485 91.565 ;
    RECT 130.775 90.845 131.285 91.565 ;
    RECT 131.955 90.845 133.505 91.565 ;
    RECT 133.855 90.845 134.205 91.565 ;
    RECT 134.86 90.845 136.4 91.565 ;
    RECT 137.2 90.845 137.52 91.565 ;
    RECT 137.8 90.845 138.26 91.565 ;
    RECT 139.06 90.845 139.6 91.565 ;
    RECT 140.07 90.845 140.785 91.565 ;
    RECT 141.075 90.845 141.28 91.565 ;
    RECT 142.28 90.845 142.44 91.565 ;
    RECT 142.79 90.845 142.96 91.565 ;
    RECT 144.03 90.845 145.765 91.565 ;
    RECT 146.505 90.845 146.695 91.565 ;
    RECT 147.045 90.845 147.17 91.565 ;
    RECT 121.21 90.125 121.33 90.845 ;
    RECT 121.62 90.125 121.97 90.845 ;
    RECT 122.555 90.125 124.12 90.845 ;
    RECT 125.39 90.125 125.545 90.845 ;
    RECT 126.005 90.125 126.63 90.845 ;
    RECT 127.1 90.125 127.25 90.845 ;
    RECT 127.6 90.125 127.995 90.845 ;
    RECT 128.285 90.125 128.605 90.845 ;
    RECT 129.035 90.125 129.315 90.845 ;
    RECT 129.785 90.125 130.485 90.845 ;
    RECT 130.775 90.125 131.285 90.845 ;
    RECT 131.955 90.125 133.505 90.845 ;
    RECT 133.855 90.125 134.205 90.845 ;
    RECT 134.86 90.125 136.4 90.845 ;
    RECT 137.2 90.125 137.52 90.845 ;
    RECT 137.8 90.125 138.26 90.845 ;
    RECT 139.06 90.125 139.6 90.845 ;
    RECT 140.07 90.125 140.785 90.845 ;
    RECT 141.075 90.125 141.28 90.845 ;
    RECT 142.28 90.125 142.44 90.845 ;
    RECT 142.79 90.125 142.96 90.845 ;
    RECT 144.03 90.125 145.765 90.845 ;
    RECT 146.505 90.125 146.695 90.845 ;
    RECT 147.045 90.125 147.17 90.845 ;
    RECT 121.21 89.405 121.33 90.125 ;
    RECT 121.62 89.405 121.97 90.125 ;
    RECT 122.555 89.405 124.12 90.125 ;
    RECT 125.39 89.405 125.545 90.125 ;
    RECT 126.005 89.405 126.63 90.125 ;
    RECT 127.1 89.405 127.25 90.125 ;
    RECT 127.6 89.405 127.995 90.125 ;
    RECT 128.285 89.405 128.605 90.125 ;
    RECT 129.035 89.405 129.315 90.125 ;
    RECT 129.785 89.405 130.485 90.125 ;
    RECT 130.775 89.405 131.285 90.125 ;
    RECT 131.955 89.405 133.505 90.125 ;
    RECT 133.855 89.405 134.205 90.125 ;
    RECT 134.86 89.405 136.4 90.125 ;
    RECT 137.2 89.405 137.52 90.125 ;
    RECT 137.8 89.405 138.26 90.125 ;
    RECT 139.06 89.405 139.6 90.125 ;
    RECT 140.07 89.405 140.785 90.125 ;
    RECT 141.075 89.405 141.28 90.125 ;
    RECT 142.28 89.405 142.44 90.125 ;
    RECT 142.79 89.405 142.96 90.125 ;
    RECT 144.03 89.405 145.765 90.125 ;
    RECT 146.505 89.405 146.695 90.125 ;
    RECT 147.045 89.405 147.17 90.125 ;
    RECT 121.21 88.685 121.33 89.405 ;
    RECT 121.62 88.685 121.97 89.405 ;
    RECT 122.555 88.685 124.12 89.405 ;
    RECT 125.39 88.685 125.545 89.405 ;
    RECT 126.005 88.685 126.63 89.405 ;
    RECT 127.1 88.685 127.25 89.405 ;
    RECT 127.6 88.685 127.995 89.405 ;
    RECT 128.285 88.685 128.605 89.405 ;
    RECT 129.035 88.685 129.315 89.405 ;
    RECT 129.785 88.685 130.485 89.405 ;
    RECT 130.775 88.685 131.285 89.405 ;
    RECT 131.955 88.685 133.505 89.405 ;
    RECT 133.855 88.685 134.205 89.405 ;
    RECT 134.86 88.685 136.4 89.405 ;
    RECT 137.2 88.685 137.52 89.405 ;
    RECT 137.8 88.685 138.26 89.405 ;
    RECT 139.06 88.685 139.6 89.405 ;
    RECT 140.07 88.685 140.785 89.405 ;
    RECT 141.075 88.685 141.28 89.405 ;
    RECT 142.28 88.685 142.44 89.405 ;
    RECT 142.79 88.685 142.96 89.405 ;
    RECT 144.03 88.685 145.765 89.405 ;
    RECT 146.505 88.685 146.695 89.405 ;
    RECT 147.045 88.685 147.17 89.405 ;
    RECT 121.21 60.585 121.33 61.325 ;
    RECT 121.62 60.585 121.97 61.325 ;
    RECT 122.555 60.585 124.12 61.325 ;
    RECT 125.39 60.585 125.545 61.325 ;
    RECT 126.005 60.585 126.63 61.325 ;
    RECT 127.1 60.585 127.25 61.325 ;
    RECT 127.6 60.585 127.995 61.325 ;
    RECT 128.285 60.585 128.605 61.325 ;
    RECT 129.035 60.585 129.315 61.325 ;
    RECT 129.785 60.585 130.485 61.325 ;
    RECT 130.775 60.585 131.285 61.325 ;
    RECT 131.755 60.585 133.505 61.325 ;
    RECT 133.855 60.585 134.205 61.325 ;
    RECT 134.86 60.585 136.4 61.325 ;
    RECT 137.2 60.585 137.52 61.325 ;
    RECT 137.8 60.585 138.26 61.325 ;
    RECT 139.06 60.585 139.6 61.325 ;
    RECT 140.07 60.585 140.785 61.325 ;
    RECT 141.075 60.585 141.28 61.325 ;
    RECT 142.28 60.585 142.44 61.325 ;
    RECT 142.79 60.585 142.96 61.325 ;
    RECT 144.03 60.585 145.765 61.325 ;
    RECT 146.505 60.585 146.695 61.325 ;
    RECT 147.045 60.585 147.17 61.325 ;
    RECT 121.21 87.965 121.33 88.685 ;
    RECT 121.62 87.965 121.97 88.685 ;
    RECT 122.555 87.965 124.12 88.685 ;
    RECT 125.39 87.965 125.545 88.685 ;
    RECT 126.005 87.965 126.63 88.685 ;
    RECT 127.1 87.965 127.25 88.685 ;
    RECT 127.6 87.965 127.995 88.685 ;
    RECT 128.285 87.965 128.605 88.685 ;
    RECT 129.035 87.965 129.315 88.685 ;
    RECT 129.785 87.965 130.485 88.685 ;
    RECT 130.775 87.965 131.285 88.685 ;
    RECT 131.955 87.965 133.505 88.685 ;
    RECT 133.855 87.965 134.205 88.685 ;
    RECT 134.86 87.965 136.4 88.685 ;
    RECT 137.2 87.965 137.52 88.685 ;
    RECT 137.8 87.965 138.26 88.685 ;
    RECT 139.06 87.965 139.6 88.685 ;
    RECT 140.07 87.965 140.785 88.685 ;
    RECT 141.075 87.965 141.28 88.685 ;
    RECT 142.28 87.965 142.44 88.685 ;
    RECT 142.79 87.965 142.96 88.685 ;
    RECT 144.03 87.965 145.765 88.685 ;
    RECT 146.505 87.965 146.695 88.685 ;
    RECT 147.045 87.965 147.17 88.685 ;
    RECT 121.21 87.245 121.33 87.965 ;
    RECT 121.62 87.245 121.97 87.965 ;
    RECT 122.555 87.245 124.12 87.965 ;
    RECT 125.39 87.245 125.545 87.965 ;
    RECT 126.005 87.245 126.63 87.965 ;
    RECT 127.1 87.245 127.25 87.965 ;
    RECT 127.6 87.245 127.995 87.965 ;
    RECT 128.285 87.245 128.605 87.965 ;
    RECT 129.035 87.245 129.315 87.965 ;
    RECT 129.785 87.245 130.485 87.965 ;
    RECT 130.775 87.245 131.285 87.965 ;
    RECT 131.955 87.245 133.505 87.965 ;
    RECT 133.855 87.245 134.205 87.965 ;
    RECT 134.86 87.245 136.4 87.965 ;
    RECT 137.2 87.245 137.52 87.965 ;
    RECT 137.8 87.245 138.26 87.965 ;
    RECT 139.06 87.245 139.6 87.965 ;
    RECT 140.07 87.245 140.785 87.965 ;
    RECT 141.075 87.245 141.28 87.965 ;
    RECT 142.28 87.245 142.44 87.965 ;
    RECT 142.79 87.245 142.96 87.965 ;
    RECT 144.03 87.245 145.765 87.965 ;
    RECT 146.505 87.245 146.695 87.965 ;
    RECT 147.045 87.245 147.17 87.965 ;
    RECT 121.21 86.525 121.33 87.245 ;
    RECT 121.62 86.525 121.97 87.245 ;
    RECT 122.555 86.525 124.12 87.245 ;
    RECT 125.39 86.525 125.545 87.245 ;
    RECT 126.005 86.525 126.63 87.245 ;
    RECT 127.1 86.525 127.25 87.245 ;
    RECT 127.6 86.525 127.995 87.245 ;
    RECT 128.285 86.525 128.605 87.245 ;
    RECT 129.035 86.525 129.315 87.245 ;
    RECT 129.785 86.525 130.485 87.245 ;
    RECT 130.775 86.525 131.285 87.245 ;
    RECT 131.955 86.525 133.505 87.245 ;
    RECT 133.855 86.525 134.205 87.245 ;
    RECT 134.86 86.525 136.4 87.245 ;
    RECT 137.2 86.525 137.52 87.245 ;
    RECT 137.8 86.525 138.26 87.245 ;
    RECT 139.06 86.525 139.6 87.245 ;
    RECT 140.07 86.525 140.785 87.245 ;
    RECT 141.075 86.525 141.28 87.245 ;
    RECT 142.28 86.525 142.44 87.245 ;
    RECT 142.79 86.525 142.96 87.245 ;
    RECT 144.03 86.525 145.765 87.245 ;
    RECT 146.505 86.525 146.695 87.245 ;
    RECT 147.045 86.525 147.17 87.245 ;
    RECT 121.21 85.805 121.33 86.525 ;
    RECT 121.62 85.805 121.97 86.525 ;
    RECT 122.555 85.805 124.12 86.525 ;
    RECT 125.39 85.805 125.545 86.525 ;
    RECT 126.005 85.805 126.63 86.525 ;
    RECT 127.1 85.805 127.25 86.525 ;
    RECT 127.6 85.805 127.995 86.525 ;
    RECT 128.285 85.805 128.605 86.525 ;
    RECT 129.035 85.805 129.315 86.525 ;
    RECT 129.785 85.805 130.485 86.525 ;
    RECT 130.775 85.805 131.285 86.525 ;
    RECT 131.955 85.805 133.505 86.525 ;
    RECT 133.855 85.805 134.205 86.525 ;
    RECT 134.86 85.805 136.4 86.525 ;
    RECT 137.2 85.805 137.52 86.525 ;
    RECT 137.8 85.805 138.26 86.525 ;
    RECT 139.06 85.805 139.6 86.525 ;
    RECT 140.07 85.805 140.785 86.525 ;
    RECT 141.075 85.805 141.28 86.525 ;
    RECT 142.28 85.805 142.44 86.525 ;
    RECT 142.79 85.805 142.96 86.525 ;
    RECT 144.03 85.805 145.765 86.525 ;
    RECT 146.505 85.805 146.695 86.525 ;
    RECT 147.045 85.805 147.17 86.525 ;
    RECT 121.21 85.085 121.33 85.805 ;
    RECT 121.62 85.085 121.97 85.805 ;
    RECT 122.555 85.085 124.12 85.805 ;
    RECT 125.39 85.085 125.545 85.805 ;
    RECT 126.005 85.085 126.63 85.805 ;
    RECT 127.1 85.085 127.25 85.805 ;
    RECT 127.6 85.085 127.995 85.805 ;
    RECT 128.285 85.085 128.605 85.805 ;
    RECT 129.035 85.085 129.315 85.805 ;
    RECT 129.785 85.085 130.485 85.805 ;
    RECT 130.775 85.085 131.285 85.805 ;
    RECT 131.955 85.085 133.505 85.805 ;
    RECT 133.855 85.085 134.205 85.805 ;
    RECT 134.86 85.085 136.4 85.805 ;
    RECT 137.2 85.085 137.52 85.805 ;
    RECT 137.8 85.085 138.26 85.805 ;
    RECT 139.06 85.085 139.6 85.805 ;
    RECT 140.07 85.085 140.785 85.805 ;
    RECT 141.075 85.085 141.28 85.805 ;
    RECT 142.28 85.085 142.44 85.805 ;
    RECT 142.79 85.085 142.96 85.805 ;
    RECT 144.03 85.085 145.765 85.805 ;
    RECT 146.505 85.085 146.695 85.805 ;
    RECT 147.045 85.085 147.17 85.805 ;
    RECT 121.21 84.365 121.33 85.085 ;
    RECT 121.62 84.365 121.97 85.085 ;
    RECT 122.555 84.365 124.12 85.085 ;
    RECT 125.39 84.365 125.545 85.085 ;
    RECT 126.005 84.365 126.63 85.085 ;
    RECT 127.1 84.365 127.25 85.085 ;
    RECT 127.6 84.365 127.995 85.085 ;
    RECT 128.285 84.365 128.605 85.085 ;
    RECT 129.035 84.365 129.315 85.085 ;
    RECT 129.785 84.365 130.485 85.085 ;
    RECT 130.775 84.365 131.285 85.085 ;
    RECT 131.955 84.365 133.505 85.085 ;
    RECT 133.855 84.365 134.205 85.085 ;
    RECT 134.86 84.365 136.4 85.085 ;
    RECT 137.2 84.365 137.52 85.085 ;
    RECT 137.8 84.365 138.26 85.085 ;
    RECT 139.06 84.365 139.6 85.085 ;
    RECT 140.07 84.365 140.785 85.085 ;
    RECT 141.075 84.365 141.28 85.085 ;
    RECT 142.28 84.365 142.44 85.085 ;
    RECT 142.79 84.365 142.96 85.085 ;
    RECT 144.03 84.365 145.765 85.085 ;
    RECT 146.505 84.365 146.695 85.085 ;
    RECT 147.045 84.365 147.17 85.085 ;
    RECT 121.21 83.645 121.33 84.365 ;
    RECT 121.62 83.645 121.97 84.365 ;
    RECT 122.555 83.645 124.12 84.365 ;
    RECT 125.39 83.645 125.545 84.365 ;
    RECT 126.005 83.645 126.63 84.365 ;
    RECT 127.1 83.645 127.25 84.365 ;
    RECT 127.6 83.645 127.995 84.365 ;
    RECT 128.285 83.645 128.605 84.365 ;
    RECT 129.035 83.645 129.315 84.365 ;
    RECT 129.785 83.645 130.485 84.365 ;
    RECT 130.775 83.645 131.285 84.365 ;
    RECT 131.955 83.645 133.505 84.365 ;
    RECT 133.855 83.645 134.205 84.365 ;
    RECT 134.86 83.645 136.4 84.365 ;
    RECT 137.2 83.645 137.52 84.365 ;
    RECT 137.8 83.645 138.26 84.365 ;
    RECT 139.06 83.645 139.6 84.365 ;
    RECT 140.07 83.645 140.785 84.365 ;
    RECT 141.075 83.645 141.28 84.365 ;
    RECT 142.28 83.645 142.44 84.365 ;
    RECT 142.79 83.645 142.96 84.365 ;
    RECT 144.03 83.645 145.765 84.365 ;
    RECT 146.505 83.645 146.695 84.365 ;
    RECT 147.045 83.645 147.17 84.365 ;
    RECT 121.21 82.925 121.33 83.645 ;
    RECT 121.62 82.925 121.97 83.645 ;
    RECT 122.555 82.925 124.12 83.645 ;
    RECT 125.39 82.925 125.545 83.645 ;
    RECT 126.005 82.925 126.63 83.645 ;
    RECT 127.1 82.925 127.25 83.645 ;
    RECT 127.6 82.925 127.995 83.645 ;
    RECT 128.285 82.925 128.605 83.645 ;
    RECT 129.035 82.925 129.315 83.645 ;
    RECT 129.785 82.925 130.485 83.645 ;
    RECT 130.775 82.925 131.285 83.645 ;
    RECT 131.955 82.925 133.505 83.645 ;
    RECT 133.855 82.925 134.205 83.645 ;
    RECT 134.86 82.925 136.4 83.645 ;
    RECT 137.2 82.925 137.52 83.645 ;
    RECT 137.8 82.925 138.26 83.645 ;
    RECT 139.06 82.925 139.6 83.645 ;
    RECT 140.07 82.925 140.785 83.645 ;
    RECT 141.075 82.925 141.28 83.645 ;
    RECT 142.28 82.925 142.44 83.645 ;
    RECT 142.79 82.925 142.96 83.645 ;
    RECT 144.03 82.925 145.765 83.645 ;
    RECT 146.505 82.925 146.695 83.645 ;
    RECT 147.045 82.925 147.17 83.645 ;
    RECT 121.21 82.205 121.33 82.925 ;
    RECT 121.62 82.205 121.97 82.925 ;
    RECT 122.555 82.205 124.12 82.925 ;
    RECT 125.39 82.205 125.545 82.925 ;
    RECT 126.005 82.205 126.63 82.925 ;
    RECT 127.1 82.205 127.25 82.925 ;
    RECT 127.6 82.205 127.995 82.925 ;
    RECT 128.285 82.205 128.605 82.925 ;
    RECT 129.035 82.205 129.315 82.925 ;
    RECT 129.785 82.205 130.485 82.925 ;
    RECT 130.775 82.205 131.285 82.925 ;
    RECT 131.955 82.205 133.505 82.925 ;
    RECT 133.855 82.205 134.205 82.925 ;
    RECT 134.86 82.205 136.4 82.925 ;
    RECT 137.2 82.205 137.52 82.925 ;
    RECT 137.8 82.205 138.26 82.925 ;
    RECT 139.06 82.205 139.6 82.925 ;
    RECT 140.07 82.205 140.785 82.925 ;
    RECT 141.075 82.205 141.28 82.925 ;
    RECT 142.28 82.205 142.44 82.925 ;
    RECT 142.79 82.205 142.96 82.925 ;
    RECT 144.03 82.205 145.765 82.925 ;
    RECT 146.505 82.205 146.695 82.925 ;
    RECT 147.045 82.205 147.17 82.925 ;
    RECT 121.21 81.485 121.33 82.205 ;
    RECT 121.62 81.485 121.97 82.205 ;
    RECT 122.555 81.485 124.12 82.205 ;
    RECT 125.39 81.485 125.545 82.205 ;
    RECT 126.005 81.485 126.63 82.205 ;
    RECT 127.1 81.485 127.25 82.205 ;
    RECT 127.6 81.485 127.995 82.205 ;
    RECT 128.285 81.485 128.605 82.205 ;
    RECT 129.035 81.485 129.315 82.205 ;
    RECT 129.785 81.485 130.485 82.205 ;
    RECT 130.775 81.485 131.285 82.205 ;
    RECT 131.955 81.485 133.505 82.205 ;
    RECT 133.855 81.485 134.205 82.205 ;
    RECT 134.86 81.485 136.4 82.205 ;
    RECT 137.2 81.485 137.52 82.205 ;
    RECT 137.8 81.485 138.26 82.205 ;
    RECT 139.06 81.485 139.6 82.205 ;
    RECT 140.07 81.485 140.785 82.205 ;
    RECT 141.075 81.485 141.28 82.205 ;
    RECT 142.28 81.485 142.44 82.205 ;
    RECT 142.79 81.485 142.96 82.205 ;
    RECT 144.03 81.485 145.765 82.205 ;
    RECT 146.505 81.485 146.695 82.205 ;
    RECT 147.045 81.485 147.17 82.205 ;
    RECT 121.21 80.765 121.33 81.485 ;
    RECT 121.62 80.765 121.97 81.485 ;
    RECT 122.555 80.765 124.12 81.485 ;
    RECT 125.39 80.765 125.545 81.485 ;
    RECT 126.005 80.765 126.63 81.485 ;
    RECT 127.1 80.765 127.25 81.485 ;
    RECT 127.6 80.765 127.995 81.485 ;
    RECT 128.285 80.765 128.605 81.485 ;
    RECT 129.035 80.765 129.315 81.485 ;
    RECT 129.785 80.765 130.485 81.485 ;
    RECT 130.775 80.765 131.285 81.485 ;
    RECT 131.955 80.765 133.505 81.485 ;
    RECT 133.855 80.765 134.205 81.485 ;
    RECT 134.86 80.765 136.4 81.485 ;
    RECT 137.2 80.765 137.52 81.485 ;
    RECT 137.8 80.765 138.26 81.485 ;
    RECT 139.06 80.765 139.6 81.485 ;
    RECT 140.07 80.765 140.785 81.485 ;
    RECT 141.075 80.765 141.28 81.485 ;
    RECT 142.28 80.765 142.44 81.485 ;
    RECT 142.79 80.765 142.96 81.485 ;
    RECT 144.03 80.765 145.765 81.485 ;
    RECT 146.505 80.765 146.695 81.485 ;
    RECT 147.045 80.765 147.17 81.485 ;
    RECT 121.21 80.045 121.33 80.765 ;
    RECT 121.62 80.045 121.97 80.765 ;
    RECT 122.555 80.045 124.12 80.765 ;
    RECT 125.39 80.045 125.545 80.765 ;
    RECT 126.005 80.045 126.63 80.765 ;
    RECT 127.1 80.045 127.25 80.765 ;
    RECT 127.6 80.045 127.995 80.765 ;
    RECT 128.285 80.045 128.605 80.765 ;
    RECT 129.035 80.045 129.315 80.765 ;
    RECT 129.785 80.045 130.485 80.765 ;
    RECT 130.775 80.045 131.285 80.765 ;
    RECT 131.955 80.045 133.505 80.765 ;
    RECT 133.855 80.045 134.205 80.765 ;
    RECT 134.86 80.045 136.4 80.765 ;
    RECT 137.2 80.045 137.52 80.765 ;
    RECT 137.8 80.045 138.26 80.765 ;
    RECT 139.06 80.045 139.6 80.765 ;
    RECT 140.07 80.045 140.785 80.765 ;
    RECT 141.075 80.045 141.28 80.765 ;
    RECT 142.28 80.045 142.44 80.765 ;
    RECT 142.79 80.045 142.96 80.765 ;
    RECT 144.03 80.045 145.765 80.765 ;
    RECT 146.505 80.045 146.695 80.765 ;
    RECT 147.045 80.045 147.17 80.765 ;
    RECT 121.21 79.325 121.33 80.045 ;
    RECT 121.62 79.325 121.97 80.045 ;
    RECT 122.555 79.325 124.12 80.045 ;
    RECT 125.39 79.325 125.545 80.045 ;
    RECT 126.005 79.325 126.63 80.045 ;
    RECT 127.1 79.325 127.25 80.045 ;
    RECT 127.6 79.325 127.995 80.045 ;
    RECT 128.285 79.325 128.605 80.045 ;
    RECT 129.035 79.325 129.315 80.045 ;
    RECT 129.785 79.325 130.485 80.045 ;
    RECT 130.775 79.325 131.285 80.045 ;
    RECT 131.955 79.325 133.505 80.045 ;
    RECT 133.855 79.325 134.205 80.045 ;
    RECT 134.86 79.325 136.4 80.045 ;
    RECT 137.2 79.325 137.52 80.045 ;
    RECT 137.8 79.325 138.26 80.045 ;
    RECT 139.06 79.325 139.6 80.045 ;
    RECT 140.07 79.325 140.785 80.045 ;
    RECT 141.075 79.325 141.28 80.045 ;
    RECT 142.28 79.325 142.44 80.045 ;
    RECT 142.79 79.325 142.96 80.045 ;
    RECT 144.03 79.325 145.765 80.045 ;
    RECT 146.505 79.325 146.695 80.045 ;
    RECT 147.045 79.325 147.17 80.045 ;
    RECT 121.21 78.605 121.33 79.325 ;
    RECT 121.62 78.605 121.97 79.325 ;
    RECT 122.555 78.605 124.12 79.325 ;
    RECT 125.39 78.605 125.545 79.325 ;
    RECT 126.005 78.605 126.63 79.325 ;
    RECT 127.1 78.605 127.25 79.325 ;
    RECT 127.6 78.605 127.995 79.325 ;
    RECT 128.285 78.605 128.605 79.325 ;
    RECT 129.035 78.605 129.315 79.325 ;
    RECT 129.785 78.605 130.485 79.325 ;
    RECT 130.775 78.605 131.285 79.325 ;
    RECT 131.955 78.605 133.505 79.325 ;
    RECT 133.855 78.605 134.205 79.325 ;
    RECT 134.86 78.605 136.4 79.325 ;
    RECT 137.2 78.605 137.52 79.325 ;
    RECT 137.8 78.605 138.26 79.325 ;
    RECT 139.06 78.605 139.6 79.325 ;
    RECT 140.07 78.605 140.785 79.325 ;
    RECT 141.075 78.605 141.28 79.325 ;
    RECT 142.28 78.605 142.44 79.325 ;
    RECT 142.79 78.605 142.96 79.325 ;
    RECT 144.03 78.605 145.765 79.325 ;
    RECT 146.505 78.605 146.695 79.325 ;
    RECT 147.045 78.605 147.17 79.325 ;
    RECT 121.21 77.885 121.33 78.605 ;
    RECT 121.62 77.885 121.97 78.605 ;
    RECT 122.555 77.885 124.12 78.605 ;
    RECT 125.39 77.885 125.545 78.605 ;
    RECT 126.005 77.885 126.63 78.605 ;
    RECT 127.1 77.885 127.25 78.605 ;
    RECT 127.6 77.885 127.995 78.605 ;
    RECT 128.285 77.885 128.605 78.605 ;
    RECT 129.035 77.885 129.315 78.605 ;
    RECT 129.785 77.885 130.485 78.605 ;
    RECT 130.775 77.885 131.285 78.605 ;
    RECT 131.955 77.885 133.505 78.605 ;
    RECT 133.855 77.885 134.205 78.605 ;
    RECT 134.86 77.885 136.4 78.605 ;
    RECT 137.2 77.885 137.52 78.605 ;
    RECT 137.8 77.885 138.26 78.605 ;
    RECT 139.06 77.885 139.6 78.605 ;
    RECT 140.07 77.885 140.785 78.605 ;
    RECT 141.075 77.885 141.28 78.605 ;
    RECT 142.28 77.885 142.44 78.605 ;
    RECT 142.79 77.885 142.96 78.605 ;
    RECT 144.03 77.885 145.765 78.605 ;
    RECT 146.505 77.885 146.695 78.605 ;
    RECT 147.045 77.885 147.17 78.605 ;
    RECT 121.21 77.165 121.33 77.885 ;
    RECT 121.62 77.165 121.97 77.885 ;
    RECT 122.555 77.165 124.12 77.885 ;
    RECT 125.39 77.165 125.545 77.885 ;
    RECT 126.005 77.165 126.63 77.885 ;
    RECT 127.1 77.165 127.25 77.885 ;
    RECT 127.6 77.165 127.995 77.885 ;
    RECT 128.285 77.165 128.605 77.885 ;
    RECT 129.035 77.165 129.315 77.885 ;
    RECT 129.785 77.165 130.485 77.885 ;
    RECT 130.775 77.165 131.285 77.885 ;
    RECT 131.955 77.165 133.505 77.885 ;
    RECT 133.855 77.165 134.205 77.885 ;
    RECT 134.86 77.165 136.4 77.885 ;
    RECT 137.2 77.165 137.52 77.885 ;
    RECT 137.8 77.165 138.26 77.885 ;
    RECT 139.06 77.165 139.6 77.885 ;
    RECT 140.07 77.165 140.785 77.885 ;
    RECT 141.075 77.165 141.28 77.885 ;
    RECT 142.28 77.165 142.44 77.885 ;
    RECT 142.79 77.165 142.96 77.885 ;
    RECT 144.03 77.165 145.765 77.885 ;
    RECT 146.505 77.165 146.695 77.885 ;
    RECT 147.045 77.165 147.17 77.885 ;
    RECT 121.21 76.445 121.33 77.165 ;
    RECT 121.62 76.445 121.97 77.165 ;
    RECT 122.555 76.445 124.12 77.165 ;
    RECT 125.39 76.445 125.545 77.165 ;
    RECT 126.005 76.445 126.63 77.165 ;
    RECT 127.1 76.445 127.25 77.165 ;
    RECT 127.6 76.445 127.995 77.165 ;
    RECT 128.285 76.445 128.605 77.165 ;
    RECT 129.035 76.445 129.315 77.165 ;
    RECT 129.785 76.445 130.485 77.165 ;
    RECT 130.775 76.445 131.285 77.165 ;
    RECT 131.955 76.445 133.505 77.165 ;
    RECT 133.855 76.445 134.205 77.165 ;
    RECT 134.86 76.445 136.4 77.165 ;
    RECT 137.2 76.445 137.52 77.165 ;
    RECT 137.8 76.445 138.26 77.165 ;
    RECT 139.06 76.445 139.6 77.165 ;
    RECT 140.07 76.445 140.785 77.165 ;
    RECT 141.075 76.445 141.28 77.165 ;
    RECT 142.28 76.445 142.44 77.165 ;
    RECT 142.79 76.445 142.96 77.165 ;
    RECT 144.03 76.445 145.765 77.165 ;
    RECT 146.505 76.445 146.695 77.165 ;
    RECT 147.045 76.445 147.17 77.165 ;
    RECT 121.21 75.725 121.33 76.445 ;
    RECT 121.62 75.725 121.97 76.445 ;
    RECT 122.555 75.725 124.12 76.445 ;
    RECT 125.39 75.725 125.545 76.445 ;
    RECT 126.005 75.725 126.63 76.445 ;
    RECT 127.1 75.725 127.25 76.445 ;
    RECT 127.6 75.725 127.995 76.445 ;
    RECT 128.285 75.725 128.605 76.445 ;
    RECT 129.035 75.725 129.315 76.445 ;
    RECT 129.785 75.725 130.485 76.445 ;
    RECT 130.775 75.725 131.285 76.445 ;
    RECT 131.955 75.725 133.505 76.445 ;
    RECT 133.855 75.725 134.205 76.445 ;
    RECT 134.86 75.725 136.4 76.445 ;
    RECT 137.2 75.725 137.52 76.445 ;
    RECT 137.8 75.725 138.26 76.445 ;
    RECT 139.06 75.725 139.6 76.445 ;
    RECT 140.07 75.725 140.785 76.445 ;
    RECT 141.075 75.725 141.28 76.445 ;
    RECT 142.28 75.725 142.44 76.445 ;
    RECT 142.79 75.725 142.96 76.445 ;
    RECT 144.03 75.725 145.765 76.445 ;
    RECT 146.505 75.725 146.695 76.445 ;
    RECT 147.045 75.725 147.17 76.445 ;
    RECT 121.21 75.005 121.33 75.725 ;
    RECT 121.62 75.005 121.97 75.725 ;
    RECT 122.555 75.005 124.12 75.725 ;
    RECT 125.39 75.005 125.545 75.725 ;
    RECT 126.005 75.005 126.63 75.725 ;
    RECT 127.1 75.005 127.25 75.725 ;
    RECT 127.6 75.005 127.995 75.725 ;
    RECT 128.285 75.005 128.605 75.725 ;
    RECT 129.035 75.005 129.315 75.725 ;
    RECT 129.785 75.005 130.485 75.725 ;
    RECT 130.775 75.005 131.285 75.725 ;
    RECT 131.955 75.005 133.505 75.725 ;
    RECT 133.855 75.005 134.205 75.725 ;
    RECT 134.86 75.005 136.4 75.725 ;
    RECT 137.2 75.005 137.52 75.725 ;
    RECT 137.8 75.005 138.26 75.725 ;
    RECT 139.06 75.005 139.6 75.725 ;
    RECT 140.07 75.005 140.785 75.725 ;
    RECT 141.075 75.005 141.28 75.725 ;
    RECT 142.28 75.005 142.44 75.725 ;
    RECT 142.79 75.005 142.96 75.725 ;
    RECT 144.03 75.005 145.765 75.725 ;
    RECT 146.505 75.005 146.695 75.725 ;
    RECT 147.045 75.005 147.17 75.725 ;
    RECT 121.21 74.285 121.33 75.005 ;
    RECT 121.62 74.285 121.97 75.005 ;
    RECT 122.555 74.285 124.12 75.005 ;
    RECT 125.39 74.285 125.545 75.005 ;
    RECT 126.005 74.285 126.63 75.005 ;
    RECT 127.1 74.285 127.25 75.005 ;
    RECT 127.6 74.285 127.995 75.005 ;
    RECT 128.285 74.285 128.605 75.005 ;
    RECT 129.035 74.285 129.315 75.005 ;
    RECT 129.785 74.285 130.485 75.005 ;
    RECT 130.775 74.285 131.285 75.005 ;
    RECT 131.955 74.285 133.505 75.005 ;
    RECT 133.855 74.285 134.205 75.005 ;
    RECT 134.86 74.285 136.4 75.005 ;
    RECT 137.2 74.285 137.52 75.005 ;
    RECT 137.8 74.285 138.26 75.005 ;
    RECT 139.06 74.285 139.6 75.005 ;
    RECT 140.07 74.285 140.785 75.005 ;
    RECT 141.075 74.285 141.28 75.005 ;
    RECT 142.28 74.285 142.44 75.005 ;
    RECT 142.79 74.285 142.96 75.005 ;
    RECT 144.03 74.285 145.765 75.005 ;
    RECT 146.505 74.285 146.695 75.005 ;
    RECT 147.045 74.285 147.17 75.005 ;
    RECT 121.21 73.565 121.33 74.285 ;
    RECT 121.62 73.565 121.97 74.285 ;
    RECT 122.555 73.565 124.12 74.285 ;
    RECT 125.39 73.565 125.545 74.285 ;
    RECT 126.005 73.565 126.63 74.285 ;
    RECT 127.1 73.565 127.25 74.285 ;
    RECT 127.6 73.565 127.995 74.285 ;
    RECT 128.285 73.565 128.605 74.285 ;
    RECT 129.035 73.565 129.315 74.285 ;
    RECT 129.785 73.565 130.485 74.285 ;
    RECT 130.775 73.565 131.285 74.285 ;
    RECT 131.955 73.565 133.505 74.285 ;
    RECT 133.855 73.565 134.205 74.285 ;
    RECT 134.86 73.565 136.4 74.285 ;
    RECT 137.2 73.565 137.52 74.285 ;
    RECT 137.8 73.565 138.26 74.285 ;
    RECT 139.06 73.565 139.6 74.285 ;
    RECT 140.07 73.565 140.785 74.285 ;
    RECT 141.075 73.565 141.28 74.285 ;
    RECT 142.28 73.565 142.44 74.285 ;
    RECT 142.79 73.565 142.96 74.285 ;
    RECT 144.03 73.565 145.765 74.285 ;
    RECT 146.505 73.565 146.695 74.285 ;
    RECT 147.045 73.565 147.17 74.285 ;
    RECT 121.21 72.845 121.33 73.565 ;
    RECT 121.62 72.845 121.97 73.565 ;
    RECT 122.555 72.845 124.12 73.565 ;
    RECT 125.39 72.845 125.545 73.565 ;
    RECT 126.005 72.845 126.63 73.565 ;
    RECT 127.1 72.845 127.25 73.565 ;
    RECT 127.6 72.845 127.995 73.565 ;
    RECT 128.285 72.845 128.605 73.565 ;
    RECT 129.035 72.845 129.315 73.565 ;
    RECT 129.785 72.845 130.485 73.565 ;
    RECT 130.775 72.845 131.285 73.565 ;
    RECT 131.955 72.845 133.505 73.565 ;
    RECT 133.855 72.845 134.205 73.565 ;
    RECT 134.86 72.845 136.4 73.565 ;
    RECT 137.2 72.845 137.52 73.565 ;
    RECT 137.8 72.845 138.26 73.565 ;
    RECT 139.06 72.845 139.6 73.565 ;
    RECT 140.07 72.845 140.785 73.565 ;
    RECT 141.075 72.845 141.28 73.565 ;
    RECT 142.28 72.845 142.44 73.565 ;
    RECT 142.79 72.845 142.96 73.565 ;
    RECT 144.03 72.845 145.765 73.565 ;
    RECT 146.505 72.845 146.695 73.565 ;
    RECT 147.045 72.845 147.17 73.565 ;
    RECT 121.21 72.125 121.33 72.845 ;
    RECT 121.62 72.125 121.97 72.845 ;
    RECT 122.555 72.125 124.12 72.845 ;
    RECT 125.39 72.125 125.545 72.845 ;
    RECT 126.005 72.125 126.63 72.845 ;
    RECT 127.1 72.125 127.25 72.845 ;
    RECT 127.6 72.125 127.995 72.845 ;
    RECT 128.285 72.125 128.605 72.845 ;
    RECT 129.035 72.125 129.315 72.845 ;
    RECT 129.785 72.125 130.485 72.845 ;
    RECT 130.775 72.125 131.285 72.845 ;
    RECT 131.955 72.125 133.505 72.845 ;
    RECT 133.855 72.125 134.205 72.845 ;
    RECT 134.86 72.125 136.4 72.845 ;
    RECT 137.2 72.125 137.52 72.845 ;
    RECT 137.8 72.125 138.26 72.845 ;
    RECT 139.06 72.125 139.6 72.845 ;
    RECT 140.07 72.125 140.785 72.845 ;
    RECT 141.075 72.125 141.28 72.845 ;
    RECT 142.28 72.125 142.44 72.845 ;
    RECT 142.79 72.125 142.96 72.845 ;
    RECT 144.03 72.125 145.765 72.845 ;
    RECT 146.505 72.125 146.695 72.845 ;
    RECT 147.045 72.125 147.17 72.845 ;
    RECT 121.21 71.405 121.33 72.125 ;
    RECT 121.62 71.405 121.97 72.125 ;
    RECT 122.555 71.405 124.12 72.125 ;
    RECT 125.39 71.405 125.545 72.125 ;
    RECT 126.005 71.405 126.63 72.125 ;
    RECT 127.1 71.405 127.25 72.125 ;
    RECT 127.6 71.405 127.995 72.125 ;
    RECT 128.285 71.405 128.605 72.125 ;
    RECT 129.035 71.405 129.315 72.125 ;
    RECT 129.785 71.405 130.485 72.125 ;
    RECT 130.775 71.405 131.285 72.125 ;
    RECT 131.955 71.405 133.505 72.125 ;
    RECT 133.855 71.405 134.205 72.125 ;
    RECT 134.86 71.405 136.4 72.125 ;
    RECT 137.2 71.405 137.52 72.125 ;
    RECT 137.8 71.405 138.26 72.125 ;
    RECT 139.06 71.405 139.6 72.125 ;
    RECT 140.07 71.405 140.785 72.125 ;
    RECT 141.075 71.405 141.28 72.125 ;
    RECT 142.28 71.405 142.44 72.125 ;
    RECT 142.79 71.405 142.96 72.125 ;
    RECT 144.03 71.405 145.765 72.125 ;
    RECT 146.505 71.405 146.695 72.125 ;
    RECT 147.045 71.405 147.17 72.125 ;
    RECT 121.21 70.685 121.33 71.405 ;
    RECT 121.62 70.685 121.97 71.405 ;
    RECT 122.555 70.685 124.12 71.405 ;
    RECT 125.39 70.685 125.545 71.405 ;
    RECT 126.005 70.685 126.63 71.405 ;
    RECT 127.1 70.685 127.25 71.405 ;
    RECT 127.6 70.685 127.995 71.405 ;
    RECT 128.285 70.685 128.605 71.405 ;
    RECT 129.035 70.685 129.315 71.405 ;
    RECT 129.785 70.685 130.485 71.405 ;
    RECT 130.775 70.685 131.285 71.405 ;
    RECT 131.955 70.685 133.505 71.405 ;
    RECT 133.855 70.685 134.205 71.405 ;
    RECT 134.86 70.685 136.4 71.405 ;
    RECT 137.2 70.685 137.52 71.405 ;
    RECT 137.8 70.685 138.26 71.405 ;
    RECT 139.06 70.685 139.6 71.405 ;
    RECT 140.07 70.685 140.785 71.405 ;
    RECT 141.075 70.685 141.28 71.405 ;
    RECT 142.28 70.685 142.44 71.405 ;
    RECT 142.79 70.685 142.96 71.405 ;
    RECT 144.03 70.685 145.765 71.405 ;
    RECT 146.505 70.685 146.695 71.405 ;
    RECT 147.045 70.685 147.17 71.405 ;
    RECT 121.21 69.965 121.33 70.685 ;
    RECT 121.62 69.965 121.97 70.685 ;
    RECT 122.555 69.965 124.12 70.685 ;
    RECT 125.39 69.965 125.545 70.685 ;
    RECT 126.005 69.965 126.63 70.685 ;
    RECT 127.1 69.965 127.25 70.685 ;
    RECT 127.6 69.965 127.995 70.685 ;
    RECT 128.285 69.965 128.605 70.685 ;
    RECT 129.035 69.965 129.315 70.685 ;
    RECT 129.785 69.965 130.485 70.685 ;
    RECT 130.775 69.965 131.285 70.685 ;
    RECT 131.955 69.965 133.505 70.685 ;
    RECT 133.855 69.965 134.205 70.685 ;
    RECT 134.86 69.965 136.4 70.685 ;
    RECT 137.2 69.965 137.52 70.685 ;
    RECT 137.8 69.965 138.26 70.685 ;
    RECT 139.06 69.965 139.6 70.685 ;
    RECT 140.07 69.965 140.785 70.685 ;
    RECT 141.075 69.965 141.28 70.685 ;
    RECT 142.28 69.965 142.44 70.685 ;
    RECT 142.79 69.965 142.96 70.685 ;
    RECT 144.03 69.965 145.765 70.685 ;
    RECT 146.505 69.965 146.695 70.685 ;
    RECT 147.045 69.965 147.17 70.685 ;
    RECT 121.21 69.245 121.33 69.965 ;
    RECT 121.62 69.245 121.97 69.965 ;
    RECT 122.555 69.245 124.12 69.965 ;
    RECT 125.39 69.245 125.545 69.965 ;
    RECT 126.005 69.245 126.63 69.965 ;
    RECT 127.1 69.245 127.25 69.965 ;
    RECT 127.6 69.245 127.995 69.965 ;
    RECT 128.285 69.245 128.605 69.965 ;
    RECT 129.035 69.245 129.315 69.965 ;
    RECT 129.785 69.245 130.485 69.965 ;
    RECT 130.775 69.245 131.285 69.965 ;
    RECT 131.955 69.245 133.505 69.965 ;
    RECT 133.855 69.245 134.205 69.965 ;
    RECT 134.86 69.245 136.4 69.965 ;
    RECT 137.2 69.245 137.52 69.965 ;
    RECT 137.8 69.245 138.26 69.965 ;
    RECT 139.06 69.245 139.6 69.965 ;
    RECT 140.07 69.245 140.785 69.965 ;
    RECT 141.075 69.245 141.28 69.965 ;
    RECT 142.28 69.245 142.44 69.965 ;
    RECT 142.79 69.245 142.96 69.965 ;
    RECT 144.03 69.245 145.765 69.965 ;
    RECT 146.505 69.245 146.695 69.965 ;
    RECT 147.045 69.245 147.17 69.965 ;
    RECT 121.21 68.525 121.33 69.245 ;
    RECT 121.62 68.525 121.97 69.245 ;
    RECT 122.555 68.525 124.12 69.245 ;
    RECT 125.39 68.525 125.545 69.245 ;
    RECT 126.005 68.525 126.63 69.245 ;
    RECT 127.1 68.525 127.25 69.245 ;
    RECT 127.6 68.525 127.995 69.245 ;
    RECT 128.285 68.525 128.605 69.245 ;
    RECT 129.035 68.525 129.315 69.245 ;
    RECT 129.785 68.525 130.485 69.245 ;
    RECT 130.775 68.525 131.285 69.245 ;
    RECT 131.955 68.525 133.505 69.245 ;
    RECT 133.855 68.525 134.205 69.245 ;
    RECT 134.86 68.525 136.4 69.245 ;
    RECT 137.2 68.525 137.52 69.245 ;
    RECT 137.8 68.525 138.26 69.245 ;
    RECT 139.06 68.525 139.6 69.245 ;
    RECT 140.07 68.525 140.785 69.245 ;
    RECT 141.075 68.525 141.28 69.245 ;
    RECT 142.28 68.525 142.44 69.245 ;
    RECT 142.79 68.525 142.96 69.245 ;
    RECT 144.03 68.525 145.765 69.245 ;
    RECT 146.505 68.525 146.695 69.245 ;
    RECT 147.045 68.525 147.17 69.245 ;
    RECT 121.21 67.805 121.33 68.525 ;
    RECT 121.62 67.805 121.97 68.525 ;
    RECT 122.555 67.805 124.12 68.525 ;
    RECT 125.39 67.805 125.545 68.525 ;
    RECT 126.005 67.805 126.63 68.525 ;
    RECT 127.1 67.805 127.25 68.525 ;
    RECT 127.6 67.805 127.995 68.525 ;
    RECT 128.285 67.805 128.605 68.525 ;
    RECT 129.035 67.805 129.315 68.525 ;
    RECT 129.785 67.805 130.485 68.525 ;
    RECT 130.775 67.805 131.285 68.525 ;
    RECT 131.955 67.805 133.505 68.525 ;
    RECT 133.855 67.805 134.205 68.525 ;
    RECT 134.86 67.805 136.4 68.525 ;
    RECT 137.2 67.805 137.52 68.525 ;
    RECT 137.8 67.805 138.26 68.525 ;
    RECT 139.06 67.805 139.6 68.525 ;
    RECT 140.07 67.805 140.785 68.525 ;
    RECT 141.075 67.805 141.28 68.525 ;
    RECT 142.28 67.805 142.44 68.525 ;
    RECT 142.79 67.805 142.96 68.525 ;
    RECT 144.03 67.805 145.765 68.525 ;
    RECT 146.505 67.805 146.695 68.525 ;
    RECT 147.045 67.805 147.17 68.525 ;
    RECT 121.21 67.085 121.33 67.805 ;
    RECT 121.62 67.085 121.97 67.805 ;
    RECT 122.555 67.085 124.12 67.805 ;
    RECT 125.39 67.085 125.545 67.805 ;
    RECT 126.005 67.085 126.63 67.805 ;
    RECT 127.1 67.085 127.25 67.805 ;
    RECT 127.6 67.085 127.995 67.805 ;
    RECT 128.285 67.085 128.605 67.805 ;
    RECT 129.035 67.085 129.315 67.805 ;
    RECT 129.785 67.085 130.485 67.805 ;
    RECT 130.775 67.085 131.285 67.805 ;
    RECT 131.955 67.085 133.505 67.805 ;
    RECT 133.855 67.085 134.205 67.805 ;
    RECT 134.86 67.085 136.4 67.805 ;
    RECT 137.2 67.085 137.52 67.805 ;
    RECT 137.8 67.085 138.26 67.805 ;
    RECT 139.06 67.085 139.6 67.805 ;
    RECT 140.07 67.085 140.785 67.805 ;
    RECT 141.075 67.085 141.28 67.805 ;
    RECT 142.28 67.085 142.44 67.805 ;
    RECT 142.79 67.085 142.96 67.805 ;
    RECT 144.03 67.085 145.765 67.805 ;
    RECT 146.505 67.085 146.695 67.805 ;
    RECT 147.045 67.085 147.17 67.805 ;
    RECT 121.21 66.365 121.33 67.085 ;
    RECT 121.62 66.365 121.97 67.085 ;
    RECT 122.555 66.365 124.12 67.085 ;
    RECT 125.39 66.365 125.545 67.085 ;
    RECT 126.005 66.365 126.63 67.085 ;
    RECT 127.1 66.365 127.25 67.085 ;
    RECT 127.6 66.365 127.995 67.085 ;
    RECT 128.285 66.365 128.605 67.085 ;
    RECT 129.035 66.365 129.315 67.085 ;
    RECT 129.785 66.365 130.485 67.085 ;
    RECT 130.775 66.365 131.285 67.085 ;
    RECT 131.955 66.365 133.505 67.085 ;
    RECT 133.855 66.365 134.205 67.085 ;
    RECT 134.86 66.365 136.4 67.085 ;
    RECT 137.2 66.365 137.52 67.085 ;
    RECT 137.8 66.365 138.26 67.085 ;
    RECT 139.06 66.365 139.6 67.085 ;
    RECT 140.07 66.365 140.785 67.085 ;
    RECT 141.075 66.365 141.28 67.085 ;
    RECT 142.28 66.365 142.44 67.085 ;
    RECT 142.79 66.365 142.96 67.085 ;
    RECT 144.03 66.365 145.765 67.085 ;
    RECT 146.505 66.365 146.695 67.085 ;
    RECT 147.045 66.365 147.17 67.085 ;
    RECT 121.21 65.645 121.33 66.365 ;
    RECT 121.62 65.645 121.97 66.365 ;
    RECT 122.555 65.645 124.12 66.365 ;
    RECT 125.39 65.645 125.545 66.365 ;
    RECT 126.005 65.645 126.63 66.365 ;
    RECT 127.1 65.645 127.25 66.365 ;
    RECT 127.6 65.645 127.995 66.365 ;
    RECT 128.285 65.645 128.605 66.365 ;
    RECT 129.035 65.645 129.315 66.365 ;
    RECT 129.785 65.645 130.485 66.365 ;
    RECT 130.775 65.645 131.285 66.365 ;
    RECT 131.955 65.645 133.505 66.365 ;
    RECT 133.855 65.645 134.205 66.365 ;
    RECT 134.86 65.645 136.4 66.365 ;
    RECT 137.2 65.645 137.52 66.365 ;
    RECT 137.8 65.645 138.26 66.365 ;
    RECT 139.06 65.645 139.6 66.365 ;
    RECT 140.07 65.645 140.785 66.365 ;
    RECT 141.075 65.645 141.28 66.365 ;
    RECT 142.28 65.645 142.44 66.365 ;
    RECT 142.79 65.645 142.96 66.365 ;
    RECT 144.03 65.645 145.765 66.365 ;
    RECT 146.505 65.645 146.695 66.365 ;
    RECT 147.045 65.645 147.17 66.365 ;
    RECT 121.21 64.925 121.33 65.645 ;
    RECT 121.62 64.925 121.97 65.645 ;
    RECT 122.555 64.925 124.12 65.645 ;
    RECT 125.39 64.925 125.545 65.645 ;
    RECT 126.005 64.925 126.63 65.645 ;
    RECT 127.1 64.925 127.25 65.645 ;
    RECT 127.6 64.925 127.995 65.645 ;
    RECT 128.285 64.925 128.605 65.645 ;
    RECT 129.035 64.925 129.315 65.645 ;
    RECT 129.785 64.925 130.485 65.645 ;
    RECT 130.775 64.925 131.285 65.645 ;
    RECT 131.955 64.925 133.505 65.645 ;
    RECT 133.855 64.925 134.205 65.645 ;
    RECT 134.86 64.925 136.4 65.645 ;
    RECT 137.2 64.925 137.52 65.645 ;
    RECT 137.8 64.925 138.26 65.645 ;
    RECT 139.06 64.925 139.6 65.645 ;
    RECT 140.07 64.925 140.785 65.645 ;
    RECT 141.075 64.925 141.28 65.645 ;
    RECT 142.28 64.925 142.44 65.645 ;
    RECT 142.79 64.925 142.96 65.645 ;
    RECT 144.03 64.925 145.765 65.645 ;
    RECT 146.505 64.925 146.695 65.645 ;
    RECT 147.045 64.925 147.17 65.645 ;
    RECT 121.21 64.205 121.33 64.925 ;
    RECT 121.62 64.205 121.97 64.925 ;
    RECT 122.555 64.205 124.12 64.925 ;
    RECT 125.39 64.205 125.545 64.925 ;
    RECT 126.005 64.205 126.63 64.925 ;
    RECT 127.1 64.205 127.25 64.925 ;
    RECT 127.6 64.205 127.995 64.925 ;
    RECT 128.285 64.205 128.605 64.925 ;
    RECT 129.035 64.205 129.315 64.925 ;
    RECT 129.785 64.205 130.485 64.925 ;
    RECT 130.775 64.205 131.285 64.925 ;
    RECT 131.955 64.205 133.505 64.925 ;
    RECT 133.855 64.205 134.205 64.925 ;
    RECT 134.86 64.205 136.4 64.925 ;
    RECT 137.2 64.205 137.52 64.925 ;
    RECT 137.8 64.205 138.26 64.925 ;
    RECT 139.06 64.205 139.6 64.925 ;
    RECT 140.07 64.205 140.785 64.925 ;
    RECT 141.075 64.205 141.28 64.925 ;
    RECT 142.28 64.205 142.44 64.925 ;
    RECT 142.79 64.205 142.96 64.925 ;
    RECT 144.03 64.205 145.765 64.925 ;
    RECT 146.505 64.205 146.695 64.925 ;
    RECT 147.045 64.205 147.17 64.925 ;
    RECT 121.21 63.485 121.33 64.205 ;
    RECT 121.62 63.485 121.97 64.205 ;
    RECT 122.555 63.485 124.12 64.205 ;
    RECT 125.39 63.485 125.545 64.205 ;
    RECT 126.005 63.485 126.63 64.205 ;
    RECT 127.1 63.485 127.25 64.205 ;
    RECT 127.6 63.485 127.995 64.205 ;
    RECT 128.285 63.485 128.605 64.205 ;
    RECT 129.035 63.485 129.315 64.205 ;
    RECT 129.785 63.485 130.485 64.205 ;
    RECT 130.775 63.485 131.285 64.205 ;
    RECT 131.955 63.485 133.505 64.205 ;
    RECT 133.855 63.485 134.205 64.205 ;
    RECT 134.86 63.485 136.4 64.205 ;
    RECT 137.2 63.485 137.52 64.205 ;
    RECT 137.8 63.485 138.26 64.205 ;
    RECT 139.06 63.485 139.6 64.205 ;
    RECT 140.07 63.485 140.785 64.205 ;
    RECT 141.075 63.485 141.28 64.205 ;
    RECT 142.28 63.485 142.44 64.205 ;
    RECT 142.79 63.485 142.96 64.205 ;
    RECT 144.03 63.485 145.765 64.205 ;
    RECT 146.505 63.485 146.695 64.205 ;
    RECT 147.045 63.485 147.17 64.205 ;
    RECT 121.21 62.765 121.33 63.485 ;
    RECT 121.62 62.765 121.97 63.485 ;
    RECT 122.555 62.765 124.12 63.485 ;
    RECT 125.39 62.765 125.545 63.485 ;
    RECT 126.005 62.765 126.63 63.485 ;
    RECT 127.1 62.765 127.25 63.485 ;
    RECT 127.6 62.765 127.995 63.485 ;
    RECT 128.285 62.765 128.605 63.485 ;
    RECT 129.035 62.765 129.315 63.485 ;
    RECT 129.785 62.765 130.485 63.485 ;
    RECT 130.775 62.765 131.285 63.485 ;
    RECT 131.955 62.765 133.505 63.485 ;
    RECT 133.855 62.765 134.205 63.485 ;
    RECT 134.86 62.765 136.4 63.485 ;
    RECT 137.2 62.765 137.52 63.485 ;
    RECT 137.8 62.765 138.26 63.485 ;
    RECT 139.06 62.765 139.6 63.485 ;
    RECT 140.07 62.765 140.785 63.485 ;
    RECT 141.075 62.765 141.28 63.485 ;
    RECT 142.28 62.765 142.44 63.485 ;
    RECT 142.79 62.765 142.96 63.485 ;
    RECT 144.03 62.765 145.765 63.485 ;
    RECT 146.505 62.765 146.695 63.485 ;
    RECT 147.045 62.765 147.17 63.485 ;
    RECT 121.21 62.045 121.33 62.765 ;
    RECT 121.62 62.045 121.97 62.765 ;
    RECT 122.555 62.045 124.12 62.765 ;
    RECT 125.39 62.045 125.545 62.765 ;
    RECT 126.005 62.045 126.63 62.765 ;
    RECT 127.1 62.045 127.25 62.765 ;
    RECT 127.6 62.045 127.995 62.765 ;
    RECT 128.285 62.045 128.605 62.765 ;
    RECT 129.035 62.045 129.315 62.765 ;
    RECT 129.785 62.045 130.485 62.765 ;
    RECT 130.775 62.045 131.285 62.765 ;
    RECT 131.955 62.045 133.505 62.765 ;
    RECT 133.855 62.045 134.205 62.765 ;
    RECT 134.86 62.045 136.4 62.765 ;
    RECT 137.2 62.045 137.52 62.765 ;
    RECT 137.8 62.045 138.26 62.765 ;
    RECT 139.06 62.045 139.6 62.765 ;
    RECT 140.07 62.045 140.785 62.765 ;
    RECT 141.075 62.045 141.28 62.765 ;
    RECT 142.28 62.045 142.44 62.765 ;
    RECT 142.79 62.045 142.96 62.765 ;
    RECT 144.03 62.045 145.765 62.765 ;
    RECT 146.505 62.045 146.695 62.765 ;
    RECT 147.045 62.045 147.17 62.765 ;
    RECT 121.21 61.325 121.33 62.045 ;
    RECT 121.62 61.325 121.97 62.045 ;
    RECT 122.555 61.325 124.12 62.045 ;
    RECT 125.39 61.325 125.545 62.045 ;
    RECT 126.005 61.325 126.63 62.045 ;
    RECT 127.1 61.325 127.25 62.045 ;
    RECT 127.6 61.325 127.995 62.045 ;
    RECT 128.285 61.325 128.605 62.045 ;
    RECT 129.035 61.325 129.315 62.045 ;
    RECT 129.785 61.325 130.485 62.045 ;
    RECT 130.775 61.325 131.285 62.045 ;
    RECT 131.955 61.325 133.505 62.045 ;
    RECT 133.855 61.325 134.205 62.045 ;
    RECT 134.86 61.325 136.4 62.045 ;
    RECT 137.2 61.325 137.52 62.045 ;
    RECT 137.8 61.325 138.26 62.045 ;
    RECT 139.06 61.325 139.6 62.045 ;
    RECT 140.07 61.325 140.785 62.045 ;
    RECT 141.075 61.325 141.28 62.045 ;
    RECT 142.28 61.325 142.44 62.045 ;
    RECT 142.79 61.325 142.96 62.045 ;
    RECT 144.03 61.325 145.765 62.045 ;
    RECT 146.505 61.325 146.695 62.045 ;
    RECT 147.045 61.325 147.17 62.045 ;
    RECT 121.21 59.865 121.33 60.585 ;
    RECT 121.62 59.865 121.97 60.585 ;
    RECT 122.555 59.865 124.12 60.585 ;
    RECT 125.39 59.865 125.545 60.585 ;
    RECT 126.005 59.865 126.63 60.585 ;
    RECT 127.1 59.865 127.25 60.585 ;
    RECT 127.6 59.865 127.995 60.585 ;
    RECT 128.285 59.865 128.605 60.585 ;
    RECT 129.035 59.865 129.315 60.585 ;
    RECT 129.785 59.865 130.485 60.585 ;
    RECT 130.775 59.865 131.285 60.585 ;
    RECT 131.955 59.865 133.505 60.585 ;
    RECT 133.855 59.865 134.205 60.585 ;
    RECT 134.86 59.865 136.4 60.585 ;
    RECT 137.2 59.865 137.52 60.585 ;
    RECT 137.8 59.865 138.26 60.585 ;
    RECT 139.06 59.865 139.6 60.585 ;
    RECT 140.07 59.865 140.785 60.585 ;
    RECT 141.075 59.865 141.28 60.585 ;
    RECT 142.28 59.865 142.44 60.585 ;
    RECT 142.79 59.865 142.96 60.585 ;
    RECT 144.03 59.865 145.765 60.585 ;
    RECT 146.505 59.865 146.695 60.585 ;
    RECT 147.045 59.865 147.17 60.585 ;
    RECT 121.21 59.145 121.33 59.865 ;
    RECT 121.62 59.145 121.97 59.865 ;
    RECT 122.555 59.145 124.12 59.865 ;
    RECT 125.39 59.145 125.545 59.865 ;
    RECT 126.005 59.145 126.63 59.865 ;
    RECT 127.1 59.145 127.25 59.865 ;
    RECT 127.6 59.145 127.995 59.865 ;
    RECT 128.285 59.145 128.605 59.865 ;
    RECT 129.035 59.145 129.315 59.865 ;
    RECT 129.785 59.145 130.485 59.865 ;
    RECT 130.775 59.145 131.285 59.865 ;
    RECT 131.955 59.145 133.505 59.865 ;
    RECT 133.855 59.145 134.205 59.865 ;
    RECT 134.86 59.145 136.4 59.865 ;
    RECT 137.2 59.145 137.52 59.865 ;
    RECT 137.8 59.145 138.26 59.865 ;
    RECT 139.06 59.145 139.6 59.865 ;
    RECT 140.07 59.145 140.785 59.865 ;
    RECT 141.075 59.145 141.28 59.865 ;
    RECT 142.28 59.145 142.44 59.865 ;
    RECT 142.79 59.145 142.96 59.865 ;
    RECT 144.03 59.145 145.765 59.865 ;
    RECT 146.505 59.145 146.695 59.865 ;
    RECT 147.045 59.145 147.17 59.865 ;
    RECT 121.21 58.425 121.33 59.145 ;
    RECT 121.62 58.425 121.97 59.145 ;
    RECT 122.555 58.425 124.12 59.145 ;
    RECT 125.39 58.425 125.545 59.145 ;
    RECT 126.005 58.425 126.63 59.145 ;
    RECT 127.1 58.425 127.25 59.145 ;
    RECT 127.6 58.425 127.995 59.145 ;
    RECT 128.285 58.425 128.605 59.145 ;
    RECT 129.035 58.425 129.315 59.145 ;
    RECT 129.785 58.425 130.485 59.145 ;
    RECT 130.775 58.425 131.285 59.145 ;
    RECT 131.955 58.425 133.505 59.145 ;
    RECT 133.855 58.425 134.205 59.145 ;
    RECT 134.86 58.425 136.4 59.145 ;
    RECT 137.2 58.425 137.52 59.145 ;
    RECT 137.8 58.425 138.26 59.145 ;
    RECT 139.06 58.425 139.6 59.145 ;
    RECT 140.07 58.425 140.785 59.145 ;
    RECT 141.075 58.425 141.28 59.145 ;
    RECT 142.28 58.425 142.44 59.145 ;
    RECT 142.79 58.425 142.96 59.145 ;
    RECT 144.03 58.425 145.765 59.145 ;
    RECT 146.505 58.425 146.695 59.145 ;
    RECT 147.045 58.425 147.17 59.145 ;
    RECT 121.21 57.705 121.33 58.425 ;
    RECT 121.62 57.705 121.97 58.425 ;
    RECT 122.555 57.705 124.12 58.425 ;
    RECT 125.39 57.705 125.545 58.425 ;
    RECT 126.005 57.705 126.63 58.425 ;
    RECT 127.1 57.705 127.25 58.425 ;
    RECT 127.6 57.705 127.995 58.425 ;
    RECT 128.285 57.705 128.605 58.425 ;
    RECT 129.035 57.705 129.315 58.425 ;
    RECT 129.785 57.705 130.485 58.425 ;
    RECT 130.775 57.705 131.285 58.425 ;
    RECT 131.955 57.705 133.505 58.425 ;
    RECT 133.855 57.705 134.205 58.425 ;
    RECT 134.86 57.705 136.4 58.425 ;
    RECT 137.2 57.705 137.52 58.425 ;
    RECT 137.8 57.705 138.26 58.425 ;
    RECT 139.06 57.705 139.6 58.425 ;
    RECT 140.07 57.705 140.785 58.425 ;
    RECT 141.075 57.705 141.28 58.425 ;
    RECT 142.28 57.705 142.44 58.425 ;
    RECT 142.79 57.705 142.96 58.425 ;
    RECT 144.03 57.705 145.765 58.425 ;
    RECT 146.505 57.705 146.695 58.425 ;
    RECT 147.045 57.705 147.17 58.425 ;
    RECT 121.21 56.985 121.33 57.705 ;
    RECT 121.62 56.985 121.97 57.705 ;
    RECT 122.555 56.985 124.12 57.705 ;
    RECT 125.39 56.985 125.545 57.705 ;
    RECT 126.005 56.985 126.63 57.705 ;
    RECT 127.1 56.985 127.25 57.705 ;
    RECT 127.6 56.985 127.995 57.705 ;
    RECT 128.285 56.985 128.605 57.705 ;
    RECT 129.035 56.985 129.315 57.705 ;
    RECT 129.785 56.985 130.485 57.705 ;
    RECT 130.775 56.985 131.285 57.705 ;
    RECT 131.955 56.985 133.505 57.705 ;
    RECT 133.855 56.985 134.205 57.705 ;
    RECT 134.86 56.985 136.4 57.705 ;
    RECT 137.2 56.985 137.52 57.705 ;
    RECT 137.8 56.985 138.26 57.705 ;
    RECT 139.06 56.985 139.6 57.705 ;
    RECT 140.07 56.985 140.785 57.705 ;
    RECT 141.075 56.985 141.28 57.705 ;
    RECT 142.28 56.985 142.44 57.705 ;
    RECT 142.79 56.985 142.96 57.705 ;
    RECT 144.03 56.985 145.765 57.705 ;
    RECT 146.505 56.985 146.695 57.705 ;
    RECT 147.045 56.985 147.17 57.705 ;
    RECT 121.21 56.265 121.33 56.985 ;
    RECT 121.62 56.265 121.97 56.985 ;
    RECT 122.555 56.265 124.12 56.985 ;
    RECT 125.39 56.265 125.545 56.985 ;
    RECT 126.005 56.265 126.63 56.985 ;
    RECT 127.1 56.265 127.25 56.985 ;
    RECT 127.6 56.265 127.995 56.985 ;
    RECT 128.285 56.265 128.605 56.985 ;
    RECT 129.035 56.265 129.315 56.985 ;
    RECT 129.785 56.265 130.485 56.985 ;
    RECT 130.775 56.265 131.285 56.985 ;
    RECT 131.955 56.265 133.505 56.985 ;
    RECT 133.855 56.265 134.205 56.985 ;
    RECT 134.86 56.265 136.4 56.985 ;
    RECT 137.2 56.265 137.52 56.985 ;
    RECT 137.8 56.265 138.26 56.985 ;
    RECT 139.06 56.265 139.6 56.985 ;
    RECT 140.07 56.265 140.785 56.985 ;
    RECT 141.075 56.265 141.28 56.985 ;
    RECT 142.28 56.265 142.44 56.985 ;
    RECT 142.79 56.265 142.96 56.985 ;
    RECT 144.03 56.265 145.765 56.985 ;
    RECT 146.505 56.265 146.695 56.985 ;
    RECT 147.045 56.265 147.17 56.985 ;
    RECT 121.21 55.545 121.33 56.265 ;
    RECT 121.62 55.545 121.97 56.265 ;
    RECT 122.555 55.545 124.12 56.265 ;
    RECT 125.39 55.545 125.545 56.265 ;
    RECT 126.005 55.545 126.63 56.265 ;
    RECT 127.1 55.545 127.25 56.265 ;
    RECT 127.6 55.545 127.995 56.265 ;
    RECT 128.285 55.545 128.605 56.265 ;
    RECT 129.035 55.545 129.315 56.265 ;
    RECT 129.785 55.545 130.485 56.265 ;
    RECT 130.775 55.545 131.285 56.265 ;
    RECT 131.955 55.545 133.505 56.265 ;
    RECT 133.855 55.545 134.205 56.265 ;
    RECT 134.86 55.545 136.4 56.265 ;
    RECT 137.2 55.545 137.52 56.265 ;
    RECT 137.8 55.545 138.26 56.265 ;
    RECT 139.06 55.545 139.6 56.265 ;
    RECT 140.07 55.545 140.785 56.265 ;
    RECT 141.075 55.545 141.28 56.265 ;
    RECT 142.28 55.545 142.44 56.265 ;
    RECT 142.79 55.545 142.96 56.265 ;
    RECT 144.03 55.545 145.765 56.265 ;
    RECT 146.505 55.545 146.695 56.265 ;
    RECT 147.045 55.545 147.17 56.265 ;
    RECT 121.21 54.825 121.33 55.545 ;
    RECT 121.62 54.825 121.97 55.545 ;
    RECT 122.555 54.825 124.12 55.545 ;
    RECT 125.39 54.825 125.545 55.545 ;
    RECT 126.005 54.825 126.63 55.545 ;
    RECT 127.1 54.825 127.25 55.545 ;
    RECT 127.6 54.825 127.995 55.545 ;
    RECT 128.285 54.825 128.605 55.545 ;
    RECT 129.035 54.825 129.315 55.545 ;
    RECT 129.785 54.825 130.485 55.545 ;
    RECT 130.775 54.825 131.285 55.545 ;
    RECT 131.955 54.825 133.505 55.545 ;
    RECT 133.855 54.825 134.205 55.545 ;
    RECT 134.86 54.825 136.4 55.545 ;
    RECT 137.2 54.825 137.52 55.545 ;
    RECT 137.8 54.825 138.26 55.545 ;
    RECT 139.06 54.825 139.6 55.545 ;
    RECT 140.07 54.825 140.785 55.545 ;
    RECT 141.075 54.825 141.28 55.545 ;
    RECT 142.28 54.825 142.44 55.545 ;
    RECT 142.79 54.825 142.96 55.545 ;
    RECT 144.03 54.825 145.765 55.545 ;
    RECT 146.505 54.825 146.695 55.545 ;
    RECT 147.045 54.825 147.17 55.545 ;
    RECT 121.21 54.105 121.33 54.825 ;
    RECT 121.62 54.105 121.97 54.825 ;
    RECT 122.555 54.105 124.12 54.825 ;
    RECT 125.39 54.105 125.545 54.825 ;
    RECT 126.005 54.105 126.63 54.825 ;
    RECT 127.1 54.105 127.25 54.825 ;
    RECT 127.6 54.105 127.995 54.825 ;
    RECT 128.285 54.105 128.605 54.825 ;
    RECT 129.035 54.105 129.315 54.825 ;
    RECT 129.785 54.105 130.485 54.825 ;
    RECT 130.775 54.105 131.285 54.825 ;
    RECT 131.955 54.105 133.505 54.825 ;
    RECT 133.855 54.105 134.205 54.825 ;
    RECT 134.86 54.105 136.4 54.825 ;
    RECT 137.2 54.105 137.52 54.825 ;
    RECT 137.8 54.105 138.26 54.825 ;
    RECT 139.06 54.105 139.6 54.825 ;
    RECT 140.07 54.105 140.785 54.825 ;
    RECT 141.075 54.105 141.28 54.825 ;
    RECT 142.28 54.105 142.44 54.825 ;
    RECT 142.79 54.105 142.96 54.825 ;
    RECT 144.03 54.105 145.765 54.825 ;
    RECT 146.505 54.105 146.695 54.825 ;
    RECT 147.045 54.105 147.17 54.825 ;
    RECT 121.21 53.385 121.33 54.105 ;
    RECT 121.62 53.385 121.97 54.105 ;
    RECT 122.555 53.385 124.12 54.105 ;
    RECT 125.39 53.385 125.545 54.105 ;
    RECT 126.005 53.385 126.63 54.105 ;
    RECT 127.1 53.385 127.25 54.105 ;
    RECT 127.6 53.385 127.995 54.105 ;
    RECT 128.285 53.385 128.605 54.105 ;
    RECT 129.035 53.385 129.315 54.105 ;
    RECT 129.785 53.385 130.485 54.105 ;
    RECT 130.775 53.385 131.285 54.105 ;
    RECT 131.955 53.385 133.505 54.105 ;
    RECT 133.855 53.385 134.205 54.105 ;
    RECT 134.86 53.385 136.4 54.105 ;
    RECT 137.2 53.385 137.52 54.105 ;
    RECT 137.8 53.385 138.26 54.105 ;
    RECT 139.06 53.385 139.6 54.105 ;
    RECT 140.07 53.385 140.785 54.105 ;
    RECT 141.075 53.385 141.28 54.105 ;
    RECT 142.28 53.385 142.44 54.105 ;
    RECT 142.79 53.385 142.96 54.105 ;
    RECT 144.03 53.385 145.765 54.105 ;
    RECT 146.505 53.385 146.695 54.105 ;
    RECT 147.045 53.385 147.17 54.105 ;
    RECT 121.21 52.665 121.33 53.385 ;
    RECT 121.62 52.665 121.97 53.385 ;
    RECT 122.555 52.665 124.12 53.385 ;
    RECT 125.39 52.665 125.545 53.385 ;
    RECT 126.005 52.665 126.63 53.385 ;
    RECT 127.1 52.665 127.25 53.385 ;
    RECT 127.6 52.665 127.995 53.385 ;
    RECT 128.285 52.665 128.605 53.385 ;
    RECT 129.035 52.665 129.315 53.385 ;
    RECT 129.785 52.665 130.485 53.385 ;
    RECT 130.775 52.665 131.285 53.385 ;
    RECT 131.955 52.665 133.505 53.385 ;
    RECT 133.855 52.665 134.205 53.385 ;
    RECT 134.86 52.665 136.4 53.385 ;
    RECT 137.2 52.665 137.52 53.385 ;
    RECT 137.8 52.665 138.26 53.385 ;
    RECT 139.06 52.665 139.6 53.385 ;
    RECT 140.07 52.665 140.785 53.385 ;
    RECT 141.075 52.665 141.28 53.385 ;
    RECT 142.28 52.665 142.44 53.385 ;
    RECT 142.79 52.665 142.96 53.385 ;
    RECT 144.03 52.665 145.765 53.385 ;
    RECT 146.505 52.665 146.695 53.385 ;
    RECT 147.045 52.665 147.17 53.385 ;
    RECT 121.21 51.945 121.33 52.665 ;
    RECT 121.62 51.945 121.97 52.665 ;
    RECT 122.555 51.945 124.12 52.665 ;
    RECT 125.39 51.945 125.545 52.665 ;
    RECT 126.005 51.945 126.63 52.665 ;
    RECT 127.1 51.945 127.25 52.665 ;
    RECT 127.6 51.945 127.995 52.665 ;
    RECT 128.285 51.945 128.605 52.665 ;
    RECT 129.035 51.945 129.315 52.665 ;
    RECT 129.785 51.945 130.485 52.665 ;
    RECT 130.775 51.945 131.285 52.665 ;
    RECT 131.955 51.945 133.505 52.665 ;
    RECT 133.855 51.945 134.205 52.665 ;
    RECT 134.86 51.945 136.4 52.665 ;
    RECT 137.2 51.945 137.52 52.665 ;
    RECT 137.8 51.945 138.26 52.665 ;
    RECT 139.06 51.945 139.6 52.665 ;
    RECT 140.07 51.945 140.785 52.665 ;
    RECT 141.075 51.945 141.28 52.665 ;
    RECT 142.28 51.945 142.44 52.665 ;
    RECT 142.79 51.945 142.96 52.665 ;
    RECT 144.03 51.945 145.765 52.665 ;
    RECT 146.505 51.945 146.695 52.665 ;
    RECT 147.045 51.945 147.17 52.665 ;
    RECT 121.21 51.225 121.33 51.945 ;
    RECT 121.62 51.225 121.97 51.945 ;
    RECT 122.555 51.225 124.12 51.945 ;
    RECT 125.39 51.225 125.545 51.945 ;
    RECT 126.005 51.225 126.63 51.945 ;
    RECT 127.1 51.225 127.25 51.945 ;
    RECT 127.6 51.225 127.995 51.945 ;
    RECT 128.285 51.225 128.605 51.945 ;
    RECT 129.035 51.225 129.315 51.945 ;
    RECT 129.785 51.225 130.485 51.945 ;
    RECT 130.775 51.225 131.285 51.945 ;
    RECT 131.955 51.225 133.505 51.945 ;
    RECT 133.855 51.225 134.205 51.945 ;
    RECT 134.86 51.225 136.4 51.945 ;
    RECT 137.2 51.225 137.52 51.945 ;
    RECT 137.8 51.225 138.26 51.945 ;
    RECT 139.06 51.225 139.6 51.945 ;
    RECT 140.07 51.225 140.785 51.945 ;
    RECT 141.075 51.225 141.28 51.945 ;
    RECT 142.28 51.225 142.44 51.945 ;
    RECT 142.79 51.225 142.96 51.945 ;
    RECT 144.03 51.225 145.765 51.945 ;
    RECT 146.505 51.225 146.695 51.945 ;
    RECT 147.045 51.225 147.17 51.945 ;
    RECT 121.21 50.505 121.33 51.225 ;
    RECT 121.62 50.505 121.97 51.225 ;
    RECT 122.555 50.505 124.12 51.225 ;
    RECT 125.39 50.505 125.545 51.225 ;
    RECT 126.005 50.505 126.63 51.225 ;
    RECT 127.1 50.505 127.25 51.225 ;
    RECT 127.6 50.505 127.995 51.225 ;
    RECT 128.285 50.505 128.605 51.225 ;
    RECT 129.035 50.505 129.315 51.225 ;
    RECT 129.785 50.505 130.485 51.225 ;
    RECT 130.775 50.505 131.285 51.225 ;
    RECT 131.955 50.505 133.505 51.225 ;
    RECT 133.855 50.505 134.205 51.225 ;
    RECT 134.86 50.505 136.4 51.225 ;
    RECT 137.2 50.505 137.52 51.225 ;
    RECT 137.8 50.505 138.26 51.225 ;
    RECT 139.06 50.505 139.6 51.225 ;
    RECT 140.07 50.505 140.785 51.225 ;
    RECT 141.075 50.505 141.28 51.225 ;
    RECT 142.28 50.505 142.44 51.225 ;
    RECT 142.79 50.505 142.96 51.225 ;
    RECT 144.03 50.505 145.765 51.225 ;
    RECT 146.505 50.505 146.695 51.225 ;
    RECT 147.045 50.505 147.17 51.225 ;
    RECT 180.59 2.9 180.66 6.45 ;
    RECT 180.59 6.685 180.66 12.485 ;
    RECT 180.39 8.225 180.46 10.34 ;
    RECT 178.915 2.135 179.195 12.49 ;
    RECT 177.27 2.9 177.34 6.45 ;
    RECT 177.27 6.685 177.34 12.485 ;
    RECT 177.07 8.225 177.14 10.34 ;
    RECT 175.595 2.135 175.875 12.49 ;
    RECT 173.95 2.9 174.02 6.45 ;
    RECT 173.95 6.685 174.02 12.485 ;
    RECT 173.75 8.225 173.82 10.34 ;
    RECT 172.275 2.135 172.555 12.49 ;
    RECT 170.63 2.9 170.7 6.45 ;
    RECT 170.63 6.685 170.7 12.485 ;
    RECT 170.43 8.225 170.5 10.34 ;
    RECT 168.955 2.135 169.235 12.49 ;
    RECT 167.31 2.9 167.38 6.45 ;
    RECT 167.31 6.685 167.38 12.485 ;
    RECT 167.11 8.225 167.18 10.34 ;
    RECT 165.635 2.135 165.915 12.49 ;
    RECT 163.99 2.9 164.06 6.45 ;
    RECT 163.99 6.685 164.06 12.485 ;
    RECT 163.79 8.225 163.86 10.34 ;
    RECT 162.315 2.135 162.595 12.49 ;
    RECT 160.67 2.9 160.74 6.45 ;
    RECT 160.67 6.685 160.74 12.485 ;
    RECT 160.47 8.225 160.54 10.34 ;
    RECT 158.995 2.135 159.275 12.49 ;
    RECT 157.35 2.9 157.42 6.45 ;
    RECT 157.35 6.685 157.42 12.485 ;
    RECT 157.15 8.225 157.22 10.34 ;
    RECT 155.675 2.135 155.955 12.49 ;
    RECT 154.03 2.9 154.1 6.45 ;
    RECT 154.03 6.685 154.1 12.485 ;
    RECT 153.83 8.225 153.9 10.34 ;
    RECT 152.355 2.135 152.635 12.49 ;
    RECT 266.91 2.9 266.98 6.45 ;
    RECT 266.91 6.685 266.98 12.485 ;
    RECT 266.71 8.225 266.78 10.34 ;
    RECT 265.235 2.135 265.515 12.49 ;
    RECT 150.71 2.9 150.78 6.45 ;
    RECT 150.71 6.685 150.78 12.485 ;
    RECT 150.51 8.225 150.58 10.34 ;
    RECT 149.035 2.135 149.315 12.49 ;
    RECT 263.59 2.9 263.66 6.45 ;
    RECT 263.59 6.685 263.66 12.485 ;
    RECT 263.39 8.225 263.46 10.34 ;
    RECT 261.915 2.135 262.195 12.49 ;
    RECT 260.27 2.9 260.34 6.45 ;
    RECT 260.27 6.685 260.34 12.485 ;
    RECT 260.07 8.225 260.14 10.34 ;
    RECT 258.595 2.135 258.875 12.49 ;
    RECT 256.95 2.9 257.02 6.45 ;
    RECT 256.95 6.685 257.02 12.485 ;
    RECT 256.75 8.225 256.82 10.34 ;
    RECT 255.275 2.135 255.555 12.49 ;
    RECT 253.63 2.9 253.7 6.45 ;
    RECT 253.63 6.685 253.7 12.485 ;
    RECT 253.43 8.225 253.5 10.34 ;
    RECT 251.955 2.135 252.235 12.49 ;
    RECT 250.31 2.9 250.38 6.45 ;
    RECT 250.31 6.685 250.38 12.485 ;
    RECT 250.11 8.225 250.18 10.34 ;
    RECT 248.635 2.135 248.915 12.49 ;
    RECT 246.99 2.9 247.06 6.45 ;
    RECT 246.99 6.685 247.06 12.485 ;
    RECT 246.79 8.225 246.86 10.34 ;
    RECT 245.315 2.135 245.595 12.49 ;
    RECT 243.67 2.9 243.74 6.45 ;
    RECT 243.67 6.685 243.74 12.485 ;
    RECT 243.47 8.225 243.54 10.34 ;
    RECT 241.995 2.135 242.275 12.49 ;
    RECT 240.35 2.9 240.42 6.45 ;
    RECT 240.35 6.685 240.42 12.485 ;
    RECT 240.15 8.225 240.22 10.34 ;
    RECT 238.675 2.135 238.955 12.49 ;
    RECT 237.03 2.9 237.1 6.45 ;
    RECT 237.03 6.685 237.1 12.485 ;
    RECT 236.83 8.225 236.9 10.34 ;
    RECT 235.355 2.135 235.635 12.49 ;
    RECT 233.71 2.9 233.78 6.45 ;
    RECT 233.71 6.685 233.78 12.485 ;
    RECT 233.51 8.225 233.58 10.34 ;
    RECT 232.035 2.135 232.315 12.49 ;
    RECT 230.39 2.9 230.46 6.45 ;
    RECT 230.39 6.685 230.46 12.485 ;
    RECT 230.19 8.225 230.26 10.34 ;
    RECT 228.715 2.135 228.995 12.49 ;
    RECT 227.07 2.9 227.14 6.45 ;
    RECT 227.07 6.685 227.14 12.485 ;
    RECT 226.87 8.225 226.94 10.34 ;
    RECT 225.395 2.135 225.675 12.49 ;
    RECT 223.75 2.9 223.82 6.45 ;
    RECT 223.75 6.685 223.82 12.485 ;
    RECT 223.55 8.225 223.62 10.34 ;
    RECT 222.075 2.135 222.355 12.49 ;
    RECT 220.43 2.9 220.5 6.45 ;
    RECT 220.43 6.685 220.5 12.485 ;
    RECT 220.23 8.225 220.3 10.34 ;
    RECT 218.755 2.135 219.035 12.49 ;
    RECT 217.11 2.9 217.18 6.45 ;
    RECT 217.11 6.685 217.18 12.485 ;
    RECT 216.91 8.225 216.98 10.34 ;
    RECT 215.435 2.135 215.715 12.49 ;
    RECT 213.79 2.9 213.86 6.45 ;
    RECT 213.79 6.685 213.86 12.485 ;
    RECT 213.59 8.225 213.66 10.34 ;
    RECT 212.115 2.135 212.395 12.49 ;
    RECT 210.47 2.9 210.54 6.45 ;
    RECT 210.47 6.685 210.54 12.485 ;
    RECT 210.27 8.225 210.34 10.34 ;
    RECT 208.795 2.135 209.075 12.49 ;
    RECT 207.15 2.9 207.22 6.45 ;
    RECT 207.15 6.685 207.22 12.485 ;
    RECT 206.95 8.225 207.02 10.34 ;
    RECT 205.475 2.135 205.755 12.49 ;
    RECT 203.83 2.9 203.9 6.45 ;
    RECT 203.83 6.685 203.9 12.485 ;
    RECT 203.63 8.225 203.7 10.34 ;
    RECT 202.155 2.135 202.435 12.49 ;
    RECT 200.51 2.9 200.58 6.45 ;
    RECT 200.51 6.685 200.58 12.485 ;
    RECT 200.31 8.225 200.38 10.34 ;
    RECT 198.835 2.135 199.115 12.49 ;
    RECT 197.19 2.9 197.26 6.45 ;
    RECT 197.19 6.685 197.26 12.485 ;
    RECT 196.99 8.225 197.06 10.34 ;
    RECT 195.515 2.135 195.795 12.49 ;
    RECT 193.87 2.9 193.94 6.45 ;
    RECT 193.87 6.685 193.94 12.485 ;
    RECT 193.67 8.225 193.74 10.34 ;
    RECT 192.195 2.135 192.475 12.49 ;
    RECT 190.55 2.9 190.62 6.45 ;
    RECT 190.55 6.685 190.62 12.485 ;
    RECT 190.35 8.225 190.42 10.34 ;
    RECT 188.875 2.135 189.155 12.49 ;
    RECT 187.23 2.9 187.3 6.45 ;
    RECT 187.23 6.685 187.3 12.485 ;
    RECT 187.03 8.225 187.1 10.34 ;
    RECT 185.555 2.135 185.835 12.49 ;
    RECT 183.91 2.9 183.98 6.45 ;
    RECT 183.91 6.685 183.98 12.485 ;
    RECT 183.71 8.225 183.78 10.34 ;
    RECT 182.235 2.135 182.515 12.49 ;
    RECT 263.4 0.695 263.47 1.11 ;
    RECT 261.915 0.695 262.195 2.135 ;
    RECT 260.08 0.695 260.15 1.11 ;
    RECT 258.595 0.695 258.875 2.135 ;
    RECT 256.76 0.695 256.83 1.11 ;
    RECT 255.275 0.695 255.555 2.135 ;
    RECT 253.44 0.695 253.51 1.11 ;
    RECT 251.955 0.695 252.235 2.135 ;
    RECT 250.12 0.695 250.19 1.11 ;
    RECT 248.635 0.695 248.915 2.135 ;
    RECT 266.72 0.695 266.79 1.11 ;
    RECT 265.235 0.695 265.515 2.135 ;
    RECT 150.52 0.695 150.59 1.11 ;
    RECT 149.035 0.695 149.315 2.135 ;
    RECT 246.8 0.695 246.87 1.11 ;
    RECT 245.315 0.695 245.595 2.135 ;
    RECT 243.48 0.695 243.55 1.11 ;
    RECT 241.995 0.695 242.275 2.135 ;
    RECT 240.16 0.695 240.23 1.11 ;
    RECT 238.675 0.695 238.955 2.135 ;
    RECT 236.84 0.695 236.91 1.11 ;
    RECT 235.355 0.695 235.635 2.135 ;
    RECT 233.52 0.695 233.59 1.11 ;
    RECT 232.035 0.695 232.315 2.135 ;
    RECT 230.2 0.695 230.27 1.11 ;
    RECT 228.715 0.695 228.995 2.135 ;
    RECT 226.88 0.695 226.95 1.11 ;
    RECT 225.395 0.695 225.675 2.135 ;
    RECT 223.56 0.695 223.63 1.11 ;
    RECT 222.075 0.695 222.355 2.135 ;
    RECT 220.24 0.695 220.31 1.11 ;
    RECT 218.755 0.695 219.035 2.135 ;
    RECT 216.92 0.695 216.99 1.11 ;
    RECT 215.435 0.695 215.715 2.135 ;
    RECT 180.4 0.695 180.47 1.11 ;
    RECT 178.915 0.695 179.195 2.135 ;
    RECT 177.08 0.695 177.15 1.11 ;
    RECT 175.595 0.695 175.875 2.135 ;
    RECT 173.76 0.695 173.83 1.11 ;
    RECT 172.275 0.695 172.555 2.135 ;
    RECT 170.44 0.695 170.51 1.11 ;
    RECT 168.955 0.695 169.235 2.135 ;
    RECT 167.12 0.695 167.19 1.11 ;
    RECT 165.635 0.695 165.915 2.135 ;
    RECT 163.8 0.695 163.87 1.11 ;
    RECT 162.315 0.695 162.595 2.135 ;
    RECT 160.48 0.695 160.55 1.11 ;
    RECT 158.995 0.695 159.275 2.135 ;
    RECT 157.16 0.695 157.23 1.11 ;
    RECT 155.675 0.695 155.955 2.135 ;
    RECT 153.84 0.695 153.91 1.11 ;
    RECT 152.355 0.695 152.635 2.135 ;
    RECT 213.6 0.695 213.67 1.11 ;
    RECT 212.115 0.695 212.395 2.135 ;
    RECT 210.28 0.695 210.35 1.11 ;
    RECT 208.795 0.695 209.075 2.135 ;
    RECT 206.96 0.695 207.03 1.11 ;
    RECT 205.475 0.695 205.755 2.135 ;
    RECT 203.64 0.695 203.71 1.11 ;
    RECT 202.155 0.695 202.435 2.135 ;
    RECT 200.32 0.695 200.39 1.11 ;
    RECT 198.835 0.695 199.115 2.135 ;
    RECT 197.0 0.695 197.07 1.11 ;
    RECT 195.515 0.695 195.795 2.135 ;
    RECT 193.68 0.695 193.75 1.11 ;
    RECT 192.195 0.695 192.475 2.135 ;
    RECT 190.36 0.695 190.43 1.11 ;
    RECT 188.875 0.695 189.155 2.135 ;
    RECT 187.04 0.695 187.11 1.11 ;
    RECT 185.555 0.695 185.835 2.135 ;
    RECT 183.72 0.695 183.79 1.11 ;
    RECT 182.235 0.695 182.515 2.135 ;
    RECT 120.445 0.695 120.525 14.505 ;
    RECT 121.195 0.695 121.33 14.505 ;
    RECT 121.62 0.695 121.97 14.505 ;
    RECT 122.555 0.695 124.12 14.505 ;
    RECT 125.39 0.695 125.545 14.505 ;
    RECT 126.005 0.695 126.63 14.505 ;
    RECT 127.1 0.695 127.25 14.505 ;
    RECT 127.6 0.695 127.995 14.505 ;
    RECT 128.285 0.695 128.605 6.55 ;
    RECT 129.035 0.695 129.315 14.505 ;
    RECT 129.785 0.695 130.485 14.505 ;
    RECT 130.775 0.695 131.285 14.505 ;
    RECT 131.955 0.695 133.505 14.505 ;
    RECT 133.855 0.695 134.205 14.505 ;
    RECT 134.685 0.695 136.4 14.505 ;
    RECT 137.2 0.695 137.52 14.505 ;
    RECT 137.8 0.695 138.26 14.505 ;
    RECT 139.06 0.695 139.6 14.505 ;
    RECT 139.6 0.695 140.07 0.915 ;
    RECT 140.07 0.695 140.785 14.505 ;
    RECT 141.075 0.695 141.28 14.505 ;
    RECT 142.28 0.695 142.44 14.505 ;
    RECT 142.79 0.695 142.96 14.505 ;
    RECT 144.03 0.695 145.765 14.505 ;
    RECT 146.505 0.695 146.695 14.505 ;
    RECT 147.045 0.695 147.185 14.505 ;
    RECT 147.855 0.695 147.935 14.505 ;
    RECT 117.79 0.695 117.86 1.11 ;
    RECT 119.065 0.695 119.345 2.135 ;
    RECT 1.59 0.695 1.66 1.11 ;
    RECT 2.865 0.695 3.145 2.135 ;
    RECT 31.47 0.695 31.54 1.11 ;
    RECT 32.745 0.695 33.025 2.135 ;
    RECT 28.15 0.695 28.22 1.11 ;
    RECT 29.425 0.695 29.705 2.135 ;
    RECT 24.83 0.695 24.9 1.11 ;
    RECT 26.105 0.695 26.385 2.135 ;
    RECT 21.51 0.695 21.58 1.11 ;
    RECT 22.785 0.695 23.065 2.135 ;
    RECT 18.19 0.695 18.26 1.11 ;
    RECT 19.465 0.695 19.745 2.135 ;
    RECT 14.87 0.695 14.94 1.11 ;
    RECT 16.145 0.695 16.425 2.135 ;
    RECT 11.55 0.695 11.62 1.11 ;
    RECT 12.825 0.695 13.105 2.135 ;
    RECT 8.23 0.695 8.3 1.11 ;
    RECT 9.505 0.695 9.785 2.135 ;
    RECT 4.91 0.695 4.98 1.11 ;
    RECT 6.185 0.695 6.465 2.135 ;
    RECT 114.47 0.695 114.54 1.11 ;
    RECT 115.745 0.695 116.025 2.135 ;
    RECT 111.15 0.695 111.22 1.11 ;
    RECT 112.425 0.695 112.705 2.135 ;
    RECT 107.83 0.695 107.9 1.11 ;
    RECT 109.105 0.695 109.385 2.135 ;
    RECT 104.51 0.695 104.58 1.11 ;
    RECT 105.785 0.695 106.065 2.135 ;
    RECT 101.19 0.695 101.26 1.11 ;
    RECT 102.465 0.695 102.745 2.135 ;
    RECT 97.87 0.695 97.94 1.11 ;
    RECT 99.145 0.695 99.425 2.135 ;
    RECT 94.55 0.695 94.62 1.11 ;
    RECT 95.825 0.695 96.105 2.135 ;
    RECT 91.23 0.695 91.3 1.11 ;
    RECT 92.505 0.695 92.785 2.135 ;
    RECT 87.91 0.695 87.98 1.11 ;
    RECT 89.185 0.695 89.465 2.135 ;
    RECT 84.59 0.695 84.66 1.11 ;
    RECT 85.865 0.695 86.145 2.135 ;
    RECT 81.27 0.695 81.34 1.11 ;
    RECT 82.545 0.695 82.825 2.135 ;
    RECT 77.95 0.695 78.02 1.11 ;
    RECT 79.225 0.695 79.505 2.135 ;
    RECT 74.63 0.695 74.7 1.11 ;
    RECT 75.905 0.695 76.185 2.135 ;
    RECT 71.31 0.695 71.38 1.11 ;
    RECT 72.585 0.695 72.865 2.135 ;
    RECT 67.99 0.695 68.06 1.11 ;
    RECT 69.265 0.695 69.545 2.135 ;
    RECT 64.67 0.695 64.74 1.11 ;
    RECT 65.945 0.695 66.225 2.135 ;
    RECT 61.35 0.695 61.42 1.11 ;
    RECT 62.625 0.695 62.905 2.135 ;
    RECT 58.03 0.695 58.1 1.11 ;
    RECT 59.305 0.695 59.585 2.135 ;
    RECT 54.71 0.695 54.78 1.11 ;
    RECT 55.985 0.695 56.265 2.135 ;
    RECT 51.39 0.695 51.46 1.11 ;
    RECT 52.665 0.695 52.945 2.135 ;
    RECT 48.07 0.695 48.14 1.11 ;
    RECT 49.345 0.695 49.625 2.135 ;
    RECT 44.75 0.695 44.82 1.11 ;
    RECT 46.025 0.695 46.305 2.135 ;
    RECT 41.43 0.695 41.5 1.11 ;
    RECT 42.705 0.695 42.985 2.135 ;
    RECT 38.11 0.695 38.18 1.11 ;
    RECT 39.385 0.695 39.665 2.135 ;
    RECT 34.79 0.695 34.86 1.11 ;
    RECT 36.065 0.695 36.345 2.135 ;
    RECT 117.6 2.9 117.67 6.45 ;
    RECT 117.6 6.685 117.67 12.485 ;
    RECT 117.8 8.225 117.87 10.34 ;
    RECT 119.065 2.135 119.345 12.49 ;
    RECT 1.4 2.9 1.47 6.45 ;
    RECT 1.4 6.685 1.47 12.485 ;
    RECT 1.6 8.225 1.67 10.34 ;
    RECT 2.865 2.135 3.145 12.49 ;
    RECT 31.28 2.9 31.35 6.45 ;
    RECT 31.28 6.685 31.35 12.485 ;
    RECT 31.48 8.225 31.55 10.34 ;
    RECT 32.745 2.135 33.025 12.49 ;
    RECT 27.96 2.9 28.03 6.45 ;
    RECT 27.96 6.685 28.03 12.485 ;
    RECT 28.16 8.225 28.23 10.34 ;
    RECT 29.425 2.135 29.705 12.49 ;
    RECT 24.64 2.9 24.71 6.45 ;
    RECT 24.64 6.685 24.71 12.485 ;
    RECT 24.84 8.225 24.91 10.34 ;
    RECT 26.105 2.135 26.385 12.49 ;
    RECT 21.32 2.9 21.39 6.45 ;
    RECT 21.32 6.685 21.39 12.485 ;
    RECT 21.52 8.225 21.59 10.34 ;
    RECT 22.785 2.135 23.065 12.49 ;
    RECT 18.0 2.9 18.07 6.45 ;
    RECT 18.0 6.685 18.07 12.485 ;
    RECT 18.2 8.225 18.27 10.34 ;
    RECT 19.465 2.135 19.745 12.49 ;
    RECT 14.68 2.9 14.75 6.45 ;
    RECT 14.68 6.685 14.75 12.485 ;
    RECT 14.88 8.225 14.95 10.34 ;
    RECT 16.145 2.135 16.425 12.49 ;
    RECT 11.36 2.9 11.43 6.45 ;
    RECT 11.36 6.685 11.43 12.485 ;
    RECT 11.56 8.225 11.63 10.34 ;
    RECT 12.825 2.135 13.105 12.49 ;
    RECT 8.04 2.9 8.11 6.45 ;
    RECT 8.04 6.685 8.11 12.485 ;
    RECT 8.24 8.225 8.31 10.34 ;
    RECT 9.505 2.135 9.785 12.49 ;
    RECT 4.72 2.9 4.79 6.45 ;
    RECT 4.72 6.685 4.79 12.485 ;
    RECT 4.92 8.225 4.99 10.34 ;
    RECT 6.185 2.135 6.465 12.49 ;
    RECT 114.28 2.9 114.35 6.45 ;
    RECT 114.28 6.685 114.35 12.485 ;
    RECT 114.48 8.225 114.55 10.34 ;
    RECT 115.745 2.135 116.025 12.49 ;
    RECT 110.96 2.9 111.03 6.45 ;
    RECT 110.96 6.685 111.03 12.485 ;
    RECT 111.16 8.225 111.23 10.34 ;
    RECT 112.425 2.135 112.705 12.49 ;
    RECT 107.64 2.9 107.71 6.45 ;
    RECT 107.64 6.685 107.71 12.485 ;
    RECT 107.84 8.225 107.91 10.34 ;
    RECT 109.105 2.135 109.385 12.49 ;
    RECT 104.32 2.9 104.39 6.45 ;
    RECT 104.32 6.685 104.39 12.485 ;
    RECT 104.52 8.225 104.59 10.34 ;
    RECT 105.785 2.135 106.065 12.49 ;
    RECT 101.0 2.9 101.07 6.45 ;
    RECT 101.0 6.685 101.07 12.485 ;
    RECT 101.2 8.225 101.27 10.34 ;
    RECT 102.465 2.135 102.745 12.49 ;
    RECT 97.68 2.9 97.75 6.45 ;
    RECT 97.68 6.685 97.75 12.485 ;
    RECT 97.88 8.225 97.95 10.34 ;
    RECT 99.145 2.135 99.425 12.49 ;
    RECT 94.36 2.9 94.43 6.45 ;
    RECT 94.36 6.685 94.43 12.485 ;
    RECT 94.56 8.225 94.63 10.34 ;
    RECT 95.825 2.135 96.105 12.49 ;
    RECT 91.04 2.9 91.11 6.45 ;
    RECT 91.04 6.685 91.11 12.485 ;
    RECT 91.24 8.225 91.31 10.34 ;
    RECT 92.505 2.135 92.785 12.49 ;
    RECT 87.72 2.9 87.79 6.45 ;
    RECT 87.72 6.685 87.79 12.485 ;
    RECT 87.92 8.225 87.99 10.34 ;
    RECT 89.185 2.135 89.465 12.49 ;
    RECT 84.4 2.9 84.47 6.45 ;
    RECT 84.4 6.685 84.47 12.485 ;
    RECT 84.6 8.225 84.67 10.34 ;
    RECT 85.865 2.135 86.145 12.49 ;
    RECT 81.08 2.9 81.15 6.45 ;
    RECT 81.08 6.685 81.15 12.485 ;
    RECT 81.28 8.225 81.35 10.34 ;
    RECT 82.545 2.135 82.825 12.49 ;
    RECT 77.76 2.9 77.83 6.45 ;
    RECT 77.76 6.685 77.83 12.485 ;
    RECT 77.96 8.225 78.03 10.34 ;
    RECT 79.225 2.135 79.505 12.49 ;
    RECT 74.44 2.9 74.51 6.45 ;
    RECT 74.44 6.685 74.51 12.485 ;
    RECT 74.64 8.225 74.71 10.34 ;
    RECT 75.905 2.135 76.185 12.49 ;
    RECT 71.12 2.9 71.19 6.45 ;
    RECT 71.12 6.685 71.19 12.485 ;
    RECT 71.32 8.225 71.39 10.34 ;
    RECT 72.585 2.135 72.865 12.49 ;
    RECT 67.8 2.9 67.87 6.45 ;
    RECT 67.8 6.685 67.87 12.485 ;
    RECT 68.0 8.225 68.07 10.34 ;
    RECT 69.265 2.135 69.545 12.49 ;
    RECT 64.48 2.9 64.55 6.45 ;
    RECT 64.48 6.685 64.55 12.485 ;
    RECT 64.68 8.225 64.75 10.34 ;
    RECT 65.945 2.135 66.225 12.49 ;
    RECT 61.16 2.9 61.23 6.45 ;
    RECT 61.16 6.685 61.23 12.485 ;
    RECT 61.36 8.225 61.43 10.34 ;
    RECT 62.625 2.135 62.905 12.49 ;
    RECT 57.84 2.9 57.91 6.45 ;
    RECT 57.84 6.685 57.91 12.485 ;
    RECT 58.04 8.225 58.11 10.34 ;
    RECT 59.305 2.135 59.585 12.49 ;
    RECT 54.52 2.9 54.59 6.45 ;
    RECT 54.52 6.685 54.59 12.485 ;
    RECT 54.72 8.225 54.79 10.34 ;
    RECT 55.985 2.135 56.265 12.49 ;
    RECT 51.2 2.9 51.27 6.45 ;
    RECT 51.2 6.685 51.27 12.485 ;
    RECT 51.4 8.225 51.47 10.34 ;
    RECT 52.665 2.135 52.945 12.49 ;
    RECT 47.88 2.9 47.95 6.45 ;
    RECT 47.88 6.685 47.95 12.485 ;
    RECT 48.08 8.225 48.15 10.34 ;
    RECT 49.345 2.135 49.625 12.49 ;
    RECT 44.56 2.9 44.63 6.45 ;
    RECT 44.56 6.685 44.63 12.485 ;
    RECT 44.76 8.225 44.83 10.34 ;
    RECT 46.025 2.135 46.305 12.49 ;
    RECT 41.24 2.9 41.31 6.45 ;
    RECT 41.24 6.685 41.31 12.485 ;
    RECT 41.44 8.225 41.51 10.34 ;
    RECT 42.705 2.135 42.985 12.49 ;
    RECT 37.92 2.9 37.99 6.45 ;
    RECT 37.92 6.685 37.99 12.485 ;
    RECT 38.12 8.225 38.19 10.34 ;
    RECT 39.385 2.135 39.665 12.49 ;
    RECT 34.6 2.9 34.67 6.45 ;
    RECT 34.6 6.685 34.67 12.485 ;
    RECT 34.8 8.225 34.87 10.34 ;
    RECT 36.065 2.135 36.345 12.49 ;
    RECT 120.445 100.295 120.525 100.88 ;
    RECT 121.195 100.295 121.33 100.88 ;
    RECT 121.62 100.685 121.97 100.88 ;
    RECT 122.555 100.295 124.12 100.88 ;
    RECT 125.39 100.295 125.545 100.88 ;
    RECT 126.005 100.295 126.63 100.88 ;
    RECT 127.1 100.295 127.25 100.88 ;
    RECT 127.6 100.295 127.995 100.88 ;
    RECT 128.285 100.295 128.605 100.88 ;
    RECT 129.035 100.295 129.315 100.88 ;
    RECT 129.785 100.295 130.485 100.88 ;
    RECT 130.775 100.295 131.285 100.88 ;
    RECT 131.955 100.295 133.505 100.88 ;
    RECT 133.855 100.295 134.205 100.88 ;
    RECT 134.685 100.295 136.4 100.88 ;
    RECT 137.2 100.295 137.52 100.88 ;
    RECT 137.8 100.295 138.26 100.88 ;
    RECT 139.06 100.295 139.6 100.88 ;
    RECT 140.07 100.295 140.785 100.88 ;
    RECT 141.075 100.295 141.28 100.88 ;
    RECT 142.28 100.295 142.44 100.88 ;
    RECT 142.79 100.295 142.96 100.88 ;
    RECT 144.03 100.295 145.765 100.88 ;
    RECT 146.505 100.295 146.695 100.88 ;
    RECT 147.045 100.295 147.185 100.88 ;
    RECT 147.855 100.295 147.935 100.88 ;
    #obstructions of filtered out pwrgnd shapes
    RECT 250.045 36.025 250.325 36.905 ;
    RECT 246.725 36.025 247.005 36.905 ;
    RECT 243.405 36.025 243.685 36.905 ;
    RECT 240.085 36.025 240.365 36.905 ;
    RECT 236.765 36.025 237.045 36.905 ;
    RECT 233.445 36.025 233.725 36.905 ;
    RECT 230.125 36.025 230.405 36.905 ;
    RECT 226.805 36.025 227.085 36.905 ;
    RECT 223.485 36.025 223.765 36.905 ;
    RECT 220.165 36.025 220.445 36.905 ;
    RECT 216.845 36.025 217.125 36.905 ;
    RECT 180.325 36.025 180.605 36.905 ;
    RECT 177.005 36.025 177.285 36.905 ;
    RECT 173.685 36.025 173.965 36.905 ;
    RECT 170.365 36.025 170.645 36.905 ;
    RECT 167.045 36.025 167.325 36.905 ;
    RECT 163.725 36.025 164.005 36.905 ;
    RECT 160.405 36.025 160.685 36.905 ;
    RECT 157.085 36.025 157.365 36.905 ;
    RECT 153.765 36.025 154.045 36.905 ;
    RECT 150.445 36.025 150.725 36.905 ;
    RECT 213.525 36.025 213.805 36.905 ;
    RECT 210.205 36.025 210.485 36.905 ;
    RECT 206.885 36.025 207.165 36.905 ;
    RECT 203.565 36.025 203.845 36.905 ;
    RECT 200.245 36.025 200.525 36.905 ;
    RECT 196.925 36.025 197.205 36.905 ;
    RECT 193.605 36.025 193.885 36.905 ;
    RECT 190.285 36.025 190.565 36.905 ;
    RECT 186.965 36.025 187.245 36.905 ;
    RECT 183.645 36.025 183.925 36.905 ;
    RECT 266.645 36.025 266.925 36.905 ;
    RECT 263.325 36.025 263.605 36.905 ;
    RECT 260.005 36.025 260.285 36.905 ;
    RECT 256.685 36.025 256.965 36.905 ;
    RECT 253.365 36.025 253.645 36.905 ;
    RECT 250.045 75.645 250.325 76.525 ;
    RECT 246.725 75.645 247.005 76.525 ;
    RECT 243.405 75.645 243.685 76.525 ;
    RECT 240.085 75.645 240.365 76.525 ;
    RECT 236.765 75.645 237.045 76.525 ;
    RECT 233.445 75.645 233.725 76.525 ;
    RECT 230.125 75.645 230.405 76.525 ;
    RECT 226.805 75.645 227.085 76.525 ;
    RECT 223.485 75.645 223.765 76.525 ;
    RECT 220.165 75.645 220.445 76.525 ;
    RECT 216.845 75.645 217.125 76.525 ;
    RECT 180.325 75.645 180.605 76.525 ;
    RECT 177.005 75.645 177.285 76.525 ;
    RECT 173.685 75.645 173.965 76.525 ;
    RECT 170.365 75.645 170.645 76.525 ;
    RECT 167.045 75.645 167.325 76.525 ;
    RECT 163.725 75.645 164.005 76.525 ;
    RECT 160.405 75.645 160.685 76.525 ;
    RECT 157.085 75.645 157.365 76.525 ;
    RECT 153.765 75.645 154.045 76.525 ;
    RECT 150.445 75.645 150.725 76.525 ;
    RECT 213.525 75.645 213.805 76.525 ;
    RECT 210.205 75.645 210.485 76.525 ;
    RECT 206.885 75.645 207.165 76.525 ;
    RECT 203.565 75.645 203.845 76.525 ;
    RECT 200.245 75.645 200.525 76.525 ;
    RECT 196.925 75.645 197.205 76.525 ;
    RECT 193.605 75.645 193.885 76.525 ;
    RECT 190.285 75.645 190.565 76.525 ;
    RECT 186.965 75.645 187.245 76.525 ;
    RECT 183.645 75.645 183.925 76.525 ;
    RECT 266.645 75.645 266.925 76.525 ;
    RECT 263.325 75.645 263.605 76.525 ;
    RECT 260.005 75.645 260.285 76.525 ;
    RECT 256.685 75.645 256.965 76.525 ;
    RECT 253.365 75.645 253.645 76.525 ;
    RECT 250.045 74.925 250.325 75.805 ;
    RECT 246.725 74.925 247.005 75.805 ;
    RECT 243.405 74.925 243.685 75.805 ;
    RECT 240.085 74.925 240.365 75.805 ;
    RECT 236.765 74.925 237.045 75.805 ;
    RECT 233.445 74.925 233.725 75.805 ;
    RECT 230.125 74.925 230.405 75.805 ;
    RECT 226.805 74.925 227.085 75.805 ;
    RECT 223.485 74.925 223.765 75.805 ;
    RECT 220.165 74.925 220.445 75.805 ;
    RECT 216.845 74.925 217.125 75.805 ;
    RECT 180.325 74.925 180.605 75.805 ;
    RECT 177.005 74.925 177.285 75.805 ;
    RECT 173.685 74.925 173.965 75.805 ;
    RECT 170.365 74.925 170.645 75.805 ;
    RECT 167.045 74.925 167.325 75.805 ;
    RECT 163.725 74.925 164.005 75.805 ;
    RECT 160.405 74.925 160.685 75.805 ;
    RECT 157.085 74.925 157.365 75.805 ;
    RECT 153.765 74.925 154.045 75.805 ;
    RECT 150.445 74.925 150.725 75.805 ;
    RECT 213.525 74.925 213.805 75.805 ;
    RECT 210.205 74.925 210.485 75.805 ;
    RECT 206.885 74.925 207.165 75.805 ;
    RECT 203.565 74.925 203.845 75.805 ;
    RECT 200.245 74.925 200.525 75.805 ;
    RECT 196.925 74.925 197.205 75.805 ;
    RECT 193.605 74.925 193.885 75.805 ;
    RECT 190.285 74.925 190.565 75.805 ;
    RECT 186.965 74.925 187.245 75.805 ;
    RECT 183.645 74.925 183.925 75.805 ;
    RECT 266.645 74.925 266.925 75.805 ;
    RECT 263.325 74.925 263.605 75.805 ;
    RECT 260.005 74.925 260.285 75.805 ;
    RECT 256.685 74.925 256.965 75.805 ;
    RECT 253.365 74.925 253.645 75.805 ;
    RECT 250.045 74.205 250.325 75.085 ;
    RECT 246.725 74.205 247.005 75.085 ;
    RECT 243.405 74.205 243.685 75.085 ;
    RECT 240.085 74.205 240.365 75.085 ;
    RECT 236.765 74.205 237.045 75.085 ;
    RECT 233.445 74.205 233.725 75.085 ;
    RECT 230.125 74.205 230.405 75.085 ;
    RECT 226.805 74.205 227.085 75.085 ;
    RECT 223.485 74.205 223.765 75.085 ;
    RECT 220.165 74.205 220.445 75.085 ;
    RECT 216.845 74.205 217.125 75.085 ;
    RECT 180.325 74.205 180.605 75.085 ;
    RECT 177.005 74.205 177.285 75.085 ;
    RECT 173.685 74.205 173.965 75.085 ;
    RECT 170.365 74.205 170.645 75.085 ;
    RECT 167.045 74.205 167.325 75.085 ;
    RECT 163.725 74.205 164.005 75.085 ;
    RECT 160.405 74.205 160.685 75.085 ;
    RECT 157.085 74.205 157.365 75.085 ;
    RECT 153.765 74.205 154.045 75.085 ;
    RECT 150.445 74.205 150.725 75.085 ;
    RECT 213.525 74.205 213.805 75.085 ;
    RECT 210.205 74.205 210.485 75.085 ;
    RECT 206.885 74.205 207.165 75.085 ;
    RECT 203.565 74.205 203.845 75.085 ;
    RECT 200.245 74.205 200.525 75.085 ;
    RECT 196.925 74.205 197.205 75.085 ;
    RECT 193.605 74.205 193.885 75.085 ;
    RECT 190.285 74.205 190.565 75.085 ;
    RECT 186.965 74.205 187.245 75.085 ;
    RECT 183.645 74.205 183.925 75.085 ;
    RECT 266.645 74.205 266.925 75.085 ;
    RECT 263.325 74.205 263.605 75.085 ;
    RECT 260.005 74.205 260.285 75.085 ;
    RECT 256.685 74.205 256.965 75.085 ;
    RECT 253.365 74.205 253.645 75.085 ;
    RECT 250.045 73.485 250.325 74.365 ;
    RECT 246.725 73.485 247.005 74.365 ;
    RECT 243.405 73.485 243.685 74.365 ;
    RECT 240.085 73.485 240.365 74.365 ;
    RECT 236.765 73.485 237.045 74.365 ;
    RECT 233.445 73.485 233.725 74.365 ;
    RECT 230.125 73.485 230.405 74.365 ;
    RECT 226.805 73.485 227.085 74.365 ;
    RECT 223.485 73.485 223.765 74.365 ;
    RECT 220.165 73.485 220.445 74.365 ;
    RECT 216.845 73.485 217.125 74.365 ;
    RECT 180.325 73.485 180.605 74.365 ;
    RECT 177.005 73.485 177.285 74.365 ;
    RECT 173.685 73.485 173.965 74.365 ;
    RECT 170.365 73.485 170.645 74.365 ;
    RECT 167.045 73.485 167.325 74.365 ;
    RECT 163.725 73.485 164.005 74.365 ;
    RECT 160.405 73.485 160.685 74.365 ;
    RECT 157.085 73.485 157.365 74.365 ;
    RECT 153.765 73.485 154.045 74.365 ;
    RECT 150.445 73.485 150.725 74.365 ;
    RECT 213.525 73.485 213.805 74.365 ;
    RECT 210.205 73.485 210.485 74.365 ;
    RECT 206.885 73.485 207.165 74.365 ;
    RECT 203.565 73.485 203.845 74.365 ;
    RECT 200.245 73.485 200.525 74.365 ;
    RECT 196.925 73.485 197.205 74.365 ;
    RECT 193.605 73.485 193.885 74.365 ;
    RECT 190.285 73.485 190.565 74.365 ;
    RECT 186.965 73.485 187.245 74.365 ;
    RECT 183.645 73.485 183.925 74.365 ;
    RECT 266.645 73.485 266.925 74.365 ;
    RECT 263.325 73.485 263.605 74.365 ;
    RECT 260.005 73.485 260.285 74.365 ;
    RECT 256.685 73.485 256.965 74.365 ;
    RECT 253.365 73.485 253.645 74.365 ;
    RECT 250.045 72.765 250.325 73.645 ;
    RECT 246.725 72.765 247.005 73.645 ;
    RECT 243.405 72.765 243.685 73.645 ;
    RECT 240.085 72.765 240.365 73.645 ;
    RECT 236.765 72.765 237.045 73.645 ;
    RECT 233.445 72.765 233.725 73.645 ;
    RECT 230.125 72.765 230.405 73.645 ;
    RECT 226.805 72.765 227.085 73.645 ;
    RECT 223.485 72.765 223.765 73.645 ;
    RECT 220.165 72.765 220.445 73.645 ;
    RECT 216.845 72.765 217.125 73.645 ;
    RECT 180.325 72.765 180.605 73.645 ;
    RECT 177.005 72.765 177.285 73.645 ;
    RECT 173.685 72.765 173.965 73.645 ;
    RECT 170.365 72.765 170.645 73.645 ;
    RECT 167.045 72.765 167.325 73.645 ;
    RECT 163.725 72.765 164.005 73.645 ;
    RECT 160.405 72.765 160.685 73.645 ;
    RECT 157.085 72.765 157.365 73.645 ;
    RECT 153.765 72.765 154.045 73.645 ;
    RECT 150.445 72.765 150.725 73.645 ;
    RECT 213.525 72.765 213.805 73.645 ;
    RECT 210.205 72.765 210.485 73.645 ;
    RECT 206.885 72.765 207.165 73.645 ;
    RECT 203.565 72.765 203.845 73.645 ;
    RECT 200.245 72.765 200.525 73.645 ;
    RECT 196.925 72.765 197.205 73.645 ;
    RECT 193.605 72.765 193.885 73.645 ;
    RECT 190.285 72.765 190.565 73.645 ;
    RECT 186.965 72.765 187.245 73.645 ;
    RECT 183.645 72.765 183.925 73.645 ;
    RECT 266.645 72.765 266.925 73.645 ;
    RECT 263.325 72.765 263.605 73.645 ;
    RECT 260.005 72.765 260.285 73.645 ;
    RECT 256.685 72.765 256.965 73.645 ;
    RECT 253.365 72.765 253.645 73.645 ;
    RECT 250.045 20.905 250.325 21.785 ;
    RECT 246.725 20.905 247.005 21.785 ;
    RECT 243.405 20.905 243.685 21.785 ;
    RECT 240.085 20.905 240.365 21.785 ;
    RECT 236.765 20.905 237.045 21.785 ;
    RECT 233.445 20.905 233.725 21.785 ;
    RECT 230.125 20.905 230.405 21.785 ;
    RECT 226.805 20.905 227.085 21.785 ;
    RECT 223.485 20.905 223.765 21.785 ;
    RECT 220.165 20.905 220.445 21.785 ;
    RECT 216.845 20.905 217.125 21.785 ;
    RECT 180.325 20.905 180.605 21.785 ;
    RECT 177.005 20.905 177.285 21.785 ;
    RECT 173.685 20.905 173.965 21.785 ;
    RECT 170.365 20.905 170.645 21.785 ;
    RECT 167.045 20.905 167.325 21.785 ;
    RECT 163.725 20.905 164.005 21.785 ;
    RECT 160.405 20.905 160.685 21.785 ;
    RECT 157.085 20.905 157.365 21.785 ;
    RECT 153.765 20.905 154.045 21.785 ;
    RECT 150.445 20.905 150.725 21.785 ;
    RECT 213.525 20.905 213.805 21.785 ;
    RECT 210.205 20.905 210.485 21.785 ;
    RECT 206.885 20.905 207.165 21.785 ;
    RECT 203.565 20.905 203.845 21.785 ;
    RECT 200.245 20.905 200.525 21.785 ;
    RECT 196.925 20.905 197.205 21.785 ;
    RECT 193.605 20.905 193.885 21.785 ;
    RECT 190.285 20.905 190.565 21.785 ;
    RECT 186.965 20.905 187.245 21.785 ;
    RECT 183.645 20.905 183.925 21.785 ;
    RECT 266.645 20.905 266.925 21.785 ;
    RECT 263.325 20.905 263.605 21.785 ;
    RECT 260.005 20.905 260.285 21.785 ;
    RECT 256.685 20.905 256.965 21.785 ;
    RECT 253.365 20.905 253.645 21.785 ;
    RECT 250.045 20.185 250.325 21.065 ;
    RECT 246.725 20.185 247.005 21.065 ;
    RECT 243.405 20.185 243.685 21.065 ;
    RECT 240.085 20.185 240.365 21.065 ;
    RECT 236.765 20.185 237.045 21.065 ;
    RECT 233.445 20.185 233.725 21.065 ;
    RECT 230.125 20.185 230.405 21.065 ;
    RECT 226.805 20.185 227.085 21.065 ;
    RECT 223.485 20.185 223.765 21.065 ;
    RECT 220.165 20.185 220.445 21.065 ;
    RECT 216.845 20.185 217.125 21.065 ;
    RECT 180.325 20.185 180.605 21.065 ;
    RECT 177.005 20.185 177.285 21.065 ;
    RECT 173.685 20.185 173.965 21.065 ;
    RECT 170.365 20.185 170.645 21.065 ;
    RECT 167.045 20.185 167.325 21.065 ;
    RECT 163.725 20.185 164.005 21.065 ;
    RECT 160.405 20.185 160.685 21.065 ;
    RECT 157.085 20.185 157.365 21.065 ;
    RECT 153.765 20.185 154.045 21.065 ;
    RECT 150.445 20.185 150.725 21.065 ;
    RECT 213.525 20.185 213.805 21.065 ;
    RECT 210.205 20.185 210.485 21.065 ;
    RECT 206.885 20.185 207.165 21.065 ;
    RECT 203.565 20.185 203.845 21.065 ;
    RECT 200.245 20.185 200.525 21.065 ;
    RECT 196.925 20.185 197.205 21.065 ;
    RECT 193.605 20.185 193.885 21.065 ;
    RECT 190.285 20.185 190.565 21.065 ;
    RECT 186.965 20.185 187.245 21.065 ;
    RECT 183.645 20.185 183.925 21.065 ;
    RECT 266.645 20.185 266.925 21.065 ;
    RECT 263.325 20.185 263.605 21.065 ;
    RECT 260.005 20.185 260.285 21.065 ;
    RECT 256.685 20.185 256.965 21.065 ;
    RECT 253.365 20.185 253.645 21.065 ;
    RECT 250.045 19.465 250.325 20.345 ;
    RECT 246.725 19.465 247.005 20.345 ;
    RECT 243.405 19.465 243.685 20.345 ;
    RECT 240.085 19.465 240.365 20.345 ;
    RECT 236.765 19.465 237.045 20.345 ;
    RECT 233.445 19.465 233.725 20.345 ;
    RECT 230.125 19.465 230.405 20.345 ;
    RECT 226.805 19.465 227.085 20.345 ;
    RECT 223.485 19.465 223.765 20.345 ;
    RECT 220.165 19.465 220.445 20.345 ;
    RECT 216.845 19.465 217.125 20.345 ;
    RECT 180.325 19.465 180.605 20.345 ;
    RECT 177.005 19.465 177.285 20.345 ;
    RECT 173.685 19.465 173.965 20.345 ;
    RECT 170.365 19.465 170.645 20.345 ;
    RECT 167.045 19.465 167.325 20.345 ;
    RECT 163.725 19.465 164.005 20.345 ;
    RECT 160.405 19.465 160.685 20.345 ;
    RECT 157.085 19.465 157.365 20.345 ;
    RECT 153.765 19.465 154.045 20.345 ;
    RECT 150.445 19.465 150.725 20.345 ;
    RECT 213.525 19.465 213.805 20.345 ;
    RECT 210.205 19.465 210.485 20.345 ;
    RECT 206.885 19.465 207.165 20.345 ;
    RECT 203.565 19.465 203.845 20.345 ;
    RECT 200.245 19.465 200.525 20.345 ;
    RECT 196.925 19.465 197.205 20.345 ;
    RECT 193.605 19.465 193.885 20.345 ;
    RECT 190.285 19.465 190.565 20.345 ;
    RECT 186.965 19.465 187.245 20.345 ;
    RECT 183.645 19.465 183.925 20.345 ;
    RECT 266.645 19.465 266.925 20.345 ;
    RECT 263.325 19.465 263.605 20.345 ;
    RECT 260.005 19.465 260.285 20.345 ;
    RECT 256.685 19.465 256.965 20.345 ;
    RECT 253.365 19.465 253.645 20.345 ;
    RECT 250.045 35.305 250.325 36.185 ;
    RECT 246.725 35.305 247.005 36.185 ;
    RECT 243.405 35.305 243.685 36.185 ;
    RECT 240.085 35.305 240.365 36.185 ;
    RECT 236.765 35.305 237.045 36.185 ;
    RECT 233.445 35.305 233.725 36.185 ;
    RECT 230.125 35.305 230.405 36.185 ;
    RECT 226.805 35.305 227.085 36.185 ;
    RECT 223.485 35.305 223.765 36.185 ;
    RECT 220.165 35.305 220.445 36.185 ;
    RECT 216.845 35.305 217.125 36.185 ;
    RECT 180.325 35.305 180.605 36.185 ;
    RECT 177.005 35.305 177.285 36.185 ;
    RECT 173.685 35.305 173.965 36.185 ;
    RECT 170.365 35.305 170.645 36.185 ;
    RECT 167.045 35.305 167.325 36.185 ;
    RECT 163.725 35.305 164.005 36.185 ;
    RECT 160.405 35.305 160.685 36.185 ;
    RECT 157.085 35.305 157.365 36.185 ;
    RECT 153.765 35.305 154.045 36.185 ;
    RECT 150.445 35.305 150.725 36.185 ;
    RECT 213.525 35.305 213.805 36.185 ;
    RECT 210.205 35.305 210.485 36.185 ;
    RECT 206.885 35.305 207.165 36.185 ;
    RECT 203.565 35.305 203.845 36.185 ;
    RECT 200.245 35.305 200.525 36.185 ;
    RECT 196.925 35.305 197.205 36.185 ;
    RECT 193.605 35.305 193.885 36.185 ;
    RECT 190.285 35.305 190.565 36.185 ;
    RECT 186.965 35.305 187.245 36.185 ;
    RECT 183.645 35.305 183.925 36.185 ;
    RECT 266.645 35.305 266.925 36.185 ;
    RECT 263.325 35.305 263.605 36.185 ;
    RECT 260.005 35.305 260.285 36.185 ;
    RECT 256.685 35.305 256.965 36.185 ;
    RECT 253.365 35.305 253.645 36.185 ;
    RECT 250.045 18.745 250.325 19.625 ;
    RECT 246.725 18.745 247.005 19.625 ;
    RECT 243.405 18.745 243.685 19.625 ;
    RECT 240.085 18.745 240.365 19.625 ;
    RECT 236.765 18.745 237.045 19.625 ;
    RECT 233.445 18.745 233.725 19.625 ;
    RECT 230.125 18.745 230.405 19.625 ;
    RECT 226.805 18.745 227.085 19.625 ;
    RECT 223.485 18.745 223.765 19.625 ;
    RECT 220.165 18.745 220.445 19.625 ;
    RECT 216.845 18.745 217.125 19.625 ;
    RECT 180.325 18.745 180.605 19.625 ;
    RECT 177.005 18.745 177.285 19.625 ;
    RECT 173.685 18.745 173.965 19.625 ;
    RECT 170.365 18.745 170.645 19.625 ;
    RECT 167.045 18.745 167.325 19.625 ;
    RECT 163.725 18.745 164.005 19.625 ;
    RECT 160.405 18.745 160.685 19.625 ;
    RECT 157.085 18.745 157.365 19.625 ;
    RECT 153.765 18.745 154.045 19.625 ;
    RECT 150.445 18.745 150.725 19.625 ;
    RECT 213.525 18.745 213.805 19.625 ;
    RECT 210.205 18.745 210.485 19.625 ;
    RECT 206.885 18.745 207.165 19.625 ;
    RECT 203.565 18.745 203.845 19.625 ;
    RECT 200.245 18.745 200.525 19.625 ;
    RECT 196.925 18.745 197.205 19.625 ;
    RECT 193.605 18.745 193.885 19.625 ;
    RECT 190.285 18.745 190.565 19.625 ;
    RECT 186.965 18.745 187.245 19.625 ;
    RECT 183.645 18.745 183.925 19.625 ;
    RECT 266.645 18.745 266.925 19.625 ;
    RECT 263.325 18.745 263.605 19.625 ;
    RECT 260.005 18.745 260.285 19.625 ;
    RECT 256.685 18.745 256.965 19.625 ;
    RECT 253.365 18.745 253.645 19.625 ;
    RECT 250.045 34.585 250.325 35.465 ;
    RECT 246.725 34.585 247.005 35.465 ;
    RECT 243.405 34.585 243.685 35.465 ;
    RECT 240.085 34.585 240.365 35.465 ;
    RECT 236.765 34.585 237.045 35.465 ;
    RECT 233.445 34.585 233.725 35.465 ;
    RECT 230.125 34.585 230.405 35.465 ;
    RECT 226.805 34.585 227.085 35.465 ;
    RECT 223.485 34.585 223.765 35.465 ;
    RECT 220.165 34.585 220.445 35.465 ;
    RECT 216.845 34.585 217.125 35.465 ;
    RECT 180.325 34.585 180.605 35.465 ;
    RECT 177.005 34.585 177.285 35.465 ;
    RECT 173.685 34.585 173.965 35.465 ;
    RECT 170.365 34.585 170.645 35.465 ;
    RECT 167.045 34.585 167.325 35.465 ;
    RECT 163.725 34.585 164.005 35.465 ;
    RECT 160.405 34.585 160.685 35.465 ;
    RECT 157.085 34.585 157.365 35.465 ;
    RECT 153.765 34.585 154.045 35.465 ;
    RECT 150.445 34.585 150.725 35.465 ;
    RECT 213.525 34.585 213.805 35.465 ;
    RECT 210.205 34.585 210.485 35.465 ;
    RECT 206.885 34.585 207.165 35.465 ;
    RECT 203.565 34.585 203.845 35.465 ;
    RECT 200.245 34.585 200.525 35.465 ;
    RECT 196.925 34.585 197.205 35.465 ;
    RECT 193.605 34.585 193.885 35.465 ;
    RECT 190.285 34.585 190.565 35.465 ;
    RECT 186.965 34.585 187.245 35.465 ;
    RECT 183.645 34.585 183.925 35.465 ;
    RECT 266.645 34.585 266.925 35.465 ;
    RECT 263.325 34.585 263.605 35.465 ;
    RECT 260.005 34.585 260.285 35.465 ;
    RECT 256.685 34.585 256.965 35.465 ;
    RECT 253.365 34.585 253.645 35.465 ;
    RECT 250.045 18.025 250.325 18.905 ;
    RECT 246.725 18.025 247.005 18.905 ;
    RECT 243.405 18.025 243.685 18.905 ;
    RECT 240.085 18.025 240.365 18.905 ;
    RECT 236.765 18.025 237.045 18.905 ;
    RECT 233.445 18.025 233.725 18.905 ;
    RECT 230.125 18.025 230.405 18.905 ;
    RECT 226.805 18.025 227.085 18.905 ;
    RECT 223.485 18.025 223.765 18.905 ;
    RECT 220.165 18.025 220.445 18.905 ;
    RECT 216.845 18.025 217.125 18.905 ;
    RECT 180.325 18.025 180.605 18.905 ;
    RECT 177.005 18.025 177.285 18.905 ;
    RECT 173.685 18.025 173.965 18.905 ;
    RECT 170.365 18.025 170.645 18.905 ;
    RECT 167.045 18.025 167.325 18.905 ;
    RECT 163.725 18.025 164.005 18.905 ;
    RECT 160.405 18.025 160.685 18.905 ;
    RECT 157.085 18.025 157.365 18.905 ;
    RECT 153.765 18.025 154.045 18.905 ;
    RECT 150.445 18.025 150.725 18.905 ;
    RECT 213.525 18.025 213.805 18.905 ;
    RECT 210.205 18.025 210.485 18.905 ;
    RECT 206.885 18.025 207.165 18.905 ;
    RECT 203.565 18.025 203.845 18.905 ;
    RECT 200.245 18.025 200.525 18.905 ;
    RECT 196.925 18.025 197.205 18.905 ;
    RECT 193.605 18.025 193.885 18.905 ;
    RECT 190.285 18.025 190.565 18.905 ;
    RECT 186.965 18.025 187.245 18.905 ;
    RECT 183.645 18.025 183.925 18.905 ;
    RECT 266.645 18.025 266.925 18.905 ;
    RECT 263.325 18.025 263.605 18.905 ;
    RECT 260.005 18.025 260.285 18.905 ;
    RECT 256.685 18.025 256.965 18.905 ;
    RECT 253.365 18.025 253.645 18.905 ;
    RECT 250.045 33.865 250.325 34.745 ;
    RECT 246.725 33.865 247.005 34.745 ;
    RECT 243.405 33.865 243.685 34.745 ;
    RECT 240.085 33.865 240.365 34.745 ;
    RECT 236.765 33.865 237.045 34.745 ;
    RECT 233.445 33.865 233.725 34.745 ;
    RECT 230.125 33.865 230.405 34.745 ;
    RECT 226.805 33.865 227.085 34.745 ;
    RECT 223.485 33.865 223.765 34.745 ;
    RECT 220.165 33.865 220.445 34.745 ;
    RECT 216.845 33.865 217.125 34.745 ;
    RECT 180.325 33.865 180.605 34.745 ;
    RECT 177.005 33.865 177.285 34.745 ;
    RECT 173.685 33.865 173.965 34.745 ;
    RECT 170.365 33.865 170.645 34.745 ;
    RECT 167.045 33.865 167.325 34.745 ;
    RECT 163.725 33.865 164.005 34.745 ;
    RECT 160.405 33.865 160.685 34.745 ;
    RECT 157.085 33.865 157.365 34.745 ;
    RECT 153.765 33.865 154.045 34.745 ;
    RECT 150.445 33.865 150.725 34.745 ;
    RECT 213.525 33.865 213.805 34.745 ;
    RECT 210.205 33.865 210.485 34.745 ;
    RECT 206.885 33.865 207.165 34.745 ;
    RECT 203.565 33.865 203.845 34.745 ;
    RECT 200.245 33.865 200.525 34.745 ;
    RECT 196.925 33.865 197.205 34.745 ;
    RECT 193.605 33.865 193.885 34.745 ;
    RECT 190.285 33.865 190.565 34.745 ;
    RECT 186.965 33.865 187.245 34.745 ;
    RECT 183.645 33.865 183.925 34.745 ;
    RECT 266.645 33.865 266.925 34.745 ;
    RECT 263.325 33.865 263.605 34.745 ;
    RECT 260.005 33.865 260.285 34.745 ;
    RECT 256.685 33.865 256.965 34.745 ;
    RECT 253.365 33.865 253.645 34.745 ;
    RECT 250.045 17.305 250.325 18.185 ;
    RECT 246.725 17.305 247.005 18.185 ;
    RECT 243.405 17.305 243.685 18.185 ;
    RECT 240.085 17.305 240.365 18.185 ;
    RECT 236.765 17.305 237.045 18.185 ;
    RECT 233.445 17.305 233.725 18.185 ;
    RECT 230.125 17.305 230.405 18.185 ;
    RECT 226.805 17.305 227.085 18.185 ;
    RECT 223.485 17.305 223.765 18.185 ;
    RECT 220.165 17.305 220.445 18.185 ;
    RECT 216.845 17.305 217.125 18.185 ;
    RECT 180.325 17.305 180.605 18.185 ;
    RECT 177.005 17.305 177.285 18.185 ;
    RECT 173.685 17.305 173.965 18.185 ;
    RECT 170.365 17.305 170.645 18.185 ;
    RECT 167.045 17.305 167.325 18.185 ;
    RECT 163.725 17.305 164.005 18.185 ;
    RECT 160.405 17.305 160.685 18.185 ;
    RECT 157.085 17.305 157.365 18.185 ;
    RECT 153.765 17.305 154.045 18.185 ;
    RECT 150.445 17.305 150.725 18.185 ;
    RECT 213.525 17.305 213.805 18.185 ;
    RECT 210.205 17.305 210.485 18.185 ;
    RECT 206.885 17.305 207.165 18.185 ;
    RECT 203.565 17.305 203.845 18.185 ;
    RECT 200.245 17.305 200.525 18.185 ;
    RECT 196.925 17.305 197.205 18.185 ;
    RECT 193.605 17.305 193.885 18.185 ;
    RECT 190.285 17.305 190.565 18.185 ;
    RECT 186.965 17.305 187.245 18.185 ;
    RECT 183.645 17.305 183.925 18.185 ;
    RECT 266.645 17.305 266.925 18.185 ;
    RECT 263.325 17.305 263.605 18.185 ;
    RECT 260.005 17.305 260.285 18.185 ;
    RECT 256.685 17.305 256.965 18.185 ;
    RECT 253.365 17.305 253.645 18.185 ;
    RECT 250.045 33.145 250.325 34.025 ;
    RECT 246.725 33.145 247.005 34.025 ;
    RECT 243.405 33.145 243.685 34.025 ;
    RECT 240.085 33.145 240.365 34.025 ;
    RECT 236.765 33.145 237.045 34.025 ;
    RECT 233.445 33.145 233.725 34.025 ;
    RECT 230.125 33.145 230.405 34.025 ;
    RECT 226.805 33.145 227.085 34.025 ;
    RECT 223.485 33.145 223.765 34.025 ;
    RECT 220.165 33.145 220.445 34.025 ;
    RECT 216.845 33.145 217.125 34.025 ;
    RECT 180.325 33.145 180.605 34.025 ;
    RECT 177.005 33.145 177.285 34.025 ;
    RECT 173.685 33.145 173.965 34.025 ;
    RECT 170.365 33.145 170.645 34.025 ;
    RECT 167.045 33.145 167.325 34.025 ;
    RECT 163.725 33.145 164.005 34.025 ;
    RECT 160.405 33.145 160.685 34.025 ;
    RECT 157.085 33.145 157.365 34.025 ;
    RECT 153.765 33.145 154.045 34.025 ;
    RECT 150.445 33.145 150.725 34.025 ;
    RECT 213.525 33.145 213.805 34.025 ;
    RECT 210.205 33.145 210.485 34.025 ;
    RECT 206.885 33.145 207.165 34.025 ;
    RECT 203.565 33.145 203.845 34.025 ;
    RECT 200.245 33.145 200.525 34.025 ;
    RECT 196.925 33.145 197.205 34.025 ;
    RECT 193.605 33.145 193.885 34.025 ;
    RECT 190.285 33.145 190.565 34.025 ;
    RECT 186.965 33.145 187.245 34.025 ;
    RECT 183.645 33.145 183.925 34.025 ;
    RECT 266.645 33.145 266.925 34.025 ;
    RECT 263.325 33.145 263.605 34.025 ;
    RECT 260.005 33.145 260.285 34.025 ;
    RECT 256.685 33.145 256.965 34.025 ;
    RECT 253.365 33.145 253.645 34.025 ;
    RECT 250.045 16.585 250.325 17.465 ;
    RECT 246.725 16.585 247.005 17.465 ;
    RECT 243.405 16.585 243.685 17.465 ;
    RECT 240.085 16.585 240.365 17.465 ;
    RECT 236.765 16.585 237.045 17.465 ;
    RECT 233.445 16.585 233.725 17.465 ;
    RECT 230.125 16.585 230.405 17.465 ;
    RECT 226.805 16.585 227.085 17.465 ;
    RECT 223.485 16.585 223.765 17.465 ;
    RECT 220.165 16.585 220.445 17.465 ;
    RECT 216.845 16.585 217.125 17.465 ;
    RECT 180.325 16.585 180.605 17.465 ;
    RECT 177.005 16.585 177.285 17.465 ;
    RECT 173.685 16.585 173.965 17.465 ;
    RECT 170.365 16.585 170.645 17.465 ;
    RECT 167.045 16.585 167.325 17.465 ;
    RECT 163.725 16.585 164.005 17.465 ;
    RECT 160.405 16.585 160.685 17.465 ;
    RECT 157.085 16.585 157.365 17.465 ;
    RECT 153.765 16.585 154.045 17.465 ;
    RECT 150.445 16.585 150.725 17.465 ;
    RECT 213.525 16.585 213.805 17.465 ;
    RECT 210.205 16.585 210.485 17.465 ;
    RECT 206.885 16.585 207.165 17.465 ;
    RECT 203.565 16.585 203.845 17.465 ;
    RECT 200.245 16.585 200.525 17.465 ;
    RECT 196.925 16.585 197.205 17.465 ;
    RECT 193.605 16.585 193.885 17.465 ;
    RECT 190.285 16.585 190.565 17.465 ;
    RECT 186.965 16.585 187.245 17.465 ;
    RECT 183.645 16.585 183.925 17.465 ;
    RECT 266.645 16.585 266.925 17.465 ;
    RECT 263.325 16.585 263.605 17.465 ;
    RECT 260.005 16.585 260.285 17.465 ;
    RECT 256.685 16.585 256.965 17.465 ;
    RECT 253.365 16.585 253.645 17.465 ;
    RECT 250.045 32.425 250.325 33.305 ;
    RECT 246.725 32.425 247.005 33.305 ;
    RECT 243.405 32.425 243.685 33.305 ;
    RECT 240.085 32.425 240.365 33.305 ;
    RECT 236.765 32.425 237.045 33.305 ;
    RECT 233.445 32.425 233.725 33.305 ;
    RECT 230.125 32.425 230.405 33.305 ;
    RECT 226.805 32.425 227.085 33.305 ;
    RECT 223.485 32.425 223.765 33.305 ;
    RECT 220.165 32.425 220.445 33.305 ;
    RECT 216.845 32.425 217.125 33.305 ;
    RECT 180.325 32.425 180.605 33.305 ;
    RECT 177.005 32.425 177.285 33.305 ;
    RECT 173.685 32.425 173.965 33.305 ;
    RECT 170.365 32.425 170.645 33.305 ;
    RECT 167.045 32.425 167.325 33.305 ;
    RECT 163.725 32.425 164.005 33.305 ;
    RECT 160.405 32.425 160.685 33.305 ;
    RECT 157.085 32.425 157.365 33.305 ;
    RECT 153.765 32.425 154.045 33.305 ;
    RECT 150.445 32.425 150.725 33.305 ;
    RECT 213.525 32.425 213.805 33.305 ;
    RECT 210.205 32.425 210.485 33.305 ;
    RECT 206.885 32.425 207.165 33.305 ;
    RECT 203.565 32.425 203.845 33.305 ;
    RECT 200.245 32.425 200.525 33.305 ;
    RECT 196.925 32.425 197.205 33.305 ;
    RECT 193.605 32.425 193.885 33.305 ;
    RECT 190.285 32.425 190.565 33.305 ;
    RECT 186.965 32.425 187.245 33.305 ;
    RECT 183.645 32.425 183.925 33.305 ;
    RECT 266.645 32.425 266.925 33.305 ;
    RECT 263.325 32.425 263.605 33.305 ;
    RECT 260.005 32.425 260.285 33.305 ;
    RECT 256.685 32.425 256.965 33.305 ;
    RECT 253.365 32.425 253.645 33.305 ;
    RECT 250.045 72.045 250.325 72.925 ;
    RECT 246.725 72.045 247.005 72.925 ;
    RECT 243.405 72.045 243.685 72.925 ;
    RECT 240.085 72.045 240.365 72.925 ;
    RECT 236.765 72.045 237.045 72.925 ;
    RECT 233.445 72.045 233.725 72.925 ;
    RECT 230.125 72.045 230.405 72.925 ;
    RECT 226.805 72.045 227.085 72.925 ;
    RECT 223.485 72.045 223.765 72.925 ;
    RECT 220.165 72.045 220.445 72.925 ;
    RECT 216.845 72.045 217.125 72.925 ;
    RECT 180.325 72.045 180.605 72.925 ;
    RECT 177.005 72.045 177.285 72.925 ;
    RECT 173.685 72.045 173.965 72.925 ;
    RECT 170.365 72.045 170.645 72.925 ;
    RECT 167.045 72.045 167.325 72.925 ;
    RECT 163.725 72.045 164.005 72.925 ;
    RECT 160.405 72.045 160.685 72.925 ;
    RECT 157.085 72.045 157.365 72.925 ;
    RECT 153.765 72.045 154.045 72.925 ;
    RECT 150.445 72.045 150.725 72.925 ;
    RECT 213.525 72.045 213.805 72.925 ;
    RECT 210.205 72.045 210.485 72.925 ;
    RECT 206.885 72.045 207.165 72.925 ;
    RECT 203.565 72.045 203.845 72.925 ;
    RECT 200.245 72.045 200.525 72.925 ;
    RECT 196.925 72.045 197.205 72.925 ;
    RECT 193.605 72.045 193.885 72.925 ;
    RECT 190.285 72.045 190.565 72.925 ;
    RECT 186.965 72.045 187.245 72.925 ;
    RECT 183.645 72.045 183.925 72.925 ;
    RECT 266.645 72.045 266.925 72.925 ;
    RECT 263.325 72.045 263.605 72.925 ;
    RECT 260.005 72.045 260.285 72.925 ;
    RECT 256.685 72.045 256.965 72.925 ;
    RECT 253.365 72.045 253.645 72.925 ;
    RECT 250.045 15.865 250.325 16.745 ;
    RECT 246.725 15.865 247.005 16.745 ;
    RECT 243.405 15.865 243.685 16.745 ;
    RECT 240.085 15.865 240.365 16.745 ;
    RECT 236.765 15.865 237.045 16.745 ;
    RECT 233.445 15.865 233.725 16.745 ;
    RECT 230.125 15.865 230.405 16.745 ;
    RECT 226.805 15.865 227.085 16.745 ;
    RECT 223.485 15.865 223.765 16.745 ;
    RECT 220.165 15.865 220.445 16.745 ;
    RECT 216.845 15.865 217.125 16.745 ;
    RECT 180.325 15.865 180.605 16.745 ;
    RECT 177.005 15.865 177.285 16.745 ;
    RECT 173.685 15.865 173.965 16.745 ;
    RECT 170.365 15.865 170.645 16.745 ;
    RECT 167.045 15.865 167.325 16.745 ;
    RECT 163.725 15.865 164.005 16.745 ;
    RECT 160.405 15.865 160.685 16.745 ;
    RECT 157.085 15.865 157.365 16.745 ;
    RECT 153.765 15.865 154.045 16.745 ;
    RECT 150.445 15.865 150.725 16.745 ;
    RECT 213.525 15.865 213.805 16.745 ;
    RECT 210.205 15.865 210.485 16.745 ;
    RECT 206.885 15.865 207.165 16.745 ;
    RECT 203.565 15.865 203.845 16.745 ;
    RECT 200.245 15.865 200.525 16.745 ;
    RECT 196.925 15.865 197.205 16.745 ;
    RECT 193.605 15.865 193.885 16.745 ;
    RECT 190.285 15.865 190.565 16.745 ;
    RECT 186.965 15.865 187.245 16.745 ;
    RECT 183.645 15.865 183.925 16.745 ;
    RECT 266.645 15.865 266.925 16.745 ;
    RECT 263.325 15.865 263.605 16.745 ;
    RECT 260.005 15.865 260.285 16.745 ;
    RECT 256.685 15.865 256.965 16.745 ;
    RECT 253.365 15.865 253.645 16.745 ;
    RECT 250.045 31.705 250.325 32.585 ;
    RECT 246.725 31.705 247.005 32.585 ;
    RECT 243.405 31.705 243.685 32.585 ;
    RECT 240.085 31.705 240.365 32.585 ;
    RECT 236.765 31.705 237.045 32.585 ;
    RECT 233.445 31.705 233.725 32.585 ;
    RECT 230.125 31.705 230.405 32.585 ;
    RECT 226.805 31.705 227.085 32.585 ;
    RECT 223.485 31.705 223.765 32.585 ;
    RECT 220.165 31.705 220.445 32.585 ;
    RECT 216.845 31.705 217.125 32.585 ;
    RECT 180.325 31.705 180.605 32.585 ;
    RECT 177.005 31.705 177.285 32.585 ;
    RECT 173.685 31.705 173.965 32.585 ;
    RECT 170.365 31.705 170.645 32.585 ;
    RECT 167.045 31.705 167.325 32.585 ;
    RECT 163.725 31.705 164.005 32.585 ;
    RECT 160.405 31.705 160.685 32.585 ;
    RECT 157.085 31.705 157.365 32.585 ;
    RECT 153.765 31.705 154.045 32.585 ;
    RECT 150.445 31.705 150.725 32.585 ;
    RECT 213.525 31.705 213.805 32.585 ;
    RECT 210.205 31.705 210.485 32.585 ;
    RECT 206.885 31.705 207.165 32.585 ;
    RECT 203.565 31.705 203.845 32.585 ;
    RECT 200.245 31.705 200.525 32.585 ;
    RECT 196.925 31.705 197.205 32.585 ;
    RECT 193.605 31.705 193.885 32.585 ;
    RECT 190.285 31.705 190.565 32.585 ;
    RECT 186.965 31.705 187.245 32.585 ;
    RECT 183.645 31.705 183.925 32.585 ;
    RECT 266.645 31.705 266.925 32.585 ;
    RECT 263.325 31.705 263.605 32.585 ;
    RECT 260.005 31.705 260.285 32.585 ;
    RECT 256.685 31.705 256.965 32.585 ;
    RECT 253.365 31.705 253.645 32.585 ;
    RECT 250.045 71.325 250.325 72.205 ;
    RECT 246.725 71.325 247.005 72.205 ;
    RECT 243.405 71.325 243.685 72.205 ;
    RECT 240.085 71.325 240.365 72.205 ;
    RECT 236.765 71.325 237.045 72.205 ;
    RECT 233.445 71.325 233.725 72.205 ;
    RECT 230.125 71.325 230.405 72.205 ;
    RECT 226.805 71.325 227.085 72.205 ;
    RECT 223.485 71.325 223.765 72.205 ;
    RECT 220.165 71.325 220.445 72.205 ;
    RECT 216.845 71.325 217.125 72.205 ;
    RECT 180.325 71.325 180.605 72.205 ;
    RECT 177.005 71.325 177.285 72.205 ;
    RECT 173.685 71.325 173.965 72.205 ;
    RECT 170.365 71.325 170.645 72.205 ;
    RECT 167.045 71.325 167.325 72.205 ;
    RECT 163.725 71.325 164.005 72.205 ;
    RECT 160.405 71.325 160.685 72.205 ;
    RECT 157.085 71.325 157.365 72.205 ;
    RECT 153.765 71.325 154.045 72.205 ;
    RECT 150.445 71.325 150.725 72.205 ;
    RECT 213.525 71.325 213.805 72.205 ;
    RECT 210.205 71.325 210.485 72.205 ;
    RECT 206.885 71.325 207.165 72.205 ;
    RECT 203.565 71.325 203.845 72.205 ;
    RECT 200.245 71.325 200.525 72.205 ;
    RECT 196.925 71.325 197.205 72.205 ;
    RECT 193.605 71.325 193.885 72.205 ;
    RECT 190.285 71.325 190.565 72.205 ;
    RECT 186.965 71.325 187.245 72.205 ;
    RECT 183.645 71.325 183.925 72.205 ;
    RECT 266.645 71.325 266.925 72.205 ;
    RECT 263.325 71.325 263.605 72.205 ;
    RECT 260.005 71.325 260.285 72.205 ;
    RECT 256.685 71.325 256.965 72.205 ;
    RECT 253.365 71.325 253.645 72.205 ;
    RECT 250.045 15.145 250.325 16.025 ;
    RECT 246.725 15.145 247.005 16.025 ;
    RECT 243.405 15.145 243.685 16.025 ;
    RECT 240.085 15.145 240.365 16.025 ;
    RECT 236.765 15.145 237.045 16.025 ;
    RECT 233.445 15.145 233.725 16.025 ;
    RECT 230.125 15.145 230.405 16.025 ;
    RECT 226.805 15.145 227.085 16.025 ;
    RECT 223.485 15.145 223.765 16.025 ;
    RECT 220.165 15.145 220.445 16.025 ;
    RECT 216.845 15.145 217.125 16.025 ;
    RECT 180.325 15.145 180.605 16.025 ;
    RECT 177.005 15.145 177.285 16.025 ;
    RECT 173.685 15.145 173.965 16.025 ;
    RECT 170.365 15.145 170.645 16.025 ;
    RECT 167.045 15.145 167.325 16.025 ;
    RECT 163.725 15.145 164.005 16.025 ;
    RECT 160.405 15.145 160.685 16.025 ;
    RECT 157.085 15.145 157.365 16.025 ;
    RECT 153.765 15.145 154.045 16.025 ;
    RECT 150.445 15.145 150.725 16.025 ;
    RECT 213.525 15.145 213.805 16.025 ;
    RECT 210.205 15.145 210.485 16.025 ;
    RECT 206.885 15.145 207.165 16.025 ;
    RECT 203.565 15.145 203.845 16.025 ;
    RECT 200.245 15.145 200.525 16.025 ;
    RECT 196.925 15.145 197.205 16.025 ;
    RECT 193.605 15.145 193.885 16.025 ;
    RECT 190.285 15.145 190.565 16.025 ;
    RECT 186.965 15.145 187.245 16.025 ;
    RECT 183.645 15.145 183.925 16.025 ;
    RECT 266.645 15.145 266.925 16.025 ;
    RECT 263.325 15.145 263.605 16.025 ;
    RECT 260.005 15.145 260.285 16.025 ;
    RECT 256.685 15.145 256.965 16.025 ;
    RECT 253.365 15.145 253.645 16.025 ;
    RECT 250.045 30.985 250.325 31.865 ;
    RECT 246.725 30.985 247.005 31.865 ;
    RECT 243.405 30.985 243.685 31.865 ;
    RECT 240.085 30.985 240.365 31.865 ;
    RECT 236.765 30.985 237.045 31.865 ;
    RECT 233.445 30.985 233.725 31.865 ;
    RECT 230.125 30.985 230.405 31.865 ;
    RECT 226.805 30.985 227.085 31.865 ;
    RECT 223.485 30.985 223.765 31.865 ;
    RECT 220.165 30.985 220.445 31.865 ;
    RECT 216.845 30.985 217.125 31.865 ;
    RECT 180.325 30.985 180.605 31.865 ;
    RECT 177.005 30.985 177.285 31.865 ;
    RECT 173.685 30.985 173.965 31.865 ;
    RECT 170.365 30.985 170.645 31.865 ;
    RECT 167.045 30.985 167.325 31.865 ;
    RECT 163.725 30.985 164.005 31.865 ;
    RECT 160.405 30.985 160.685 31.865 ;
    RECT 157.085 30.985 157.365 31.865 ;
    RECT 153.765 30.985 154.045 31.865 ;
    RECT 150.445 30.985 150.725 31.865 ;
    RECT 213.525 30.985 213.805 31.865 ;
    RECT 210.205 30.985 210.485 31.865 ;
    RECT 206.885 30.985 207.165 31.865 ;
    RECT 203.565 30.985 203.845 31.865 ;
    RECT 200.245 30.985 200.525 31.865 ;
    RECT 196.925 30.985 197.205 31.865 ;
    RECT 193.605 30.985 193.885 31.865 ;
    RECT 190.285 30.985 190.565 31.865 ;
    RECT 186.965 30.985 187.245 31.865 ;
    RECT 183.645 30.985 183.925 31.865 ;
    RECT 266.645 30.985 266.925 31.865 ;
    RECT 263.325 30.985 263.605 31.865 ;
    RECT 260.005 30.985 260.285 31.865 ;
    RECT 256.685 30.985 256.965 31.865 ;
    RECT 253.365 30.985 253.645 31.865 ;
    RECT 250.045 70.605 250.325 71.485 ;
    RECT 246.725 70.605 247.005 71.485 ;
    RECT 243.405 70.605 243.685 71.485 ;
    RECT 240.085 70.605 240.365 71.485 ;
    RECT 236.765 70.605 237.045 71.485 ;
    RECT 233.445 70.605 233.725 71.485 ;
    RECT 230.125 70.605 230.405 71.485 ;
    RECT 226.805 70.605 227.085 71.485 ;
    RECT 223.485 70.605 223.765 71.485 ;
    RECT 220.165 70.605 220.445 71.485 ;
    RECT 216.845 70.605 217.125 71.485 ;
    RECT 180.325 70.605 180.605 71.485 ;
    RECT 177.005 70.605 177.285 71.485 ;
    RECT 173.685 70.605 173.965 71.485 ;
    RECT 170.365 70.605 170.645 71.485 ;
    RECT 167.045 70.605 167.325 71.485 ;
    RECT 163.725 70.605 164.005 71.485 ;
    RECT 160.405 70.605 160.685 71.485 ;
    RECT 157.085 70.605 157.365 71.485 ;
    RECT 153.765 70.605 154.045 71.485 ;
    RECT 150.445 70.605 150.725 71.485 ;
    RECT 213.525 70.605 213.805 71.485 ;
    RECT 210.205 70.605 210.485 71.485 ;
    RECT 206.885 70.605 207.165 71.485 ;
    RECT 203.565 70.605 203.845 71.485 ;
    RECT 200.245 70.605 200.525 71.485 ;
    RECT 196.925 70.605 197.205 71.485 ;
    RECT 193.605 70.605 193.885 71.485 ;
    RECT 190.285 70.605 190.565 71.485 ;
    RECT 186.965 70.605 187.245 71.485 ;
    RECT 183.645 70.605 183.925 71.485 ;
    RECT 266.645 70.605 266.925 71.485 ;
    RECT 263.325 70.605 263.605 71.485 ;
    RECT 260.005 70.605 260.285 71.485 ;
    RECT 256.685 70.605 256.965 71.485 ;
    RECT 253.365 70.605 253.645 71.485 ;
    RECT 250.045 30.265 250.325 31.145 ;
    RECT 246.725 30.265 247.005 31.145 ;
    RECT 243.405 30.265 243.685 31.145 ;
    RECT 240.085 30.265 240.365 31.145 ;
    RECT 236.765 30.265 237.045 31.145 ;
    RECT 233.445 30.265 233.725 31.145 ;
    RECT 230.125 30.265 230.405 31.145 ;
    RECT 226.805 30.265 227.085 31.145 ;
    RECT 223.485 30.265 223.765 31.145 ;
    RECT 220.165 30.265 220.445 31.145 ;
    RECT 216.845 30.265 217.125 31.145 ;
    RECT 180.325 30.265 180.605 31.145 ;
    RECT 177.005 30.265 177.285 31.145 ;
    RECT 173.685 30.265 173.965 31.145 ;
    RECT 170.365 30.265 170.645 31.145 ;
    RECT 167.045 30.265 167.325 31.145 ;
    RECT 163.725 30.265 164.005 31.145 ;
    RECT 160.405 30.265 160.685 31.145 ;
    RECT 157.085 30.265 157.365 31.145 ;
    RECT 153.765 30.265 154.045 31.145 ;
    RECT 150.445 30.265 150.725 31.145 ;
    RECT 213.525 30.265 213.805 31.145 ;
    RECT 210.205 30.265 210.485 31.145 ;
    RECT 206.885 30.265 207.165 31.145 ;
    RECT 203.565 30.265 203.845 31.145 ;
    RECT 200.245 30.265 200.525 31.145 ;
    RECT 196.925 30.265 197.205 31.145 ;
    RECT 193.605 30.265 193.885 31.145 ;
    RECT 190.285 30.265 190.565 31.145 ;
    RECT 186.965 30.265 187.245 31.145 ;
    RECT 183.645 30.265 183.925 31.145 ;
    RECT 266.645 30.265 266.925 31.145 ;
    RECT 263.325 30.265 263.605 31.145 ;
    RECT 260.005 30.265 260.285 31.145 ;
    RECT 256.685 30.265 256.965 31.145 ;
    RECT 253.365 30.265 253.645 31.145 ;
    RECT 250.045 69.885 250.325 70.765 ;
    RECT 246.725 69.885 247.005 70.765 ;
    RECT 243.405 69.885 243.685 70.765 ;
    RECT 240.085 69.885 240.365 70.765 ;
    RECT 236.765 69.885 237.045 70.765 ;
    RECT 233.445 69.885 233.725 70.765 ;
    RECT 230.125 69.885 230.405 70.765 ;
    RECT 226.805 69.885 227.085 70.765 ;
    RECT 223.485 69.885 223.765 70.765 ;
    RECT 220.165 69.885 220.445 70.765 ;
    RECT 216.845 69.885 217.125 70.765 ;
    RECT 180.325 69.885 180.605 70.765 ;
    RECT 177.005 69.885 177.285 70.765 ;
    RECT 173.685 69.885 173.965 70.765 ;
    RECT 170.365 69.885 170.645 70.765 ;
    RECT 167.045 69.885 167.325 70.765 ;
    RECT 163.725 69.885 164.005 70.765 ;
    RECT 160.405 69.885 160.685 70.765 ;
    RECT 157.085 69.885 157.365 70.765 ;
    RECT 153.765 69.885 154.045 70.765 ;
    RECT 150.445 69.885 150.725 70.765 ;
    RECT 213.525 69.885 213.805 70.765 ;
    RECT 210.205 69.885 210.485 70.765 ;
    RECT 206.885 69.885 207.165 70.765 ;
    RECT 203.565 69.885 203.845 70.765 ;
    RECT 200.245 69.885 200.525 70.765 ;
    RECT 196.925 69.885 197.205 70.765 ;
    RECT 193.605 69.885 193.885 70.765 ;
    RECT 190.285 69.885 190.565 70.765 ;
    RECT 186.965 69.885 187.245 70.765 ;
    RECT 183.645 69.885 183.925 70.765 ;
    RECT 266.645 69.885 266.925 70.765 ;
    RECT 263.325 69.885 263.605 70.765 ;
    RECT 260.005 69.885 260.285 70.765 ;
    RECT 256.685 69.885 256.965 70.765 ;
    RECT 253.365 69.885 253.645 70.765 ;
    RECT 250.045 29.545 250.325 30.425 ;
    RECT 246.725 29.545 247.005 30.425 ;
    RECT 243.405 29.545 243.685 30.425 ;
    RECT 240.085 29.545 240.365 30.425 ;
    RECT 236.765 29.545 237.045 30.425 ;
    RECT 233.445 29.545 233.725 30.425 ;
    RECT 230.125 29.545 230.405 30.425 ;
    RECT 226.805 29.545 227.085 30.425 ;
    RECT 223.485 29.545 223.765 30.425 ;
    RECT 220.165 29.545 220.445 30.425 ;
    RECT 216.845 29.545 217.125 30.425 ;
    RECT 180.325 29.545 180.605 30.425 ;
    RECT 177.005 29.545 177.285 30.425 ;
    RECT 173.685 29.545 173.965 30.425 ;
    RECT 170.365 29.545 170.645 30.425 ;
    RECT 167.045 29.545 167.325 30.425 ;
    RECT 163.725 29.545 164.005 30.425 ;
    RECT 160.405 29.545 160.685 30.425 ;
    RECT 157.085 29.545 157.365 30.425 ;
    RECT 153.765 29.545 154.045 30.425 ;
    RECT 150.445 29.545 150.725 30.425 ;
    RECT 213.525 29.545 213.805 30.425 ;
    RECT 210.205 29.545 210.485 30.425 ;
    RECT 206.885 29.545 207.165 30.425 ;
    RECT 203.565 29.545 203.845 30.425 ;
    RECT 200.245 29.545 200.525 30.425 ;
    RECT 196.925 29.545 197.205 30.425 ;
    RECT 193.605 29.545 193.885 30.425 ;
    RECT 190.285 29.545 190.565 30.425 ;
    RECT 186.965 29.545 187.245 30.425 ;
    RECT 183.645 29.545 183.925 30.425 ;
    RECT 266.645 29.545 266.925 30.425 ;
    RECT 263.325 29.545 263.605 30.425 ;
    RECT 260.005 29.545 260.285 30.425 ;
    RECT 256.685 29.545 256.965 30.425 ;
    RECT 253.365 29.545 253.645 30.425 ;
    RECT 250.045 69.165 250.325 70.045 ;
    RECT 246.725 69.165 247.005 70.045 ;
    RECT 243.405 69.165 243.685 70.045 ;
    RECT 240.085 69.165 240.365 70.045 ;
    RECT 236.765 69.165 237.045 70.045 ;
    RECT 233.445 69.165 233.725 70.045 ;
    RECT 230.125 69.165 230.405 70.045 ;
    RECT 226.805 69.165 227.085 70.045 ;
    RECT 223.485 69.165 223.765 70.045 ;
    RECT 220.165 69.165 220.445 70.045 ;
    RECT 216.845 69.165 217.125 70.045 ;
    RECT 180.325 69.165 180.605 70.045 ;
    RECT 177.005 69.165 177.285 70.045 ;
    RECT 173.685 69.165 173.965 70.045 ;
    RECT 170.365 69.165 170.645 70.045 ;
    RECT 167.045 69.165 167.325 70.045 ;
    RECT 163.725 69.165 164.005 70.045 ;
    RECT 160.405 69.165 160.685 70.045 ;
    RECT 157.085 69.165 157.365 70.045 ;
    RECT 153.765 69.165 154.045 70.045 ;
    RECT 150.445 69.165 150.725 70.045 ;
    RECT 213.525 69.165 213.805 70.045 ;
    RECT 210.205 69.165 210.485 70.045 ;
    RECT 206.885 69.165 207.165 70.045 ;
    RECT 203.565 69.165 203.845 70.045 ;
    RECT 200.245 69.165 200.525 70.045 ;
    RECT 196.925 69.165 197.205 70.045 ;
    RECT 193.605 69.165 193.885 70.045 ;
    RECT 190.285 69.165 190.565 70.045 ;
    RECT 186.965 69.165 187.245 70.045 ;
    RECT 183.645 69.165 183.925 70.045 ;
    RECT 266.645 69.165 266.925 70.045 ;
    RECT 263.325 69.165 263.605 70.045 ;
    RECT 260.005 69.165 260.285 70.045 ;
    RECT 256.685 69.165 256.965 70.045 ;
    RECT 253.365 69.165 253.645 70.045 ;
    RECT 250.045 28.825 250.325 29.705 ;
    RECT 246.725 28.825 247.005 29.705 ;
    RECT 243.405 28.825 243.685 29.705 ;
    RECT 240.085 28.825 240.365 29.705 ;
    RECT 236.765 28.825 237.045 29.705 ;
    RECT 233.445 28.825 233.725 29.705 ;
    RECT 230.125 28.825 230.405 29.705 ;
    RECT 226.805 28.825 227.085 29.705 ;
    RECT 223.485 28.825 223.765 29.705 ;
    RECT 220.165 28.825 220.445 29.705 ;
    RECT 216.845 28.825 217.125 29.705 ;
    RECT 180.325 28.825 180.605 29.705 ;
    RECT 177.005 28.825 177.285 29.705 ;
    RECT 173.685 28.825 173.965 29.705 ;
    RECT 170.365 28.825 170.645 29.705 ;
    RECT 167.045 28.825 167.325 29.705 ;
    RECT 163.725 28.825 164.005 29.705 ;
    RECT 160.405 28.825 160.685 29.705 ;
    RECT 157.085 28.825 157.365 29.705 ;
    RECT 153.765 28.825 154.045 29.705 ;
    RECT 150.445 28.825 150.725 29.705 ;
    RECT 213.525 28.825 213.805 29.705 ;
    RECT 210.205 28.825 210.485 29.705 ;
    RECT 206.885 28.825 207.165 29.705 ;
    RECT 203.565 28.825 203.845 29.705 ;
    RECT 200.245 28.825 200.525 29.705 ;
    RECT 196.925 28.825 197.205 29.705 ;
    RECT 193.605 28.825 193.885 29.705 ;
    RECT 190.285 28.825 190.565 29.705 ;
    RECT 186.965 28.825 187.245 29.705 ;
    RECT 183.645 28.825 183.925 29.705 ;
    RECT 266.645 28.825 266.925 29.705 ;
    RECT 263.325 28.825 263.605 29.705 ;
    RECT 260.005 28.825 260.285 29.705 ;
    RECT 256.685 28.825 256.965 29.705 ;
    RECT 253.365 28.825 253.645 29.705 ;
    RECT 250.045 68.445 250.325 69.325 ;
    RECT 246.725 68.445 247.005 69.325 ;
    RECT 243.405 68.445 243.685 69.325 ;
    RECT 240.085 68.445 240.365 69.325 ;
    RECT 236.765 68.445 237.045 69.325 ;
    RECT 233.445 68.445 233.725 69.325 ;
    RECT 230.125 68.445 230.405 69.325 ;
    RECT 226.805 68.445 227.085 69.325 ;
    RECT 223.485 68.445 223.765 69.325 ;
    RECT 220.165 68.445 220.445 69.325 ;
    RECT 216.845 68.445 217.125 69.325 ;
    RECT 180.325 68.445 180.605 69.325 ;
    RECT 177.005 68.445 177.285 69.325 ;
    RECT 173.685 68.445 173.965 69.325 ;
    RECT 170.365 68.445 170.645 69.325 ;
    RECT 167.045 68.445 167.325 69.325 ;
    RECT 163.725 68.445 164.005 69.325 ;
    RECT 160.405 68.445 160.685 69.325 ;
    RECT 157.085 68.445 157.365 69.325 ;
    RECT 153.765 68.445 154.045 69.325 ;
    RECT 150.445 68.445 150.725 69.325 ;
    RECT 213.525 68.445 213.805 69.325 ;
    RECT 210.205 68.445 210.485 69.325 ;
    RECT 206.885 68.445 207.165 69.325 ;
    RECT 203.565 68.445 203.845 69.325 ;
    RECT 200.245 68.445 200.525 69.325 ;
    RECT 196.925 68.445 197.205 69.325 ;
    RECT 193.605 68.445 193.885 69.325 ;
    RECT 190.285 68.445 190.565 69.325 ;
    RECT 186.965 68.445 187.245 69.325 ;
    RECT 183.645 68.445 183.925 69.325 ;
    RECT 266.645 68.445 266.925 69.325 ;
    RECT 263.325 68.445 263.605 69.325 ;
    RECT 260.005 68.445 260.285 69.325 ;
    RECT 256.685 68.445 256.965 69.325 ;
    RECT 253.365 68.445 253.645 69.325 ;
    RECT 250.045 67.725 250.325 68.605 ;
    RECT 246.725 67.725 247.005 68.605 ;
    RECT 243.405 67.725 243.685 68.605 ;
    RECT 240.085 67.725 240.365 68.605 ;
    RECT 236.765 67.725 237.045 68.605 ;
    RECT 233.445 67.725 233.725 68.605 ;
    RECT 230.125 67.725 230.405 68.605 ;
    RECT 226.805 67.725 227.085 68.605 ;
    RECT 223.485 67.725 223.765 68.605 ;
    RECT 220.165 67.725 220.445 68.605 ;
    RECT 216.845 67.725 217.125 68.605 ;
    RECT 180.325 67.725 180.605 68.605 ;
    RECT 177.005 67.725 177.285 68.605 ;
    RECT 173.685 67.725 173.965 68.605 ;
    RECT 170.365 67.725 170.645 68.605 ;
    RECT 167.045 67.725 167.325 68.605 ;
    RECT 163.725 67.725 164.005 68.605 ;
    RECT 160.405 67.725 160.685 68.605 ;
    RECT 157.085 67.725 157.365 68.605 ;
    RECT 153.765 67.725 154.045 68.605 ;
    RECT 150.445 67.725 150.725 68.605 ;
    RECT 213.525 67.725 213.805 68.605 ;
    RECT 210.205 67.725 210.485 68.605 ;
    RECT 206.885 67.725 207.165 68.605 ;
    RECT 203.565 67.725 203.845 68.605 ;
    RECT 200.245 67.725 200.525 68.605 ;
    RECT 196.925 67.725 197.205 68.605 ;
    RECT 193.605 67.725 193.885 68.605 ;
    RECT 190.285 67.725 190.565 68.605 ;
    RECT 186.965 67.725 187.245 68.605 ;
    RECT 183.645 67.725 183.925 68.605 ;
    RECT 266.645 67.725 266.925 68.605 ;
    RECT 263.325 67.725 263.605 68.605 ;
    RECT 260.005 67.725 260.285 68.605 ;
    RECT 256.685 67.725 256.965 68.605 ;
    RECT 253.365 67.725 253.645 68.605 ;
    RECT 250.045 67.005 250.325 67.885 ;
    RECT 246.725 67.005 247.005 67.885 ;
    RECT 243.405 67.005 243.685 67.885 ;
    RECT 240.085 67.005 240.365 67.885 ;
    RECT 236.765 67.005 237.045 67.885 ;
    RECT 233.445 67.005 233.725 67.885 ;
    RECT 230.125 67.005 230.405 67.885 ;
    RECT 226.805 67.005 227.085 67.885 ;
    RECT 223.485 67.005 223.765 67.885 ;
    RECT 220.165 67.005 220.445 67.885 ;
    RECT 216.845 67.005 217.125 67.885 ;
    RECT 180.325 67.005 180.605 67.885 ;
    RECT 177.005 67.005 177.285 67.885 ;
    RECT 173.685 67.005 173.965 67.885 ;
    RECT 170.365 67.005 170.645 67.885 ;
    RECT 167.045 67.005 167.325 67.885 ;
    RECT 163.725 67.005 164.005 67.885 ;
    RECT 160.405 67.005 160.685 67.885 ;
    RECT 157.085 67.005 157.365 67.885 ;
    RECT 153.765 67.005 154.045 67.885 ;
    RECT 150.445 67.005 150.725 67.885 ;
    RECT 213.525 67.005 213.805 67.885 ;
    RECT 210.205 67.005 210.485 67.885 ;
    RECT 206.885 67.005 207.165 67.885 ;
    RECT 203.565 67.005 203.845 67.885 ;
    RECT 200.245 67.005 200.525 67.885 ;
    RECT 196.925 67.005 197.205 67.885 ;
    RECT 193.605 67.005 193.885 67.885 ;
    RECT 190.285 67.005 190.565 67.885 ;
    RECT 186.965 67.005 187.245 67.885 ;
    RECT 183.645 67.005 183.925 67.885 ;
    RECT 266.645 67.005 266.925 67.885 ;
    RECT 263.325 67.005 263.605 67.885 ;
    RECT 260.005 67.005 260.285 67.885 ;
    RECT 256.685 67.005 256.965 67.885 ;
    RECT 253.365 67.005 253.645 67.885 ;
    RECT 250.045 66.285 250.325 67.165 ;
    RECT 246.725 66.285 247.005 67.165 ;
    RECT 243.405 66.285 243.685 67.165 ;
    RECT 240.085 66.285 240.365 67.165 ;
    RECT 236.765 66.285 237.045 67.165 ;
    RECT 233.445 66.285 233.725 67.165 ;
    RECT 230.125 66.285 230.405 67.165 ;
    RECT 226.805 66.285 227.085 67.165 ;
    RECT 223.485 66.285 223.765 67.165 ;
    RECT 220.165 66.285 220.445 67.165 ;
    RECT 216.845 66.285 217.125 67.165 ;
    RECT 180.325 66.285 180.605 67.165 ;
    RECT 177.005 66.285 177.285 67.165 ;
    RECT 173.685 66.285 173.965 67.165 ;
    RECT 170.365 66.285 170.645 67.165 ;
    RECT 167.045 66.285 167.325 67.165 ;
    RECT 163.725 66.285 164.005 67.165 ;
    RECT 160.405 66.285 160.685 67.165 ;
    RECT 157.085 66.285 157.365 67.165 ;
    RECT 153.765 66.285 154.045 67.165 ;
    RECT 150.445 66.285 150.725 67.165 ;
    RECT 213.525 66.285 213.805 67.165 ;
    RECT 210.205 66.285 210.485 67.165 ;
    RECT 206.885 66.285 207.165 67.165 ;
    RECT 203.565 66.285 203.845 67.165 ;
    RECT 200.245 66.285 200.525 67.165 ;
    RECT 196.925 66.285 197.205 67.165 ;
    RECT 193.605 66.285 193.885 67.165 ;
    RECT 190.285 66.285 190.565 67.165 ;
    RECT 186.965 66.285 187.245 67.165 ;
    RECT 183.645 66.285 183.925 67.165 ;
    RECT 266.645 66.285 266.925 67.165 ;
    RECT 263.325 66.285 263.605 67.165 ;
    RECT 260.005 66.285 260.285 67.165 ;
    RECT 256.685 66.285 256.965 67.165 ;
    RECT 253.365 66.285 253.645 67.165 ;
    RECT 250.045 65.565 250.325 66.445 ;
    RECT 246.725 65.565 247.005 66.445 ;
    RECT 243.405 65.565 243.685 66.445 ;
    RECT 240.085 65.565 240.365 66.445 ;
    RECT 236.765 65.565 237.045 66.445 ;
    RECT 233.445 65.565 233.725 66.445 ;
    RECT 230.125 65.565 230.405 66.445 ;
    RECT 226.805 65.565 227.085 66.445 ;
    RECT 223.485 65.565 223.765 66.445 ;
    RECT 220.165 65.565 220.445 66.445 ;
    RECT 216.845 65.565 217.125 66.445 ;
    RECT 180.325 65.565 180.605 66.445 ;
    RECT 177.005 65.565 177.285 66.445 ;
    RECT 173.685 65.565 173.965 66.445 ;
    RECT 170.365 65.565 170.645 66.445 ;
    RECT 167.045 65.565 167.325 66.445 ;
    RECT 163.725 65.565 164.005 66.445 ;
    RECT 160.405 65.565 160.685 66.445 ;
    RECT 157.085 65.565 157.365 66.445 ;
    RECT 153.765 65.565 154.045 66.445 ;
    RECT 150.445 65.565 150.725 66.445 ;
    RECT 213.525 65.565 213.805 66.445 ;
    RECT 210.205 65.565 210.485 66.445 ;
    RECT 206.885 65.565 207.165 66.445 ;
    RECT 203.565 65.565 203.845 66.445 ;
    RECT 200.245 65.565 200.525 66.445 ;
    RECT 196.925 65.565 197.205 66.445 ;
    RECT 193.605 65.565 193.885 66.445 ;
    RECT 190.285 65.565 190.565 66.445 ;
    RECT 186.965 65.565 187.245 66.445 ;
    RECT 183.645 65.565 183.925 66.445 ;
    RECT 266.645 65.565 266.925 66.445 ;
    RECT 263.325 65.565 263.605 66.445 ;
    RECT 260.005 65.565 260.285 66.445 ;
    RECT 256.685 65.565 256.965 66.445 ;
    RECT 253.365 65.565 253.645 66.445 ;
    RECT 250.045 56.185 250.325 57.065 ;
    RECT 246.725 56.185 247.005 57.065 ;
    RECT 243.405 56.185 243.685 57.065 ;
    RECT 240.085 56.185 240.365 57.065 ;
    RECT 236.765 56.185 237.045 57.065 ;
    RECT 233.445 56.185 233.725 57.065 ;
    RECT 230.125 56.185 230.405 57.065 ;
    RECT 226.805 56.185 227.085 57.065 ;
    RECT 223.485 56.185 223.765 57.065 ;
    RECT 220.165 56.185 220.445 57.065 ;
    RECT 216.845 56.185 217.125 57.065 ;
    RECT 180.325 56.185 180.605 57.065 ;
    RECT 177.005 56.185 177.285 57.065 ;
    RECT 173.685 56.185 173.965 57.065 ;
    RECT 170.365 56.185 170.645 57.065 ;
    RECT 167.045 56.185 167.325 57.065 ;
    RECT 163.725 56.185 164.005 57.065 ;
    RECT 160.405 56.185 160.685 57.065 ;
    RECT 157.085 56.185 157.365 57.065 ;
    RECT 153.765 56.185 154.045 57.065 ;
    RECT 150.445 56.185 150.725 57.065 ;
    RECT 213.525 56.185 213.805 57.065 ;
    RECT 210.205 56.185 210.485 57.065 ;
    RECT 206.885 56.185 207.165 57.065 ;
    RECT 203.565 56.185 203.845 57.065 ;
    RECT 200.245 56.185 200.525 57.065 ;
    RECT 196.925 56.185 197.205 57.065 ;
    RECT 193.605 56.185 193.885 57.065 ;
    RECT 190.285 56.185 190.565 57.065 ;
    RECT 186.965 56.185 187.245 57.065 ;
    RECT 183.645 56.185 183.925 57.065 ;
    RECT 266.645 56.185 266.925 57.065 ;
    RECT 263.325 56.185 263.605 57.065 ;
    RECT 260.005 56.185 260.285 57.065 ;
    RECT 256.685 56.185 256.965 57.065 ;
    RECT 253.365 56.185 253.645 57.065 ;
    RECT 266.645 98.765 266.925 100.295 ;
    RECT 263.325 98.765 263.605 100.295 ;
    RECT 260.005 98.765 260.285 100.295 ;
    RECT 256.685 98.765 256.965 100.295 ;
    RECT 253.365 98.765 253.645 100.295 ;
    RECT 250.045 98.765 250.325 100.295 ;
    RECT 246.725 98.765 247.005 100.295 ;
    RECT 243.405 98.765 243.685 100.295 ;
    RECT 240.085 98.765 240.365 100.295 ;
    RECT 236.765 98.765 237.045 100.295 ;
    RECT 233.445 98.765 233.725 100.295 ;
    RECT 230.125 98.765 230.405 100.295 ;
    RECT 226.805 98.765 227.085 100.295 ;
    RECT 223.485 98.765 223.765 100.295 ;
    RECT 220.165 98.765 220.445 100.295 ;
    RECT 216.845 98.765 217.125 100.295 ;
    RECT 213.525 98.765 213.805 100.295 ;
    RECT 210.205 98.765 210.485 100.295 ;
    RECT 206.885 98.765 207.165 100.295 ;
    RECT 203.565 98.765 203.845 100.295 ;
    RECT 200.245 98.765 200.525 100.295 ;
    RECT 196.925 98.765 197.205 100.295 ;
    RECT 193.605 98.765 193.885 100.295 ;
    RECT 190.285 98.765 190.565 100.295 ;
    RECT 186.965 98.765 187.245 100.295 ;
    RECT 183.645 98.765 183.925 100.295 ;
    RECT 180.325 98.765 180.605 100.295 ;
    RECT 177.005 98.765 177.285 100.295 ;
    RECT 173.685 98.765 173.965 100.295 ;
    RECT 170.365 98.765 170.645 100.295 ;
    RECT 167.045 98.765 167.325 100.295 ;
    RECT 163.725 98.765 164.005 100.295 ;
    RECT 160.405 98.765 160.685 100.295 ;
    RECT 157.085 98.765 157.365 100.295 ;
    RECT 153.765 98.765 154.045 100.295 ;
    RECT 150.445 98.765 150.725 100.295 ;
    RECT 250.045 28.105 250.325 28.985 ;
    RECT 246.725 28.105 247.005 28.985 ;
    RECT 243.405 28.105 243.685 28.985 ;
    RECT 240.085 28.105 240.365 28.985 ;
    RECT 236.765 28.105 237.045 28.985 ;
    RECT 233.445 28.105 233.725 28.985 ;
    RECT 230.125 28.105 230.405 28.985 ;
    RECT 226.805 28.105 227.085 28.985 ;
    RECT 223.485 28.105 223.765 28.985 ;
    RECT 220.165 28.105 220.445 28.985 ;
    RECT 216.845 28.105 217.125 28.985 ;
    RECT 180.325 28.105 180.605 28.985 ;
    RECT 177.005 28.105 177.285 28.985 ;
    RECT 173.685 28.105 173.965 28.985 ;
    RECT 170.365 28.105 170.645 28.985 ;
    RECT 167.045 28.105 167.325 28.985 ;
    RECT 163.725 28.105 164.005 28.985 ;
    RECT 160.405 28.105 160.685 28.985 ;
    RECT 157.085 28.105 157.365 28.985 ;
    RECT 153.765 28.105 154.045 28.985 ;
    RECT 150.445 28.105 150.725 28.985 ;
    RECT 213.525 28.105 213.805 28.985 ;
    RECT 210.205 28.105 210.485 28.985 ;
    RECT 206.885 28.105 207.165 28.985 ;
    RECT 203.565 28.105 203.845 28.985 ;
    RECT 200.245 28.105 200.525 28.985 ;
    RECT 196.925 28.105 197.205 28.985 ;
    RECT 193.605 28.105 193.885 28.985 ;
    RECT 190.285 28.105 190.565 28.985 ;
    RECT 186.965 28.105 187.245 28.985 ;
    RECT 183.645 28.105 183.925 28.985 ;
    RECT 266.645 28.105 266.925 28.985 ;
    RECT 263.325 28.105 263.605 28.985 ;
    RECT 260.005 28.105 260.285 28.985 ;
    RECT 256.685 28.105 256.965 28.985 ;
    RECT 253.365 28.105 253.645 28.985 ;
    RECT 250.045 27.385 250.325 28.265 ;
    RECT 246.725 27.385 247.005 28.265 ;
    RECT 243.405 27.385 243.685 28.265 ;
    RECT 240.085 27.385 240.365 28.265 ;
    RECT 236.765 27.385 237.045 28.265 ;
    RECT 233.445 27.385 233.725 28.265 ;
    RECT 230.125 27.385 230.405 28.265 ;
    RECT 226.805 27.385 227.085 28.265 ;
    RECT 223.485 27.385 223.765 28.265 ;
    RECT 220.165 27.385 220.445 28.265 ;
    RECT 216.845 27.385 217.125 28.265 ;
    RECT 180.325 27.385 180.605 28.265 ;
    RECT 177.005 27.385 177.285 28.265 ;
    RECT 173.685 27.385 173.965 28.265 ;
    RECT 170.365 27.385 170.645 28.265 ;
    RECT 167.045 27.385 167.325 28.265 ;
    RECT 163.725 27.385 164.005 28.265 ;
    RECT 160.405 27.385 160.685 28.265 ;
    RECT 157.085 27.385 157.365 28.265 ;
    RECT 153.765 27.385 154.045 28.265 ;
    RECT 150.445 27.385 150.725 28.265 ;
    RECT 213.525 27.385 213.805 28.265 ;
    RECT 210.205 27.385 210.485 28.265 ;
    RECT 206.885 27.385 207.165 28.265 ;
    RECT 203.565 27.385 203.845 28.265 ;
    RECT 200.245 27.385 200.525 28.265 ;
    RECT 196.925 27.385 197.205 28.265 ;
    RECT 193.605 27.385 193.885 28.265 ;
    RECT 190.285 27.385 190.565 28.265 ;
    RECT 186.965 27.385 187.245 28.265 ;
    RECT 183.645 27.385 183.925 28.265 ;
    RECT 266.645 27.385 266.925 28.265 ;
    RECT 263.325 27.385 263.605 28.265 ;
    RECT 260.005 27.385 260.285 28.265 ;
    RECT 256.685 27.385 256.965 28.265 ;
    RECT 253.365 27.385 253.645 28.265 ;
    RECT 250.045 26.665 250.325 27.545 ;
    RECT 246.725 26.665 247.005 27.545 ;
    RECT 243.405 26.665 243.685 27.545 ;
    RECT 240.085 26.665 240.365 27.545 ;
    RECT 236.765 26.665 237.045 27.545 ;
    RECT 233.445 26.665 233.725 27.545 ;
    RECT 230.125 26.665 230.405 27.545 ;
    RECT 226.805 26.665 227.085 27.545 ;
    RECT 223.485 26.665 223.765 27.545 ;
    RECT 220.165 26.665 220.445 27.545 ;
    RECT 216.845 26.665 217.125 27.545 ;
    RECT 180.325 26.665 180.605 27.545 ;
    RECT 177.005 26.665 177.285 27.545 ;
    RECT 173.685 26.665 173.965 27.545 ;
    RECT 170.365 26.665 170.645 27.545 ;
    RECT 167.045 26.665 167.325 27.545 ;
    RECT 163.725 26.665 164.005 27.545 ;
    RECT 160.405 26.665 160.685 27.545 ;
    RECT 157.085 26.665 157.365 27.545 ;
    RECT 153.765 26.665 154.045 27.545 ;
    RECT 150.445 26.665 150.725 27.545 ;
    RECT 213.525 26.665 213.805 27.545 ;
    RECT 210.205 26.665 210.485 27.545 ;
    RECT 206.885 26.665 207.165 27.545 ;
    RECT 203.565 26.665 203.845 27.545 ;
    RECT 200.245 26.665 200.525 27.545 ;
    RECT 196.925 26.665 197.205 27.545 ;
    RECT 193.605 26.665 193.885 27.545 ;
    RECT 190.285 26.665 190.565 27.545 ;
    RECT 186.965 26.665 187.245 27.545 ;
    RECT 183.645 26.665 183.925 27.545 ;
    RECT 266.645 26.665 266.925 27.545 ;
    RECT 263.325 26.665 263.605 27.545 ;
    RECT 260.005 26.665 260.285 27.545 ;
    RECT 256.685 26.665 256.965 27.545 ;
    RECT 253.365 26.665 253.645 27.545 ;
    RECT 250.045 25.945 250.325 26.825 ;
    RECT 246.725 25.945 247.005 26.825 ;
    RECT 243.405 25.945 243.685 26.825 ;
    RECT 240.085 25.945 240.365 26.825 ;
    RECT 236.765 25.945 237.045 26.825 ;
    RECT 233.445 25.945 233.725 26.825 ;
    RECT 230.125 25.945 230.405 26.825 ;
    RECT 226.805 25.945 227.085 26.825 ;
    RECT 223.485 25.945 223.765 26.825 ;
    RECT 220.165 25.945 220.445 26.825 ;
    RECT 216.845 25.945 217.125 26.825 ;
    RECT 180.325 25.945 180.605 26.825 ;
    RECT 177.005 25.945 177.285 26.825 ;
    RECT 173.685 25.945 173.965 26.825 ;
    RECT 170.365 25.945 170.645 26.825 ;
    RECT 167.045 25.945 167.325 26.825 ;
    RECT 163.725 25.945 164.005 26.825 ;
    RECT 160.405 25.945 160.685 26.825 ;
    RECT 157.085 25.945 157.365 26.825 ;
    RECT 153.765 25.945 154.045 26.825 ;
    RECT 150.445 25.945 150.725 26.825 ;
    RECT 213.525 25.945 213.805 26.825 ;
    RECT 210.205 25.945 210.485 26.825 ;
    RECT 206.885 25.945 207.165 26.825 ;
    RECT 203.565 25.945 203.845 26.825 ;
    RECT 200.245 25.945 200.525 26.825 ;
    RECT 196.925 25.945 197.205 26.825 ;
    RECT 193.605 25.945 193.885 26.825 ;
    RECT 190.285 25.945 190.565 26.825 ;
    RECT 186.965 25.945 187.245 26.825 ;
    RECT 183.645 25.945 183.925 26.825 ;
    RECT 266.645 25.945 266.925 26.825 ;
    RECT 263.325 25.945 263.605 26.825 ;
    RECT 260.005 25.945 260.285 26.825 ;
    RECT 256.685 25.945 256.965 26.825 ;
    RECT 253.365 25.945 253.645 26.825 ;
    RECT 250.045 25.225 250.325 26.105 ;
    RECT 246.725 25.225 247.005 26.105 ;
    RECT 243.405 25.225 243.685 26.105 ;
    RECT 240.085 25.225 240.365 26.105 ;
    RECT 236.765 25.225 237.045 26.105 ;
    RECT 233.445 25.225 233.725 26.105 ;
    RECT 230.125 25.225 230.405 26.105 ;
    RECT 226.805 25.225 227.085 26.105 ;
    RECT 223.485 25.225 223.765 26.105 ;
    RECT 220.165 25.225 220.445 26.105 ;
    RECT 216.845 25.225 217.125 26.105 ;
    RECT 180.325 25.225 180.605 26.105 ;
    RECT 177.005 25.225 177.285 26.105 ;
    RECT 173.685 25.225 173.965 26.105 ;
    RECT 170.365 25.225 170.645 26.105 ;
    RECT 167.045 25.225 167.325 26.105 ;
    RECT 163.725 25.225 164.005 26.105 ;
    RECT 160.405 25.225 160.685 26.105 ;
    RECT 157.085 25.225 157.365 26.105 ;
    RECT 153.765 25.225 154.045 26.105 ;
    RECT 150.445 25.225 150.725 26.105 ;
    RECT 213.525 25.225 213.805 26.105 ;
    RECT 210.205 25.225 210.485 26.105 ;
    RECT 206.885 25.225 207.165 26.105 ;
    RECT 203.565 25.225 203.845 26.105 ;
    RECT 200.245 25.225 200.525 26.105 ;
    RECT 196.925 25.225 197.205 26.105 ;
    RECT 193.605 25.225 193.885 26.105 ;
    RECT 190.285 25.225 190.565 26.105 ;
    RECT 186.965 25.225 187.245 26.105 ;
    RECT 183.645 25.225 183.925 26.105 ;
    RECT 266.645 25.225 266.925 26.105 ;
    RECT 263.325 25.225 263.605 26.105 ;
    RECT 260.005 25.225 260.285 26.105 ;
    RECT 256.685 25.225 256.965 26.105 ;
    RECT 253.365 25.225 253.645 26.105 ;
    RECT 250.045 64.845 250.325 65.725 ;
    RECT 246.725 64.845 247.005 65.725 ;
    RECT 243.405 64.845 243.685 65.725 ;
    RECT 240.085 64.845 240.365 65.725 ;
    RECT 236.765 64.845 237.045 65.725 ;
    RECT 233.445 64.845 233.725 65.725 ;
    RECT 230.125 64.845 230.405 65.725 ;
    RECT 226.805 64.845 227.085 65.725 ;
    RECT 223.485 64.845 223.765 65.725 ;
    RECT 220.165 64.845 220.445 65.725 ;
    RECT 216.845 64.845 217.125 65.725 ;
    RECT 180.325 64.845 180.605 65.725 ;
    RECT 177.005 64.845 177.285 65.725 ;
    RECT 173.685 64.845 173.965 65.725 ;
    RECT 170.365 64.845 170.645 65.725 ;
    RECT 167.045 64.845 167.325 65.725 ;
    RECT 163.725 64.845 164.005 65.725 ;
    RECT 160.405 64.845 160.685 65.725 ;
    RECT 157.085 64.845 157.365 65.725 ;
    RECT 153.765 64.845 154.045 65.725 ;
    RECT 150.445 64.845 150.725 65.725 ;
    RECT 213.525 64.845 213.805 65.725 ;
    RECT 210.205 64.845 210.485 65.725 ;
    RECT 206.885 64.845 207.165 65.725 ;
    RECT 203.565 64.845 203.845 65.725 ;
    RECT 200.245 64.845 200.525 65.725 ;
    RECT 196.925 64.845 197.205 65.725 ;
    RECT 193.605 64.845 193.885 65.725 ;
    RECT 190.285 64.845 190.565 65.725 ;
    RECT 186.965 64.845 187.245 65.725 ;
    RECT 183.645 64.845 183.925 65.725 ;
    RECT 266.645 64.845 266.925 65.725 ;
    RECT 263.325 64.845 263.605 65.725 ;
    RECT 260.005 64.845 260.285 65.725 ;
    RECT 256.685 64.845 256.965 65.725 ;
    RECT 253.365 64.845 253.645 65.725 ;
    RECT 250.045 24.505 250.325 25.385 ;
    RECT 246.725 24.505 247.005 25.385 ;
    RECT 243.405 24.505 243.685 25.385 ;
    RECT 240.085 24.505 240.365 25.385 ;
    RECT 236.765 24.505 237.045 25.385 ;
    RECT 233.445 24.505 233.725 25.385 ;
    RECT 230.125 24.505 230.405 25.385 ;
    RECT 226.805 24.505 227.085 25.385 ;
    RECT 223.485 24.505 223.765 25.385 ;
    RECT 220.165 24.505 220.445 25.385 ;
    RECT 216.845 24.505 217.125 25.385 ;
    RECT 180.325 24.505 180.605 25.385 ;
    RECT 177.005 24.505 177.285 25.385 ;
    RECT 173.685 24.505 173.965 25.385 ;
    RECT 170.365 24.505 170.645 25.385 ;
    RECT 167.045 24.505 167.325 25.385 ;
    RECT 163.725 24.505 164.005 25.385 ;
    RECT 160.405 24.505 160.685 25.385 ;
    RECT 157.085 24.505 157.365 25.385 ;
    RECT 153.765 24.505 154.045 25.385 ;
    RECT 150.445 24.505 150.725 25.385 ;
    RECT 213.525 24.505 213.805 25.385 ;
    RECT 210.205 24.505 210.485 25.385 ;
    RECT 206.885 24.505 207.165 25.385 ;
    RECT 203.565 24.505 203.845 25.385 ;
    RECT 200.245 24.505 200.525 25.385 ;
    RECT 196.925 24.505 197.205 25.385 ;
    RECT 193.605 24.505 193.885 25.385 ;
    RECT 190.285 24.505 190.565 25.385 ;
    RECT 186.965 24.505 187.245 25.385 ;
    RECT 183.645 24.505 183.925 25.385 ;
    RECT 266.645 24.505 266.925 25.385 ;
    RECT 263.325 24.505 263.605 25.385 ;
    RECT 260.005 24.505 260.285 25.385 ;
    RECT 256.685 24.505 256.965 25.385 ;
    RECT 253.365 24.505 253.645 25.385 ;
    RECT 250.045 64.125 250.325 65.005 ;
    RECT 246.725 64.125 247.005 65.005 ;
    RECT 243.405 64.125 243.685 65.005 ;
    RECT 240.085 64.125 240.365 65.005 ;
    RECT 236.765 64.125 237.045 65.005 ;
    RECT 233.445 64.125 233.725 65.005 ;
    RECT 230.125 64.125 230.405 65.005 ;
    RECT 226.805 64.125 227.085 65.005 ;
    RECT 223.485 64.125 223.765 65.005 ;
    RECT 220.165 64.125 220.445 65.005 ;
    RECT 216.845 64.125 217.125 65.005 ;
    RECT 180.325 64.125 180.605 65.005 ;
    RECT 177.005 64.125 177.285 65.005 ;
    RECT 173.685 64.125 173.965 65.005 ;
    RECT 170.365 64.125 170.645 65.005 ;
    RECT 167.045 64.125 167.325 65.005 ;
    RECT 163.725 64.125 164.005 65.005 ;
    RECT 160.405 64.125 160.685 65.005 ;
    RECT 157.085 64.125 157.365 65.005 ;
    RECT 153.765 64.125 154.045 65.005 ;
    RECT 150.445 64.125 150.725 65.005 ;
    RECT 213.525 64.125 213.805 65.005 ;
    RECT 210.205 64.125 210.485 65.005 ;
    RECT 206.885 64.125 207.165 65.005 ;
    RECT 203.565 64.125 203.845 65.005 ;
    RECT 200.245 64.125 200.525 65.005 ;
    RECT 196.925 64.125 197.205 65.005 ;
    RECT 193.605 64.125 193.885 65.005 ;
    RECT 190.285 64.125 190.565 65.005 ;
    RECT 186.965 64.125 187.245 65.005 ;
    RECT 183.645 64.125 183.925 65.005 ;
    RECT 266.645 64.125 266.925 65.005 ;
    RECT 263.325 64.125 263.605 65.005 ;
    RECT 260.005 64.125 260.285 65.005 ;
    RECT 256.685 64.125 256.965 65.005 ;
    RECT 253.365 64.125 253.645 65.005 ;
    RECT 250.045 23.785 250.325 24.665 ;
    RECT 246.725 23.785 247.005 24.665 ;
    RECT 243.405 23.785 243.685 24.665 ;
    RECT 240.085 23.785 240.365 24.665 ;
    RECT 236.765 23.785 237.045 24.665 ;
    RECT 233.445 23.785 233.725 24.665 ;
    RECT 230.125 23.785 230.405 24.665 ;
    RECT 226.805 23.785 227.085 24.665 ;
    RECT 223.485 23.785 223.765 24.665 ;
    RECT 220.165 23.785 220.445 24.665 ;
    RECT 216.845 23.785 217.125 24.665 ;
    RECT 180.325 23.785 180.605 24.665 ;
    RECT 177.005 23.785 177.285 24.665 ;
    RECT 173.685 23.785 173.965 24.665 ;
    RECT 170.365 23.785 170.645 24.665 ;
    RECT 167.045 23.785 167.325 24.665 ;
    RECT 163.725 23.785 164.005 24.665 ;
    RECT 160.405 23.785 160.685 24.665 ;
    RECT 157.085 23.785 157.365 24.665 ;
    RECT 153.765 23.785 154.045 24.665 ;
    RECT 150.445 23.785 150.725 24.665 ;
    RECT 213.525 23.785 213.805 24.665 ;
    RECT 210.205 23.785 210.485 24.665 ;
    RECT 206.885 23.785 207.165 24.665 ;
    RECT 203.565 23.785 203.845 24.665 ;
    RECT 200.245 23.785 200.525 24.665 ;
    RECT 196.925 23.785 197.205 24.665 ;
    RECT 193.605 23.785 193.885 24.665 ;
    RECT 190.285 23.785 190.565 24.665 ;
    RECT 186.965 23.785 187.245 24.665 ;
    RECT 183.645 23.785 183.925 24.665 ;
    RECT 266.645 23.785 266.925 24.665 ;
    RECT 263.325 23.785 263.605 24.665 ;
    RECT 260.005 23.785 260.285 24.665 ;
    RECT 256.685 23.785 256.965 24.665 ;
    RECT 253.365 23.785 253.645 24.665 ;
    RECT 250.045 63.405 250.325 64.285 ;
    RECT 246.725 63.405 247.005 64.285 ;
    RECT 243.405 63.405 243.685 64.285 ;
    RECT 240.085 63.405 240.365 64.285 ;
    RECT 236.765 63.405 237.045 64.285 ;
    RECT 233.445 63.405 233.725 64.285 ;
    RECT 230.125 63.405 230.405 64.285 ;
    RECT 226.805 63.405 227.085 64.285 ;
    RECT 223.485 63.405 223.765 64.285 ;
    RECT 220.165 63.405 220.445 64.285 ;
    RECT 216.845 63.405 217.125 64.285 ;
    RECT 180.325 63.405 180.605 64.285 ;
    RECT 177.005 63.405 177.285 64.285 ;
    RECT 173.685 63.405 173.965 64.285 ;
    RECT 170.365 63.405 170.645 64.285 ;
    RECT 167.045 63.405 167.325 64.285 ;
    RECT 163.725 63.405 164.005 64.285 ;
    RECT 160.405 63.405 160.685 64.285 ;
    RECT 157.085 63.405 157.365 64.285 ;
    RECT 153.765 63.405 154.045 64.285 ;
    RECT 150.445 63.405 150.725 64.285 ;
    RECT 213.525 63.405 213.805 64.285 ;
    RECT 210.205 63.405 210.485 64.285 ;
    RECT 206.885 63.405 207.165 64.285 ;
    RECT 203.565 63.405 203.845 64.285 ;
    RECT 200.245 63.405 200.525 64.285 ;
    RECT 196.925 63.405 197.205 64.285 ;
    RECT 193.605 63.405 193.885 64.285 ;
    RECT 190.285 63.405 190.565 64.285 ;
    RECT 186.965 63.405 187.245 64.285 ;
    RECT 183.645 63.405 183.925 64.285 ;
    RECT 266.645 63.405 266.925 64.285 ;
    RECT 263.325 63.405 263.605 64.285 ;
    RECT 260.005 63.405 260.285 64.285 ;
    RECT 256.685 63.405 256.965 64.285 ;
    RECT 253.365 63.405 253.645 64.285 ;
    RECT 250.045 55.465 250.325 56.345 ;
    RECT 246.725 55.465 247.005 56.345 ;
    RECT 243.405 55.465 243.685 56.345 ;
    RECT 240.085 55.465 240.365 56.345 ;
    RECT 236.765 55.465 237.045 56.345 ;
    RECT 233.445 55.465 233.725 56.345 ;
    RECT 230.125 55.465 230.405 56.345 ;
    RECT 226.805 55.465 227.085 56.345 ;
    RECT 223.485 55.465 223.765 56.345 ;
    RECT 220.165 55.465 220.445 56.345 ;
    RECT 216.845 55.465 217.125 56.345 ;
    RECT 180.325 55.465 180.605 56.345 ;
    RECT 177.005 55.465 177.285 56.345 ;
    RECT 173.685 55.465 173.965 56.345 ;
    RECT 170.365 55.465 170.645 56.345 ;
    RECT 167.045 55.465 167.325 56.345 ;
    RECT 163.725 55.465 164.005 56.345 ;
    RECT 160.405 55.465 160.685 56.345 ;
    RECT 157.085 55.465 157.365 56.345 ;
    RECT 153.765 55.465 154.045 56.345 ;
    RECT 150.445 55.465 150.725 56.345 ;
    RECT 213.525 55.465 213.805 56.345 ;
    RECT 210.205 55.465 210.485 56.345 ;
    RECT 206.885 55.465 207.165 56.345 ;
    RECT 203.565 55.465 203.845 56.345 ;
    RECT 200.245 55.465 200.525 56.345 ;
    RECT 196.925 55.465 197.205 56.345 ;
    RECT 193.605 55.465 193.885 56.345 ;
    RECT 190.285 55.465 190.565 56.345 ;
    RECT 186.965 55.465 187.245 56.345 ;
    RECT 183.645 55.465 183.925 56.345 ;
    RECT 266.645 55.465 266.925 56.345 ;
    RECT 263.325 55.465 263.605 56.345 ;
    RECT 260.005 55.465 260.285 56.345 ;
    RECT 256.685 55.465 256.965 56.345 ;
    RECT 253.365 55.465 253.645 56.345 ;
    RECT 250.045 23.065 250.325 23.945 ;
    RECT 246.725 23.065 247.005 23.945 ;
    RECT 243.405 23.065 243.685 23.945 ;
    RECT 240.085 23.065 240.365 23.945 ;
    RECT 236.765 23.065 237.045 23.945 ;
    RECT 233.445 23.065 233.725 23.945 ;
    RECT 230.125 23.065 230.405 23.945 ;
    RECT 226.805 23.065 227.085 23.945 ;
    RECT 223.485 23.065 223.765 23.945 ;
    RECT 220.165 23.065 220.445 23.945 ;
    RECT 216.845 23.065 217.125 23.945 ;
    RECT 180.325 23.065 180.605 23.945 ;
    RECT 177.005 23.065 177.285 23.945 ;
    RECT 173.685 23.065 173.965 23.945 ;
    RECT 170.365 23.065 170.645 23.945 ;
    RECT 167.045 23.065 167.325 23.945 ;
    RECT 163.725 23.065 164.005 23.945 ;
    RECT 160.405 23.065 160.685 23.945 ;
    RECT 157.085 23.065 157.365 23.945 ;
    RECT 153.765 23.065 154.045 23.945 ;
    RECT 150.445 23.065 150.725 23.945 ;
    RECT 213.525 23.065 213.805 23.945 ;
    RECT 210.205 23.065 210.485 23.945 ;
    RECT 206.885 23.065 207.165 23.945 ;
    RECT 203.565 23.065 203.845 23.945 ;
    RECT 200.245 23.065 200.525 23.945 ;
    RECT 196.925 23.065 197.205 23.945 ;
    RECT 193.605 23.065 193.885 23.945 ;
    RECT 190.285 23.065 190.565 23.945 ;
    RECT 186.965 23.065 187.245 23.945 ;
    RECT 183.645 23.065 183.925 23.945 ;
    RECT 266.645 23.065 266.925 23.945 ;
    RECT 263.325 23.065 263.605 23.945 ;
    RECT 260.005 23.065 260.285 23.945 ;
    RECT 256.685 23.065 256.965 23.945 ;
    RECT 253.365 23.065 253.645 23.945 ;
    RECT 250.045 62.685 250.325 63.565 ;
    RECT 246.725 62.685 247.005 63.565 ;
    RECT 243.405 62.685 243.685 63.565 ;
    RECT 240.085 62.685 240.365 63.565 ;
    RECT 236.765 62.685 237.045 63.565 ;
    RECT 233.445 62.685 233.725 63.565 ;
    RECT 230.125 62.685 230.405 63.565 ;
    RECT 226.805 62.685 227.085 63.565 ;
    RECT 223.485 62.685 223.765 63.565 ;
    RECT 220.165 62.685 220.445 63.565 ;
    RECT 216.845 62.685 217.125 63.565 ;
    RECT 180.325 62.685 180.605 63.565 ;
    RECT 177.005 62.685 177.285 63.565 ;
    RECT 173.685 62.685 173.965 63.565 ;
    RECT 170.365 62.685 170.645 63.565 ;
    RECT 167.045 62.685 167.325 63.565 ;
    RECT 163.725 62.685 164.005 63.565 ;
    RECT 160.405 62.685 160.685 63.565 ;
    RECT 157.085 62.685 157.365 63.565 ;
    RECT 153.765 62.685 154.045 63.565 ;
    RECT 150.445 62.685 150.725 63.565 ;
    RECT 213.525 62.685 213.805 63.565 ;
    RECT 210.205 62.685 210.485 63.565 ;
    RECT 206.885 62.685 207.165 63.565 ;
    RECT 203.565 62.685 203.845 63.565 ;
    RECT 200.245 62.685 200.525 63.565 ;
    RECT 196.925 62.685 197.205 63.565 ;
    RECT 193.605 62.685 193.885 63.565 ;
    RECT 190.285 62.685 190.565 63.565 ;
    RECT 186.965 62.685 187.245 63.565 ;
    RECT 183.645 62.685 183.925 63.565 ;
    RECT 266.645 62.685 266.925 63.565 ;
    RECT 263.325 62.685 263.605 63.565 ;
    RECT 260.005 62.685 260.285 63.565 ;
    RECT 256.685 62.685 256.965 63.565 ;
    RECT 253.365 62.685 253.645 63.565 ;
    RECT 250.045 54.745 250.325 55.625 ;
    RECT 246.725 54.745 247.005 55.625 ;
    RECT 243.405 54.745 243.685 55.625 ;
    RECT 240.085 54.745 240.365 55.625 ;
    RECT 236.765 54.745 237.045 55.625 ;
    RECT 233.445 54.745 233.725 55.625 ;
    RECT 230.125 54.745 230.405 55.625 ;
    RECT 226.805 54.745 227.085 55.625 ;
    RECT 223.485 54.745 223.765 55.625 ;
    RECT 220.165 54.745 220.445 55.625 ;
    RECT 216.845 54.745 217.125 55.625 ;
    RECT 180.325 54.745 180.605 55.625 ;
    RECT 177.005 54.745 177.285 55.625 ;
    RECT 173.685 54.745 173.965 55.625 ;
    RECT 170.365 54.745 170.645 55.625 ;
    RECT 167.045 54.745 167.325 55.625 ;
    RECT 163.725 54.745 164.005 55.625 ;
    RECT 160.405 54.745 160.685 55.625 ;
    RECT 157.085 54.745 157.365 55.625 ;
    RECT 153.765 54.745 154.045 55.625 ;
    RECT 150.445 54.745 150.725 55.625 ;
    RECT 213.525 54.745 213.805 55.625 ;
    RECT 210.205 54.745 210.485 55.625 ;
    RECT 206.885 54.745 207.165 55.625 ;
    RECT 203.565 54.745 203.845 55.625 ;
    RECT 200.245 54.745 200.525 55.625 ;
    RECT 196.925 54.745 197.205 55.625 ;
    RECT 193.605 54.745 193.885 55.625 ;
    RECT 190.285 54.745 190.565 55.625 ;
    RECT 186.965 54.745 187.245 55.625 ;
    RECT 183.645 54.745 183.925 55.625 ;
    RECT 266.645 54.745 266.925 55.625 ;
    RECT 263.325 54.745 263.605 55.625 ;
    RECT 260.005 54.745 260.285 55.625 ;
    RECT 256.685 54.745 256.965 55.625 ;
    RECT 253.365 54.745 253.645 55.625 ;
    RECT 250.045 22.345 250.325 23.225 ;
    RECT 246.725 22.345 247.005 23.225 ;
    RECT 243.405 22.345 243.685 23.225 ;
    RECT 240.085 22.345 240.365 23.225 ;
    RECT 236.765 22.345 237.045 23.225 ;
    RECT 233.445 22.345 233.725 23.225 ;
    RECT 230.125 22.345 230.405 23.225 ;
    RECT 226.805 22.345 227.085 23.225 ;
    RECT 223.485 22.345 223.765 23.225 ;
    RECT 220.165 22.345 220.445 23.225 ;
    RECT 216.845 22.345 217.125 23.225 ;
    RECT 180.325 22.345 180.605 23.225 ;
    RECT 177.005 22.345 177.285 23.225 ;
    RECT 173.685 22.345 173.965 23.225 ;
    RECT 170.365 22.345 170.645 23.225 ;
    RECT 167.045 22.345 167.325 23.225 ;
    RECT 163.725 22.345 164.005 23.225 ;
    RECT 160.405 22.345 160.685 23.225 ;
    RECT 157.085 22.345 157.365 23.225 ;
    RECT 153.765 22.345 154.045 23.225 ;
    RECT 150.445 22.345 150.725 23.225 ;
    RECT 213.525 22.345 213.805 23.225 ;
    RECT 210.205 22.345 210.485 23.225 ;
    RECT 206.885 22.345 207.165 23.225 ;
    RECT 203.565 22.345 203.845 23.225 ;
    RECT 200.245 22.345 200.525 23.225 ;
    RECT 196.925 22.345 197.205 23.225 ;
    RECT 193.605 22.345 193.885 23.225 ;
    RECT 190.285 22.345 190.565 23.225 ;
    RECT 186.965 22.345 187.245 23.225 ;
    RECT 183.645 22.345 183.925 23.225 ;
    RECT 266.645 22.345 266.925 23.225 ;
    RECT 263.325 22.345 263.605 23.225 ;
    RECT 260.005 22.345 260.285 23.225 ;
    RECT 256.685 22.345 256.965 23.225 ;
    RECT 253.365 22.345 253.645 23.225 ;
    RECT 250.045 61.965 250.325 62.845 ;
    RECT 246.725 61.965 247.005 62.845 ;
    RECT 243.405 61.965 243.685 62.845 ;
    RECT 240.085 61.965 240.365 62.845 ;
    RECT 236.765 61.965 237.045 62.845 ;
    RECT 233.445 61.965 233.725 62.845 ;
    RECT 230.125 61.965 230.405 62.845 ;
    RECT 226.805 61.965 227.085 62.845 ;
    RECT 223.485 61.965 223.765 62.845 ;
    RECT 220.165 61.965 220.445 62.845 ;
    RECT 216.845 61.965 217.125 62.845 ;
    RECT 180.325 61.965 180.605 62.845 ;
    RECT 177.005 61.965 177.285 62.845 ;
    RECT 173.685 61.965 173.965 62.845 ;
    RECT 170.365 61.965 170.645 62.845 ;
    RECT 167.045 61.965 167.325 62.845 ;
    RECT 163.725 61.965 164.005 62.845 ;
    RECT 160.405 61.965 160.685 62.845 ;
    RECT 157.085 61.965 157.365 62.845 ;
    RECT 153.765 61.965 154.045 62.845 ;
    RECT 150.445 61.965 150.725 62.845 ;
    RECT 213.525 61.965 213.805 62.845 ;
    RECT 210.205 61.965 210.485 62.845 ;
    RECT 206.885 61.965 207.165 62.845 ;
    RECT 203.565 61.965 203.845 62.845 ;
    RECT 200.245 61.965 200.525 62.845 ;
    RECT 196.925 61.965 197.205 62.845 ;
    RECT 193.605 61.965 193.885 62.845 ;
    RECT 190.285 61.965 190.565 62.845 ;
    RECT 186.965 61.965 187.245 62.845 ;
    RECT 183.645 61.965 183.925 62.845 ;
    RECT 266.645 61.965 266.925 62.845 ;
    RECT 263.325 61.965 263.605 62.845 ;
    RECT 260.005 61.965 260.285 62.845 ;
    RECT 256.685 61.965 256.965 62.845 ;
    RECT 253.365 61.965 253.645 62.845 ;
    RECT 250.045 97.245 250.325 98.125 ;
    RECT 246.725 97.245 247.005 98.125 ;
    RECT 243.405 97.245 243.685 98.125 ;
    RECT 240.085 97.245 240.365 98.125 ;
    RECT 236.765 97.245 237.045 98.125 ;
    RECT 233.445 97.245 233.725 98.125 ;
    RECT 230.125 97.245 230.405 98.125 ;
    RECT 226.805 97.245 227.085 98.125 ;
    RECT 223.485 97.245 223.765 98.125 ;
    RECT 220.165 97.245 220.445 98.125 ;
    RECT 216.845 97.245 217.125 98.125 ;
    RECT 180.325 97.245 180.605 98.125 ;
    RECT 177.005 97.245 177.285 98.125 ;
    RECT 173.685 97.245 173.965 98.125 ;
    RECT 170.365 97.245 170.645 98.125 ;
    RECT 167.045 97.245 167.325 98.125 ;
    RECT 163.725 97.245 164.005 98.125 ;
    RECT 160.405 97.245 160.685 98.125 ;
    RECT 157.085 97.245 157.365 98.125 ;
    RECT 153.765 97.245 154.045 98.125 ;
    RECT 150.445 97.245 150.725 98.125 ;
    RECT 213.525 97.245 213.805 98.125 ;
    RECT 210.205 97.245 210.485 98.125 ;
    RECT 206.885 97.245 207.165 98.125 ;
    RECT 203.565 97.245 203.845 98.125 ;
    RECT 200.245 97.245 200.525 98.125 ;
    RECT 196.925 97.245 197.205 98.125 ;
    RECT 193.605 97.245 193.885 98.125 ;
    RECT 190.285 97.245 190.565 98.125 ;
    RECT 186.965 97.245 187.245 98.125 ;
    RECT 183.645 97.245 183.925 98.125 ;
    RECT 266.645 97.245 266.925 98.125 ;
    RECT 263.325 97.245 263.605 98.125 ;
    RECT 260.005 97.245 260.285 98.125 ;
    RECT 256.685 97.245 256.965 98.125 ;
    RECT 253.365 97.245 253.645 98.125 ;
    RECT 250.045 21.625 250.325 22.505 ;
    RECT 246.725 21.625 247.005 22.505 ;
    RECT 243.405 21.625 243.685 22.505 ;
    RECT 240.085 21.625 240.365 22.505 ;
    RECT 236.765 21.625 237.045 22.505 ;
    RECT 233.445 21.625 233.725 22.505 ;
    RECT 230.125 21.625 230.405 22.505 ;
    RECT 226.805 21.625 227.085 22.505 ;
    RECT 223.485 21.625 223.765 22.505 ;
    RECT 220.165 21.625 220.445 22.505 ;
    RECT 216.845 21.625 217.125 22.505 ;
    RECT 180.325 21.625 180.605 22.505 ;
    RECT 177.005 21.625 177.285 22.505 ;
    RECT 173.685 21.625 173.965 22.505 ;
    RECT 170.365 21.625 170.645 22.505 ;
    RECT 167.045 21.625 167.325 22.505 ;
    RECT 163.725 21.625 164.005 22.505 ;
    RECT 160.405 21.625 160.685 22.505 ;
    RECT 157.085 21.625 157.365 22.505 ;
    RECT 153.765 21.625 154.045 22.505 ;
    RECT 150.445 21.625 150.725 22.505 ;
    RECT 213.525 21.625 213.805 22.505 ;
    RECT 210.205 21.625 210.485 22.505 ;
    RECT 206.885 21.625 207.165 22.505 ;
    RECT 203.565 21.625 203.845 22.505 ;
    RECT 200.245 21.625 200.525 22.505 ;
    RECT 196.925 21.625 197.205 22.505 ;
    RECT 193.605 21.625 193.885 22.505 ;
    RECT 190.285 21.625 190.565 22.505 ;
    RECT 186.965 21.625 187.245 22.505 ;
    RECT 183.645 21.625 183.925 22.505 ;
    RECT 266.645 21.625 266.925 22.505 ;
    RECT 263.325 21.625 263.605 22.505 ;
    RECT 260.005 21.625 260.285 22.505 ;
    RECT 256.685 21.625 256.965 22.505 ;
    RECT 253.365 21.625 253.645 22.505 ;
    RECT 250.045 61.245 250.325 62.125 ;
    RECT 246.725 61.245 247.005 62.125 ;
    RECT 243.405 61.245 243.685 62.125 ;
    RECT 240.085 61.245 240.365 62.125 ;
    RECT 236.765 61.245 237.045 62.125 ;
    RECT 233.445 61.245 233.725 62.125 ;
    RECT 230.125 61.245 230.405 62.125 ;
    RECT 226.805 61.245 227.085 62.125 ;
    RECT 223.485 61.245 223.765 62.125 ;
    RECT 220.165 61.245 220.445 62.125 ;
    RECT 216.845 61.245 217.125 62.125 ;
    RECT 180.325 61.245 180.605 62.125 ;
    RECT 177.005 61.245 177.285 62.125 ;
    RECT 173.685 61.245 173.965 62.125 ;
    RECT 170.365 61.245 170.645 62.125 ;
    RECT 167.045 61.245 167.325 62.125 ;
    RECT 163.725 61.245 164.005 62.125 ;
    RECT 160.405 61.245 160.685 62.125 ;
    RECT 157.085 61.245 157.365 62.125 ;
    RECT 153.765 61.245 154.045 62.125 ;
    RECT 150.445 61.245 150.725 62.125 ;
    RECT 213.525 61.245 213.805 62.125 ;
    RECT 210.205 61.245 210.485 62.125 ;
    RECT 206.885 61.245 207.165 62.125 ;
    RECT 203.565 61.245 203.845 62.125 ;
    RECT 200.245 61.245 200.525 62.125 ;
    RECT 196.925 61.245 197.205 62.125 ;
    RECT 193.605 61.245 193.885 62.125 ;
    RECT 190.285 61.245 190.565 62.125 ;
    RECT 186.965 61.245 187.245 62.125 ;
    RECT 183.645 61.245 183.925 62.125 ;
    RECT 266.645 61.245 266.925 62.125 ;
    RECT 263.325 61.245 263.605 62.125 ;
    RECT 260.005 61.245 260.285 62.125 ;
    RECT 256.685 61.245 256.965 62.125 ;
    RECT 253.365 61.245 253.645 62.125 ;
    RECT 180.325 60.585 180.605 61.325 ;
    RECT 177.005 60.585 177.285 61.325 ;
    RECT 173.685 60.585 173.965 61.325 ;
    RECT 170.365 60.585 170.645 61.325 ;
    RECT 167.045 60.585 167.325 61.325 ;
    RECT 163.725 60.585 164.005 61.325 ;
    RECT 160.405 60.585 160.685 61.325 ;
    RECT 157.085 60.585 157.365 61.325 ;
    RECT 153.765 60.585 154.045 61.325 ;
    RECT 150.445 60.585 150.725 61.325 ;
    RECT 266.645 60.585 266.925 61.325 ;
    RECT 263.325 60.585 263.605 61.325 ;
    RECT 260.005 60.585 260.285 61.325 ;
    RECT 256.685 60.585 256.965 61.325 ;
    RECT 253.365 60.585 253.645 61.325 ;
    RECT 250.045 60.585 250.325 61.325 ;
    RECT 246.725 60.585 247.005 61.325 ;
    RECT 243.405 60.585 243.685 61.325 ;
    RECT 240.085 60.585 240.365 61.325 ;
    RECT 236.765 60.585 237.045 61.325 ;
    RECT 233.445 60.585 233.725 61.325 ;
    RECT 230.125 60.585 230.405 61.325 ;
    RECT 226.805 60.585 227.085 61.325 ;
    RECT 223.485 60.585 223.765 61.325 ;
    RECT 220.165 60.585 220.445 61.325 ;
    RECT 216.845 60.585 217.125 61.325 ;
    RECT 213.525 60.585 213.805 61.325 ;
    RECT 210.205 60.585 210.485 61.325 ;
    RECT 206.885 60.585 207.165 61.325 ;
    RECT 203.565 60.585 203.845 61.325 ;
    RECT 200.245 60.585 200.525 61.325 ;
    RECT 196.925 60.585 197.205 61.325 ;
    RECT 193.605 60.585 193.885 61.325 ;
    RECT 190.285 60.585 190.565 61.325 ;
    RECT 186.965 60.585 187.245 61.325 ;
    RECT 183.645 60.585 183.925 61.325 ;
    RECT 250.045 96.525 250.325 97.405 ;
    RECT 246.725 96.525 247.005 97.405 ;
    RECT 243.405 96.525 243.685 97.405 ;
    RECT 240.085 96.525 240.365 97.405 ;
    RECT 236.765 96.525 237.045 97.405 ;
    RECT 233.445 96.525 233.725 97.405 ;
    RECT 230.125 96.525 230.405 97.405 ;
    RECT 226.805 96.525 227.085 97.405 ;
    RECT 223.485 96.525 223.765 97.405 ;
    RECT 220.165 96.525 220.445 97.405 ;
    RECT 216.845 96.525 217.125 97.405 ;
    RECT 180.325 96.525 180.605 97.405 ;
    RECT 177.005 96.525 177.285 97.405 ;
    RECT 173.685 96.525 173.965 97.405 ;
    RECT 170.365 96.525 170.645 97.405 ;
    RECT 167.045 96.525 167.325 97.405 ;
    RECT 163.725 96.525 164.005 97.405 ;
    RECT 160.405 96.525 160.685 97.405 ;
    RECT 157.085 96.525 157.365 97.405 ;
    RECT 153.765 96.525 154.045 97.405 ;
    RECT 150.445 96.525 150.725 97.405 ;
    RECT 213.525 96.525 213.805 97.405 ;
    RECT 210.205 96.525 210.485 97.405 ;
    RECT 206.885 96.525 207.165 97.405 ;
    RECT 203.565 96.525 203.845 97.405 ;
    RECT 200.245 96.525 200.525 97.405 ;
    RECT 196.925 96.525 197.205 97.405 ;
    RECT 193.605 96.525 193.885 97.405 ;
    RECT 190.285 96.525 190.565 97.405 ;
    RECT 186.965 96.525 187.245 97.405 ;
    RECT 183.645 96.525 183.925 97.405 ;
    RECT 266.645 96.525 266.925 97.405 ;
    RECT 263.325 96.525 263.605 97.405 ;
    RECT 260.005 96.525 260.285 97.405 ;
    RECT 256.685 96.525 256.965 97.405 ;
    RECT 253.365 96.525 253.645 97.405 ;
    RECT 250.045 59.785 250.325 60.665 ;
    RECT 246.725 59.785 247.005 60.665 ;
    RECT 243.405 59.785 243.685 60.665 ;
    RECT 240.085 59.785 240.365 60.665 ;
    RECT 236.765 59.785 237.045 60.665 ;
    RECT 233.445 59.785 233.725 60.665 ;
    RECT 230.125 59.785 230.405 60.665 ;
    RECT 226.805 59.785 227.085 60.665 ;
    RECT 223.485 59.785 223.765 60.665 ;
    RECT 220.165 59.785 220.445 60.665 ;
    RECT 216.845 59.785 217.125 60.665 ;
    RECT 180.325 59.785 180.605 60.665 ;
    RECT 177.005 59.785 177.285 60.665 ;
    RECT 173.685 59.785 173.965 60.665 ;
    RECT 170.365 59.785 170.645 60.665 ;
    RECT 167.045 59.785 167.325 60.665 ;
    RECT 163.725 59.785 164.005 60.665 ;
    RECT 160.405 59.785 160.685 60.665 ;
    RECT 157.085 59.785 157.365 60.665 ;
    RECT 153.765 59.785 154.045 60.665 ;
    RECT 150.445 59.785 150.725 60.665 ;
    RECT 213.525 59.785 213.805 60.665 ;
    RECT 210.205 59.785 210.485 60.665 ;
    RECT 206.885 59.785 207.165 60.665 ;
    RECT 203.565 59.785 203.845 60.665 ;
    RECT 200.245 59.785 200.525 60.665 ;
    RECT 196.925 59.785 197.205 60.665 ;
    RECT 193.605 59.785 193.885 60.665 ;
    RECT 190.285 59.785 190.565 60.665 ;
    RECT 186.965 59.785 187.245 60.665 ;
    RECT 183.645 59.785 183.925 60.665 ;
    RECT 266.645 59.785 266.925 60.665 ;
    RECT 263.325 59.785 263.605 60.665 ;
    RECT 260.005 59.785 260.285 60.665 ;
    RECT 256.685 59.785 256.965 60.665 ;
    RECT 253.365 59.785 253.645 60.665 ;
    RECT 250.045 95.805 250.325 96.685 ;
    RECT 246.725 95.805 247.005 96.685 ;
    RECT 243.405 95.805 243.685 96.685 ;
    RECT 240.085 95.805 240.365 96.685 ;
    RECT 236.765 95.805 237.045 96.685 ;
    RECT 233.445 95.805 233.725 96.685 ;
    RECT 230.125 95.805 230.405 96.685 ;
    RECT 226.805 95.805 227.085 96.685 ;
    RECT 223.485 95.805 223.765 96.685 ;
    RECT 220.165 95.805 220.445 96.685 ;
    RECT 216.845 95.805 217.125 96.685 ;
    RECT 180.325 95.805 180.605 96.685 ;
    RECT 177.005 95.805 177.285 96.685 ;
    RECT 173.685 95.805 173.965 96.685 ;
    RECT 170.365 95.805 170.645 96.685 ;
    RECT 167.045 95.805 167.325 96.685 ;
    RECT 163.725 95.805 164.005 96.685 ;
    RECT 160.405 95.805 160.685 96.685 ;
    RECT 157.085 95.805 157.365 96.685 ;
    RECT 153.765 95.805 154.045 96.685 ;
    RECT 150.445 95.805 150.725 96.685 ;
    RECT 213.525 95.805 213.805 96.685 ;
    RECT 210.205 95.805 210.485 96.685 ;
    RECT 206.885 95.805 207.165 96.685 ;
    RECT 203.565 95.805 203.845 96.685 ;
    RECT 200.245 95.805 200.525 96.685 ;
    RECT 196.925 95.805 197.205 96.685 ;
    RECT 193.605 95.805 193.885 96.685 ;
    RECT 190.285 95.805 190.565 96.685 ;
    RECT 186.965 95.805 187.245 96.685 ;
    RECT 183.645 95.805 183.925 96.685 ;
    RECT 266.645 95.805 266.925 96.685 ;
    RECT 263.325 95.805 263.605 96.685 ;
    RECT 260.005 95.805 260.285 96.685 ;
    RECT 256.685 95.805 256.965 96.685 ;
    RECT 253.365 95.805 253.645 96.685 ;
    RECT 250.045 59.065 250.325 59.945 ;
    RECT 246.725 59.065 247.005 59.945 ;
    RECT 243.405 59.065 243.685 59.945 ;
    RECT 240.085 59.065 240.365 59.945 ;
    RECT 236.765 59.065 237.045 59.945 ;
    RECT 233.445 59.065 233.725 59.945 ;
    RECT 230.125 59.065 230.405 59.945 ;
    RECT 226.805 59.065 227.085 59.945 ;
    RECT 223.485 59.065 223.765 59.945 ;
    RECT 220.165 59.065 220.445 59.945 ;
    RECT 216.845 59.065 217.125 59.945 ;
    RECT 180.325 59.065 180.605 59.945 ;
    RECT 177.005 59.065 177.285 59.945 ;
    RECT 173.685 59.065 173.965 59.945 ;
    RECT 170.365 59.065 170.645 59.945 ;
    RECT 167.045 59.065 167.325 59.945 ;
    RECT 163.725 59.065 164.005 59.945 ;
    RECT 160.405 59.065 160.685 59.945 ;
    RECT 157.085 59.065 157.365 59.945 ;
    RECT 153.765 59.065 154.045 59.945 ;
    RECT 150.445 59.065 150.725 59.945 ;
    RECT 213.525 59.065 213.805 59.945 ;
    RECT 210.205 59.065 210.485 59.945 ;
    RECT 206.885 59.065 207.165 59.945 ;
    RECT 203.565 59.065 203.845 59.945 ;
    RECT 200.245 59.065 200.525 59.945 ;
    RECT 196.925 59.065 197.205 59.945 ;
    RECT 193.605 59.065 193.885 59.945 ;
    RECT 190.285 59.065 190.565 59.945 ;
    RECT 186.965 59.065 187.245 59.945 ;
    RECT 183.645 59.065 183.925 59.945 ;
    RECT 266.645 59.065 266.925 59.945 ;
    RECT 263.325 59.065 263.605 59.945 ;
    RECT 260.005 59.065 260.285 59.945 ;
    RECT 256.685 59.065 256.965 59.945 ;
    RECT 253.365 59.065 253.645 59.945 ;
    RECT 250.045 95.085 250.325 95.965 ;
    RECT 246.725 95.085 247.005 95.965 ;
    RECT 243.405 95.085 243.685 95.965 ;
    RECT 240.085 95.085 240.365 95.965 ;
    RECT 236.765 95.085 237.045 95.965 ;
    RECT 233.445 95.085 233.725 95.965 ;
    RECT 230.125 95.085 230.405 95.965 ;
    RECT 226.805 95.085 227.085 95.965 ;
    RECT 223.485 95.085 223.765 95.965 ;
    RECT 220.165 95.085 220.445 95.965 ;
    RECT 216.845 95.085 217.125 95.965 ;
    RECT 180.325 95.085 180.605 95.965 ;
    RECT 177.005 95.085 177.285 95.965 ;
    RECT 173.685 95.085 173.965 95.965 ;
    RECT 170.365 95.085 170.645 95.965 ;
    RECT 167.045 95.085 167.325 95.965 ;
    RECT 163.725 95.085 164.005 95.965 ;
    RECT 160.405 95.085 160.685 95.965 ;
    RECT 157.085 95.085 157.365 95.965 ;
    RECT 153.765 95.085 154.045 95.965 ;
    RECT 150.445 95.085 150.725 95.965 ;
    RECT 213.525 95.085 213.805 95.965 ;
    RECT 210.205 95.085 210.485 95.965 ;
    RECT 206.885 95.085 207.165 95.965 ;
    RECT 203.565 95.085 203.845 95.965 ;
    RECT 200.245 95.085 200.525 95.965 ;
    RECT 196.925 95.085 197.205 95.965 ;
    RECT 193.605 95.085 193.885 95.965 ;
    RECT 190.285 95.085 190.565 95.965 ;
    RECT 186.965 95.085 187.245 95.965 ;
    RECT 183.645 95.085 183.925 95.965 ;
    RECT 266.645 95.085 266.925 95.965 ;
    RECT 263.325 95.085 263.605 95.965 ;
    RECT 260.005 95.085 260.285 95.965 ;
    RECT 256.685 95.085 256.965 95.965 ;
    RECT 253.365 95.085 253.645 95.965 ;
    RECT 250.045 58.345 250.325 59.225 ;
    RECT 246.725 58.345 247.005 59.225 ;
    RECT 243.405 58.345 243.685 59.225 ;
    RECT 240.085 58.345 240.365 59.225 ;
    RECT 236.765 58.345 237.045 59.225 ;
    RECT 233.445 58.345 233.725 59.225 ;
    RECT 230.125 58.345 230.405 59.225 ;
    RECT 226.805 58.345 227.085 59.225 ;
    RECT 223.485 58.345 223.765 59.225 ;
    RECT 220.165 58.345 220.445 59.225 ;
    RECT 216.845 58.345 217.125 59.225 ;
    RECT 180.325 58.345 180.605 59.225 ;
    RECT 177.005 58.345 177.285 59.225 ;
    RECT 173.685 58.345 173.965 59.225 ;
    RECT 170.365 58.345 170.645 59.225 ;
    RECT 167.045 58.345 167.325 59.225 ;
    RECT 163.725 58.345 164.005 59.225 ;
    RECT 160.405 58.345 160.685 59.225 ;
    RECT 157.085 58.345 157.365 59.225 ;
    RECT 153.765 58.345 154.045 59.225 ;
    RECT 150.445 58.345 150.725 59.225 ;
    RECT 213.525 58.345 213.805 59.225 ;
    RECT 210.205 58.345 210.485 59.225 ;
    RECT 206.885 58.345 207.165 59.225 ;
    RECT 203.565 58.345 203.845 59.225 ;
    RECT 200.245 58.345 200.525 59.225 ;
    RECT 196.925 58.345 197.205 59.225 ;
    RECT 193.605 58.345 193.885 59.225 ;
    RECT 190.285 58.345 190.565 59.225 ;
    RECT 186.965 58.345 187.245 59.225 ;
    RECT 183.645 58.345 183.925 59.225 ;
    RECT 266.645 58.345 266.925 59.225 ;
    RECT 263.325 58.345 263.605 59.225 ;
    RECT 260.005 58.345 260.285 59.225 ;
    RECT 256.685 58.345 256.965 59.225 ;
    RECT 253.365 58.345 253.645 59.225 ;
    RECT 250.045 94.365 250.325 95.245 ;
    RECT 246.725 94.365 247.005 95.245 ;
    RECT 243.405 94.365 243.685 95.245 ;
    RECT 240.085 94.365 240.365 95.245 ;
    RECT 236.765 94.365 237.045 95.245 ;
    RECT 233.445 94.365 233.725 95.245 ;
    RECT 230.125 94.365 230.405 95.245 ;
    RECT 226.805 94.365 227.085 95.245 ;
    RECT 223.485 94.365 223.765 95.245 ;
    RECT 220.165 94.365 220.445 95.245 ;
    RECT 216.845 94.365 217.125 95.245 ;
    RECT 180.325 94.365 180.605 95.245 ;
    RECT 177.005 94.365 177.285 95.245 ;
    RECT 173.685 94.365 173.965 95.245 ;
    RECT 170.365 94.365 170.645 95.245 ;
    RECT 167.045 94.365 167.325 95.245 ;
    RECT 163.725 94.365 164.005 95.245 ;
    RECT 160.405 94.365 160.685 95.245 ;
    RECT 157.085 94.365 157.365 95.245 ;
    RECT 153.765 94.365 154.045 95.245 ;
    RECT 150.445 94.365 150.725 95.245 ;
    RECT 213.525 94.365 213.805 95.245 ;
    RECT 210.205 94.365 210.485 95.245 ;
    RECT 206.885 94.365 207.165 95.245 ;
    RECT 203.565 94.365 203.845 95.245 ;
    RECT 200.245 94.365 200.525 95.245 ;
    RECT 196.925 94.365 197.205 95.245 ;
    RECT 193.605 94.365 193.885 95.245 ;
    RECT 190.285 94.365 190.565 95.245 ;
    RECT 186.965 94.365 187.245 95.245 ;
    RECT 183.645 94.365 183.925 95.245 ;
    RECT 266.645 94.365 266.925 95.245 ;
    RECT 263.325 94.365 263.605 95.245 ;
    RECT 260.005 94.365 260.285 95.245 ;
    RECT 256.685 94.365 256.965 95.245 ;
    RECT 253.365 94.365 253.645 95.245 ;
    RECT 250.045 57.625 250.325 58.505 ;
    RECT 246.725 57.625 247.005 58.505 ;
    RECT 243.405 57.625 243.685 58.505 ;
    RECT 240.085 57.625 240.365 58.505 ;
    RECT 236.765 57.625 237.045 58.505 ;
    RECT 233.445 57.625 233.725 58.505 ;
    RECT 230.125 57.625 230.405 58.505 ;
    RECT 226.805 57.625 227.085 58.505 ;
    RECT 223.485 57.625 223.765 58.505 ;
    RECT 220.165 57.625 220.445 58.505 ;
    RECT 216.845 57.625 217.125 58.505 ;
    RECT 180.325 57.625 180.605 58.505 ;
    RECT 177.005 57.625 177.285 58.505 ;
    RECT 173.685 57.625 173.965 58.505 ;
    RECT 170.365 57.625 170.645 58.505 ;
    RECT 167.045 57.625 167.325 58.505 ;
    RECT 163.725 57.625 164.005 58.505 ;
    RECT 160.405 57.625 160.685 58.505 ;
    RECT 157.085 57.625 157.365 58.505 ;
    RECT 153.765 57.625 154.045 58.505 ;
    RECT 150.445 57.625 150.725 58.505 ;
    RECT 213.525 57.625 213.805 58.505 ;
    RECT 210.205 57.625 210.485 58.505 ;
    RECT 206.885 57.625 207.165 58.505 ;
    RECT 203.565 57.625 203.845 58.505 ;
    RECT 200.245 57.625 200.525 58.505 ;
    RECT 196.925 57.625 197.205 58.505 ;
    RECT 193.605 57.625 193.885 58.505 ;
    RECT 190.285 57.625 190.565 58.505 ;
    RECT 186.965 57.625 187.245 58.505 ;
    RECT 183.645 57.625 183.925 58.505 ;
    RECT 266.645 57.625 266.925 58.505 ;
    RECT 263.325 57.625 263.605 58.505 ;
    RECT 260.005 57.625 260.285 58.505 ;
    RECT 256.685 57.625 256.965 58.505 ;
    RECT 253.365 57.625 253.645 58.505 ;
    RECT 250.045 93.645 250.325 94.525 ;
    RECT 246.725 93.645 247.005 94.525 ;
    RECT 243.405 93.645 243.685 94.525 ;
    RECT 240.085 93.645 240.365 94.525 ;
    RECT 236.765 93.645 237.045 94.525 ;
    RECT 233.445 93.645 233.725 94.525 ;
    RECT 230.125 93.645 230.405 94.525 ;
    RECT 226.805 93.645 227.085 94.525 ;
    RECT 223.485 93.645 223.765 94.525 ;
    RECT 220.165 93.645 220.445 94.525 ;
    RECT 216.845 93.645 217.125 94.525 ;
    RECT 180.325 93.645 180.605 94.525 ;
    RECT 177.005 93.645 177.285 94.525 ;
    RECT 173.685 93.645 173.965 94.525 ;
    RECT 170.365 93.645 170.645 94.525 ;
    RECT 167.045 93.645 167.325 94.525 ;
    RECT 163.725 93.645 164.005 94.525 ;
    RECT 160.405 93.645 160.685 94.525 ;
    RECT 157.085 93.645 157.365 94.525 ;
    RECT 153.765 93.645 154.045 94.525 ;
    RECT 150.445 93.645 150.725 94.525 ;
    RECT 213.525 93.645 213.805 94.525 ;
    RECT 210.205 93.645 210.485 94.525 ;
    RECT 206.885 93.645 207.165 94.525 ;
    RECT 203.565 93.645 203.845 94.525 ;
    RECT 200.245 93.645 200.525 94.525 ;
    RECT 196.925 93.645 197.205 94.525 ;
    RECT 193.605 93.645 193.885 94.525 ;
    RECT 190.285 93.645 190.565 94.525 ;
    RECT 186.965 93.645 187.245 94.525 ;
    RECT 183.645 93.645 183.925 94.525 ;
    RECT 266.645 93.645 266.925 94.525 ;
    RECT 263.325 93.645 263.605 94.525 ;
    RECT 260.005 93.645 260.285 94.525 ;
    RECT 256.685 93.645 256.965 94.525 ;
    RECT 253.365 93.645 253.645 94.525 ;
    RECT 250.045 56.905 250.325 57.785 ;
    RECT 246.725 56.905 247.005 57.785 ;
    RECT 243.405 56.905 243.685 57.785 ;
    RECT 240.085 56.905 240.365 57.785 ;
    RECT 236.765 56.905 237.045 57.785 ;
    RECT 233.445 56.905 233.725 57.785 ;
    RECT 230.125 56.905 230.405 57.785 ;
    RECT 226.805 56.905 227.085 57.785 ;
    RECT 223.485 56.905 223.765 57.785 ;
    RECT 220.165 56.905 220.445 57.785 ;
    RECT 216.845 56.905 217.125 57.785 ;
    RECT 180.325 56.905 180.605 57.785 ;
    RECT 177.005 56.905 177.285 57.785 ;
    RECT 173.685 56.905 173.965 57.785 ;
    RECT 170.365 56.905 170.645 57.785 ;
    RECT 167.045 56.905 167.325 57.785 ;
    RECT 163.725 56.905 164.005 57.785 ;
    RECT 160.405 56.905 160.685 57.785 ;
    RECT 157.085 56.905 157.365 57.785 ;
    RECT 153.765 56.905 154.045 57.785 ;
    RECT 150.445 56.905 150.725 57.785 ;
    RECT 213.525 56.905 213.805 57.785 ;
    RECT 210.205 56.905 210.485 57.785 ;
    RECT 206.885 56.905 207.165 57.785 ;
    RECT 203.565 56.905 203.845 57.785 ;
    RECT 200.245 56.905 200.525 57.785 ;
    RECT 196.925 56.905 197.205 57.785 ;
    RECT 193.605 56.905 193.885 57.785 ;
    RECT 190.285 56.905 190.565 57.785 ;
    RECT 186.965 56.905 187.245 57.785 ;
    RECT 183.645 56.905 183.925 57.785 ;
    RECT 266.645 56.905 266.925 57.785 ;
    RECT 263.325 56.905 263.605 57.785 ;
    RECT 260.005 56.905 260.285 57.785 ;
    RECT 256.685 56.905 256.965 57.785 ;
    RECT 253.365 56.905 253.645 57.785 ;
    RECT 250.045 92.925 250.325 93.805 ;
    RECT 246.725 92.925 247.005 93.805 ;
    RECT 243.405 92.925 243.685 93.805 ;
    RECT 240.085 92.925 240.365 93.805 ;
    RECT 236.765 92.925 237.045 93.805 ;
    RECT 233.445 92.925 233.725 93.805 ;
    RECT 230.125 92.925 230.405 93.805 ;
    RECT 226.805 92.925 227.085 93.805 ;
    RECT 223.485 92.925 223.765 93.805 ;
    RECT 220.165 92.925 220.445 93.805 ;
    RECT 216.845 92.925 217.125 93.805 ;
    RECT 180.325 92.925 180.605 93.805 ;
    RECT 177.005 92.925 177.285 93.805 ;
    RECT 173.685 92.925 173.965 93.805 ;
    RECT 170.365 92.925 170.645 93.805 ;
    RECT 167.045 92.925 167.325 93.805 ;
    RECT 163.725 92.925 164.005 93.805 ;
    RECT 160.405 92.925 160.685 93.805 ;
    RECT 157.085 92.925 157.365 93.805 ;
    RECT 153.765 92.925 154.045 93.805 ;
    RECT 150.445 92.925 150.725 93.805 ;
    RECT 213.525 92.925 213.805 93.805 ;
    RECT 210.205 92.925 210.485 93.805 ;
    RECT 206.885 92.925 207.165 93.805 ;
    RECT 203.565 92.925 203.845 93.805 ;
    RECT 200.245 92.925 200.525 93.805 ;
    RECT 196.925 92.925 197.205 93.805 ;
    RECT 193.605 92.925 193.885 93.805 ;
    RECT 190.285 92.925 190.565 93.805 ;
    RECT 186.965 92.925 187.245 93.805 ;
    RECT 183.645 92.925 183.925 93.805 ;
    RECT 266.645 92.925 266.925 93.805 ;
    RECT 263.325 92.925 263.605 93.805 ;
    RECT 260.005 92.925 260.285 93.805 ;
    RECT 256.685 92.925 256.965 93.805 ;
    RECT 253.365 92.925 253.645 93.805 ;
    RECT 250.045 92.205 250.325 93.085 ;
    RECT 246.725 92.205 247.005 93.085 ;
    RECT 243.405 92.205 243.685 93.085 ;
    RECT 240.085 92.205 240.365 93.085 ;
    RECT 236.765 92.205 237.045 93.085 ;
    RECT 233.445 92.205 233.725 93.085 ;
    RECT 230.125 92.205 230.405 93.085 ;
    RECT 226.805 92.205 227.085 93.085 ;
    RECT 223.485 92.205 223.765 93.085 ;
    RECT 220.165 92.205 220.445 93.085 ;
    RECT 216.845 92.205 217.125 93.085 ;
    RECT 180.325 92.205 180.605 93.085 ;
    RECT 177.005 92.205 177.285 93.085 ;
    RECT 173.685 92.205 173.965 93.085 ;
    RECT 170.365 92.205 170.645 93.085 ;
    RECT 167.045 92.205 167.325 93.085 ;
    RECT 163.725 92.205 164.005 93.085 ;
    RECT 160.405 92.205 160.685 93.085 ;
    RECT 157.085 92.205 157.365 93.085 ;
    RECT 153.765 92.205 154.045 93.085 ;
    RECT 150.445 92.205 150.725 93.085 ;
    RECT 213.525 92.205 213.805 93.085 ;
    RECT 210.205 92.205 210.485 93.085 ;
    RECT 206.885 92.205 207.165 93.085 ;
    RECT 203.565 92.205 203.845 93.085 ;
    RECT 200.245 92.205 200.525 93.085 ;
    RECT 196.925 92.205 197.205 93.085 ;
    RECT 193.605 92.205 193.885 93.085 ;
    RECT 190.285 92.205 190.565 93.085 ;
    RECT 186.965 92.205 187.245 93.085 ;
    RECT 183.645 92.205 183.925 93.085 ;
    RECT 266.645 92.205 266.925 93.085 ;
    RECT 263.325 92.205 263.605 93.085 ;
    RECT 260.005 92.205 260.285 93.085 ;
    RECT 256.685 92.205 256.965 93.085 ;
    RECT 253.365 92.205 253.645 93.085 ;
    RECT 250.045 91.485 250.325 92.365 ;
    RECT 246.725 91.485 247.005 92.365 ;
    RECT 243.405 91.485 243.685 92.365 ;
    RECT 240.085 91.485 240.365 92.365 ;
    RECT 236.765 91.485 237.045 92.365 ;
    RECT 233.445 91.485 233.725 92.365 ;
    RECT 230.125 91.485 230.405 92.365 ;
    RECT 226.805 91.485 227.085 92.365 ;
    RECT 223.485 91.485 223.765 92.365 ;
    RECT 220.165 91.485 220.445 92.365 ;
    RECT 216.845 91.485 217.125 92.365 ;
    RECT 180.325 91.485 180.605 92.365 ;
    RECT 177.005 91.485 177.285 92.365 ;
    RECT 173.685 91.485 173.965 92.365 ;
    RECT 170.365 91.485 170.645 92.365 ;
    RECT 167.045 91.485 167.325 92.365 ;
    RECT 163.725 91.485 164.005 92.365 ;
    RECT 160.405 91.485 160.685 92.365 ;
    RECT 157.085 91.485 157.365 92.365 ;
    RECT 153.765 91.485 154.045 92.365 ;
    RECT 150.445 91.485 150.725 92.365 ;
    RECT 213.525 91.485 213.805 92.365 ;
    RECT 210.205 91.485 210.485 92.365 ;
    RECT 206.885 91.485 207.165 92.365 ;
    RECT 203.565 91.485 203.845 92.365 ;
    RECT 200.245 91.485 200.525 92.365 ;
    RECT 196.925 91.485 197.205 92.365 ;
    RECT 193.605 91.485 193.885 92.365 ;
    RECT 190.285 91.485 190.565 92.365 ;
    RECT 186.965 91.485 187.245 92.365 ;
    RECT 183.645 91.485 183.925 92.365 ;
    RECT 266.645 91.485 266.925 92.365 ;
    RECT 263.325 91.485 263.605 92.365 ;
    RECT 260.005 91.485 260.285 92.365 ;
    RECT 256.685 91.485 256.965 92.365 ;
    RECT 253.365 91.485 253.645 92.365 ;
    RECT 250.045 90.765 250.325 91.645 ;
    RECT 246.725 90.765 247.005 91.645 ;
    RECT 243.405 90.765 243.685 91.645 ;
    RECT 240.085 90.765 240.365 91.645 ;
    RECT 236.765 90.765 237.045 91.645 ;
    RECT 233.445 90.765 233.725 91.645 ;
    RECT 230.125 90.765 230.405 91.645 ;
    RECT 226.805 90.765 227.085 91.645 ;
    RECT 223.485 90.765 223.765 91.645 ;
    RECT 220.165 90.765 220.445 91.645 ;
    RECT 216.845 90.765 217.125 91.645 ;
    RECT 180.325 90.765 180.605 91.645 ;
    RECT 177.005 90.765 177.285 91.645 ;
    RECT 173.685 90.765 173.965 91.645 ;
    RECT 170.365 90.765 170.645 91.645 ;
    RECT 167.045 90.765 167.325 91.645 ;
    RECT 163.725 90.765 164.005 91.645 ;
    RECT 160.405 90.765 160.685 91.645 ;
    RECT 157.085 90.765 157.365 91.645 ;
    RECT 153.765 90.765 154.045 91.645 ;
    RECT 150.445 90.765 150.725 91.645 ;
    RECT 213.525 90.765 213.805 91.645 ;
    RECT 210.205 90.765 210.485 91.645 ;
    RECT 206.885 90.765 207.165 91.645 ;
    RECT 203.565 90.765 203.845 91.645 ;
    RECT 200.245 90.765 200.525 91.645 ;
    RECT 196.925 90.765 197.205 91.645 ;
    RECT 193.605 90.765 193.885 91.645 ;
    RECT 190.285 90.765 190.565 91.645 ;
    RECT 186.965 90.765 187.245 91.645 ;
    RECT 183.645 90.765 183.925 91.645 ;
    RECT 266.645 90.765 266.925 91.645 ;
    RECT 263.325 90.765 263.605 91.645 ;
    RECT 260.005 90.765 260.285 91.645 ;
    RECT 256.685 90.765 256.965 91.645 ;
    RECT 253.365 90.765 253.645 91.645 ;
    RECT 250.045 54.025 250.325 54.905 ;
    RECT 246.725 54.025 247.005 54.905 ;
    RECT 243.405 54.025 243.685 54.905 ;
    RECT 240.085 54.025 240.365 54.905 ;
    RECT 236.765 54.025 237.045 54.905 ;
    RECT 233.445 54.025 233.725 54.905 ;
    RECT 230.125 54.025 230.405 54.905 ;
    RECT 226.805 54.025 227.085 54.905 ;
    RECT 223.485 54.025 223.765 54.905 ;
    RECT 220.165 54.025 220.445 54.905 ;
    RECT 216.845 54.025 217.125 54.905 ;
    RECT 180.325 54.025 180.605 54.905 ;
    RECT 177.005 54.025 177.285 54.905 ;
    RECT 173.685 54.025 173.965 54.905 ;
    RECT 170.365 54.025 170.645 54.905 ;
    RECT 167.045 54.025 167.325 54.905 ;
    RECT 163.725 54.025 164.005 54.905 ;
    RECT 160.405 54.025 160.685 54.905 ;
    RECT 157.085 54.025 157.365 54.905 ;
    RECT 153.765 54.025 154.045 54.905 ;
    RECT 150.445 54.025 150.725 54.905 ;
    RECT 213.525 54.025 213.805 54.905 ;
    RECT 210.205 54.025 210.485 54.905 ;
    RECT 206.885 54.025 207.165 54.905 ;
    RECT 203.565 54.025 203.845 54.905 ;
    RECT 200.245 54.025 200.525 54.905 ;
    RECT 196.925 54.025 197.205 54.905 ;
    RECT 193.605 54.025 193.885 54.905 ;
    RECT 190.285 54.025 190.565 54.905 ;
    RECT 186.965 54.025 187.245 54.905 ;
    RECT 183.645 54.025 183.925 54.905 ;
    RECT 266.645 54.025 266.925 54.905 ;
    RECT 263.325 54.025 263.605 54.905 ;
    RECT 260.005 54.025 260.285 54.905 ;
    RECT 256.685 54.025 256.965 54.905 ;
    RECT 253.365 54.025 253.645 54.905 ;
    RECT 250.045 90.045 250.325 90.925 ;
    RECT 246.725 90.045 247.005 90.925 ;
    RECT 243.405 90.045 243.685 90.925 ;
    RECT 240.085 90.045 240.365 90.925 ;
    RECT 236.765 90.045 237.045 90.925 ;
    RECT 233.445 90.045 233.725 90.925 ;
    RECT 230.125 90.045 230.405 90.925 ;
    RECT 226.805 90.045 227.085 90.925 ;
    RECT 223.485 90.045 223.765 90.925 ;
    RECT 220.165 90.045 220.445 90.925 ;
    RECT 216.845 90.045 217.125 90.925 ;
    RECT 180.325 90.045 180.605 90.925 ;
    RECT 177.005 90.045 177.285 90.925 ;
    RECT 173.685 90.045 173.965 90.925 ;
    RECT 170.365 90.045 170.645 90.925 ;
    RECT 167.045 90.045 167.325 90.925 ;
    RECT 163.725 90.045 164.005 90.925 ;
    RECT 160.405 90.045 160.685 90.925 ;
    RECT 157.085 90.045 157.365 90.925 ;
    RECT 153.765 90.045 154.045 90.925 ;
    RECT 150.445 90.045 150.725 90.925 ;
    RECT 213.525 90.045 213.805 90.925 ;
    RECT 210.205 90.045 210.485 90.925 ;
    RECT 206.885 90.045 207.165 90.925 ;
    RECT 203.565 90.045 203.845 90.925 ;
    RECT 200.245 90.045 200.525 90.925 ;
    RECT 196.925 90.045 197.205 90.925 ;
    RECT 193.605 90.045 193.885 90.925 ;
    RECT 190.285 90.045 190.565 90.925 ;
    RECT 186.965 90.045 187.245 90.925 ;
    RECT 183.645 90.045 183.925 90.925 ;
    RECT 266.645 90.045 266.925 90.925 ;
    RECT 263.325 90.045 263.605 90.925 ;
    RECT 260.005 90.045 260.285 90.925 ;
    RECT 256.685 90.045 256.965 90.925 ;
    RECT 253.365 90.045 253.645 90.925 ;
    RECT 250.045 53.305 250.325 54.185 ;
    RECT 246.725 53.305 247.005 54.185 ;
    RECT 243.405 53.305 243.685 54.185 ;
    RECT 240.085 53.305 240.365 54.185 ;
    RECT 236.765 53.305 237.045 54.185 ;
    RECT 233.445 53.305 233.725 54.185 ;
    RECT 230.125 53.305 230.405 54.185 ;
    RECT 226.805 53.305 227.085 54.185 ;
    RECT 223.485 53.305 223.765 54.185 ;
    RECT 220.165 53.305 220.445 54.185 ;
    RECT 216.845 53.305 217.125 54.185 ;
    RECT 180.325 53.305 180.605 54.185 ;
    RECT 177.005 53.305 177.285 54.185 ;
    RECT 173.685 53.305 173.965 54.185 ;
    RECT 170.365 53.305 170.645 54.185 ;
    RECT 167.045 53.305 167.325 54.185 ;
    RECT 163.725 53.305 164.005 54.185 ;
    RECT 160.405 53.305 160.685 54.185 ;
    RECT 157.085 53.305 157.365 54.185 ;
    RECT 153.765 53.305 154.045 54.185 ;
    RECT 150.445 53.305 150.725 54.185 ;
    RECT 213.525 53.305 213.805 54.185 ;
    RECT 210.205 53.305 210.485 54.185 ;
    RECT 206.885 53.305 207.165 54.185 ;
    RECT 203.565 53.305 203.845 54.185 ;
    RECT 200.245 53.305 200.525 54.185 ;
    RECT 196.925 53.305 197.205 54.185 ;
    RECT 193.605 53.305 193.885 54.185 ;
    RECT 190.285 53.305 190.565 54.185 ;
    RECT 186.965 53.305 187.245 54.185 ;
    RECT 183.645 53.305 183.925 54.185 ;
    RECT 266.645 53.305 266.925 54.185 ;
    RECT 263.325 53.305 263.605 54.185 ;
    RECT 260.005 53.305 260.285 54.185 ;
    RECT 256.685 53.305 256.965 54.185 ;
    RECT 253.365 53.305 253.645 54.185 ;
    RECT 250.045 14.425 250.325 15.305 ;
    RECT 246.725 14.425 247.005 15.305 ;
    RECT 243.405 14.425 243.685 15.305 ;
    RECT 240.085 14.425 240.365 15.305 ;
    RECT 236.765 14.425 237.045 15.305 ;
    RECT 233.445 14.425 233.725 15.305 ;
    RECT 230.125 14.425 230.405 15.305 ;
    RECT 226.805 14.425 227.085 15.305 ;
    RECT 223.485 14.425 223.765 15.305 ;
    RECT 220.165 14.425 220.445 15.305 ;
    RECT 216.845 14.425 217.125 15.305 ;
    RECT 180.325 14.425 180.605 15.305 ;
    RECT 177.005 14.425 177.285 15.305 ;
    RECT 173.685 14.425 173.965 15.305 ;
    RECT 170.365 14.425 170.645 15.305 ;
    RECT 167.045 14.425 167.325 15.305 ;
    RECT 163.725 14.425 164.005 15.305 ;
    RECT 160.405 14.425 160.685 15.305 ;
    RECT 157.085 14.425 157.365 15.305 ;
    RECT 153.765 14.425 154.045 15.305 ;
    RECT 213.525 14.425 213.805 15.305 ;
    RECT 210.205 14.425 210.485 15.305 ;
    RECT 266.645 14.425 266.925 15.305 ;
    RECT 206.885 14.425 207.165 15.305 ;
    RECT 203.565 14.425 203.845 15.305 ;
    RECT 200.245 14.425 200.525 15.305 ;
    RECT 196.925 14.425 197.205 15.305 ;
    RECT 193.605 14.425 193.885 15.305 ;
    RECT 190.285 14.425 190.565 15.305 ;
    RECT 150.445 14.425 150.725 15.305 ;
    RECT 186.965 14.425 187.245 15.305 ;
    RECT 183.645 14.425 183.925 15.305 ;
    RECT 263.325 14.425 263.605 15.305 ;
    RECT 260.005 14.425 260.285 15.305 ;
    RECT 256.685 14.425 256.965 15.305 ;
    RECT 253.365 14.425 253.645 15.305 ;
    RECT 250.045 89.325 250.325 90.205 ;
    RECT 246.725 89.325 247.005 90.205 ;
    RECT 243.405 89.325 243.685 90.205 ;
    RECT 240.085 89.325 240.365 90.205 ;
    RECT 236.765 89.325 237.045 90.205 ;
    RECT 233.445 89.325 233.725 90.205 ;
    RECT 230.125 89.325 230.405 90.205 ;
    RECT 226.805 89.325 227.085 90.205 ;
    RECT 223.485 89.325 223.765 90.205 ;
    RECT 220.165 89.325 220.445 90.205 ;
    RECT 216.845 89.325 217.125 90.205 ;
    RECT 180.325 89.325 180.605 90.205 ;
    RECT 177.005 89.325 177.285 90.205 ;
    RECT 173.685 89.325 173.965 90.205 ;
    RECT 170.365 89.325 170.645 90.205 ;
    RECT 167.045 89.325 167.325 90.205 ;
    RECT 163.725 89.325 164.005 90.205 ;
    RECT 160.405 89.325 160.685 90.205 ;
    RECT 157.085 89.325 157.365 90.205 ;
    RECT 153.765 89.325 154.045 90.205 ;
    RECT 150.445 89.325 150.725 90.205 ;
    RECT 213.525 89.325 213.805 90.205 ;
    RECT 210.205 89.325 210.485 90.205 ;
    RECT 206.885 89.325 207.165 90.205 ;
    RECT 203.565 89.325 203.845 90.205 ;
    RECT 200.245 89.325 200.525 90.205 ;
    RECT 196.925 89.325 197.205 90.205 ;
    RECT 193.605 89.325 193.885 90.205 ;
    RECT 190.285 89.325 190.565 90.205 ;
    RECT 186.965 89.325 187.245 90.205 ;
    RECT 183.645 89.325 183.925 90.205 ;
    RECT 266.645 89.325 266.925 90.205 ;
    RECT 263.325 89.325 263.605 90.205 ;
    RECT 260.005 89.325 260.285 90.205 ;
    RECT 256.685 89.325 256.965 90.205 ;
    RECT 253.365 89.325 253.645 90.205 ;
    RECT 250.045 52.585 250.325 53.465 ;
    RECT 246.725 52.585 247.005 53.465 ;
    RECT 243.405 52.585 243.685 53.465 ;
    RECT 240.085 52.585 240.365 53.465 ;
    RECT 236.765 52.585 237.045 53.465 ;
    RECT 233.445 52.585 233.725 53.465 ;
    RECT 230.125 52.585 230.405 53.465 ;
    RECT 226.805 52.585 227.085 53.465 ;
    RECT 223.485 52.585 223.765 53.465 ;
    RECT 220.165 52.585 220.445 53.465 ;
    RECT 216.845 52.585 217.125 53.465 ;
    RECT 180.325 52.585 180.605 53.465 ;
    RECT 177.005 52.585 177.285 53.465 ;
    RECT 173.685 52.585 173.965 53.465 ;
    RECT 170.365 52.585 170.645 53.465 ;
    RECT 167.045 52.585 167.325 53.465 ;
    RECT 163.725 52.585 164.005 53.465 ;
    RECT 160.405 52.585 160.685 53.465 ;
    RECT 157.085 52.585 157.365 53.465 ;
    RECT 153.765 52.585 154.045 53.465 ;
    RECT 150.445 52.585 150.725 53.465 ;
    RECT 213.525 52.585 213.805 53.465 ;
    RECT 210.205 52.585 210.485 53.465 ;
    RECT 206.885 52.585 207.165 53.465 ;
    RECT 203.565 52.585 203.845 53.465 ;
    RECT 200.245 52.585 200.525 53.465 ;
    RECT 196.925 52.585 197.205 53.465 ;
    RECT 193.605 52.585 193.885 53.465 ;
    RECT 190.285 52.585 190.565 53.465 ;
    RECT 186.965 52.585 187.245 53.465 ;
    RECT 183.645 52.585 183.925 53.465 ;
    RECT 266.645 52.585 266.925 53.465 ;
    RECT 263.325 52.585 263.605 53.465 ;
    RECT 260.005 52.585 260.285 53.465 ;
    RECT 256.685 52.585 256.965 53.465 ;
    RECT 253.365 52.585 253.645 53.465 ;
    RECT 250.045 88.605 250.325 89.485 ;
    RECT 246.725 88.605 247.005 89.485 ;
    RECT 243.405 88.605 243.685 89.485 ;
    RECT 240.085 88.605 240.365 89.485 ;
    RECT 236.765 88.605 237.045 89.485 ;
    RECT 233.445 88.605 233.725 89.485 ;
    RECT 230.125 88.605 230.405 89.485 ;
    RECT 226.805 88.605 227.085 89.485 ;
    RECT 223.485 88.605 223.765 89.485 ;
    RECT 220.165 88.605 220.445 89.485 ;
    RECT 216.845 88.605 217.125 89.485 ;
    RECT 180.325 88.605 180.605 89.485 ;
    RECT 177.005 88.605 177.285 89.485 ;
    RECT 173.685 88.605 173.965 89.485 ;
    RECT 170.365 88.605 170.645 89.485 ;
    RECT 167.045 88.605 167.325 89.485 ;
    RECT 163.725 88.605 164.005 89.485 ;
    RECT 160.405 88.605 160.685 89.485 ;
    RECT 157.085 88.605 157.365 89.485 ;
    RECT 153.765 88.605 154.045 89.485 ;
    RECT 150.445 88.605 150.725 89.485 ;
    RECT 213.525 88.605 213.805 89.485 ;
    RECT 210.205 88.605 210.485 89.485 ;
    RECT 206.885 88.605 207.165 89.485 ;
    RECT 203.565 88.605 203.845 89.485 ;
    RECT 200.245 88.605 200.525 89.485 ;
    RECT 196.925 88.605 197.205 89.485 ;
    RECT 193.605 88.605 193.885 89.485 ;
    RECT 190.285 88.605 190.565 89.485 ;
    RECT 186.965 88.605 187.245 89.485 ;
    RECT 183.645 88.605 183.925 89.485 ;
    RECT 266.645 88.605 266.925 89.485 ;
    RECT 263.325 88.605 263.605 89.485 ;
    RECT 260.005 88.605 260.285 89.485 ;
    RECT 256.685 88.605 256.965 89.485 ;
    RECT 253.365 88.605 253.645 89.485 ;
    RECT 250.045 51.865 250.325 52.745 ;
    RECT 246.725 51.865 247.005 52.745 ;
    RECT 243.405 51.865 243.685 52.745 ;
    RECT 240.085 51.865 240.365 52.745 ;
    RECT 236.765 51.865 237.045 52.745 ;
    RECT 233.445 51.865 233.725 52.745 ;
    RECT 230.125 51.865 230.405 52.745 ;
    RECT 226.805 51.865 227.085 52.745 ;
    RECT 223.485 51.865 223.765 52.745 ;
    RECT 220.165 51.865 220.445 52.745 ;
    RECT 216.845 51.865 217.125 52.745 ;
    RECT 180.325 51.865 180.605 52.745 ;
    RECT 177.005 51.865 177.285 52.745 ;
    RECT 173.685 51.865 173.965 52.745 ;
    RECT 170.365 51.865 170.645 52.745 ;
    RECT 167.045 51.865 167.325 52.745 ;
    RECT 163.725 51.865 164.005 52.745 ;
    RECT 160.405 51.865 160.685 52.745 ;
    RECT 157.085 51.865 157.365 52.745 ;
    RECT 153.765 51.865 154.045 52.745 ;
    RECT 150.445 51.865 150.725 52.745 ;
    RECT 213.525 51.865 213.805 52.745 ;
    RECT 210.205 51.865 210.485 52.745 ;
    RECT 206.885 51.865 207.165 52.745 ;
    RECT 203.565 51.865 203.845 52.745 ;
    RECT 200.245 51.865 200.525 52.745 ;
    RECT 196.925 51.865 197.205 52.745 ;
    RECT 193.605 51.865 193.885 52.745 ;
    RECT 190.285 51.865 190.565 52.745 ;
    RECT 186.965 51.865 187.245 52.745 ;
    RECT 183.645 51.865 183.925 52.745 ;
    RECT 266.645 51.865 266.925 52.745 ;
    RECT 263.325 51.865 263.605 52.745 ;
    RECT 260.005 51.865 260.285 52.745 ;
    RECT 256.685 51.865 256.965 52.745 ;
    RECT 253.365 51.865 253.645 52.745 ;
    RECT 250.045 87.885 250.325 88.765 ;
    RECT 246.725 87.885 247.005 88.765 ;
    RECT 243.405 87.885 243.685 88.765 ;
    RECT 240.085 87.885 240.365 88.765 ;
    RECT 236.765 87.885 237.045 88.765 ;
    RECT 233.445 87.885 233.725 88.765 ;
    RECT 230.125 87.885 230.405 88.765 ;
    RECT 226.805 87.885 227.085 88.765 ;
    RECT 223.485 87.885 223.765 88.765 ;
    RECT 220.165 87.885 220.445 88.765 ;
    RECT 216.845 87.885 217.125 88.765 ;
    RECT 180.325 87.885 180.605 88.765 ;
    RECT 177.005 87.885 177.285 88.765 ;
    RECT 173.685 87.885 173.965 88.765 ;
    RECT 170.365 87.885 170.645 88.765 ;
    RECT 167.045 87.885 167.325 88.765 ;
    RECT 163.725 87.885 164.005 88.765 ;
    RECT 160.405 87.885 160.685 88.765 ;
    RECT 157.085 87.885 157.365 88.765 ;
    RECT 153.765 87.885 154.045 88.765 ;
    RECT 150.445 87.885 150.725 88.765 ;
    RECT 213.525 87.885 213.805 88.765 ;
    RECT 210.205 87.885 210.485 88.765 ;
    RECT 206.885 87.885 207.165 88.765 ;
    RECT 203.565 87.885 203.845 88.765 ;
    RECT 200.245 87.885 200.525 88.765 ;
    RECT 196.925 87.885 197.205 88.765 ;
    RECT 193.605 87.885 193.885 88.765 ;
    RECT 190.285 87.885 190.565 88.765 ;
    RECT 186.965 87.885 187.245 88.765 ;
    RECT 183.645 87.885 183.925 88.765 ;
    RECT 266.645 87.885 266.925 88.765 ;
    RECT 263.325 87.885 263.605 88.765 ;
    RECT 260.005 87.885 260.285 88.765 ;
    RECT 256.685 87.885 256.965 88.765 ;
    RECT 253.365 87.885 253.645 88.765 ;
    RECT 250.045 51.145 250.325 52.025 ;
    RECT 246.725 51.145 247.005 52.025 ;
    RECT 243.405 51.145 243.685 52.025 ;
    RECT 240.085 51.145 240.365 52.025 ;
    RECT 236.765 51.145 237.045 52.025 ;
    RECT 233.445 51.145 233.725 52.025 ;
    RECT 230.125 51.145 230.405 52.025 ;
    RECT 226.805 51.145 227.085 52.025 ;
    RECT 223.485 51.145 223.765 52.025 ;
    RECT 220.165 51.145 220.445 52.025 ;
    RECT 216.845 51.145 217.125 52.025 ;
    RECT 180.325 51.145 180.605 52.025 ;
    RECT 177.005 51.145 177.285 52.025 ;
    RECT 173.685 51.145 173.965 52.025 ;
    RECT 170.365 51.145 170.645 52.025 ;
    RECT 167.045 51.145 167.325 52.025 ;
    RECT 163.725 51.145 164.005 52.025 ;
    RECT 160.405 51.145 160.685 52.025 ;
    RECT 157.085 51.145 157.365 52.025 ;
    RECT 153.765 51.145 154.045 52.025 ;
    RECT 150.445 51.145 150.725 52.025 ;
    RECT 213.525 51.145 213.805 52.025 ;
    RECT 210.205 51.145 210.485 52.025 ;
    RECT 206.885 51.145 207.165 52.025 ;
    RECT 203.565 51.145 203.845 52.025 ;
    RECT 200.245 51.145 200.525 52.025 ;
    RECT 196.925 51.145 197.205 52.025 ;
    RECT 193.605 51.145 193.885 52.025 ;
    RECT 190.285 51.145 190.565 52.025 ;
    RECT 186.965 51.145 187.245 52.025 ;
    RECT 183.645 51.145 183.925 52.025 ;
    RECT 266.645 51.145 266.925 52.025 ;
    RECT 263.325 51.145 263.605 52.025 ;
    RECT 260.005 51.145 260.285 52.025 ;
    RECT 256.685 51.145 256.965 52.025 ;
    RECT 253.365 51.145 253.645 52.025 ;
    RECT 250.045 87.165 250.325 88.045 ;
    RECT 246.725 87.165 247.005 88.045 ;
    RECT 243.405 87.165 243.685 88.045 ;
    RECT 240.085 87.165 240.365 88.045 ;
    RECT 236.765 87.165 237.045 88.045 ;
    RECT 233.445 87.165 233.725 88.045 ;
    RECT 230.125 87.165 230.405 88.045 ;
    RECT 226.805 87.165 227.085 88.045 ;
    RECT 223.485 87.165 223.765 88.045 ;
    RECT 220.165 87.165 220.445 88.045 ;
    RECT 216.845 87.165 217.125 88.045 ;
    RECT 180.325 87.165 180.605 88.045 ;
    RECT 177.005 87.165 177.285 88.045 ;
    RECT 173.685 87.165 173.965 88.045 ;
    RECT 170.365 87.165 170.645 88.045 ;
    RECT 167.045 87.165 167.325 88.045 ;
    RECT 163.725 87.165 164.005 88.045 ;
    RECT 160.405 87.165 160.685 88.045 ;
    RECT 157.085 87.165 157.365 88.045 ;
    RECT 153.765 87.165 154.045 88.045 ;
    RECT 150.445 87.165 150.725 88.045 ;
    RECT 213.525 87.165 213.805 88.045 ;
    RECT 210.205 87.165 210.485 88.045 ;
    RECT 206.885 87.165 207.165 88.045 ;
    RECT 203.565 87.165 203.845 88.045 ;
    RECT 200.245 87.165 200.525 88.045 ;
    RECT 196.925 87.165 197.205 88.045 ;
    RECT 193.605 87.165 193.885 88.045 ;
    RECT 190.285 87.165 190.565 88.045 ;
    RECT 186.965 87.165 187.245 88.045 ;
    RECT 183.645 87.165 183.925 88.045 ;
    RECT 266.645 87.165 266.925 88.045 ;
    RECT 263.325 87.165 263.605 88.045 ;
    RECT 260.005 87.165 260.285 88.045 ;
    RECT 256.685 87.165 256.965 88.045 ;
    RECT 253.365 87.165 253.645 88.045 ;
    RECT 250.045 50.425 250.325 51.305 ;
    RECT 246.725 50.425 247.005 51.305 ;
    RECT 243.405 50.425 243.685 51.305 ;
    RECT 240.085 50.425 240.365 51.305 ;
    RECT 236.765 50.425 237.045 51.305 ;
    RECT 233.445 50.425 233.725 51.305 ;
    RECT 230.125 50.425 230.405 51.305 ;
    RECT 226.805 50.425 227.085 51.305 ;
    RECT 223.485 50.425 223.765 51.305 ;
    RECT 220.165 50.425 220.445 51.305 ;
    RECT 216.845 50.425 217.125 51.305 ;
    RECT 180.325 50.425 180.605 51.305 ;
    RECT 177.005 50.425 177.285 51.305 ;
    RECT 173.685 50.425 173.965 51.305 ;
    RECT 170.365 50.425 170.645 51.305 ;
    RECT 167.045 50.425 167.325 51.305 ;
    RECT 163.725 50.425 164.005 51.305 ;
    RECT 160.405 50.425 160.685 51.305 ;
    RECT 157.085 50.425 157.365 51.305 ;
    RECT 153.765 50.425 154.045 51.305 ;
    RECT 150.445 50.425 150.725 51.305 ;
    RECT 213.525 50.425 213.805 51.305 ;
    RECT 210.205 50.425 210.485 51.305 ;
    RECT 206.885 50.425 207.165 51.305 ;
    RECT 203.565 50.425 203.845 51.305 ;
    RECT 200.245 50.425 200.525 51.305 ;
    RECT 196.925 50.425 197.205 51.305 ;
    RECT 193.605 50.425 193.885 51.305 ;
    RECT 190.285 50.425 190.565 51.305 ;
    RECT 186.965 50.425 187.245 51.305 ;
    RECT 183.645 50.425 183.925 51.305 ;
    RECT 266.645 50.425 266.925 51.305 ;
    RECT 263.325 50.425 263.605 51.305 ;
    RECT 260.005 50.425 260.285 51.305 ;
    RECT 256.685 50.425 256.965 51.305 ;
    RECT 253.365 50.425 253.645 51.305 ;
    RECT 250.045 49.705 250.325 50.585 ;
    RECT 246.725 49.705 247.005 50.585 ;
    RECT 243.405 49.705 243.685 50.585 ;
    RECT 240.085 49.705 240.365 50.585 ;
    RECT 236.765 49.705 237.045 50.585 ;
    RECT 233.445 49.705 233.725 50.585 ;
    RECT 230.125 49.705 230.405 50.585 ;
    RECT 226.805 49.705 227.085 50.585 ;
    RECT 223.485 49.705 223.765 50.585 ;
    RECT 220.165 49.705 220.445 50.585 ;
    RECT 216.845 49.705 217.125 50.585 ;
    RECT 180.325 49.705 180.605 50.585 ;
    RECT 177.005 49.705 177.285 50.585 ;
    RECT 173.685 49.705 173.965 50.585 ;
    RECT 170.365 49.705 170.645 50.585 ;
    RECT 167.045 49.705 167.325 50.585 ;
    RECT 163.725 49.705 164.005 50.585 ;
    RECT 160.405 49.705 160.685 50.585 ;
    RECT 157.085 49.705 157.365 50.585 ;
    RECT 153.765 49.705 154.045 50.585 ;
    RECT 150.445 49.705 150.725 50.585 ;
    RECT 213.525 49.705 213.805 50.585 ;
    RECT 210.205 49.705 210.485 50.585 ;
    RECT 206.885 49.705 207.165 50.585 ;
    RECT 203.565 49.705 203.845 50.585 ;
    RECT 200.245 49.705 200.525 50.585 ;
    RECT 196.925 49.705 197.205 50.585 ;
    RECT 193.605 49.705 193.885 50.585 ;
    RECT 190.285 49.705 190.565 50.585 ;
    RECT 186.965 49.705 187.245 50.585 ;
    RECT 183.645 49.705 183.925 50.585 ;
    RECT 266.645 49.705 266.925 50.585 ;
    RECT 263.325 49.705 263.605 50.585 ;
    RECT 260.005 49.705 260.285 50.585 ;
    RECT 256.685 49.705 256.965 50.585 ;
    RECT 253.365 49.705 253.645 50.585 ;
    RECT 250.045 48.985 250.325 49.865 ;
    RECT 246.725 48.985 247.005 49.865 ;
    RECT 243.405 48.985 243.685 49.865 ;
    RECT 240.085 48.985 240.365 49.865 ;
    RECT 236.765 48.985 237.045 49.865 ;
    RECT 233.445 48.985 233.725 49.865 ;
    RECT 230.125 48.985 230.405 49.865 ;
    RECT 226.805 48.985 227.085 49.865 ;
    RECT 223.485 48.985 223.765 49.865 ;
    RECT 220.165 48.985 220.445 49.865 ;
    RECT 216.845 48.985 217.125 49.865 ;
    RECT 180.325 48.985 180.605 49.865 ;
    RECT 177.005 48.985 177.285 49.865 ;
    RECT 173.685 48.985 173.965 49.865 ;
    RECT 170.365 48.985 170.645 49.865 ;
    RECT 167.045 48.985 167.325 49.865 ;
    RECT 163.725 48.985 164.005 49.865 ;
    RECT 160.405 48.985 160.685 49.865 ;
    RECT 157.085 48.985 157.365 49.865 ;
    RECT 153.765 48.985 154.045 49.865 ;
    RECT 150.445 48.985 150.725 49.865 ;
    RECT 213.525 48.985 213.805 49.865 ;
    RECT 210.205 48.985 210.485 49.865 ;
    RECT 206.885 48.985 207.165 49.865 ;
    RECT 203.565 48.985 203.845 49.865 ;
    RECT 200.245 48.985 200.525 49.865 ;
    RECT 196.925 48.985 197.205 49.865 ;
    RECT 193.605 48.985 193.885 49.865 ;
    RECT 190.285 48.985 190.565 49.865 ;
    RECT 186.965 48.985 187.245 49.865 ;
    RECT 183.645 48.985 183.925 49.865 ;
    RECT 266.645 48.985 266.925 49.865 ;
    RECT 263.325 48.985 263.605 49.865 ;
    RECT 260.005 48.985 260.285 49.865 ;
    RECT 256.685 48.985 256.965 49.865 ;
    RECT 253.365 48.985 253.645 49.865 ;
    RECT 250.045 48.265 250.325 49.145 ;
    RECT 246.725 48.265 247.005 49.145 ;
    RECT 243.405 48.265 243.685 49.145 ;
    RECT 240.085 48.265 240.365 49.145 ;
    RECT 236.765 48.265 237.045 49.145 ;
    RECT 233.445 48.265 233.725 49.145 ;
    RECT 230.125 48.265 230.405 49.145 ;
    RECT 226.805 48.265 227.085 49.145 ;
    RECT 223.485 48.265 223.765 49.145 ;
    RECT 220.165 48.265 220.445 49.145 ;
    RECT 216.845 48.265 217.125 49.145 ;
    RECT 180.325 48.265 180.605 49.145 ;
    RECT 177.005 48.265 177.285 49.145 ;
    RECT 173.685 48.265 173.965 49.145 ;
    RECT 170.365 48.265 170.645 49.145 ;
    RECT 167.045 48.265 167.325 49.145 ;
    RECT 163.725 48.265 164.005 49.145 ;
    RECT 160.405 48.265 160.685 49.145 ;
    RECT 157.085 48.265 157.365 49.145 ;
    RECT 153.765 48.265 154.045 49.145 ;
    RECT 150.445 48.265 150.725 49.145 ;
    RECT 213.525 48.265 213.805 49.145 ;
    RECT 210.205 48.265 210.485 49.145 ;
    RECT 206.885 48.265 207.165 49.145 ;
    RECT 203.565 48.265 203.845 49.145 ;
    RECT 200.245 48.265 200.525 49.145 ;
    RECT 196.925 48.265 197.205 49.145 ;
    RECT 193.605 48.265 193.885 49.145 ;
    RECT 190.285 48.265 190.565 49.145 ;
    RECT 186.965 48.265 187.245 49.145 ;
    RECT 183.645 48.265 183.925 49.145 ;
    RECT 266.645 48.265 266.925 49.145 ;
    RECT 263.325 48.265 263.605 49.145 ;
    RECT 260.005 48.265 260.285 49.145 ;
    RECT 256.685 48.265 256.965 49.145 ;
    RECT 253.365 48.265 253.645 49.145 ;
    RECT 250.045 47.545 250.325 48.425 ;
    RECT 246.725 47.545 247.005 48.425 ;
    RECT 243.405 47.545 243.685 48.425 ;
    RECT 240.085 47.545 240.365 48.425 ;
    RECT 236.765 47.545 237.045 48.425 ;
    RECT 233.445 47.545 233.725 48.425 ;
    RECT 230.125 47.545 230.405 48.425 ;
    RECT 226.805 47.545 227.085 48.425 ;
    RECT 223.485 47.545 223.765 48.425 ;
    RECT 220.165 47.545 220.445 48.425 ;
    RECT 216.845 47.545 217.125 48.425 ;
    RECT 180.325 47.545 180.605 48.425 ;
    RECT 177.005 47.545 177.285 48.425 ;
    RECT 173.685 47.545 173.965 48.425 ;
    RECT 170.365 47.545 170.645 48.425 ;
    RECT 167.045 47.545 167.325 48.425 ;
    RECT 163.725 47.545 164.005 48.425 ;
    RECT 160.405 47.545 160.685 48.425 ;
    RECT 157.085 47.545 157.365 48.425 ;
    RECT 153.765 47.545 154.045 48.425 ;
    RECT 150.445 47.545 150.725 48.425 ;
    RECT 213.525 47.545 213.805 48.425 ;
    RECT 210.205 47.545 210.485 48.425 ;
    RECT 206.885 47.545 207.165 48.425 ;
    RECT 203.565 47.545 203.845 48.425 ;
    RECT 200.245 47.545 200.525 48.425 ;
    RECT 196.925 47.545 197.205 48.425 ;
    RECT 193.605 47.545 193.885 48.425 ;
    RECT 190.285 47.545 190.565 48.425 ;
    RECT 186.965 47.545 187.245 48.425 ;
    RECT 183.645 47.545 183.925 48.425 ;
    RECT 266.645 47.545 266.925 48.425 ;
    RECT 263.325 47.545 263.605 48.425 ;
    RECT 260.005 47.545 260.285 48.425 ;
    RECT 256.685 47.545 256.965 48.425 ;
    RECT 253.365 47.545 253.645 48.425 ;
    RECT 250.045 46.825 250.325 47.705 ;
    RECT 246.725 46.825 247.005 47.705 ;
    RECT 243.405 46.825 243.685 47.705 ;
    RECT 240.085 46.825 240.365 47.705 ;
    RECT 236.765 46.825 237.045 47.705 ;
    RECT 233.445 46.825 233.725 47.705 ;
    RECT 230.125 46.825 230.405 47.705 ;
    RECT 226.805 46.825 227.085 47.705 ;
    RECT 223.485 46.825 223.765 47.705 ;
    RECT 220.165 46.825 220.445 47.705 ;
    RECT 216.845 46.825 217.125 47.705 ;
    RECT 180.325 46.825 180.605 47.705 ;
    RECT 177.005 46.825 177.285 47.705 ;
    RECT 173.685 46.825 173.965 47.705 ;
    RECT 170.365 46.825 170.645 47.705 ;
    RECT 167.045 46.825 167.325 47.705 ;
    RECT 163.725 46.825 164.005 47.705 ;
    RECT 160.405 46.825 160.685 47.705 ;
    RECT 157.085 46.825 157.365 47.705 ;
    RECT 153.765 46.825 154.045 47.705 ;
    RECT 150.445 46.825 150.725 47.705 ;
    RECT 213.525 46.825 213.805 47.705 ;
    RECT 210.205 46.825 210.485 47.705 ;
    RECT 206.885 46.825 207.165 47.705 ;
    RECT 203.565 46.825 203.845 47.705 ;
    RECT 200.245 46.825 200.525 47.705 ;
    RECT 196.925 46.825 197.205 47.705 ;
    RECT 193.605 46.825 193.885 47.705 ;
    RECT 190.285 46.825 190.565 47.705 ;
    RECT 186.965 46.825 187.245 47.705 ;
    RECT 183.645 46.825 183.925 47.705 ;
    RECT 266.645 46.825 266.925 47.705 ;
    RECT 263.325 46.825 263.605 47.705 ;
    RECT 260.005 46.825 260.285 47.705 ;
    RECT 256.685 46.825 256.965 47.705 ;
    RECT 253.365 46.825 253.645 47.705 ;
    RECT 250.045 86.445 250.325 87.325 ;
    RECT 246.725 86.445 247.005 87.325 ;
    RECT 243.405 86.445 243.685 87.325 ;
    RECT 240.085 86.445 240.365 87.325 ;
    RECT 236.765 86.445 237.045 87.325 ;
    RECT 233.445 86.445 233.725 87.325 ;
    RECT 230.125 86.445 230.405 87.325 ;
    RECT 226.805 86.445 227.085 87.325 ;
    RECT 223.485 86.445 223.765 87.325 ;
    RECT 220.165 86.445 220.445 87.325 ;
    RECT 216.845 86.445 217.125 87.325 ;
    RECT 180.325 86.445 180.605 87.325 ;
    RECT 177.005 86.445 177.285 87.325 ;
    RECT 173.685 86.445 173.965 87.325 ;
    RECT 170.365 86.445 170.645 87.325 ;
    RECT 167.045 86.445 167.325 87.325 ;
    RECT 163.725 86.445 164.005 87.325 ;
    RECT 160.405 86.445 160.685 87.325 ;
    RECT 157.085 86.445 157.365 87.325 ;
    RECT 153.765 86.445 154.045 87.325 ;
    RECT 150.445 86.445 150.725 87.325 ;
    RECT 213.525 86.445 213.805 87.325 ;
    RECT 210.205 86.445 210.485 87.325 ;
    RECT 206.885 86.445 207.165 87.325 ;
    RECT 203.565 86.445 203.845 87.325 ;
    RECT 200.245 86.445 200.525 87.325 ;
    RECT 196.925 86.445 197.205 87.325 ;
    RECT 193.605 86.445 193.885 87.325 ;
    RECT 190.285 86.445 190.565 87.325 ;
    RECT 186.965 86.445 187.245 87.325 ;
    RECT 183.645 86.445 183.925 87.325 ;
    RECT 266.645 86.445 266.925 87.325 ;
    RECT 263.325 86.445 263.605 87.325 ;
    RECT 260.005 86.445 260.285 87.325 ;
    RECT 256.685 86.445 256.965 87.325 ;
    RECT 253.365 86.445 253.645 87.325 ;
    RECT 250.045 46.105 250.325 46.985 ;
    RECT 246.725 46.105 247.005 46.985 ;
    RECT 243.405 46.105 243.685 46.985 ;
    RECT 240.085 46.105 240.365 46.985 ;
    RECT 236.765 46.105 237.045 46.985 ;
    RECT 233.445 46.105 233.725 46.985 ;
    RECT 230.125 46.105 230.405 46.985 ;
    RECT 226.805 46.105 227.085 46.985 ;
    RECT 223.485 46.105 223.765 46.985 ;
    RECT 220.165 46.105 220.445 46.985 ;
    RECT 216.845 46.105 217.125 46.985 ;
    RECT 180.325 46.105 180.605 46.985 ;
    RECT 177.005 46.105 177.285 46.985 ;
    RECT 173.685 46.105 173.965 46.985 ;
    RECT 170.365 46.105 170.645 46.985 ;
    RECT 167.045 46.105 167.325 46.985 ;
    RECT 163.725 46.105 164.005 46.985 ;
    RECT 160.405 46.105 160.685 46.985 ;
    RECT 157.085 46.105 157.365 46.985 ;
    RECT 153.765 46.105 154.045 46.985 ;
    RECT 150.445 46.105 150.725 46.985 ;
    RECT 213.525 46.105 213.805 46.985 ;
    RECT 210.205 46.105 210.485 46.985 ;
    RECT 206.885 46.105 207.165 46.985 ;
    RECT 203.565 46.105 203.845 46.985 ;
    RECT 200.245 46.105 200.525 46.985 ;
    RECT 196.925 46.105 197.205 46.985 ;
    RECT 193.605 46.105 193.885 46.985 ;
    RECT 190.285 46.105 190.565 46.985 ;
    RECT 186.965 46.105 187.245 46.985 ;
    RECT 183.645 46.105 183.925 46.985 ;
    RECT 266.645 46.105 266.925 46.985 ;
    RECT 263.325 46.105 263.605 46.985 ;
    RECT 260.005 46.105 260.285 46.985 ;
    RECT 256.685 46.105 256.965 46.985 ;
    RECT 253.365 46.105 253.645 46.985 ;
    RECT 250.045 85.725 250.325 86.605 ;
    RECT 246.725 85.725 247.005 86.605 ;
    RECT 243.405 85.725 243.685 86.605 ;
    RECT 240.085 85.725 240.365 86.605 ;
    RECT 236.765 85.725 237.045 86.605 ;
    RECT 233.445 85.725 233.725 86.605 ;
    RECT 230.125 85.725 230.405 86.605 ;
    RECT 226.805 85.725 227.085 86.605 ;
    RECT 223.485 85.725 223.765 86.605 ;
    RECT 220.165 85.725 220.445 86.605 ;
    RECT 216.845 85.725 217.125 86.605 ;
    RECT 180.325 85.725 180.605 86.605 ;
    RECT 177.005 85.725 177.285 86.605 ;
    RECT 173.685 85.725 173.965 86.605 ;
    RECT 170.365 85.725 170.645 86.605 ;
    RECT 167.045 85.725 167.325 86.605 ;
    RECT 163.725 85.725 164.005 86.605 ;
    RECT 160.405 85.725 160.685 86.605 ;
    RECT 157.085 85.725 157.365 86.605 ;
    RECT 153.765 85.725 154.045 86.605 ;
    RECT 150.445 85.725 150.725 86.605 ;
    RECT 213.525 85.725 213.805 86.605 ;
    RECT 210.205 85.725 210.485 86.605 ;
    RECT 206.885 85.725 207.165 86.605 ;
    RECT 203.565 85.725 203.845 86.605 ;
    RECT 200.245 85.725 200.525 86.605 ;
    RECT 196.925 85.725 197.205 86.605 ;
    RECT 193.605 85.725 193.885 86.605 ;
    RECT 190.285 85.725 190.565 86.605 ;
    RECT 186.965 85.725 187.245 86.605 ;
    RECT 183.645 85.725 183.925 86.605 ;
    RECT 266.645 85.725 266.925 86.605 ;
    RECT 263.325 85.725 263.605 86.605 ;
    RECT 260.005 85.725 260.285 86.605 ;
    RECT 256.685 85.725 256.965 86.605 ;
    RECT 253.365 85.725 253.645 86.605 ;
    RECT 250.045 45.385 250.325 46.265 ;
    RECT 246.725 45.385 247.005 46.265 ;
    RECT 243.405 45.385 243.685 46.265 ;
    RECT 240.085 45.385 240.365 46.265 ;
    RECT 236.765 45.385 237.045 46.265 ;
    RECT 233.445 45.385 233.725 46.265 ;
    RECT 230.125 45.385 230.405 46.265 ;
    RECT 226.805 45.385 227.085 46.265 ;
    RECT 223.485 45.385 223.765 46.265 ;
    RECT 220.165 45.385 220.445 46.265 ;
    RECT 216.845 45.385 217.125 46.265 ;
    RECT 180.325 45.385 180.605 46.265 ;
    RECT 177.005 45.385 177.285 46.265 ;
    RECT 173.685 45.385 173.965 46.265 ;
    RECT 170.365 45.385 170.645 46.265 ;
    RECT 167.045 45.385 167.325 46.265 ;
    RECT 163.725 45.385 164.005 46.265 ;
    RECT 160.405 45.385 160.685 46.265 ;
    RECT 157.085 45.385 157.365 46.265 ;
    RECT 153.765 45.385 154.045 46.265 ;
    RECT 150.445 45.385 150.725 46.265 ;
    RECT 213.525 45.385 213.805 46.265 ;
    RECT 210.205 45.385 210.485 46.265 ;
    RECT 206.885 45.385 207.165 46.265 ;
    RECT 203.565 45.385 203.845 46.265 ;
    RECT 200.245 45.385 200.525 46.265 ;
    RECT 196.925 45.385 197.205 46.265 ;
    RECT 193.605 45.385 193.885 46.265 ;
    RECT 190.285 45.385 190.565 46.265 ;
    RECT 186.965 45.385 187.245 46.265 ;
    RECT 183.645 45.385 183.925 46.265 ;
    RECT 266.645 45.385 266.925 46.265 ;
    RECT 263.325 45.385 263.605 46.265 ;
    RECT 260.005 45.385 260.285 46.265 ;
    RECT 256.685 45.385 256.965 46.265 ;
    RECT 253.365 45.385 253.645 46.265 ;
    RECT 250.045 85.005 250.325 85.885 ;
    RECT 246.725 85.005 247.005 85.885 ;
    RECT 243.405 85.005 243.685 85.885 ;
    RECT 240.085 85.005 240.365 85.885 ;
    RECT 236.765 85.005 237.045 85.885 ;
    RECT 233.445 85.005 233.725 85.885 ;
    RECT 230.125 85.005 230.405 85.885 ;
    RECT 226.805 85.005 227.085 85.885 ;
    RECT 223.485 85.005 223.765 85.885 ;
    RECT 220.165 85.005 220.445 85.885 ;
    RECT 216.845 85.005 217.125 85.885 ;
    RECT 180.325 85.005 180.605 85.885 ;
    RECT 177.005 85.005 177.285 85.885 ;
    RECT 173.685 85.005 173.965 85.885 ;
    RECT 170.365 85.005 170.645 85.885 ;
    RECT 167.045 85.005 167.325 85.885 ;
    RECT 163.725 85.005 164.005 85.885 ;
    RECT 160.405 85.005 160.685 85.885 ;
    RECT 157.085 85.005 157.365 85.885 ;
    RECT 153.765 85.005 154.045 85.885 ;
    RECT 150.445 85.005 150.725 85.885 ;
    RECT 213.525 85.005 213.805 85.885 ;
    RECT 210.205 85.005 210.485 85.885 ;
    RECT 206.885 85.005 207.165 85.885 ;
    RECT 203.565 85.005 203.845 85.885 ;
    RECT 200.245 85.005 200.525 85.885 ;
    RECT 196.925 85.005 197.205 85.885 ;
    RECT 193.605 85.005 193.885 85.885 ;
    RECT 190.285 85.005 190.565 85.885 ;
    RECT 186.965 85.005 187.245 85.885 ;
    RECT 183.645 85.005 183.925 85.885 ;
    RECT 266.645 85.005 266.925 85.885 ;
    RECT 263.325 85.005 263.605 85.885 ;
    RECT 260.005 85.005 260.285 85.885 ;
    RECT 256.685 85.005 256.965 85.885 ;
    RECT 253.365 85.005 253.645 85.885 ;
    RECT 250.045 44.665 250.325 45.545 ;
    RECT 246.725 44.665 247.005 45.545 ;
    RECT 243.405 44.665 243.685 45.545 ;
    RECT 240.085 44.665 240.365 45.545 ;
    RECT 236.765 44.665 237.045 45.545 ;
    RECT 233.445 44.665 233.725 45.545 ;
    RECT 230.125 44.665 230.405 45.545 ;
    RECT 226.805 44.665 227.085 45.545 ;
    RECT 223.485 44.665 223.765 45.545 ;
    RECT 220.165 44.665 220.445 45.545 ;
    RECT 216.845 44.665 217.125 45.545 ;
    RECT 180.325 44.665 180.605 45.545 ;
    RECT 177.005 44.665 177.285 45.545 ;
    RECT 173.685 44.665 173.965 45.545 ;
    RECT 170.365 44.665 170.645 45.545 ;
    RECT 167.045 44.665 167.325 45.545 ;
    RECT 163.725 44.665 164.005 45.545 ;
    RECT 160.405 44.665 160.685 45.545 ;
    RECT 157.085 44.665 157.365 45.545 ;
    RECT 153.765 44.665 154.045 45.545 ;
    RECT 150.445 44.665 150.725 45.545 ;
    RECT 213.525 44.665 213.805 45.545 ;
    RECT 210.205 44.665 210.485 45.545 ;
    RECT 206.885 44.665 207.165 45.545 ;
    RECT 203.565 44.665 203.845 45.545 ;
    RECT 200.245 44.665 200.525 45.545 ;
    RECT 196.925 44.665 197.205 45.545 ;
    RECT 193.605 44.665 193.885 45.545 ;
    RECT 190.285 44.665 190.565 45.545 ;
    RECT 186.965 44.665 187.245 45.545 ;
    RECT 183.645 44.665 183.925 45.545 ;
    RECT 266.645 44.665 266.925 45.545 ;
    RECT 263.325 44.665 263.605 45.545 ;
    RECT 260.005 44.665 260.285 45.545 ;
    RECT 256.685 44.665 256.965 45.545 ;
    RECT 253.365 44.665 253.645 45.545 ;
    RECT 250.045 84.285 250.325 85.165 ;
    RECT 246.725 84.285 247.005 85.165 ;
    RECT 243.405 84.285 243.685 85.165 ;
    RECT 240.085 84.285 240.365 85.165 ;
    RECT 236.765 84.285 237.045 85.165 ;
    RECT 233.445 84.285 233.725 85.165 ;
    RECT 230.125 84.285 230.405 85.165 ;
    RECT 226.805 84.285 227.085 85.165 ;
    RECT 223.485 84.285 223.765 85.165 ;
    RECT 220.165 84.285 220.445 85.165 ;
    RECT 216.845 84.285 217.125 85.165 ;
    RECT 180.325 84.285 180.605 85.165 ;
    RECT 177.005 84.285 177.285 85.165 ;
    RECT 173.685 84.285 173.965 85.165 ;
    RECT 170.365 84.285 170.645 85.165 ;
    RECT 167.045 84.285 167.325 85.165 ;
    RECT 163.725 84.285 164.005 85.165 ;
    RECT 160.405 84.285 160.685 85.165 ;
    RECT 157.085 84.285 157.365 85.165 ;
    RECT 153.765 84.285 154.045 85.165 ;
    RECT 150.445 84.285 150.725 85.165 ;
    RECT 213.525 84.285 213.805 85.165 ;
    RECT 210.205 84.285 210.485 85.165 ;
    RECT 206.885 84.285 207.165 85.165 ;
    RECT 203.565 84.285 203.845 85.165 ;
    RECT 200.245 84.285 200.525 85.165 ;
    RECT 196.925 84.285 197.205 85.165 ;
    RECT 193.605 84.285 193.885 85.165 ;
    RECT 190.285 84.285 190.565 85.165 ;
    RECT 186.965 84.285 187.245 85.165 ;
    RECT 183.645 84.285 183.925 85.165 ;
    RECT 266.645 84.285 266.925 85.165 ;
    RECT 263.325 84.285 263.605 85.165 ;
    RECT 260.005 84.285 260.285 85.165 ;
    RECT 256.685 84.285 256.965 85.165 ;
    RECT 253.365 84.285 253.645 85.165 ;
    RECT 250.045 43.945 250.325 44.825 ;
    RECT 246.725 43.945 247.005 44.825 ;
    RECT 243.405 43.945 243.685 44.825 ;
    RECT 240.085 43.945 240.365 44.825 ;
    RECT 236.765 43.945 237.045 44.825 ;
    RECT 233.445 43.945 233.725 44.825 ;
    RECT 230.125 43.945 230.405 44.825 ;
    RECT 226.805 43.945 227.085 44.825 ;
    RECT 223.485 43.945 223.765 44.825 ;
    RECT 220.165 43.945 220.445 44.825 ;
    RECT 216.845 43.945 217.125 44.825 ;
    RECT 180.325 43.945 180.605 44.825 ;
    RECT 177.005 43.945 177.285 44.825 ;
    RECT 173.685 43.945 173.965 44.825 ;
    RECT 170.365 43.945 170.645 44.825 ;
    RECT 167.045 43.945 167.325 44.825 ;
    RECT 163.725 43.945 164.005 44.825 ;
    RECT 160.405 43.945 160.685 44.825 ;
    RECT 157.085 43.945 157.365 44.825 ;
    RECT 153.765 43.945 154.045 44.825 ;
    RECT 150.445 43.945 150.725 44.825 ;
    RECT 213.525 43.945 213.805 44.825 ;
    RECT 210.205 43.945 210.485 44.825 ;
    RECT 206.885 43.945 207.165 44.825 ;
    RECT 203.565 43.945 203.845 44.825 ;
    RECT 200.245 43.945 200.525 44.825 ;
    RECT 196.925 43.945 197.205 44.825 ;
    RECT 193.605 43.945 193.885 44.825 ;
    RECT 190.285 43.945 190.565 44.825 ;
    RECT 186.965 43.945 187.245 44.825 ;
    RECT 183.645 43.945 183.925 44.825 ;
    RECT 266.645 43.945 266.925 44.825 ;
    RECT 263.325 43.945 263.605 44.825 ;
    RECT 260.005 43.945 260.285 44.825 ;
    RECT 256.685 43.945 256.965 44.825 ;
    RECT 253.365 43.945 253.645 44.825 ;
    RECT 250.045 83.565 250.325 84.445 ;
    RECT 246.725 83.565 247.005 84.445 ;
    RECT 243.405 83.565 243.685 84.445 ;
    RECT 240.085 83.565 240.365 84.445 ;
    RECT 236.765 83.565 237.045 84.445 ;
    RECT 233.445 83.565 233.725 84.445 ;
    RECT 230.125 83.565 230.405 84.445 ;
    RECT 226.805 83.565 227.085 84.445 ;
    RECT 223.485 83.565 223.765 84.445 ;
    RECT 220.165 83.565 220.445 84.445 ;
    RECT 216.845 83.565 217.125 84.445 ;
    RECT 180.325 83.565 180.605 84.445 ;
    RECT 177.005 83.565 177.285 84.445 ;
    RECT 173.685 83.565 173.965 84.445 ;
    RECT 170.365 83.565 170.645 84.445 ;
    RECT 167.045 83.565 167.325 84.445 ;
    RECT 163.725 83.565 164.005 84.445 ;
    RECT 160.405 83.565 160.685 84.445 ;
    RECT 157.085 83.565 157.365 84.445 ;
    RECT 153.765 83.565 154.045 84.445 ;
    RECT 150.445 83.565 150.725 84.445 ;
    RECT 213.525 83.565 213.805 84.445 ;
    RECT 210.205 83.565 210.485 84.445 ;
    RECT 206.885 83.565 207.165 84.445 ;
    RECT 203.565 83.565 203.845 84.445 ;
    RECT 200.245 83.565 200.525 84.445 ;
    RECT 196.925 83.565 197.205 84.445 ;
    RECT 193.605 83.565 193.885 84.445 ;
    RECT 190.285 83.565 190.565 84.445 ;
    RECT 186.965 83.565 187.245 84.445 ;
    RECT 183.645 83.565 183.925 84.445 ;
    RECT 266.645 83.565 266.925 84.445 ;
    RECT 263.325 83.565 263.605 84.445 ;
    RECT 260.005 83.565 260.285 84.445 ;
    RECT 256.685 83.565 256.965 84.445 ;
    RECT 253.365 83.565 253.645 84.445 ;
    RECT 250.045 43.225 250.325 44.105 ;
    RECT 246.725 43.225 247.005 44.105 ;
    RECT 243.405 43.225 243.685 44.105 ;
    RECT 240.085 43.225 240.365 44.105 ;
    RECT 236.765 43.225 237.045 44.105 ;
    RECT 233.445 43.225 233.725 44.105 ;
    RECT 230.125 43.225 230.405 44.105 ;
    RECT 226.805 43.225 227.085 44.105 ;
    RECT 223.485 43.225 223.765 44.105 ;
    RECT 220.165 43.225 220.445 44.105 ;
    RECT 216.845 43.225 217.125 44.105 ;
    RECT 180.325 43.225 180.605 44.105 ;
    RECT 177.005 43.225 177.285 44.105 ;
    RECT 173.685 43.225 173.965 44.105 ;
    RECT 170.365 43.225 170.645 44.105 ;
    RECT 167.045 43.225 167.325 44.105 ;
    RECT 163.725 43.225 164.005 44.105 ;
    RECT 160.405 43.225 160.685 44.105 ;
    RECT 157.085 43.225 157.365 44.105 ;
    RECT 153.765 43.225 154.045 44.105 ;
    RECT 150.445 43.225 150.725 44.105 ;
    RECT 213.525 43.225 213.805 44.105 ;
    RECT 210.205 43.225 210.485 44.105 ;
    RECT 206.885 43.225 207.165 44.105 ;
    RECT 203.565 43.225 203.845 44.105 ;
    RECT 200.245 43.225 200.525 44.105 ;
    RECT 196.925 43.225 197.205 44.105 ;
    RECT 193.605 43.225 193.885 44.105 ;
    RECT 190.285 43.225 190.565 44.105 ;
    RECT 186.965 43.225 187.245 44.105 ;
    RECT 183.645 43.225 183.925 44.105 ;
    RECT 266.645 43.225 266.925 44.105 ;
    RECT 263.325 43.225 263.605 44.105 ;
    RECT 260.005 43.225 260.285 44.105 ;
    RECT 256.685 43.225 256.965 44.105 ;
    RECT 253.365 43.225 253.645 44.105 ;
    RECT 250.045 82.845 250.325 83.725 ;
    RECT 246.725 82.845 247.005 83.725 ;
    RECT 243.405 82.845 243.685 83.725 ;
    RECT 240.085 82.845 240.365 83.725 ;
    RECT 236.765 82.845 237.045 83.725 ;
    RECT 233.445 82.845 233.725 83.725 ;
    RECT 230.125 82.845 230.405 83.725 ;
    RECT 226.805 82.845 227.085 83.725 ;
    RECT 223.485 82.845 223.765 83.725 ;
    RECT 220.165 82.845 220.445 83.725 ;
    RECT 216.845 82.845 217.125 83.725 ;
    RECT 180.325 82.845 180.605 83.725 ;
    RECT 177.005 82.845 177.285 83.725 ;
    RECT 173.685 82.845 173.965 83.725 ;
    RECT 170.365 82.845 170.645 83.725 ;
    RECT 167.045 82.845 167.325 83.725 ;
    RECT 163.725 82.845 164.005 83.725 ;
    RECT 160.405 82.845 160.685 83.725 ;
    RECT 157.085 82.845 157.365 83.725 ;
    RECT 153.765 82.845 154.045 83.725 ;
    RECT 150.445 82.845 150.725 83.725 ;
    RECT 213.525 82.845 213.805 83.725 ;
    RECT 210.205 82.845 210.485 83.725 ;
    RECT 206.885 82.845 207.165 83.725 ;
    RECT 203.565 82.845 203.845 83.725 ;
    RECT 200.245 82.845 200.525 83.725 ;
    RECT 196.925 82.845 197.205 83.725 ;
    RECT 193.605 82.845 193.885 83.725 ;
    RECT 190.285 82.845 190.565 83.725 ;
    RECT 186.965 82.845 187.245 83.725 ;
    RECT 183.645 82.845 183.925 83.725 ;
    RECT 266.645 82.845 266.925 83.725 ;
    RECT 263.325 82.845 263.605 83.725 ;
    RECT 260.005 82.845 260.285 83.725 ;
    RECT 256.685 82.845 256.965 83.725 ;
    RECT 253.365 82.845 253.645 83.725 ;
    RECT 250.045 82.125 250.325 83.005 ;
    RECT 246.725 82.125 247.005 83.005 ;
    RECT 243.405 82.125 243.685 83.005 ;
    RECT 240.085 82.125 240.365 83.005 ;
    RECT 236.765 82.125 237.045 83.005 ;
    RECT 233.445 82.125 233.725 83.005 ;
    RECT 230.125 82.125 230.405 83.005 ;
    RECT 226.805 82.125 227.085 83.005 ;
    RECT 223.485 82.125 223.765 83.005 ;
    RECT 220.165 82.125 220.445 83.005 ;
    RECT 216.845 82.125 217.125 83.005 ;
    RECT 180.325 82.125 180.605 83.005 ;
    RECT 177.005 82.125 177.285 83.005 ;
    RECT 173.685 82.125 173.965 83.005 ;
    RECT 170.365 82.125 170.645 83.005 ;
    RECT 167.045 82.125 167.325 83.005 ;
    RECT 163.725 82.125 164.005 83.005 ;
    RECT 160.405 82.125 160.685 83.005 ;
    RECT 157.085 82.125 157.365 83.005 ;
    RECT 153.765 82.125 154.045 83.005 ;
    RECT 150.445 82.125 150.725 83.005 ;
    RECT 213.525 82.125 213.805 83.005 ;
    RECT 210.205 82.125 210.485 83.005 ;
    RECT 206.885 82.125 207.165 83.005 ;
    RECT 203.565 82.125 203.845 83.005 ;
    RECT 200.245 82.125 200.525 83.005 ;
    RECT 196.925 82.125 197.205 83.005 ;
    RECT 193.605 82.125 193.885 83.005 ;
    RECT 190.285 82.125 190.565 83.005 ;
    RECT 186.965 82.125 187.245 83.005 ;
    RECT 183.645 82.125 183.925 83.005 ;
    RECT 266.645 82.125 266.925 83.005 ;
    RECT 263.325 82.125 263.605 83.005 ;
    RECT 260.005 82.125 260.285 83.005 ;
    RECT 256.685 82.125 256.965 83.005 ;
    RECT 253.365 82.125 253.645 83.005 ;
    RECT 250.045 81.405 250.325 82.285 ;
    RECT 246.725 81.405 247.005 82.285 ;
    RECT 243.405 81.405 243.685 82.285 ;
    RECT 240.085 81.405 240.365 82.285 ;
    RECT 236.765 81.405 237.045 82.285 ;
    RECT 233.445 81.405 233.725 82.285 ;
    RECT 230.125 81.405 230.405 82.285 ;
    RECT 226.805 81.405 227.085 82.285 ;
    RECT 223.485 81.405 223.765 82.285 ;
    RECT 220.165 81.405 220.445 82.285 ;
    RECT 216.845 81.405 217.125 82.285 ;
    RECT 180.325 81.405 180.605 82.285 ;
    RECT 177.005 81.405 177.285 82.285 ;
    RECT 173.685 81.405 173.965 82.285 ;
    RECT 170.365 81.405 170.645 82.285 ;
    RECT 167.045 81.405 167.325 82.285 ;
    RECT 163.725 81.405 164.005 82.285 ;
    RECT 160.405 81.405 160.685 82.285 ;
    RECT 157.085 81.405 157.365 82.285 ;
    RECT 153.765 81.405 154.045 82.285 ;
    RECT 150.445 81.405 150.725 82.285 ;
    RECT 213.525 81.405 213.805 82.285 ;
    RECT 210.205 81.405 210.485 82.285 ;
    RECT 206.885 81.405 207.165 82.285 ;
    RECT 203.565 81.405 203.845 82.285 ;
    RECT 200.245 81.405 200.525 82.285 ;
    RECT 196.925 81.405 197.205 82.285 ;
    RECT 193.605 81.405 193.885 82.285 ;
    RECT 190.285 81.405 190.565 82.285 ;
    RECT 186.965 81.405 187.245 82.285 ;
    RECT 183.645 81.405 183.925 82.285 ;
    RECT 266.645 81.405 266.925 82.285 ;
    RECT 263.325 81.405 263.605 82.285 ;
    RECT 260.005 81.405 260.285 82.285 ;
    RECT 256.685 81.405 256.965 82.285 ;
    RECT 253.365 81.405 253.645 82.285 ;
    RECT 250.045 97.965 250.325 98.845 ;
    RECT 246.725 97.965 247.005 98.845 ;
    RECT 243.405 97.965 243.685 98.845 ;
    RECT 240.085 97.965 240.365 98.845 ;
    RECT 236.765 97.965 237.045 98.845 ;
    RECT 233.445 97.965 233.725 98.845 ;
    RECT 230.125 97.965 230.405 98.845 ;
    RECT 226.805 97.965 227.085 98.845 ;
    RECT 223.485 97.965 223.765 98.845 ;
    RECT 220.165 97.965 220.445 98.845 ;
    RECT 216.845 97.965 217.125 98.845 ;
    RECT 180.325 97.965 180.605 98.845 ;
    RECT 177.005 97.965 177.285 98.845 ;
    RECT 173.685 97.965 173.965 98.845 ;
    RECT 170.365 97.965 170.645 98.845 ;
    RECT 167.045 97.965 167.325 98.845 ;
    RECT 163.725 97.965 164.005 98.845 ;
    RECT 160.405 97.965 160.685 98.845 ;
    RECT 157.085 97.965 157.365 98.845 ;
    RECT 153.765 97.965 154.045 98.845 ;
    RECT 213.525 97.965 213.805 98.845 ;
    RECT 210.205 97.965 210.485 98.845 ;
    RECT 206.885 97.965 207.165 98.845 ;
    RECT 203.565 97.965 203.845 98.845 ;
    RECT 200.245 97.965 200.525 98.845 ;
    RECT 196.925 97.965 197.205 98.845 ;
    RECT 193.605 97.965 193.885 98.845 ;
    RECT 190.285 97.965 190.565 98.845 ;
    RECT 186.965 97.965 187.245 98.845 ;
    RECT 183.645 97.965 183.925 98.845 ;
    RECT 266.645 97.965 266.925 98.845 ;
    RECT 150.445 97.965 150.725 98.845 ;
    RECT 263.325 97.965 263.605 98.845 ;
    RECT 260.005 97.965 260.285 98.845 ;
    RECT 256.685 97.965 256.965 98.845 ;
    RECT 253.365 97.965 253.645 98.845 ;
    RECT 250.045 80.685 250.325 81.565 ;
    RECT 246.725 80.685 247.005 81.565 ;
    RECT 243.405 80.685 243.685 81.565 ;
    RECT 240.085 80.685 240.365 81.565 ;
    RECT 236.765 80.685 237.045 81.565 ;
    RECT 233.445 80.685 233.725 81.565 ;
    RECT 230.125 80.685 230.405 81.565 ;
    RECT 226.805 80.685 227.085 81.565 ;
    RECT 223.485 80.685 223.765 81.565 ;
    RECT 220.165 80.685 220.445 81.565 ;
    RECT 216.845 80.685 217.125 81.565 ;
    RECT 180.325 80.685 180.605 81.565 ;
    RECT 177.005 80.685 177.285 81.565 ;
    RECT 173.685 80.685 173.965 81.565 ;
    RECT 170.365 80.685 170.645 81.565 ;
    RECT 167.045 80.685 167.325 81.565 ;
    RECT 163.725 80.685 164.005 81.565 ;
    RECT 160.405 80.685 160.685 81.565 ;
    RECT 157.085 80.685 157.365 81.565 ;
    RECT 153.765 80.685 154.045 81.565 ;
    RECT 150.445 80.685 150.725 81.565 ;
    RECT 213.525 80.685 213.805 81.565 ;
    RECT 210.205 80.685 210.485 81.565 ;
    RECT 206.885 80.685 207.165 81.565 ;
    RECT 203.565 80.685 203.845 81.565 ;
    RECT 200.245 80.685 200.525 81.565 ;
    RECT 196.925 80.685 197.205 81.565 ;
    RECT 193.605 80.685 193.885 81.565 ;
    RECT 190.285 80.685 190.565 81.565 ;
    RECT 186.965 80.685 187.245 81.565 ;
    RECT 183.645 80.685 183.925 81.565 ;
    RECT 266.645 80.685 266.925 81.565 ;
    RECT 263.325 80.685 263.605 81.565 ;
    RECT 260.005 80.685 260.285 81.565 ;
    RECT 256.685 80.685 256.965 81.565 ;
    RECT 253.365 80.685 253.645 81.565 ;
    RECT 250.045 79.965 250.325 80.845 ;
    RECT 246.725 79.965 247.005 80.845 ;
    RECT 243.405 79.965 243.685 80.845 ;
    RECT 240.085 79.965 240.365 80.845 ;
    RECT 236.765 79.965 237.045 80.845 ;
    RECT 233.445 79.965 233.725 80.845 ;
    RECT 230.125 79.965 230.405 80.845 ;
    RECT 226.805 79.965 227.085 80.845 ;
    RECT 223.485 79.965 223.765 80.845 ;
    RECT 220.165 79.965 220.445 80.845 ;
    RECT 216.845 79.965 217.125 80.845 ;
    RECT 180.325 79.965 180.605 80.845 ;
    RECT 177.005 79.965 177.285 80.845 ;
    RECT 173.685 79.965 173.965 80.845 ;
    RECT 170.365 79.965 170.645 80.845 ;
    RECT 167.045 79.965 167.325 80.845 ;
    RECT 163.725 79.965 164.005 80.845 ;
    RECT 160.405 79.965 160.685 80.845 ;
    RECT 157.085 79.965 157.365 80.845 ;
    RECT 153.765 79.965 154.045 80.845 ;
    RECT 150.445 79.965 150.725 80.845 ;
    RECT 213.525 79.965 213.805 80.845 ;
    RECT 210.205 79.965 210.485 80.845 ;
    RECT 206.885 79.965 207.165 80.845 ;
    RECT 203.565 79.965 203.845 80.845 ;
    RECT 200.245 79.965 200.525 80.845 ;
    RECT 196.925 79.965 197.205 80.845 ;
    RECT 193.605 79.965 193.885 80.845 ;
    RECT 190.285 79.965 190.565 80.845 ;
    RECT 186.965 79.965 187.245 80.845 ;
    RECT 183.645 79.965 183.925 80.845 ;
    RECT 266.645 79.965 266.925 80.845 ;
    RECT 263.325 79.965 263.605 80.845 ;
    RECT 260.005 79.965 260.285 80.845 ;
    RECT 256.685 79.965 256.965 80.845 ;
    RECT 253.365 79.965 253.645 80.845 ;
    RECT 250.045 42.505 250.325 43.385 ;
    RECT 246.725 42.505 247.005 43.385 ;
    RECT 243.405 42.505 243.685 43.385 ;
    RECT 240.085 42.505 240.365 43.385 ;
    RECT 236.765 42.505 237.045 43.385 ;
    RECT 233.445 42.505 233.725 43.385 ;
    RECT 230.125 42.505 230.405 43.385 ;
    RECT 226.805 42.505 227.085 43.385 ;
    RECT 223.485 42.505 223.765 43.385 ;
    RECT 220.165 42.505 220.445 43.385 ;
    RECT 216.845 42.505 217.125 43.385 ;
    RECT 180.325 42.505 180.605 43.385 ;
    RECT 177.005 42.505 177.285 43.385 ;
    RECT 173.685 42.505 173.965 43.385 ;
    RECT 170.365 42.505 170.645 43.385 ;
    RECT 167.045 42.505 167.325 43.385 ;
    RECT 163.725 42.505 164.005 43.385 ;
    RECT 160.405 42.505 160.685 43.385 ;
    RECT 157.085 42.505 157.365 43.385 ;
    RECT 153.765 42.505 154.045 43.385 ;
    RECT 150.445 42.505 150.725 43.385 ;
    RECT 213.525 42.505 213.805 43.385 ;
    RECT 210.205 42.505 210.485 43.385 ;
    RECT 206.885 42.505 207.165 43.385 ;
    RECT 203.565 42.505 203.845 43.385 ;
    RECT 200.245 42.505 200.525 43.385 ;
    RECT 196.925 42.505 197.205 43.385 ;
    RECT 193.605 42.505 193.885 43.385 ;
    RECT 190.285 42.505 190.565 43.385 ;
    RECT 186.965 42.505 187.245 43.385 ;
    RECT 183.645 42.505 183.925 43.385 ;
    RECT 266.645 42.505 266.925 43.385 ;
    RECT 263.325 42.505 263.605 43.385 ;
    RECT 260.005 42.505 260.285 43.385 ;
    RECT 256.685 42.505 256.965 43.385 ;
    RECT 253.365 42.505 253.645 43.385 ;
    RECT 250.045 41.785 250.325 42.665 ;
    RECT 246.725 41.785 247.005 42.665 ;
    RECT 243.405 41.785 243.685 42.665 ;
    RECT 240.085 41.785 240.365 42.665 ;
    RECT 236.765 41.785 237.045 42.665 ;
    RECT 233.445 41.785 233.725 42.665 ;
    RECT 230.125 41.785 230.405 42.665 ;
    RECT 226.805 41.785 227.085 42.665 ;
    RECT 223.485 41.785 223.765 42.665 ;
    RECT 220.165 41.785 220.445 42.665 ;
    RECT 216.845 41.785 217.125 42.665 ;
    RECT 180.325 41.785 180.605 42.665 ;
    RECT 177.005 41.785 177.285 42.665 ;
    RECT 173.685 41.785 173.965 42.665 ;
    RECT 170.365 41.785 170.645 42.665 ;
    RECT 167.045 41.785 167.325 42.665 ;
    RECT 163.725 41.785 164.005 42.665 ;
    RECT 160.405 41.785 160.685 42.665 ;
    RECT 157.085 41.785 157.365 42.665 ;
    RECT 153.765 41.785 154.045 42.665 ;
    RECT 150.445 41.785 150.725 42.665 ;
    RECT 213.525 41.785 213.805 42.665 ;
    RECT 210.205 41.785 210.485 42.665 ;
    RECT 206.885 41.785 207.165 42.665 ;
    RECT 203.565 41.785 203.845 42.665 ;
    RECT 200.245 41.785 200.525 42.665 ;
    RECT 196.925 41.785 197.205 42.665 ;
    RECT 193.605 41.785 193.885 42.665 ;
    RECT 190.285 41.785 190.565 42.665 ;
    RECT 186.965 41.785 187.245 42.665 ;
    RECT 183.645 41.785 183.925 42.665 ;
    RECT 266.645 41.785 266.925 42.665 ;
    RECT 263.325 41.785 263.605 42.665 ;
    RECT 260.005 41.785 260.285 42.665 ;
    RECT 256.685 41.785 256.965 42.665 ;
    RECT 253.365 41.785 253.645 42.665 ;
    RECT 250.045 41.065 250.325 41.945 ;
    RECT 246.725 41.065 247.005 41.945 ;
    RECT 243.405 41.065 243.685 41.945 ;
    RECT 240.085 41.065 240.365 41.945 ;
    RECT 236.765 41.065 237.045 41.945 ;
    RECT 233.445 41.065 233.725 41.945 ;
    RECT 230.125 41.065 230.405 41.945 ;
    RECT 226.805 41.065 227.085 41.945 ;
    RECT 223.485 41.065 223.765 41.945 ;
    RECT 220.165 41.065 220.445 41.945 ;
    RECT 216.845 41.065 217.125 41.945 ;
    RECT 180.325 41.065 180.605 41.945 ;
    RECT 177.005 41.065 177.285 41.945 ;
    RECT 173.685 41.065 173.965 41.945 ;
    RECT 170.365 41.065 170.645 41.945 ;
    RECT 167.045 41.065 167.325 41.945 ;
    RECT 163.725 41.065 164.005 41.945 ;
    RECT 160.405 41.065 160.685 41.945 ;
    RECT 157.085 41.065 157.365 41.945 ;
    RECT 153.765 41.065 154.045 41.945 ;
    RECT 150.445 41.065 150.725 41.945 ;
    RECT 213.525 41.065 213.805 41.945 ;
    RECT 210.205 41.065 210.485 41.945 ;
    RECT 206.885 41.065 207.165 41.945 ;
    RECT 203.565 41.065 203.845 41.945 ;
    RECT 200.245 41.065 200.525 41.945 ;
    RECT 196.925 41.065 197.205 41.945 ;
    RECT 193.605 41.065 193.885 41.945 ;
    RECT 190.285 41.065 190.565 41.945 ;
    RECT 186.965 41.065 187.245 41.945 ;
    RECT 183.645 41.065 183.925 41.945 ;
    RECT 266.645 41.065 266.925 41.945 ;
    RECT 263.325 41.065 263.605 41.945 ;
    RECT 260.005 41.065 260.285 41.945 ;
    RECT 256.685 41.065 256.965 41.945 ;
    RECT 253.365 41.065 253.645 41.945 ;
    RECT 250.045 40.345 250.325 41.225 ;
    RECT 246.725 40.345 247.005 41.225 ;
    RECT 243.405 40.345 243.685 41.225 ;
    RECT 240.085 40.345 240.365 41.225 ;
    RECT 236.765 40.345 237.045 41.225 ;
    RECT 233.445 40.345 233.725 41.225 ;
    RECT 230.125 40.345 230.405 41.225 ;
    RECT 226.805 40.345 227.085 41.225 ;
    RECT 223.485 40.345 223.765 41.225 ;
    RECT 220.165 40.345 220.445 41.225 ;
    RECT 216.845 40.345 217.125 41.225 ;
    RECT 180.325 40.345 180.605 41.225 ;
    RECT 177.005 40.345 177.285 41.225 ;
    RECT 173.685 40.345 173.965 41.225 ;
    RECT 170.365 40.345 170.645 41.225 ;
    RECT 167.045 40.345 167.325 41.225 ;
    RECT 163.725 40.345 164.005 41.225 ;
    RECT 160.405 40.345 160.685 41.225 ;
    RECT 157.085 40.345 157.365 41.225 ;
    RECT 153.765 40.345 154.045 41.225 ;
    RECT 150.445 40.345 150.725 41.225 ;
    RECT 213.525 40.345 213.805 41.225 ;
    RECT 210.205 40.345 210.485 41.225 ;
    RECT 206.885 40.345 207.165 41.225 ;
    RECT 203.565 40.345 203.845 41.225 ;
    RECT 200.245 40.345 200.525 41.225 ;
    RECT 196.925 40.345 197.205 41.225 ;
    RECT 193.605 40.345 193.885 41.225 ;
    RECT 190.285 40.345 190.565 41.225 ;
    RECT 186.965 40.345 187.245 41.225 ;
    RECT 183.645 40.345 183.925 41.225 ;
    RECT 266.645 40.345 266.925 41.225 ;
    RECT 263.325 40.345 263.605 41.225 ;
    RECT 260.005 40.345 260.285 41.225 ;
    RECT 256.685 40.345 256.965 41.225 ;
    RECT 253.365 40.345 253.645 41.225 ;
    RECT 250.045 39.625 250.325 40.505 ;
    RECT 246.725 39.625 247.005 40.505 ;
    RECT 243.405 39.625 243.685 40.505 ;
    RECT 240.085 39.625 240.365 40.505 ;
    RECT 236.765 39.625 237.045 40.505 ;
    RECT 233.445 39.625 233.725 40.505 ;
    RECT 230.125 39.625 230.405 40.505 ;
    RECT 226.805 39.625 227.085 40.505 ;
    RECT 223.485 39.625 223.765 40.505 ;
    RECT 220.165 39.625 220.445 40.505 ;
    RECT 216.845 39.625 217.125 40.505 ;
    RECT 180.325 39.625 180.605 40.505 ;
    RECT 177.005 39.625 177.285 40.505 ;
    RECT 173.685 39.625 173.965 40.505 ;
    RECT 170.365 39.625 170.645 40.505 ;
    RECT 167.045 39.625 167.325 40.505 ;
    RECT 163.725 39.625 164.005 40.505 ;
    RECT 160.405 39.625 160.685 40.505 ;
    RECT 157.085 39.625 157.365 40.505 ;
    RECT 153.765 39.625 154.045 40.505 ;
    RECT 150.445 39.625 150.725 40.505 ;
    RECT 213.525 39.625 213.805 40.505 ;
    RECT 210.205 39.625 210.485 40.505 ;
    RECT 206.885 39.625 207.165 40.505 ;
    RECT 203.565 39.625 203.845 40.505 ;
    RECT 200.245 39.625 200.525 40.505 ;
    RECT 196.925 39.625 197.205 40.505 ;
    RECT 193.605 39.625 193.885 40.505 ;
    RECT 190.285 39.625 190.565 40.505 ;
    RECT 186.965 39.625 187.245 40.505 ;
    RECT 183.645 39.625 183.925 40.505 ;
    RECT 266.645 39.625 266.925 40.505 ;
    RECT 263.325 39.625 263.605 40.505 ;
    RECT 260.005 39.625 260.285 40.505 ;
    RECT 256.685 39.625 256.965 40.505 ;
    RECT 253.365 39.625 253.645 40.505 ;
    RECT 250.045 79.245 250.325 80.125 ;
    RECT 246.725 79.245 247.005 80.125 ;
    RECT 243.405 79.245 243.685 80.125 ;
    RECT 240.085 79.245 240.365 80.125 ;
    RECT 236.765 79.245 237.045 80.125 ;
    RECT 233.445 79.245 233.725 80.125 ;
    RECT 230.125 79.245 230.405 80.125 ;
    RECT 226.805 79.245 227.085 80.125 ;
    RECT 223.485 79.245 223.765 80.125 ;
    RECT 220.165 79.245 220.445 80.125 ;
    RECT 216.845 79.245 217.125 80.125 ;
    RECT 180.325 79.245 180.605 80.125 ;
    RECT 177.005 79.245 177.285 80.125 ;
    RECT 173.685 79.245 173.965 80.125 ;
    RECT 170.365 79.245 170.645 80.125 ;
    RECT 167.045 79.245 167.325 80.125 ;
    RECT 163.725 79.245 164.005 80.125 ;
    RECT 160.405 79.245 160.685 80.125 ;
    RECT 157.085 79.245 157.365 80.125 ;
    RECT 153.765 79.245 154.045 80.125 ;
    RECT 150.445 79.245 150.725 80.125 ;
    RECT 213.525 79.245 213.805 80.125 ;
    RECT 210.205 79.245 210.485 80.125 ;
    RECT 206.885 79.245 207.165 80.125 ;
    RECT 203.565 79.245 203.845 80.125 ;
    RECT 200.245 79.245 200.525 80.125 ;
    RECT 196.925 79.245 197.205 80.125 ;
    RECT 193.605 79.245 193.885 80.125 ;
    RECT 190.285 79.245 190.565 80.125 ;
    RECT 186.965 79.245 187.245 80.125 ;
    RECT 183.645 79.245 183.925 80.125 ;
    RECT 266.645 79.245 266.925 80.125 ;
    RECT 263.325 79.245 263.605 80.125 ;
    RECT 260.005 79.245 260.285 80.125 ;
    RECT 256.685 79.245 256.965 80.125 ;
    RECT 253.365 79.245 253.645 80.125 ;
    RECT 250.045 38.905 250.325 39.785 ;
    RECT 246.725 38.905 247.005 39.785 ;
    RECT 243.405 38.905 243.685 39.785 ;
    RECT 240.085 38.905 240.365 39.785 ;
    RECT 236.765 38.905 237.045 39.785 ;
    RECT 233.445 38.905 233.725 39.785 ;
    RECT 230.125 38.905 230.405 39.785 ;
    RECT 226.805 38.905 227.085 39.785 ;
    RECT 223.485 38.905 223.765 39.785 ;
    RECT 220.165 38.905 220.445 39.785 ;
    RECT 216.845 38.905 217.125 39.785 ;
    RECT 180.325 38.905 180.605 39.785 ;
    RECT 177.005 38.905 177.285 39.785 ;
    RECT 173.685 38.905 173.965 39.785 ;
    RECT 170.365 38.905 170.645 39.785 ;
    RECT 167.045 38.905 167.325 39.785 ;
    RECT 163.725 38.905 164.005 39.785 ;
    RECT 160.405 38.905 160.685 39.785 ;
    RECT 157.085 38.905 157.365 39.785 ;
    RECT 153.765 38.905 154.045 39.785 ;
    RECT 150.445 38.905 150.725 39.785 ;
    RECT 213.525 38.905 213.805 39.785 ;
    RECT 210.205 38.905 210.485 39.785 ;
    RECT 206.885 38.905 207.165 39.785 ;
    RECT 203.565 38.905 203.845 39.785 ;
    RECT 200.245 38.905 200.525 39.785 ;
    RECT 196.925 38.905 197.205 39.785 ;
    RECT 193.605 38.905 193.885 39.785 ;
    RECT 190.285 38.905 190.565 39.785 ;
    RECT 186.965 38.905 187.245 39.785 ;
    RECT 183.645 38.905 183.925 39.785 ;
    RECT 266.645 38.905 266.925 39.785 ;
    RECT 263.325 38.905 263.605 39.785 ;
    RECT 260.005 38.905 260.285 39.785 ;
    RECT 256.685 38.905 256.965 39.785 ;
    RECT 253.365 38.905 253.645 39.785 ;
    RECT 250.045 78.525 250.325 79.405 ;
    RECT 246.725 78.525 247.005 79.405 ;
    RECT 243.405 78.525 243.685 79.405 ;
    RECT 240.085 78.525 240.365 79.405 ;
    RECT 236.765 78.525 237.045 79.405 ;
    RECT 233.445 78.525 233.725 79.405 ;
    RECT 230.125 78.525 230.405 79.405 ;
    RECT 226.805 78.525 227.085 79.405 ;
    RECT 223.485 78.525 223.765 79.405 ;
    RECT 220.165 78.525 220.445 79.405 ;
    RECT 216.845 78.525 217.125 79.405 ;
    RECT 180.325 78.525 180.605 79.405 ;
    RECT 177.005 78.525 177.285 79.405 ;
    RECT 173.685 78.525 173.965 79.405 ;
    RECT 170.365 78.525 170.645 79.405 ;
    RECT 167.045 78.525 167.325 79.405 ;
    RECT 163.725 78.525 164.005 79.405 ;
    RECT 160.405 78.525 160.685 79.405 ;
    RECT 157.085 78.525 157.365 79.405 ;
    RECT 153.765 78.525 154.045 79.405 ;
    RECT 150.445 78.525 150.725 79.405 ;
    RECT 213.525 78.525 213.805 79.405 ;
    RECT 210.205 78.525 210.485 79.405 ;
    RECT 206.885 78.525 207.165 79.405 ;
    RECT 203.565 78.525 203.845 79.405 ;
    RECT 200.245 78.525 200.525 79.405 ;
    RECT 196.925 78.525 197.205 79.405 ;
    RECT 193.605 78.525 193.885 79.405 ;
    RECT 190.285 78.525 190.565 79.405 ;
    RECT 186.965 78.525 187.245 79.405 ;
    RECT 183.645 78.525 183.925 79.405 ;
    RECT 266.645 78.525 266.925 79.405 ;
    RECT 263.325 78.525 263.605 79.405 ;
    RECT 260.005 78.525 260.285 79.405 ;
    RECT 256.685 78.525 256.965 79.405 ;
    RECT 253.365 78.525 253.645 79.405 ;
    RECT 250.045 38.185 250.325 39.065 ;
    RECT 246.725 38.185 247.005 39.065 ;
    RECT 243.405 38.185 243.685 39.065 ;
    RECT 240.085 38.185 240.365 39.065 ;
    RECT 236.765 38.185 237.045 39.065 ;
    RECT 233.445 38.185 233.725 39.065 ;
    RECT 230.125 38.185 230.405 39.065 ;
    RECT 226.805 38.185 227.085 39.065 ;
    RECT 223.485 38.185 223.765 39.065 ;
    RECT 220.165 38.185 220.445 39.065 ;
    RECT 216.845 38.185 217.125 39.065 ;
    RECT 180.325 38.185 180.605 39.065 ;
    RECT 177.005 38.185 177.285 39.065 ;
    RECT 173.685 38.185 173.965 39.065 ;
    RECT 170.365 38.185 170.645 39.065 ;
    RECT 167.045 38.185 167.325 39.065 ;
    RECT 163.725 38.185 164.005 39.065 ;
    RECT 160.405 38.185 160.685 39.065 ;
    RECT 157.085 38.185 157.365 39.065 ;
    RECT 153.765 38.185 154.045 39.065 ;
    RECT 150.445 38.185 150.725 39.065 ;
    RECT 213.525 38.185 213.805 39.065 ;
    RECT 210.205 38.185 210.485 39.065 ;
    RECT 206.885 38.185 207.165 39.065 ;
    RECT 203.565 38.185 203.845 39.065 ;
    RECT 200.245 38.185 200.525 39.065 ;
    RECT 196.925 38.185 197.205 39.065 ;
    RECT 193.605 38.185 193.885 39.065 ;
    RECT 190.285 38.185 190.565 39.065 ;
    RECT 186.965 38.185 187.245 39.065 ;
    RECT 183.645 38.185 183.925 39.065 ;
    RECT 266.645 38.185 266.925 39.065 ;
    RECT 263.325 38.185 263.605 39.065 ;
    RECT 260.005 38.185 260.285 39.065 ;
    RECT 256.685 38.185 256.965 39.065 ;
    RECT 253.365 38.185 253.645 39.065 ;
    RECT 250.045 77.805 250.325 78.685 ;
    RECT 246.725 77.805 247.005 78.685 ;
    RECT 243.405 77.805 243.685 78.685 ;
    RECT 240.085 77.805 240.365 78.685 ;
    RECT 236.765 77.805 237.045 78.685 ;
    RECT 233.445 77.805 233.725 78.685 ;
    RECT 230.125 77.805 230.405 78.685 ;
    RECT 226.805 77.805 227.085 78.685 ;
    RECT 223.485 77.805 223.765 78.685 ;
    RECT 220.165 77.805 220.445 78.685 ;
    RECT 216.845 77.805 217.125 78.685 ;
    RECT 180.325 77.805 180.605 78.685 ;
    RECT 177.005 77.805 177.285 78.685 ;
    RECT 173.685 77.805 173.965 78.685 ;
    RECT 170.365 77.805 170.645 78.685 ;
    RECT 167.045 77.805 167.325 78.685 ;
    RECT 163.725 77.805 164.005 78.685 ;
    RECT 160.405 77.805 160.685 78.685 ;
    RECT 157.085 77.805 157.365 78.685 ;
    RECT 153.765 77.805 154.045 78.685 ;
    RECT 150.445 77.805 150.725 78.685 ;
    RECT 213.525 77.805 213.805 78.685 ;
    RECT 210.205 77.805 210.485 78.685 ;
    RECT 206.885 77.805 207.165 78.685 ;
    RECT 203.565 77.805 203.845 78.685 ;
    RECT 200.245 77.805 200.525 78.685 ;
    RECT 196.925 77.805 197.205 78.685 ;
    RECT 193.605 77.805 193.885 78.685 ;
    RECT 190.285 77.805 190.565 78.685 ;
    RECT 186.965 77.805 187.245 78.685 ;
    RECT 183.645 77.805 183.925 78.685 ;
    RECT 266.645 77.805 266.925 78.685 ;
    RECT 263.325 77.805 263.605 78.685 ;
    RECT 260.005 77.805 260.285 78.685 ;
    RECT 256.685 77.805 256.965 78.685 ;
    RECT 253.365 77.805 253.645 78.685 ;
    RECT 250.045 37.465 250.325 38.345 ;
    RECT 246.725 37.465 247.005 38.345 ;
    RECT 243.405 37.465 243.685 38.345 ;
    RECT 240.085 37.465 240.365 38.345 ;
    RECT 236.765 37.465 237.045 38.345 ;
    RECT 233.445 37.465 233.725 38.345 ;
    RECT 230.125 37.465 230.405 38.345 ;
    RECT 226.805 37.465 227.085 38.345 ;
    RECT 223.485 37.465 223.765 38.345 ;
    RECT 220.165 37.465 220.445 38.345 ;
    RECT 216.845 37.465 217.125 38.345 ;
    RECT 180.325 37.465 180.605 38.345 ;
    RECT 177.005 37.465 177.285 38.345 ;
    RECT 173.685 37.465 173.965 38.345 ;
    RECT 170.365 37.465 170.645 38.345 ;
    RECT 167.045 37.465 167.325 38.345 ;
    RECT 163.725 37.465 164.005 38.345 ;
    RECT 160.405 37.465 160.685 38.345 ;
    RECT 157.085 37.465 157.365 38.345 ;
    RECT 153.765 37.465 154.045 38.345 ;
    RECT 150.445 37.465 150.725 38.345 ;
    RECT 213.525 37.465 213.805 38.345 ;
    RECT 210.205 37.465 210.485 38.345 ;
    RECT 206.885 37.465 207.165 38.345 ;
    RECT 203.565 37.465 203.845 38.345 ;
    RECT 200.245 37.465 200.525 38.345 ;
    RECT 196.925 37.465 197.205 38.345 ;
    RECT 193.605 37.465 193.885 38.345 ;
    RECT 190.285 37.465 190.565 38.345 ;
    RECT 186.965 37.465 187.245 38.345 ;
    RECT 183.645 37.465 183.925 38.345 ;
    RECT 266.645 37.465 266.925 38.345 ;
    RECT 263.325 37.465 263.605 38.345 ;
    RECT 260.005 37.465 260.285 38.345 ;
    RECT 256.685 37.465 256.965 38.345 ;
    RECT 253.365 37.465 253.645 38.345 ;
    RECT 250.045 77.085 250.325 77.965 ;
    RECT 246.725 77.085 247.005 77.965 ;
    RECT 243.405 77.085 243.685 77.965 ;
    RECT 240.085 77.085 240.365 77.965 ;
    RECT 236.765 77.085 237.045 77.965 ;
    RECT 233.445 77.085 233.725 77.965 ;
    RECT 230.125 77.085 230.405 77.965 ;
    RECT 226.805 77.085 227.085 77.965 ;
    RECT 223.485 77.085 223.765 77.965 ;
    RECT 220.165 77.085 220.445 77.965 ;
    RECT 216.845 77.085 217.125 77.965 ;
    RECT 180.325 77.085 180.605 77.965 ;
    RECT 177.005 77.085 177.285 77.965 ;
    RECT 173.685 77.085 173.965 77.965 ;
    RECT 170.365 77.085 170.645 77.965 ;
    RECT 167.045 77.085 167.325 77.965 ;
    RECT 163.725 77.085 164.005 77.965 ;
    RECT 160.405 77.085 160.685 77.965 ;
    RECT 157.085 77.085 157.365 77.965 ;
    RECT 153.765 77.085 154.045 77.965 ;
    RECT 150.445 77.085 150.725 77.965 ;
    RECT 213.525 77.085 213.805 77.965 ;
    RECT 210.205 77.085 210.485 77.965 ;
    RECT 206.885 77.085 207.165 77.965 ;
    RECT 203.565 77.085 203.845 77.965 ;
    RECT 200.245 77.085 200.525 77.965 ;
    RECT 196.925 77.085 197.205 77.965 ;
    RECT 193.605 77.085 193.885 77.965 ;
    RECT 190.285 77.085 190.565 77.965 ;
    RECT 186.965 77.085 187.245 77.965 ;
    RECT 183.645 77.085 183.925 77.965 ;
    RECT 266.645 77.085 266.925 77.965 ;
    RECT 263.325 77.085 263.605 77.965 ;
    RECT 260.005 77.085 260.285 77.965 ;
    RECT 256.685 77.085 256.965 77.965 ;
    RECT 253.365 77.085 253.645 77.965 ;
    RECT 250.045 36.745 250.325 37.625 ;
    RECT 246.725 36.745 247.005 37.625 ;
    RECT 243.405 36.745 243.685 37.625 ;
    RECT 240.085 36.745 240.365 37.625 ;
    RECT 236.765 36.745 237.045 37.625 ;
    RECT 233.445 36.745 233.725 37.625 ;
    RECT 230.125 36.745 230.405 37.625 ;
    RECT 226.805 36.745 227.085 37.625 ;
    RECT 223.485 36.745 223.765 37.625 ;
    RECT 220.165 36.745 220.445 37.625 ;
    RECT 216.845 36.745 217.125 37.625 ;
    RECT 180.325 36.745 180.605 37.625 ;
    RECT 177.005 36.745 177.285 37.625 ;
    RECT 173.685 36.745 173.965 37.625 ;
    RECT 170.365 36.745 170.645 37.625 ;
    RECT 167.045 36.745 167.325 37.625 ;
    RECT 163.725 36.745 164.005 37.625 ;
    RECT 160.405 36.745 160.685 37.625 ;
    RECT 157.085 36.745 157.365 37.625 ;
    RECT 153.765 36.745 154.045 37.625 ;
    RECT 150.445 36.745 150.725 37.625 ;
    RECT 213.525 36.745 213.805 37.625 ;
    RECT 210.205 36.745 210.485 37.625 ;
    RECT 206.885 36.745 207.165 37.625 ;
    RECT 203.565 36.745 203.845 37.625 ;
    RECT 200.245 36.745 200.525 37.625 ;
    RECT 196.925 36.745 197.205 37.625 ;
    RECT 193.605 36.745 193.885 37.625 ;
    RECT 190.285 36.745 190.565 37.625 ;
    RECT 186.965 36.745 187.245 37.625 ;
    RECT 183.645 36.745 183.925 37.625 ;
    RECT 266.645 36.745 266.925 37.625 ;
    RECT 263.325 36.745 263.605 37.625 ;
    RECT 260.005 36.745 260.285 37.625 ;
    RECT 256.685 36.745 256.965 37.625 ;
    RECT 253.365 36.745 253.645 37.625 ;
    RECT 250.045 76.365 250.325 77.245 ;
    RECT 246.725 76.365 247.005 77.245 ;
    RECT 243.405 76.365 243.685 77.245 ;
    RECT 240.085 76.365 240.365 77.245 ;
    RECT 236.765 76.365 237.045 77.245 ;
    RECT 233.445 76.365 233.725 77.245 ;
    RECT 230.125 76.365 230.405 77.245 ;
    RECT 226.805 76.365 227.085 77.245 ;
    RECT 223.485 76.365 223.765 77.245 ;
    RECT 220.165 76.365 220.445 77.245 ;
    RECT 216.845 76.365 217.125 77.245 ;
    RECT 180.325 76.365 180.605 77.245 ;
    RECT 177.005 76.365 177.285 77.245 ;
    RECT 173.685 76.365 173.965 77.245 ;
    RECT 170.365 76.365 170.645 77.245 ;
    RECT 167.045 76.365 167.325 77.245 ;
    RECT 163.725 76.365 164.005 77.245 ;
    RECT 160.405 76.365 160.685 77.245 ;
    RECT 157.085 76.365 157.365 77.245 ;
    RECT 153.765 76.365 154.045 77.245 ;
    RECT 150.445 76.365 150.725 77.245 ;
    RECT 213.525 76.365 213.805 77.245 ;
    RECT 210.205 76.365 210.485 77.245 ;
    RECT 206.885 76.365 207.165 77.245 ;
    RECT 203.565 76.365 203.845 77.245 ;
    RECT 200.245 76.365 200.525 77.245 ;
    RECT 196.925 76.365 197.205 77.245 ;
    RECT 193.605 76.365 193.885 77.245 ;
    RECT 190.285 76.365 190.565 77.245 ;
    RECT 186.965 76.365 187.245 77.245 ;
    RECT 183.645 76.365 183.925 77.245 ;
    RECT 266.645 76.365 266.925 77.245 ;
    RECT 263.325 76.365 263.605 77.245 ;
    RECT 260.005 76.365 260.285 77.245 ;
    RECT 256.685 76.365 256.965 77.245 ;
    RECT 253.365 76.365 253.645 77.245 ;
    RECT 61.215 52.585 61.495 53.465 ;
    RECT 57.895 52.585 58.175 53.465 ;
    RECT 54.575 52.585 54.855 53.465 ;
    RECT 51.255 52.585 51.535 53.465 ;
    RECT 47.935 52.585 48.215 53.465 ;
    RECT 44.615 52.585 44.895 53.465 ;
    RECT 41.295 52.585 41.575 53.465 ;
    RECT 37.975 52.585 38.255 53.465 ;
    RECT 34.655 52.585 34.935 53.465 ;
    RECT 117.655 52.585 117.935 53.465 ;
    RECT 114.335 52.585 114.615 53.465 ;
    RECT 111.015 52.585 111.295 53.465 ;
    RECT 107.695 52.585 107.975 53.465 ;
    RECT 104.375 52.585 104.655 53.465 ;
    RECT 101.055 52.585 101.335 53.465 ;
    RECT 97.735 52.585 98.015 53.465 ;
    RECT 94.415 52.585 94.695 53.465 ;
    RECT 91.095 52.585 91.375 53.465 ;
    RECT 87.775 52.585 88.055 53.465 ;
    RECT 84.455 52.585 84.735 53.465 ;
    RECT 81.135 52.585 81.415 53.465 ;
    RECT 77.815 52.585 78.095 53.465 ;
    RECT 74.495 52.585 74.775 53.465 ;
    RECT 71.175 52.585 71.455 53.465 ;
    RECT 31.335 52.585 31.615 53.465 ;
    RECT 67.855 52.585 68.135 53.465 ;
    RECT 28.015 52.585 28.295 53.465 ;
    RECT 24.695 52.585 24.975 53.465 ;
    RECT 21.375 52.585 21.655 53.465 ;
    RECT 18.055 52.585 18.335 53.465 ;
    RECT 14.735 52.585 15.015 53.465 ;
    RECT 11.415 52.585 11.695 53.465 ;
    RECT 8.095 52.585 8.375 53.465 ;
    RECT 4.775 52.585 5.055 53.465 ;
    RECT 1.455 52.585 1.735 53.465 ;
    RECT 64.535 52.585 64.815 53.465 ;
    RECT 61.215 51.865 61.495 52.745 ;
    RECT 57.895 51.865 58.175 52.745 ;
    RECT 54.575 51.865 54.855 52.745 ;
    RECT 51.255 51.865 51.535 52.745 ;
    RECT 47.935 51.865 48.215 52.745 ;
    RECT 44.615 51.865 44.895 52.745 ;
    RECT 41.295 51.865 41.575 52.745 ;
    RECT 37.975 51.865 38.255 52.745 ;
    RECT 34.655 51.865 34.935 52.745 ;
    RECT 117.655 51.865 117.935 52.745 ;
    RECT 114.335 51.865 114.615 52.745 ;
    RECT 111.015 51.865 111.295 52.745 ;
    RECT 107.695 51.865 107.975 52.745 ;
    RECT 104.375 51.865 104.655 52.745 ;
    RECT 101.055 51.865 101.335 52.745 ;
    RECT 97.735 51.865 98.015 52.745 ;
    RECT 94.415 51.865 94.695 52.745 ;
    RECT 91.095 51.865 91.375 52.745 ;
    RECT 87.775 51.865 88.055 52.745 ;
    RECT 84.455 51.865 84.735 52.745 ;
    RECT 81.135 51.865 81.415 52.745 ;
    RECT 77.815 51.865 78.095 52.745 ;
    RECT 74.495 51.865 74.775 52.745 ;
    RECT 71.175 51.865 71.455 52.745 ;
    RECT 31.335 51.865 31.615 52.745 ;
    RECT 67.855 51.865 68.135 52.745 ;
    RECT 28.015 51.865 28.295 52.745 ;
    RECT 24.695 51.865 24.975 52.745 ;
    RECT 21.375 51.865 21.655 52.745 ;
    RECT 18.055 51.865 18.335 52.745 ;
    RECT 14.735 51.865 15.015 52.745 ;
    RECT 11.415 51.865 11.695 52.745 ;
    RECT 8.095 51.865 8.375 52.745 ;
    RECT 4.775 51.865 5.055 52.745 ;
    RECT 1.455 51.865 1.735 52.745 ;
    RECT 64.535 51.865 64.815 52.745 ;
    RECT 61.215 51.145 61.495 52.025 ;
    RECT 57.895 51.145 58.175 52.025 ;
    RECT 54.575 51.145 54.855 52.025 ;
    RECT 51.255 51.145 51.535 52.025 ;
    RECT 47.935 51.145 48.215 52.025 ;
    RECT 44.615 51.145 44.895 52.025 ;
    RECT 41.295 51.145 41.575 52.025 ;
    RECT 37.975 51.145 38.255 52.025 ;
    RECT 34.655 51.145 34.935 52.025 ;
    RECT 117.655 51.145 117.935 52.025 ;
    RECT 114.335 51.145 114.615 52.025 ;
    RECT 111.015 51.145 111.295 52.025 ;
    RECT 107.695 51.145 107.975 52.025 ;
    RECT 104.375 51.145 104.655 52.025 ;
    RECT 101.055 51.145 101.335 52.025 ;
    RECT 97.735 51.145 98.015 52.025 ;
    RECT 94.415 51.145 94.695 52.025 ;
    RECT 91.095 51.145 91.375 52.025 ;
    RECT 87.775 51.145 88.055 52.025 ;
    RECT 84.455 51.145 84.735 52.025 ;
    RECT 81.135 51.145 81.415 52.025 ;
    RECT 77.815 51.145 78.095 52.025 ;
    RECT 74.495 51.145 74.775 52.025 ;
    RECT 71.175 51.145 71.455 52.025 ;
    RECT 31.335 51.145 31.615 52.025 ;
    RECT 67.855 51.145 68.135 52.025 ;
    RECT 28.015 51.145 28.295 52.025 ;
    RECT 24.695 51.145 24.975 52.025 ;
    RECT 21.375 51.145 21.655 52.025 ;
    RECT 18.055 51.145 18.335 52.025 ;
    RECT 14.735 51.145 15.015 52.025 ;
    RECT 11.415 51.145 11.695 52.025 ;
    RECT 8.095 51.145 8.375 52.025 ;
    RECT 4.775 51.145 5.055 52.025 ;
    RECT 1.455 51.145 1.735 52.025 ;
    RECT 64.535 51.145 64.815 52.025 ;
    RECT 61.215 50.425 61.495 51.305 ;
    RECT 57.895 50.425 58.175 51.305 ;
    RECT 54.575 50.425 54.855 51.305 ;
    RECT 51.255 50.425 51.535 51.305 ;
    RECT 47.935 50.425 48.215 51.305 ;
    RECT 44.615 50.425 44.895 51.305 ;
    RECT 41.295 50.425 41.575 51.305 ;
    RECT 37.975 50.425 38.255 51.305 ;
    RECT 34.655 50.425 34.935 51.305 ;
    RECT 117.655 50.425 117.935 51.305 ;
    RECT 114.335 50.425 114.615 51.305 ;
    RECT 111.015 50.425 111.295 51.305 ;
    RECT 107.695 50.425 107.975 51.305 ;
    RECT 104.375 50.425 104.655 51.305 ;
    RECT 101.055 50.425 101.335 51.305 ;
    RECT 97.735 50.425 98.015 51.305 ;
    RECT 94.415 50.425 94.695 51.305 ;
    RECT 91.095 50.425 91.375 51.305 ;
    RECT 87.775 50.425 88.055 51.305 ;
    RECT 84.455 50.425 84.735 51.305 ;
    RECT 81.135 50.425 81.415 51.305 ;
    RECT 77.815 50.425 78.095 51.305 ;
    RECT 74.495 50.425 74.775 51.305 ;
    RECT 71.175 50.425 71.455 51.305 ;
    RECT 31.335 50.425 31.615 51.305 ;
    RECT 67.855 50.425 68.135 51.305 ;
    RECT 28.015 50.425 28.295 51.305 ;
    RECT 24.695 50.425 24.975 51.305 ;
    RECT 21.375 50.425 21.655 51.305 ;
    RECT 18.055 50.425 18.335 51.305 ;
    RECT 14.735 50.425 15.015 51.305 ;
    RECT 11.415 50.425 11.695 51.305 ;
    RECT 8.095 50.425 8.375 51.305 ;
    RECT 4.775 50.425 5.055 51.305 ;
    RECT 1.455 50.425 1.735 51.305 ;
    RECT 64.535 50.425 64.815 51.305 ;
    RECT 61.215 93.645 61.495 94.525 ;
    RECT 57.895 93.645 58.175 94.525 ;
    RECT 54.575 93.645 54.855 94.525 ;
    RECT 51.255 93.645 51.535 94.525 ;
    RECT 47.935 93.645 48.215 94.525 ;
    RECT 44.615 93.645 44.895 94.525 ;
    RECT 41.295 93.645 41.575 94.525 ;
    RECT 37.975 93.645 38.255 94.525 ;
    RECT 34.655 93.645 34.935 94.525 ;
    RECT 117.655 93.645 117.935 94.525 ;
    RECT 114.335 93.645 114.615 94.525 ;
    RECT 111.015 93.645 111.295 94.525 ;
    RECT 107.695 93.645 107.975 94.525 ;
    RECT 104.375 93.645 104.655 94.525 ;
    RECT 101.055 93.645 101.335 94.525 ;
    RECT 97.735 93.645 98.015 94.525 ;
    RECT 94.415 93.645 94.695 94.525 ;
    RECT 91.095 93.645 91.375 94.525 ;
    RECT 87.775 93.645 88.055 94.525 ;
    RECT 84.455 93.645 84.735 94.525 ;
    RECT 81.135 93.645 81.415 94.525 ;
    RECT 77.815 93.645 78.095 94.525 ;
    RECT 74.495 93.645 74.775 94.525 ;
    RECT 71.175 93.645 71.455 94.525 ;
    RECT 31.335 93.645 31.615 94.525 ;
    RECT 67.855 93.645 68.135 94.525 ;
    RECT 28.015 93.645 28.295 94.525 ;
    RECT 24.695 93.645 24.975 94.525 ;
    RECT 21.375 93.645 21.655 94.525 ;
    RECT 18.055 93.645 18.335 94.525 ;
    RECT 14.735 93.645 15.015 94.525 ;
    RECT 11.415 93.645 11.695 94.525 ;
    RECT 8.095 93.645 8.375 94.525 ;
    RECT 4.775 93.645 5.055 94.525 ;
    RECT 1.455 93.645 1.735 94.525 ;
    RECT 64.535 93.645 64.815 94.525 ;
    RECT 61.215 92.925 61.495 93.805 ;
    RECT 57.895 92.925 58.175 93.805 ;
    RECT 54.575 92.925 54.855 93.805 ;
    RECT 51.255 92.925 51.535 93.805 ;
    RECT 47.935 92.925 48.215 93.805 ;
    RECT 44.615 92.925 44.895 93.805 ;
    RECT 41.295 92.925 41.575 93.805 ;
    RECT 37.975 92.925 38.255 93.805 ;
    RECT 34.655 92.925 34.935 93.805 ;
    RECT 117.655 92.925 117.935 93.805 ;
    RECT 114.335 92.925 114.615 93.805 ;
    RECT 111.015 92.925 111.295 93.805 ;
    RECT 107.695 92.925 107.975 93.805 ;
    RECT 104.375 92.925 104.655 93.805 ;
    RECT 101.055 92.925 101.335 93.805 ;
    RECT 97.735 92.925 98.015 93.805 ;
    RECT 94.415 92.925 94.695 93.805 ;
    RECT 91.095 92.925 91.375 93.805 ;
    RECT 87.775 92.925 88.055 93.805 ;
    RECT 84.455 92.925 84.735 93.805 ;
    RECT 81.135 92.925 81.415 93.805 ;
    RECT 77.815 92.925 78.095 93.805 ;
    RECT 74.495 92.925 74.775 93.805 ;
    RECT 71.175 92.925 71.455 93.805 ;
    RECT 31.335 92.925 31.615 93.805 ;
    RECT 67.855 92.925 68.135 93.805 ;
    RECT 28.015 92.925 28.295 93.805 ;
    RECT 24.695 92.925 24.975 93.805 ;
    RECT 21.375 92.925 21.655 93.805 ;
    RECT 18.055 92.925 18.335 93.805 ;
    RECT 14.735 92.925 15.015 93.805 ;
    RECT 11.415 92.925 11.695 93.805 ;
    RECT 8.095 92.925 8.375 93.805 ;
    RECT 4.775 92.925 5.055 93.805 ;
    RECT 1.455 92.925 1.735 93.805 ;
    RECT 64.535 92.925 64.815 93.805 ;
    RECT 61.215 92.205 61.495 93.085 ;
    RECT 57.895 92.205 58.175 93.085 ;
    RECT 54.575 92.205 54.855 93.085 ;
    RECT 51.255 92.205 51.535 93.085 ;
    RECT 47.935 92.205 48.215 93.085 ;
    RECT 44.615 92.205 44.895 93.085 ;
    RECT 41.295 92.205 41.575 93.085 ;
    RECT 37.975 92.205 38.255 93.085 ;
    RECT 34.655 92.205 34.935 93.085 ;
    RECT 117.655 92.205 117.935 93.085 ;
    RECT 114.335 92.205 114.615 93.085 ;
    RECT 111.015 92.205 111.295 93.085 ;
    RECT 107.695 92.205 107.975 93.085 ;
    RECT 104.375 92.205 104.655 93.085 ;
    RECT 101.055 92.205 101.335 93.085 ;
    RECT 97.735 92.205 98.015 93.085 ;
    RECT 94.415 92.205 94.695 93.085 ;
    RECT 91.095 92.205 91.375 93.085 ;
    RECT 87.775 92.205 88.055 93.085 ;
    RECT 84.455 92.205 84.735 93.085 ;
    RECT 81.135 92.205 81.415 93.085 ;
    RECT 77.815 92.205 78.095 93.085 ;
    RECT 74.495 92.205 74.775 93.085 ;
    RECT 71.175 92.205 71.455 93.085 ;
    RECT 31.335 92.205 31.615 93.085 ;
    RECT 67.855 92.205 68.135 93.085 ;
    RECT 28.015 92.205 28.295 93.085 ;
    RECT 24.695 92.205 24.975 93.085 ;
    RECT 21.375 92.205 21.655 93.085 ;
    RECT 18.055 92.205 18.335 93.085 ;
    RECT 14.735 92.205 15.015 93.085 ;
    RECT 11.415 92.205 11.695 93.085 ;
    RECT 8.095 92.205 8.375 93.085 ;
    RECT 4.775 92.205 5.055 93.085 ;
    RECT 1.455 92.205 1.735 93.085 ;
    RECT 64.535 92.205 64.815 93.085 ;
    RECT 61.215 91.485 61.495 92.365 ;
    RECT 57.895 91.485 58.175 92.365 ;
    RECT 54.575 91.485 54.855 92.365 ;
    RECT 51.255 91.485 51.535 92.365 ;
    RECT 47.935 91.485 48.215 92.365 ;
    RECT 44.615 91.485 44.895 92.365 ;
    RECT 41.295 91.485 41.575 92.365 ;
    RECT 37.975 91.485 38.255 92.365 ;
    RECT 34.655 91.485 34.935 92.365 ;
    RECT 117.655 91.485 117.935 92.365 ;
    RECT 114.335 91.485 114.615 92.365 ;
    RECT 111.015 91.485 111.295 92.365 ;
    RECT 107.695 91.485 107.975 92.365 ;
    RECT 104.375 91.485 104.655 92.365 ;
    RECT 101.055 91.485 101.335 92.365 ;
    RECT 97.735 91.485 98.015 92.365 ;
    RECT 94.415 91.485 94.695 92.365 ;
    RECT 91.095 91.485 91.375 92.365 ;
    RECT 87.775 91.485 88.055 92.365 ;
    RECT 84.455 91.485 84.735 92.365 ;
    RECT 81.135 91.485 81.415 92.365 ;
    RECT 77.815 91.485 78.095 92.365 ;
    RECT 74.495 91.485 74.775 92.365 ;
    RECT 71.175 91.485 71.455 92.365 ;
    RECT 31.335 91.485 31.615 92.365 ;
    RECT 67.855 91.485 68.135 92.365 ;
    RECT 28.015 91.485 28.295 92.365 ;
    RECT 24.695 91.485 24.975 92.365 ;
    RECT 21.375 91.485 21.655 92.365 ;
    RECT 18.055 91.485 18.335 92.365 ;
    RECT 14.735 91.485 15.015 92.365 ;
    RECT 11.415 91.485 11.695 92.365 ;
    RECT 8.095 91.485 8.375 92.365 ;
    RECT 4.775 91.485 5.055 92.365 ;
    RECT 1.455 91.485 1.735 92.365 ;
    RECT 64.535 91.485 64.815 92.365 ;
    RECT 61.215 90.765 61.495 91.645 ;
    RECT 57.895 90.765 58.175 91.645 ;
    RECT 54.575 90.765 54.855 91.645 ;
    RECT 51.255 90.765 51.535 91.645 ;
    RECT 47.935 90.765 48.215 91.645 ;
    RECT 44.615 90.765 44.895 91.645 ;
    RECT 41.295 90.765 41.575 91.645 ;
    RECT 37.975 90.765 38.255 91.645 ;
    RECT 34.655 90.765 34.935 91.645 ;
    RECT 117.655 90.765 117.935 91.645 ;
    RECT 114.335 90.765 114.615 91.645 ;
    RECT 111.015 90.765 111.295 91.645 ;
    RECT 107.695 90.765 107.975 91.645 ;
    RECT 104.375 90.765 104.655 91.645 ;
    RECT 101.055 90.765 101.335 91.645 ;
    RECT 97.735 90.765 98.015 91.645 ;
    RECT 94.415 90.765 94.695 91.645 ;
    RECT 91.095 90.765 91.375 91.645 ;
    RECT 87.775 90.765 88.055 91.645 ;
    RECT 84.455 90.765 84.735 91.645 ;
    RECT 81.135 90.765 81.415 91.645 ;
    RECT 77.815 90.765 78.095 91.645 ;
    RECT 74.495 90.765 74.775 91.645 ;
    RECT 71.175 90.765 71.455 91.645 ;
    RECT 31.335 90.765 31.615 91.645 ;
    RECT 67.855 90.765 68.135 91.645 ;
    RECT 28.015 90.765 28.295 91.645 ;
    RECT 24.695 90.765 24.975 91.645 ;
    RECT 21.375 90.765 21.655 91.645 ;
    RECT 18.055 90.765 18.335 91.645 ;
    RECT 14.735 90.765 15.015 91.645 ;
    RECT 11.415 90.765 11.695 91.645 ;
    RECT 8.095 90.765 8.375 91.645 ;
    RECT 4.775 90.765 5.055 91.645 ;
    RECT 1.455 90.765 1.735 91.645 ;
    RECT 64.535 90.765 64.815 91.645 ;
    RECT 61.215 90.045 61.495 90.925 ;
    RECT 57.895 90.045 58.175 90.925 ;
    RECT 54.575 90.045 54.855 90.925 ;
    RECT 51.255 90.045 51.535 90.925 ;
    RECT 47.935 90.045 48.215 90.925 ;
    RECT 44.615 90.045 44.895 90.925 ;
    RECT 41.295 90.045 41.575 90.925 ;
    RECT 37.975 90.045 38.255 90.925 ;
    RECT 34.655 90.045 34.935 90.925 ;
    RECT 117.655 90.045 117.935 90.925 ;
    RECT 114.335 90.045 114.615 90.925 ;
    RECT 111.015 90.045 111.295 90.925 ;
    RECT 107.695 90.045 107.975 90.925 ;
    RECT 104.375 90.045 104.655 90.925 ;
    RECT 101.055 90.045 101.335 90.925 ;
    RECT 97.735 90.045 98.015 90.925 ;
    RECT 94.415 90.045 94.695 90.925 ;
    RECT 91.095 90.045 91.375 90.925 ;
    RECT 87.775 90.045 88.055 90.925 ;
    RECT 84.455 90.045 84.735 90.925 ;
    RECT 81.135 90.045 81.415 90.925 ;
    RECT 77.815 90.045 78.095 90.925 ;
    RECT 74.495 90.045 74.775 90.925 ;
    RECT 71.175 90.045 71.455 90.925 ;
    RECT 31.335 90.045 31.615 90.925 ;
    RECT 67.855 90.045 68.135 90.925 ;
    RECT 28.015 90.045 28.295 90.925 ;
    RECT 24.695 90.045 24.975 90.925 ;
    RECT 21.375 90.045 21.655 90.925 ;
    RECT 18.055 90.045 18.335 90.925 ;
    RECT 14.735 90.045 15.015 90.925 ;
    RECT 11.415 90.045 11.695 90.925 ;
    RECT 8.095 90.045 8.375 90.925 ;
    RECT 4.775 90.045 5.055 90.925 ;
    RECT 1.455 90.045 1.735 90.925 ;
    RECT 64.535 90.045 64.815 90.925 ;
    RECT 61.215 89.325 61.495 90.205 ;
    RECT 57.895 89.325 58.175 90.205 ;
    RECT 54.575 89.325 54.855 90.205 ;
    RECT 51.255 89.325 51.535 90.205 ;
    RECT 47.935 89.325 48.215 90.205 ;
    RECT 44.615 89.325 44.895 90.205 ;
    RECT 41.295 89.325 41.575 90.205 ;
    RECT 37.975 89.325 38.255 90.205 ;
    RECT 34.655 89.325 34.935 90.205 ;
    RECT 117.655 89.325 117.935 90.205 ;
    RECT 114.335 89.325 114.615 90.205 ;
    RECT 111.015 89.325 111.295 90.205 ;
    RECT 107.695 89.325 107.975 90.205 ;
    RECT 104.375 89.325 104.655 90.205 ;
    RECT 101.055 89.325 101.335 90.205 ;
    RECT 97.735 89.325 98.015 90.205 ;
    RECT 94.415 89.325 94.695 90.205 ;
    RECT 91.095 89.325 91.375 90.205 ;
    RECT 87.775 89.325 88.055 90.205 ;
    RECT 84.455 89.325 84.735 90.205 ;
    RECT 81.135 89.325 81.415 90.205 ;
    RECT 77.815 89.325 78.095 90.205 ;
    RECT 74.495 89.325 74.775 90.205 ;
    RECT 71.175 89.325 71.455 90.205 ;
    RECT 31.335 89.325 31.615 90.205 ;
    RECT 67.855 89.325 68.135 90.205 ;
    RECT 28.015 89.325 28.295 90.205 ;
    RECT 24.695 89.325 24.975 90.205 ;
    RECT 21.375 89.325 21.655 90.205 ;
    RECT 18.055 89.325 18.335 90.205 ;
    RECT 14.735 89.325 15.015 90.205 ;
    RECT 11.415 89.325 11.695 90.205 ;
    RECT 8.095 89.325 8.375 90.205 ;
    RECT 4.775 89.325 5.055 90.205 ;
    RECT 1.455 89.325 1.735 90.205 ;
    RECT 64.535 89.325 64.815 90.205 ;
    RECT 61.215 14.425 61.495 15.305 ;
    RECT 57.895 14.425 58.175 15.305 ;
    RECT 54.575 14.425 54.855 15.305 ;
    RECT 51.255 14.425 51.535 15.305 ;
    RECT 47.935 14.425 48.215 15.305 ;
    RECT 44.615 14.425 44.895 15.305 ;
    RECT 41.295 14.425 41.575 15.305 ;
    RECT 37.975 14.425 38.255 15.305 ;
    RECT 34.655 14.425 34.935 15.305 ;
    RECT 114.335 14.425 114.615 15.305 ;
    RECT 111.015 14.425 111.295 15.305 ;
    RECT 107.695 14.425 107.975 15.305 ;
    RECT 104.375 14.425 104.655 15.305 ;
    RECT 101.055 14.425 101.335 15.305 ;
    RECT 97.735 14.425 98.015 15.305 ;
    RECT 94.415 14.425 94.695 15.305 ;
    RECT 91.095 14.425 91.375 15.305 ;
    RECT 87.775 14.425 88.055 15.305 ;
    RECT 84.455 14.425 84.735 15.305 ;
    RECT 81.135 14.425 81.415 15.305 ;
    RECT 77.815 14.425 78.095 15.305 ;
    RECT 74.495 14.425 74.775 15.305 ;
    RECT 71.175 14.425 71.455 15.305 ;
    RECT 31.335 14.425 31.615 15.305 ;
    RECT 67.855 14.425 68.135 15.305 ;
    RECT 28.015 14.425 28.295 15.305 ;
    RECT 24.695 14.425 24.975 15.305 ;
    RECT 21.375 14.425 21.655 15.305 ;
    RECT 18.055 14.425 18.335 15.305 ;
    RECT 14.735 14.425 15.015 15.305 ;
    RECT 11.415 14.425 11.695 15.305 ;
    RECT 8.095 14.425 8.375 15.305 ;
    RECT 4.775 14.425 5.055 15.305 ;
    RECT 117.655 14.425 117.935 15.305 ;
    RECT 1.455 14.425 1.735 15.305 ;
    RECT 64.535 14.425 64.815 15.305 ;
    RECT 61.215 88.605 61.495 89.485 ;
    RECT 57.895 88.605 58.175 89.485 ;
    RECT 54.575 88.605 54.855 89.485 ;
    RECT 51.255 88.605 51.535 89.485 ;
    RECT 47.935 88.605 48.215 89.485 ;
    RECT 44.615 88.605 44.895 89.485 ;
    RECT 41.295 88.605 41.575 89.485 ;
    RECT 37.975 88.605 38.255 89.485 ;
    RECT 34.655 88.605 34.935 89.485 ;
    RECT 117.655 88.605 117.935 89.485 ;
    RECT 114.335 88.605 114.615 89.485 ;
    RECT 111.015 88.605 111.295 89.485 ;
    RECT 107.695 88.605 107.975 89.485 ;
    RECT 104.375 88.605 104.655 89.485 ;
    RECT 101.055 88.605 101.335 89.485 ;
    RECT 97.735 88.605 98.015 89.485 ;
    RECT 94.415 88.605 94.695 89.485 ;
    RECT 91.095 88.605 91.375 89.485 ;
    RECT 87.775 88.605 88.055 89.485 ;
    RECT 84.455 88.605 84.735 89.485 ;
    RECT 81.135 88.605 81.415 89.485 ;
    RECT 77.815 88.605 78.095 89.485 ;
    RECT 74.495 88.605 74.775 89.485 ;
    RECT 71.175 88.605 71.455 89.485 ;
    RECT 31.335 88.605 31.615 89.485 ;
    RECT 67.855 88.605 68.135 89.485 ;
    RECT 28.015 88.605 28.295 89.485 ;
    RECT 24.695 88.605 24.975 89.485 ;
    RECT 21.375 88.605 21.655 89.485 ;
    RECT 18.055 88.605 18.335 89.485 ;
    RECT 14.735 88.605 15.015 89.485 ;
    RECT 11.415 88.605 11.695 89.485 ;
    RECT 8.095 88.605 8.375 89.485 ;
    RECT 4.775 88.605 5.055 89.485 ;
    RECT 1.455 88.605 1.735 89.485 ;
    RECT 64.535 88.605 64.815 89.485 ;
    RECT 61.215 20.905 61.495 21.785 ;
    RECT 57.895 20.905 58.175 21.785 ;
    RECT 54.575 20.905 54.855 21.785 ;
    RECT 51.255 20.905 51.535 21.785 ;
    RECT 47.935 20.905 48.215 21.785 ;
    RECT 44.615 20.905 44.895 21.785 ;
    RECT 41.295 20.905 41.575 21.785 ;
    RECT 37.975 20.905 38.255 21.785 ;
    RECT 34.655 20.905 34.935 21.785 ;
    RECT 117.655 20.905 117.935 21.785 ;
    RECT 114.335 20.905 114.615 21.785 ;
    RECT 111.015 20.905 111.295 21.785 ;
    RECT 107.695 20.905 107.975 21.785 ;
    RECT 104.375 20.905 104.655 21.785 ;
    RECT 101.055 20.905 101.335 21.785 ;
    RECT 97.735 20.905 98.015 21.785 ;
    RECT 94.415 20.905 94.695 21.785 ;
    RECT 91.095 20.905 91.375 21.785 ;
    RECT 87.775 20.905 88.055 21.785 ;
    RECT 84.455 20.905 84.735 21.785 ;
    RECT 81.135 20.905 81.415 21.785 ;
    RECT 77.815 20.905 78.095 21.785 ;
    RECT 74.495 20.905 74.775 21.785 ;
    RECT 71.175 20.905 71.455 21.785 ;
    RECT 31.335 20.905 31.615 21.785 ;
    RECT 67.855 20.905 68.135 21.785 ;
    RECT 28.015 20.905 28.295 21.785 ;
    RECT 24.695 20.905 24.975 21.785 ;
    RECT 21.375 20.905 21.655 21.785 ;
    RECT 18.055 20.905 18.335 21.785 ;
    RECT 14.735 20.905 15.015 21.785 ;
    RECT 11.415 20.905 11.695 21.785 ;
    RECT 8.095 20.905 8.375 21.785 ;
    RECT 4.775 20.905 5.055 21.785 ;
    RECT 1.455 20.905 1.735 21.785 ;
    RECT 64.535 20.905 64.815 21.785 ;
    RECT 61.215 87.885 61.495 88.765 ;
    RECT 57.895 87.885 58.175 88.765 ;
    RECT 54.575 87.885 54.855 88.765 ;
    RECT 51.255 87.885 51.535 88.765 ;
    RECT 47.935 87.885 48.215 88.765 ;
    RECT 44.615 87.885 44.895 88.765 ;
    RECT 41.295 87.885 41.575 88.765 ;
    RECT 37.975 87.885 38.255 88.765 ;
    RECT 34.655 87.885 34.935 88.765 ;
    RECT 117.655 87.885 117.935 88.765 ;
    RECT 114.335 87.885 114.615 88.765 ;
    RECT 111.015 87.885 111.295 88.765 ;
    RECT 107.695 87.885 107.975 88.765 ;
    RECT 104.375 87.885 104.655 88.765 ;
    RECT 101.055 87.885 101.335 88.765 ;
    RECT 97.735 87.885 98.015 88.765 ;
    RECT 94.415 87.885 94.695 88.765 ;
    RECT 91.095 87.885 91.375 88.765 ;
    RECT 87.775 87.885 88.055 88.765 ;
    RECT 84.455 87.885 84.735 88.765 ;
    RECT 81.135 87.885 81.415 88.765 ;
    RECT 77.815 87.885 78.095 88.765 ;
    RECT 74.495 87.885 74.775 88.765 ;
    RECT 71.175 87.885 71.455 88.765 ;
    RECT 31.335 87.885 31.615 88.765 ;
    RECT 67.855 87.885 68.135 88.765 ;
    RECT 28.015 87.885 28.295 88.765 ;
    RECT 24.695 87.885 24.975 88.765 ;
    RECT 21.375 87.885 21.655 88.765 ;
    RECT 18.055 87.885 18.335 88.765 ;
    RECT 14.735 87.885 15.015 88.765 ;
    RECT 11.415 87.885 11.695 88.765 ;
    RECT 8.095 87.885 8.375 88.765 ;
    RECT 4.775 87.885 5.055 88.765 ;
    RECT 1.455 87.885 1.735 88.765 ;
    RECT 64.535 87.885 64.815 88.765 ;
    RECT 61.215 20.185 61.495 21.065 ;
    RECT 57.895 20.185 58.175 21.065 ;
    RECT 54.575 20.185 54.855 21.065 ;
    RECT 51.255 20.185 51.535 21.065 ;
    RECT 47.935 20.185 48.215 21.065 ;
    RECT 44.615 20.185 44.895 21.065 ;
    RECT 41.295 20.185 41.575 21.065 ;
    RECT 37.975 20.185 38.255 21.065 ;
    RECT 34.655 20.185 34.935 21.065 ;
    RECT 117.655 20.185 117.935 21.065 ;
    RECT 114.335 20.185 114.615 21.065 ;
    RECT 111.015 20.185 111.295 21.065 ;
    RECT 107.695 20.185 107.975 21.065 ;
    RECT 104.375 20.185 104.655 21.065 ;
    RECT 101.055 20.185 101.335 21.065 ;
    RECT 97.735 20.185 98.015 21.065 ;
    RECT 94.415 20.185 94.695 21.065 ;
    RECT 91.095 20.185 91.375 21.065 ;
    RECT 87.775 20.185 88.055 21.065 ;
    RECT 84.455 20.185 84.735 21.065 ;
    RECT 81.135 20.185 81.415 21.065 ;
    RECT 77.815 20.185 78.095 21.065 ;
    RECT 74.495 20.185 74.775 21.065 ;
    RECT 71.175 20.185 71.455 21.065 ;
    RECT 31.335 20.185 31.615 21.065 ;
    RECT 67.855 20.185 68.135 21.065 ;
    RECT 28.015 20.185 28.295 21.065 ;
    RECT 24.695 20.185 24.975 21.065 ;
    RECT 21.375 20.185 21.655 21.065 ;
    RECT 18.055 20.185 18.335 21.065 ;
    RECT 14.735 20.185 15.015 21.065 ;
    RECT 11.415 20.185 11.695 21.065 ;
    RECT 8.095 20.185 8.375 21.065 ;
    RECT 4.775 20.185 5.055 21.065 ;
    RECT 1.455 20.185 1.735 21.065 ;
    RECT 64.535 20.185 64.815 21.065 ;
    RECT 61.215 87.165 61.495 88.045 ;
    RECT 57.895 87.165 58.175 88.045 ;
    RECT 54.575 87.165 54.855 88.045 ;
    RECT 51.255 87.165 51.535 88.045 ;
    RECT 47.935 87.165 48.215 88.045 ;
    RECT 44.615 87.165 44.895 88.045 ;
    RECT 41.295 87.165 41.575 88.045 ;
    RECT 37.975 87.165 38.255 88.045 ;
    RECT 34.655 87.165 34.935 88.045 ;
    RECT 117.655 87.165 117.935 88.045 ;
    RECT 114.335 87.165 114.615 88.045 ;
    RECT 111.015 87.165 111.295 88.045 ;
    RECT 107.695 87.165 107.975 88.045 ;
    RECT 104.375 87.165 104.655 88.045 ;
    RECT 101.055 87.165 101.335 88.045 ;
    RECT 97.735 87.165 98.015 88.045 ;
    RECT 94.415 87.165 94.695 88.045 ;
    RECT 91.095 87.165 91.375 88.045 ;
    RECT 87.775 87.165 88.055 88.045 ;
    RECT 84.455 87.165 84.735 88.045 ;
    RECT 81.135 87.165 81.415 88.045 ;
    RECT 77.815 87.165 78.095 88.045 ;
    RECT 74.495 87.165 74.775 88.045 ;
    RECT 71.175 87.165 71.455 88.045 ;
    RECT 31.335 87.165 31.615 88.045 ;
    RECT 67.855 87.165 68.135 88.045 ;
    RECT 28.015 87.165 28.295 88.045 ;
    RECT 24.695 87.165 24.975 88.045 ;
    RECT 21.375 87.165 21.655 88.045 ;
    RECT 18.055 87.165 18.335 88.045 ;
    RECT 14.735 87.165 15.015 88.045 ;
    RECT 11.415 87.165 11.695 88.045 ;
    RECT 8.095 87.165 8.375 88.045 ;
    RECT 4.775 87.165 5.055 88.045 ;
    RECT 1.455 87.165 1.735 88.045 ;
    RECT 64.535 87.165 64.815 88.045 ;
    RECT 61.215 19.465 61.495 20.345 ;
    RECT 57.895 19.465 58.175 20.345 ;
    RECT 54.575 19.465 54.855 20.345 ;
    RECT 51.255 19.465 51.535 20.345 ;
    RECT 47.935 19.465 48.215 20.345 ;
    RECT 44.615 19.465 44.895 20.345 ;
    RECT 41.295 19.465 41.575 20.345 ;
    RECT 37.975 19.465 38.255 20.345 ;
    RECT 34.655 19.465 34.935 20.345 ;
    RECT 117.655 19.465 117.935 20.345 ;
    RECT 114.335 19.465 114.615 20.345 ;
    RECT 111.015 19.465 111.295 20.345 ;
    RECT 107.695 19.465 107.975 20.345 ;
    RECT 104.375 19.465 104.655 20.345 ;
    RECT 101.055 19.465 101.335 20.345 ;
    RECT 97.735 19.465 98.015 20.345 ;
    RECT 94.415 19.465 94.695 20.345 ;
    RECT 91.095 19.465 91.375 20.345 ;
    RECT 87.775 19.465 88.055 20.345 ;
    RECT 84.455 19.465 84.735 20.345 ;
    RECT 81.135 19.465 81.415 20.345 ;
    RECT 77.815 19.465 78.095 20.345 ;
    RECT 74.495 19.465 74.775 20.345 ;
    RECT 71.175 19.465 71.455 20.345 ;
    RECT 31.335 19.465 31.615 20.345 ;
    RECT 67.855 19.465 68.135 20.345 ;
    RECT 28.015 19.465 28.295 20.345 ;
    RECT 24.695 19.465 24.975 20.345 ;
    RECT 21.375 19.465 21.655 20.345 ;
    RECT 18.055 19.465 18.335 20.345 ;
    RECT 14.735 19.465 15.015 20.345 ;
    RECT 11.415 19.465 11.695 20.345 ;
    RECT 8.095 19.465 8.375 20.345 ;
    RECT 4.775 19.465 5.055 20.345 ;
    RECT 1.455 19.465 1.735 20.345 ;
    RECT 64.535 19.465 64.815 20.345 ;
    RECT 61.215 18.745 61.495 19.625 ;
    RECT 57.895 18.745 58.175 19.625 ;
    RECT 54.575 18.745 54.855 19.625 ;
    RECT 51.255 18.745 51.535 19.625 ;
    RECT 47.935 18.745 48.215 19.625 ;
    RECT 44.615 18.745 44.895 19.625 ;
    RECT 41.295 18.745 41.575 19.625 ;
    RECT 37.975 18.745 38.255 19.625 ;
    RECT 34.655 18.745 34.935 19.625 ;
    RECT 117.655 18.745 117.935 19.625 ;
    RECT 114.335 18.745 114.615 19.625 ;
    RECT 111.015 18.745 111.295 19.625 ;
    RECT 107.695 18.745 107.975 19.625 ;
    RECT 104.375 18.745 104.655 19.625 ;
    RECT 101.055 18.745 101.335 19.625 ;
    RECT 97.735 18.745 98.015 19.625 ;
    RECT 94.415 18.745 94.695 19.625 ;
    RECT 91.095 18.745 91.375 19.625 ;
    RECT 87.775 18.745 88.055 19.625 ;
    RECT 84.455 18.745 84.735 19.625 ;
    RECT 81.135 18.745 81.415 19.625 ;
    RECT 77.815 18.745 78.095 19.625 ;
    RECT 74.495 18.745 74.775 19.625 ;
    RECT 71.175 18.745 71.455 19.625 ;
    RECT 31.335 18.745 31.615 19.625 ;
    RECT 67.855 18.745 68.135 19.625 ;
    RECT 28.015 18.745 28.295 19.625 ;
    RECT 24.695 18.745 24.975 19.625 ;
    RECT 21.375 18.745 21.655 19.625 ;
    RECT 18.055 18.745 18.335 19.625 ;
    RECT 14.735 18.745 15.015 19.625 ;
    RECT 11.415 18.745 11.695 19.625 ;
    RECT 8.095 18.745 8.375 19.625 ;
    RECT 4.775 18.745 5.055 19.625 ;
    RECT 1.455 18.745 1.735 19.625 ;
    RECT 64.535 18.745 64.815 19.625 ;
    RECT 61.215 49.705 61.495 50.585 ;
    RECT 57.895 49.705 58.175 50.585 ;
    RECT 54.575 49.705 54.855 50.585 ;
    RECT 51.255 49.705 51.535 50.585 ;
    RECT 47.935 49.705 48.215 50.585 ;
    RECT 44.615 49.705 44.895 50.585 ;
    RECT 41.295 49.705 41.575 50.585 ;
    RECT 37.975 49.705 38.255 50.585 ;
    RECT 34.655 49.705 34.935 50.585 ;
    RECT 117.655 49.705 117.935 50.585 ;
    RECT 114.335 49.705 114.615 50.585 ;
    RECT 111.015 49.705 111.295 50.585 ;
    RECT 107.695 49.705 107.975 50.585 ;
    RECT 104.375 49.705 104.655 50.585 ;
    RECT 101.055 49.705 101.335 50.585 ;
    RECT 97.735 49.705 98.015 50.585 ;
    RECT 94.415 49.705 94.695 50.585 ;
    RECT 91.095 49.705 91.375 50.585 ;
    RECT 87.775 49.705 88.055 50.585 ;
    RECT 84.455 49.705 84.735 50.585 ;
    RECT 81.135 49.705 81.415 50.585 ;
    RECT 77.815 49.705 78.095 50.585 ;
    RECT 74.495 49.705 74.775 50.585 ;
    RECT 71.175 49.705 71.455 50.585 ;
    RECT 31.335 49.705 31.615 50.585 ;
    RECT 67.855 49.705 68.135 50.585 ;
    RECT 28.015 49.705 28.295 50.585 ;
    RECT 24.695 49.705 24.975 50.585 ;
    RECT 21.375 49.705 21.655 50.585 ;
    RECT 18.055 49.705 18.335 50.585 ;
    RECT 14.735 49.705 15.015 50.585 ;
    RECT 11.415 49.705 11.695 50.585 ;
    RECT 8.095 49.705 8.375 50.585 ;
    RECT 4.775 49.705 5.055 50.585 ;
    RECT 1.455 49.705 1.735 50.585 ;
    RECT 64.535 49.705 64.815 50.585 ;
    RECT 61.215 18.025 61.495 18.905 ;
    RECT 57.895 18.025 58.175 18.905 ;
    RECT 54.575 18.025 54.855 18.905 ;
    RECT 51.255 18.025 51.535 18.905 ;
    RECT 47.935 18.025 48.215 18.905 ;
    RECT 44.615 18.025 44.895 18.905 ;
    RECT 41.295 18.025 41.575 18.905 ;
    RECT 37.975 18.025 38.255 18.905 ;
    RECT 34.655 18.025 34.935 18.905 ;
    RECT 117.655 18.025 117.935 18.905 ;
    RECT 114.335 18.025 114.615 18.905 ;
    RECT 111.015 18.025 111.295 18.905 ;
    RECT 107.695 18.025 107.975 18.905 ;
    RECT 104.375 18.025 104.655 18.905 ;
    RECT 101.055 18.025 101.335 18.905 ;
    RECT 97.735 18.025 98.015 18.905 ;
    RECT 94.415 18.025 94.695 18.905 ;
    RECT 91.095 18.025 91.375 18.905 ;
    RECT 87.775 18.025 88.055 18.905 ;
    RECT 84.455 18.025 84.735 18.905 ;
    RECT 81.135 18.025 81.415 18.905 ;
    RECT 77.815 18.025 78.095 18.905 ;
    RECT 74.495 18.025 74.775 18.905 ;
    RECT 71.175 18.025 71.455 18.905 ;
    RECT 31.335 18.025 31.615 18.905 ;
    RECT 67.855 18.025 68.135 18.905 ;
    RECT 28.015 18.025 28.295 18.905 ;
    RECT 24.695 18.025 24.975 18.905 ;
    RECT 21.375 18.025 21.655 18.905 ;
    RECT 18.055 18.025 18.335 18.905 ;
    RECT 14.735 18.025 15.015 18.905 ;
    RECT 11.415 18.025 11.695 18.905 ;
    RECT 8.095 18.025 8.375 18.905 ;
    RECT 4.775 18.025 5.055 18.905 ;
    RECT 1.455 18.025 1.735 18.905 ;
    RECT 64.535 18.025 64.815 18.905 ;
    RECT 61.215 48.985 61.495 49.865 ;
    RECT 57.895 48.985 58.175 49.865 ;
    RECT 54.575 48.985 54.855 49.865 ;
    RECT 51.255 48.985 51.535 49.865 ;
    RECT 47.935 48.985 48.215 49.865 ;
    RECT 44.615 48.985 44.895 49.865 ;
    RECT 41.295 48.985 41.575 49.865 ;
    RECT 37.975 48.985 38.255 49.865 ;
    RECT 34.655 48.985 34.935 49.865 ;
    RECT 117.655 48.985 117.935 49.865 ;
    RECT 114.335 48.985 114.615 49.865 ;
    RECT 111.015 48.985 111.295 49.865 ;
    RECT 107.695 48.985 107.975 49.865 ;
    RECT 104.375 48.985 104.655 49.865 ;
    RECT 101.055 48.985 101.335 49.865 ;
    RECT 97.735 48.985 98.015 49.865 ;
    RECT 94.415 48.985 94.695 49.865 ;
    RECT 91.095 48.985 91.375 49.865 ;
    RECT 87.775 48.985 88.055 49.865 ;
    RECT 84.455 48.985 84.735 49.865 ;
    RECT 81.135 48.985 81.415 49.865 ;
    RECT 77.815 48.985 78.095 49.865 ;
    RECT 74.495 48.985 74.775 49.865 ;
    RECT 71.175 48.985 71.455 49.865 ;
    RECT 31.335 48.985 31.615 49.865 ;
    RECT 67.855 48.985 68.135 49.865 ;
    RECT 28.015 48.985 28.295 49.865 ;
    RECT 24.695 48.985 24.975 49.865 ;
    RECT 21.375 48.985 21.655 49.865 ;
    RECT 18.055 48.985 18.335 49.865 ;
    RECT 14.735 48.985 15.015 49.865 ;
    RECT 11.415 48.985 11.695 49.865 ;
    RECT 8.095 48.985 8.375 49.865 ;
    RECT 4.775 48.985 5.055 49.865 ;
    RECT 1.455 48.985 1.735 49.865 ;
    RECT 64.535 48.985 64.815 49.865 ;
    RECT 61.215 17.305 61.495 18.185 ;
    RECT 57.895 17.305 58.175 18.185 ;
    RECT 54.575 17.305 54.855 18.185 ;
    RECT 51.255 17.305 51.535 18.185 ;
    RECT 47.935 17.305 48.215 18.185 ;
    RECT 44.615 17.305 44.895 18.185 ;
    RECT 41.295 17.305 41.575 18.185 ;
    RECT 37.975 17.305 38.255 18.185 ;
    RECT 34.655 17.305 34.935 18.185 ;
    RECT 117.655 17.305 117.935 18.185 ;
    RECT 114.335 17.305 114.615 18.185 ;
    RECT 111.015 17.305 111.295 18.185 ;
    RECT 107.695 17.305 107.975 18.185 ;
    RECT 104.375 17.305 104.655 18.185 ;
    RECT 101.055 17.305 101.335 18.185 ;
    RECT 97.735 17.305 98.015 18.185 ;
    RECT 94.415 17.305 94.695 18.185 ;
    RECT 91.095 17.305 91.375 18.185 ;
    RECT 87.775 17.305 88.055 18.185 ;
    RECT 84.455 17.305 84.735 18.185 ;
    RECT 81.135 17.305 81.415 18.185 ;
    RECT 77.815 17.305 78.095 18.185 ;
    RECT 74.495 17.305 74.775 18.185 ;
    RECT 71.175 17.305 71.455 18.185 ;
    RECT 31.335 17.305 31.615 18.185 ;
    RECT 67.855 17.305 68.135 18.185 ;
    RECT 28.015 17.305 28.295 18.185 ;
    RECT 24.695 17.305 24.975 18.185 ;
    RECT 21.375 17.305 21.655 18.185 ;
    RECT 18.055 17.305 18.335 18.185 ;
    RECT 14.735 17.305 15.015 18.185 ;
    RECT 11.415 17.305 11.695 18.185 ;
    RECT 8.095 17.305 8.375 18.185 ;
    RECT 4.775 17.305 5.055 18.185 ;
    RECT 1.455 17.305 1.735 18.185 ;
    RECT 64.535 17.305 64.815 18.185 ;
    RECT 61.215 48.265 61.495 49.145 ;
    RECT 57.895 48.265 58.175 49.145 ;
    RECT 54.575 48.265 54.855 49.145 ;
    RECT 51.255 48.265 51.535 49.145 ;
    RECT 47.935 48.265 48.215 49.145 ;
    RECT 44.615 48.265 44.895 49.145 ;
    RECT 41.295 48.265 41.575 49.145 ;
    RECT 37.975 48.265 38.255 49.145 ;
    RECT 34.655 48.265 34.935 49.145 ;
    RECT 117.655 48.265 117.935 49.145 ;
    RECT 114.335 48.265 114.615 49.145 ;
    RECT 111.015 48.265 111.295 49.145 ;
    RECT 107.695 48.265 107.975 49.145 ;
    RECT 104.375 48.265 104.655 49.145 ;
    RECT 101.055 48.265 101.335 49.145 ;
    RECT 97.735 48.265 98.015 49.145 ;
    RECT 94.415 48.265 94.695 49.145 ;
    RECT 91.095 48.265 91.375 49.145 ;
    RECT 87.775 48.265 88.055 49.145 ;
    RECT 84.455 48.265 84.735 49.145 ;
    RECT 81.135 48.265 81.415 49.145 ;
    RECT 77.815 48.265 78.095 49.145 ;
    RECT 74.495 48.265 74.775 49.145 ;
    RECT 71.175 48.265 71.455 49.145 ;
    RECT 31.335 48.265 31.615 49.145 ;
    RECT 67.855 48.265 68.135 49.145 ;
    RECT 28.015 48.265 28.295 49.145 ;
    RECT 24.695 48.265 24.975 49.145 ;
    RECT 21.375 48.265 21.655 49.145 ;
    RECT 18.055 48.265 18.335 49.145 ;
    RECT 14.735 48.265 15.015 49.145 ;
    RECT 11.415 48.265 11.695 49.145 ;
    RECT 8.095 48.265 8.375 49.145 ;
    RECT 4.775 48.265 5.055 49.145 ;
    RECT 1.455 48.265 1.735 49.145 ;
    RECT 64.535 48.265 64.815 49.145 ;
    RECT 61.215 16.585 61.495 17.465 ;
    RECT 57.895 16.585 58.175 17.465 ;
    RECT 54.575 16.585 54.855 17.465 ;
    RECT 51.255 16.585 51.535 17.465 ;
    RECT 47.935 16.585 48.215 17.465 ;
    RECT 44.615 16.585 44.895 17.465 ;
    RECT 41.295 16.585 41.575 17.465 ;
    RECT 37.975 16.585 38.255 17.465 ;
    RECT 34.655 16.585 34.935 17.465 ;
    RECT 117.655 16.585 117.935 17.465 ;
    RECT 114.335 16.585 114.615 17.465 ;
    RECT 111.015 16.585 111.295 17.465 ;
    RECT 107.695 16.585 107.975 17.465 ;
    RECT 104.375 16.585 104.655 17.465 ;
    RECT 101.055 16.585 101.335 17.465 ;
    RECT 97.735 16.585 98.015 17.465 ;
    RECT 94.415 16.585 94.695 17.465 ;
    RECT 91.095 16.585 91.375 17.465 ;
    RECT 87.775 16.585 88.055 17.465 ;
    RECT 84.455 16.585 84.735 17.465 ;
    RECT 81.135 16.585 81.415 17.465 ;
    RECT 77.815 16.585 78.095 17.465 ;
    RECT 74.495 16.585 74.775 17.465 ;
    RECT 71.175 16.585 71.455 17.465 ;
    RECT 31.335 16.585 31.615 17.465 ;
    RECT 67.855 16.585 68.135 17.465 ;
    RECT 28.015 16.585 28.295 17.465 ;
    RECT 24.695 16.585 24.975 17.465 ;
    RECT 21.375 16.585 21.655 17.465 ;
    RECT 18.055 16.585 18.335 17.465 ;
    RECT 14.735 16.585 15.015 17.465 ;
    RECT 11.415 16.585 11.695 17.465 ;
    RECT 8.095 16.585 8.375 17.465 ;
    RECT 4.775 16.585 5.055 17.465 ;
    RECT 1.455 16.585 1.735 17.465 ;
    RECT 64.535 16.585 64.815 17.465 ;
    RECT 61.215 47.545 61.495 48.425 ;
    RECT 57.895 47.545 58.175 48.425 ;
    RECT 54.575 47.545 54.855 48.425 ;
    RECT 51.255 47.545 51.535 48.425 ;
    RECT 47.935 47.545 48.215 48.425 ;
    RECT 44.615 47.545 44.895 48.425 ;
    RECT 41.295 47.545 41.575 48.425 ;
    RECT 37.975 47.545 38.255 48.425 ;
    RECT 34.655 47.545 34.935 48.425 ;
    RECT 117.655 47.545 117.935 48.425 ;
    RECT 114.335 47.545 114.615 48.425 ;
    RECT 111.015 47.545 111.295 48.425 ;
    RECT 107.695 47.545 107.975 48.425 ;
    RECT 104.375 47.545 104.655 48.425 ;
    RECT 101.055 47.545 101.335 48.425 ;
    RECT 97.735 47.545 98.015 48.425 ;
    RECT 94.415 47.545 94.695 48.425 ;
    RECT 91.095 47.545 91.375 48.425 ;
    RECT 87.775 47.545 88.055 48.425 ;
    RECT 84.455 47.545 84.735 48.425 ;
    RECT 81.135 47.545 81.415 48.425 ;
    RECT 77.815 47.545 78.095 48.425 ;
    RECT 74.495 47.545 74.775 48.425 ;
    RECT 71.175 47.545 71.455 48.425 ;
    RECT 31.335 47.545 31.615 48.425 ;
    RECT 67.855 47.545 68.135 48.425 ;
    RECT 28.015 47.545 28.295 48.425 ;
    RECT 24.695 47.545 24.975 48.425 ;
    RECT 21.375 47.545 21.655 48.425 ;
    RECT 18.055 47.545 18.335 48.425 ;
    RECT 14.735 47.545 15.015 48.425 ;
    RECT 11.415 47.545 11.695 48.425 ;
    RECT 8.095 47.545 8.375 48.425 ;
    RECT 4.775 47.545 5.055 48.425 ;
    RECT 1.455 47.545 1.735 48.425 ;
    RECT 64.535 47.545 64.815 48.425 ;
    RECT 61.215 15.865 61.495 16.745 ;
    RECT 57.895 15.865 58.175 16.745 ;
    RECT 54.575 15.865 54.855 16.745 ;
    RECT 51.255 15.865 51.535 16.745 ;
    RECT 47.935 15.865 48.215 16.745 ;
    RECT 44.615 15.865 44.895 16.745 ;
    RECT 41.295 15.865 41.575 16.745 ;
    RECT 37.975 15.865 38.255 16.745 ;
    RECT 34.655 15.865 34.935 16.745 ;
    RECT 117.655 15.865 117.935 16.745 ;
    RECT 114.335 15.865 114.615 16.745 ;
    RECT 111.015 15.865 111.295 16.745 ;
    RECT 107.695 15.865 107.975 16.745 ;
    RECT 104.375 15.865 104.655 16.745 ;
    RECT 101.055 15.865 101.335 16.745 ;
    RECT 97.735 15.865 98.015 16.745 ;
    RECT 94.415 15.865 94.695 16.745 ;
    RECT 91.095 15.865 91.375 16.745 ;
    RECT 87.775 15.865 88.055 16.745 ;
    RECT 84.455 15.865 84.735 16.745 ;
    RECT 81.135 15.865 81.415 16.745 ;
    RECT 77.815 15.865 78.095 16.745 ;
    RECT 74.495 15.865 74.775 16.745 ;
    RECT 71.175 15.865 71.455 16.745 ;
    RECT 31.335 15.865 31.615 16.745 ;
    RECT 67.855 15.865 68.135 16.745 ;
    RECT 28.015 15.865 28.295 16.745 ;
    RECT 24.695 15.865 24.975 16.745 ;
    RECT 21.375 15.865 21.655 16.745 ;
    RECT 18.055 15.865 18.335 16.745 ;
    RECT 14.735 15.865 15.015 16.745 ;
    RECT 11.415 15.865 11.695 16.745 ;
    RECT 8.095 15.865 8.375 16.745 ;
    RECT 4.775 15.865 5.055 16.745 ;
    RECT 1.455 15.865 1.735 16.745 ;
    RECT 64.535 15.865 64.815 16.745 ;
    RECT 61.215 46.825 61.495 47.705 ;
    RECT 57.895 46.825 58.175 47.705 ;
    RECT 54.575 46.825 54.855 47.705 ;
    RECT 51.255 46.825 51.535 47.705 ;
    RECT 47.935 46.825 48.215 47.705 ;
    RECT 44.615 46.825 44.895 47.705 ;
    RECT 41.295 46.825 41.575 47.705 ;
    RECT 37.975 46.825 38.255 47.705 ;
    RECT 34.655 46.825 34.935 47.705 ;
    RECT 117.655 46.825 117.935 47.705 ;
    RECT 114.335 46.825 114.615 47.705 ;
    RECT 111.015 46.825 111.295 47.705 ;
    RECT 107.695 46.825 107.975 47.705 ;
    RECT 104.375 46.825 104.655 47.705 ;
    RECT 101.055 46.825 101.335 47.705 ;
    RECT 97.735 46.825 98.015 47.705 ;
    RECT 94.415 46.825 94.695 47.705 ;
    RECT 91.095 46.825 91.375 47.705 ;
    RECT 87.775 46.825 88.055 47.705 ;
    RECT 84.455 46.825 84.735 47.705 ;
    RECT 81.135 46.825 81.415 47.705 ;
    RECT 77.815 46.825 78.095 47.705 ;
    RECT 74.495 46.825 74.775 47.705 ;
    RECT 71.175 46.825 71.455 47.705 ;
    RECT 31.335 46.825 31.615 47.705 ;
    RECT 67.855 46.825 68.135 47.705 ;
    RECT 28.015 46.825 28.295 47.705 ;
    RECT 24.695 46.825 24.975 47.705 ;
    RECT 21.375 46.825 21.655 47.705 ;
    RECT 18.055 46.825 18.335 47.705 ;
    RECT 14.735 46.825 15.015 47.705 ;
    RECT 11.415 46.825 11.695 47.705 ;
    RECT 8.095 46.825 8.375 47.705 ;
    RECT 4.775 46.825 5.055 47.705 ;
    RECT 1.455 46.825 1.735 47.705 ;
    RECT 64.535 46.825 64.815 47.705 ;
    RECT 61.215 86.445 61.495 87.325 ;
    RECT 57.895 86.445 58.175 87.325 ;
    RECT 54.575 86.445 54.855 87.325 ;
    RECT 51.255 86.445 51.535 87.325 ;
    RECT 47.935 86.445 48.215 87.325 ;
    RECT 44.615 86.445 44.895 87.325 ;
    RECT 41.295 86.445 41.575 87.325 ;
    RECT 37.975 86.445 38.255 87.325 ;
    RECT 34.655 86.445 34.935 87.325 ;
    RECT 117.655 86.445 117.935 87.325 ;
    RECT 114.335 86.445 114.615 87.325 ;
    RECT 111.015 86.445 111.295 87.325 ;
    RECT 107.695 86.445 107.975 87.325 ;
    RECT 104.375 86.445 104.655 87.325 ;
    RECT 101.055 86.445 101.335 87.325 ;
    RECT 97.735 86.445 98.015 87.325 ;
    RECT 94.415 86.445 94.695 87.325 ;
    RECT 91.095 86.445 91.375 87.325 ;
    RECT 87.775 86.445 88.055 87.325 ;
    RECT 84.455 86.445 84.735 87.325 ;
    RECT 81.135 86.445 81.415 87.325 ;
    RECT 77.815 86.445 78.095 87.325 ;
    RECT 74.495 86.445 74.775 87.325 ;
    RECT 71.175 86.445 71.455 87.325 ;
    RECT 31.335 86.445 31.615 87.325 ;
    RECT 67.855 86.445 68.135 87.325 ;
    RECT 28.015 86.445 28.295 87.325 ;
    RECT 24.695 86.445 24.975 87.325 ;
    RECT 21.375 86.445 21.655 87.325 ;
    RECT 18.055 86.445 18.335 87.325 ;
    RECT 14.735 86.445 15.015 87.325 ;
    RECT 11.415 86.445 11.695 87.325 ;
    RECT 8.095 86.445 8.375 87.325 ;
    RECT 4.775 86.445 5.055 87.325 ;
    RECT 1.455 86.445 1.735 87.325 ;
    RECT 64.535 86.445 64.815 87.325 ;
    RECT 61.215 15.145 61.495 16.025 ;
    RECT 57.895 15.145 58.175 16.025 ;
    RECT 54.575 15.145 54.855 16.025 ;
    RECT 51.255 15.145 51.535 16.025 ;
    RECT 47.935 15.145 48.215 16.025 ;
    RECT 44.615 15.145 44.895 16.025 ;
    RECT 41.295 15.145 41.575 16.025 ;
    RECT 37.975 15.145 38.255 16.025 ;
    RECT 34.655 15.145 34.935 16.025 ;
    RECT 117.655 15.145 117.935 16.025 ;
    RECT 114.335 15.145 114.615 16.025 ;
    RECT 111.015 15.145 111.295 16.025 ;
    RECT 107.695 15.145 107.975 16.025 ;
    RECT 104.375 15.145 104.655 16.025 ;
    RECT 101.055 15.145 101.335 16.025 ;
    RECT 97.735 15.145 98.015 16.025 ;
    RECT 94.415 15.145 94.695 16.025 ;
    RECT 91.095 15.145 91.375 16.025 ;
    RECT 87.775 15.145 88.055 16.025 ;
    RECT 84.455 15.145 84.735 16.025 ;
    RECT 81.135 15.145 81.415 16.025 ;
    RECT 77.815 15.145 78.095 16.025 ;
    RECT 74.495 15.145 74.775 16.025 ;
    RECT 71.175 15.145 71.455 16.025 ;
    RECT 31.335 15.145 31.615 16.025 ;
    RECT 67.855 15.145 68.135 16.025 ;
    RECT 28.015 15.145 28.295 16.025 ;
    RECT 24.695 15.145 24.975 16.025 ;
    RECT 21.375 15.145 21.655 16.025 ;
    RECT 18.055 15.145 18.335 16.025 ;
    RECT 14.735 15.145 15.015 16.025 ;
    RECT 11.415 15.145 11.695 16.025 ;
    RECT 8.095 15.145 8.375 16.025 ;
    RECT 4.775 15.145 5.055 16.025 ;
    RECT 1.455 15.145 1.735 16.025 ;
    RECT 64.535 15.145 64.815 16.025 ;
    RECT 61.215 46.105 61.495 46.985 ;
    RECT 57.895 46.105 58.175 46.985 ;
    RECT 54.575 46.105 54.855 46.985 ;
    RECT 51.255 46.105 51.535 46.985 ;
    RECT 47.935 46.105 48.215 46.985 ;
    RECT 44.615 46.105 44.895 46.985 ;
    RECT 41.295 46.105 41.575 46.985 ;
    RECT 37.975 46.105 38.255 46.985 ;
    RECT 34.655 46.105 34.935 46.985 ;
    RECT 117.655 46.105 117.935 46.985 ;
    RECT 114.335 46.105 114.615 46.985 ;
    RECT 111.015 46.105 111.295 46.985 ;
    RECT 107.695 46.105 107.975 46.985 ;
    RECT 104.375 46.105 104.655 46.985 ;
    RECT 101.055 46.105 101.335 46.985 ;
    RECT 97.735 46.105 98.015 46.985 ;
    RECT 94.415 46.105 94.695 46.985 ;
    RECT 91.095 46.105 91.375 46.985 ;
    RECT 87.775 46.105 88.055 46.985 ;
    RECT 84.455 46.105 84.735 46.985 ;
    RECT 81.135 46.105 81.415 46.985 ;
    RECT 77.815 46.105 78.095 46.985 ;
    RECT 74.495 46.105 74.775 46.985 ;
    RECT 71.175 46.105 71.455 46.985 ;
    RECT 31.335 46.105 31.615 46.985 ;
    RECT 67.855 46.105 68.135 46.985 ;
    RECT 28.015 46.105 28.295 46.985 ;
    RECT 24.695 46.105 24.975 46.985 ;
    RECT 21.375 46.105 21.655 46.985 ;
    RECT 18.055 46.105 18.335 46.985 ;
    RECT 14.735 46.105 15.015 46.985 ;
    RECT 11.415 46.105 11.695 46.985 ;
    RECT 8.095 46.105 8.375 46.985 ;
    RECT 4.775 46.105 5.055 46.985 ;
    RECT 1.455 46.105 1.735 46.985 ;
    RECT 64.535 46.105 64.815 46.985 ;
    RECT 61.215 85.725 61.495 86.605 ;
    RECT 57.895 85.725 58.175 86.605 ;
    RECT 54.575 85.725 54.855 86.605 ;
    RECT 51.255 85.725 51.535 86.605 ;
    RECT 47.935 85.725 48.215 86.605 ;
    RECT 44.615 85.725 44.895 86.605 ;
    RECT 41.295 85.725 41.575 86.605 ;
    RECT 37.975 85.725 38.255 86.605 ;
    RECT 34.655 85.725 34.935 86.605 ;
    RECT 117.655 85.725 117.935 86.605 ;
    RECT 114.335 85.725 114.615 86.605 ;
    RECT 111.015 85.725 111.295 86.605 ;
    RECT 107.695 85.725 107.975 86.605 ;
    RECT 104.375 85.725 104.655 86.605 ;
    RECT 101.055 85.725 101.335 86.605 ;
    RECT 97.735 85.725 98.015 86.605 ;
    RECT 94.415 85.725 94.695 86.605 ;
    RECT 91.095 85.725 91.375 86.605 ;
    RECT 87.775 85.725 88.055 86.605 ;
    RECT 84.455 85.725 84.735 86.605 ;
    RECT 81.135 85.725 81.415 86.605 ;
    RECT 77.815 85.725 78.095 86.605 ;
    RECT 74.495 85.725 74.775 86.605 ;
    RECT 71.175 85.725 71.455 86.605 ;
    RECT 31.335 85.725 31.615 86.605 ;
    RECT 67.855 85.725 68.135 86.605 ;
    RECT 28.015 85.725 28.295 86.605 ;
    RECT 24.695 85.725 24.975 86.605 ;
    RECT 21.375 85.725 21.655 86.605 ;
    RECT 18.055 85.725 18.335 86.605 ;
    RECT 14.735 85.725 15.015 86.605 ;
    RECT 11.415 85.725 11.695 86.605 ;
    RECT 8.095 85.725 8.375 86.605 ;
    RECT 4.775 85.725 5.055 86.605 ;
    RECT 1.455 85.725 1.735 86.605 ;
    RECT 64.535 85.725 64.815 86.605 ;
    RECT 61.215 45.385 61.495 46.265 ;
    RECT 57.895 45.385 58.175 46.265 ;
    RECT 54.575 45.385 54.855 46.265 ;
    RECT 51.255 45.385 51.535 46.265 ;
    RECT 47.935 45.385 48.215 46.265 ;
    RECT 44.615 45.385 44.895 46.265 ;
    RECT 41.295 45.385 41.575 46.265 ;
    RECT 37.975 45.385 38.255 46.265 ;
    RECT 34.655 45.385 34.935 46.265 ;
    RECT 117.655 45.385 117.935 46.265 ;
    RECT 114.335 45.385 114.615 46.265 ;
    RECT 111.015 45.385 111.295 46.265 ;
    RECT 107.695 45.385 107.975 46.265 ;
    RECT 104.375 45.385 104.655 46.265 ;
    RECT 101.055 45.385 101.335 46.265 ;
    RECT 97.735 45.385 98.015 46.265 ;
    RECT 94.415 45.385 94.695 46.265 ;
    RECT 91.095 45.385 91.375 46.265 ;
    RECT 87.775 45.385 88.055 46.265 ;
    RECT 84.455 45.385 84.735 46.265 ;
    RECT 81.135 45.385 81.415 46.265 ;
    RECT 77.815 45.385 78.095 46.265 ;
    RECT 74.495 45.385 74.775 46.265 ;
    RECT 71.175 45.385 71.455 46.265 ;
    RECT 31.335 45.385 31.615 46.265 ;
    RECT 67.855 45.385 68.135 46.265 ;
    RECT 28.015 45.385 28.295 46.265 ;
    RECT 24.695 45.385 24.975 46.265 ;
    RECT 21.375 45.385 21.655 46.265 ;
    RECT 18.055 45.385 18.335 46.265 ;
    RECT 14.735 45.385 15.015 46.265 ;
    RECT 11.415 45.385 11.695 46.265 ;
    RECT 8.095 45.385 8.375 46.265 ;
    RECT 4.775 45.385 5.055 46.265 ;
    RECT 1.455 45.385 1.735 46.265 ;
    RECT 64.535 45.385 64.815 46.265 ;
    RECT 61.215 85.005 61.495 85.885 ;
    RECT 57.895 85.005 58.175 85.885 ;
    RECT 54.575 85.005 54.855 85.885 ;
    RECT 51.255 85.005 51.535 85.885 ;
    RECT 47.935 85.005 48.215 85.885 ;
    RECT 44.615 85.005 44.895 85.885 ;
    RECT 41.295 85.005 41.575 85.885 ;
    RECT 37.975 85.005 38.255 85.885 ;
    RECT 34.655 85.005 34.935 85.885 ;
    RECT 117.655 85.005 117.935 85.885 ;
    RECT 114.335 85.005 114.615 85.885 ;
    RECT 111.015 85.005 111.295 85.885 ;
    RECT 107.695 85.005 107.975 85.885 ;
    RECT 104.375 85.005 104.655 85.885 ;
    RECT 101.055 85.005 101.335 85.885 ;
    RECT 97.735 85.005 98.015 85.885 ;
    RECT 94.415 85.005 94.695 85.885 ;
    RECT 91.095 85.005 91.375 85.885 ;
    RECT 87.775 85.005 88.055 85.885 ;
    RECT 84.455 85.005 84.735 85.885 ;
    RECT 81.135 85.005 81.415 85.885 ;
    RECT 77.815 85.005 78.095 85.885 ;
    RECT 74.495 85.005 74.775 85.885 ;
    RECT 71.175 85.005 71.455 85.885 ;
    RECT 31.335 85.005 31.615 85.885 ;
    RECT 67.855 85.005 68.135 85.885 ;
    RECT 28.015 85.005 28.295 85.885 ;
    RECT 24.695 85.005 24.975 85.885 ;
    RECT 21.375 85.005 21.655 85.885 ;
    RECT 18.055 85.005 18.335 85.885 ;
    RECT 14.735 85.005 15.015 85.885 ;
    RECT 11.415 85.005 11.695 85.885 ;
    RECT 8.095 85.005 8.375 85.885 ;
    RECT 4.775 85.005 5.055 85.885 ;
    RECT 1.455 85.005 1.735 85.885 ;
    RECT 64.535 85.005 64.815 85.885 ;
    RECT 61.215 44.665 61.495 45.545 ;
    RECT 57.895 44.665 58.175 45.545 ;
    RECT 54.575 44.665 54.855 45.545 ;
    RECT 51.255 44.665 51.535 45.545 ;
    RECT 47.935 44.665 48.215 45.545 ;
    RECT 44.615 44.665 44.895 45.545 ;
    RECT 41.295 44.665 41.575 45.545 ;
    RECT 37.975 44.665 38.255 45.545 ;
    RECT 34.655 44.665 34.935 45.545 ;
    RECT 117.655 44.665 117.935 45.545 ;
    RECT 114.335 44.665 114.615 45.545 ;
    RECT 111.015 44.665 111.295 45.545 ;
    RECT 107.695 44.665 107.975 45.545 ;
    RECT 104.375 44.665 104.655 45.545 ;
    RECT 101.055 44.665 101.335 45.545 ;
    RECT 97.735 44.665 98.015 45.545 ;
    RECT 94.415 44.665 94.695 45.545 ;
    RECT 91.095 44.665 91.375 45.545 ;
    RECT 87.775 44.665 88.055 45.545 ;
    RECT 84.455 44.665 84.735 45.545 ;
    RECT 81.135 44.665 81.415 45.545 ;
    RECT 77.815 44.665 78.095 45.545 ;
    RECT 74.495 44.665 74.775 45.545 ;
    RECT 71.175 44.665 71.455 45.545 ;
    RECT 31.335 44.665 31.615 45.545 ;
    RECT 67.855 44.665 68.135 45.545 ;
    RECT 28.015 44.665 28.295 45.545 ;
    RECT 24.695 44.665 24.975 45.545 ;
    RECT 21.375 44.665 21.655 45.545 ;
    RECT 18.055 44.665 18.335 45.545 ;
    RECT 14.735 44.665 15.015 45.545 ;
    RECT 11.415 44.665 11.695 45.545 ;
    RECT 8.095 44.665 8.375 45.545 ;
    RECT 4.775 44.665 5.055 45.545 ;
    RECT 1.455 44.665 1.735 45.545 ;
    RECT 64.535 44.665 64.815 45.545 ;
    RECT 61.215 84.285 61.495 85.165 ;
    RECT 57.895 84.285 58.175 85.165 ;
    RECT 54.575 84.285 54.855 85.165 ;
    RECT 51.255 84.285 51.535 85.165 ;
    RECT 47.935 84.285 48.215 85.165 ;
    RECT 44.615 84.285 44.895 85.165 ;
    RECT 41.295 84.285 41.575 85.165 ;
    RECT 37.975 84.285 38.255 85.165 ;
    RECT 34.655 84.285 34.935 85.165 ;
    RECT 117.655 84.285 117.935 85.165 ;
    RECT 114.335 84.285 114.615 85.165 ;
    RECT 111.015 84.285 111.295 85.165 ;
    RECT 107.695 84.285 107.975 85.165 ;
    RECT 104.375 84.285 104.655 85.165 ;
    RECT 101.055 84.285 101.335 85.165 ;
    RECT 97.735 84.285 98.015 85.165 ;
    RECT 94.415 84.285 94.695 85.165 ;
    RECT 91.095 84.285 91.375 85.165 ;
    RECT 87.775 84.285 88.055 85.165 ;
    RECT 84.455 84.285 84.735 85.165 ;
    RECT 81.135 84.285 81.415 85.165 ;
    RECT 77.815 84.285 78.095 85.165 ;
    RECT 74.495 84.285 74.775 85.165 ;
    RECT 71.175 84.285 71.455 85.165 ;
    RECT 31.335 84.285 31.615 85.165 ;
    RECT 67.855 84.285 68.135 85.165 ;
    RECT 28.015 84.285 28.295 85.165 ;
    RECT 24.695 84.285 24.975 85.165 ;
    RECT 21.375 84.285 21.655 85.165 ;
    RECT 18.055 84.285 18.335 85.165 ;
    RECT 14.735 84.285 15.015 85.165 ;
    RECT 11.415 84.285 11.695 85.165 ;
    RECT 8.095 84.285 8.375 85.165 ;
    RECT 4.775 84.285 5.055 85.165 ;
    RECT 1.455 84.285 1.735 85.165 ;
    RECT 64.535 84.285 64.815 85.165 ;
    RECT 61.215 43.945 61.495 44.825 ;
    RECT 57.895 43.945 58.175 44.825 ;
    RECT 54.575 43.945 54.855 44.825 ;
    RECT 51.255 43.945 51.535 44.825 ;
    RECT 47.935 43.945 48.215 44.825 ;
    RECT 44.615 43.945 44.895 44.825 ;
    RECT 41.295 43.945 41.575 44.825 ;
    RECT 37.975 43.945 38.255 44.825 ;
    RECT 34.655 43.945 34.935 44.825 ;
    RECT 117.655 43.945 117.935 44.825 ;
    RECT 114.335 43.945 114.615 44.825 ;
    RECT 111.015 43.945 111.295 44.825 ;
    RECT 107.695 43.945 107.975 44.825 ;
    RECT 104.375 43.945 104.655 44.825 ;
    RECT 101.055 43.945 101.335 44.825 ;
    RECT 97.735 43.945 98.015 44.825 ;
    RECT 94.415 43.945 94.695 44.825 ;
    RECT 91.095 43.945 91.375 44.825 ;
    RECT 87.775 43.945 88.055 44.825 ;
    RECT 84.455 43.945 84.735 44.825 ;
    RECT 81.135 43.945 81.415 44.825 ;
    RECT 77.815 43.945 78.095 44.825 ;
    RECT 74.495 43.945 74.775 44.825 ;
    RECT 71.175 43.945 71.455 44.825 ;
    RECT 31.335 43.945 31.615 44.825 ;
    RECT 67.855 43.945 68.135 44.825 ;
    RECT 28.015 43.945 28.295 44.825 ;
    RECT 24.695 43.945 24.975 44.825 ;
    RECT 21.375 43.945 21.655 44.825 ;
    RECT 18.055 43.945 18.335 44.825 ;
    RECT 14.735 43.945 15.015 44.825 ;
    RECT 11.415 43.945 11.695 44.825 ;
    RECT 8.095 43.945 8.375 44.825 ;
    RECT 4.775 43.945 5.055 44.825 ;
    RECT 1.455 43.945 1.735 44.825 ;
    RECT 64.535 43.945 64.815 44.825 ;
    RECT 61.215 83.565 61.495 84.445 ;
    RECT 57.895 83.565 58.175 84.445 ;
    RECT 54.575 83.565 54.855 84.445 ;
    RECT 51.255 83.565 51.535 84.445 ;
    RECT 47.935 83.565 48.215 84.445 ;
    RECT 44.615 83.565 44.895 84.445 ;
    RECT 41.295 83.565 41.575 84.445 ;
    RECT 37.975 83.565 38.255 84.445 ;
    RECT 34.655 83.565 34.935 84.445 ;
    RECT 117.655 83.565 117.935 84.445 ;
    RECT 114.335 83.565 114.615 84.445 ;
    RECT 111.015 83.565 111.295 84.445 ;
    RECT 107.695 83.565 107.975 84.445 ;
    RECT 104.375 83.565 104.655 84.445 ;
    RECT 101.055 83.565 101.335 84.445 ;
    RECT 97.735 83.565 98.015 84.445 ;
    RECT 94.415 83.565 94.695 84.445 ;
    RECT 91.095 83.565 91.375 84.445 ;
    RECT 87.775 83.565 88.055 84.445 ;
    RECT 84.455 83.565 84.735 84.445 ;
    RECT 81.135 83.565 81.415 84.445 ;
    RECT 77.815 83.565 78.095 84.445 ;
    RECT 74.495 83.565 74.775 84.445 ;
    RECT 71.175 83.565 71.455 84.445 ;
    RECT 31.335 83.565 31.615 84.445 ;
    RECT 67.855 83.565 68.135 84.445 ;
    RECT 28.015 83.565 28.295 84.445 ;
    RECT 24.695 83.565 24.975 84.445 ;
    RECT 21.375 83.565 21.655 84.445 ;
    RECT 18.055 83.565 18.335 84.445 ;
    RECT 14.735 83.565 15.015 84.445 ;
    RECT 11.415 83.565 11.695 84.445 ;
    RECT 8.095 83.565 8.375 84.445 ;
    RECT 4.775 83.565 5.055 84.445 ;
    RECT 1.455 83.565 1.735 84.445 ;
    RECT 64.535 83.565 64.815 84.445 ;
    RECT 61.215 43.225 61.495 44.105 ;
    RECT 57.895 43.225 58.175 44.105 ;
    RECT 54.575 43.225 54.855 44.105 ;
    RECT 51.255 43.225 51.535 44.105 ;
    RECT 47.935 43.225 48.215 44.105 ;
    RECT 44.615 43.225 44.895 44.105 ;
    RECT 41.295 43.225 41.575 44.105 ;
    RECT 37.975 43.225 38.255 44.105 ;
    RECT 34.655 43.225 34.935 44.105 ;
    RECT 117.655 43.225 117.935 44.105 ;
    RECT 114.335 43.225 114.615 44.105 ;
    RECT 111.015 43.225 111.295 44.105 ;
    RECT 107.695 43.225 107.975 44.105 ;
    RECT 104.375 43.225 104.655 44.105 ;
    RECT 101.055 43.225 101.335 44.105 ;
    RECT 97.735 43.225 98.015 44.105 ;
    RECT 94.415 43.225 94.695 44.105 ;
    RECT 91.095 43.225 91.375 44.105 ;
    RECT 87.775 43.225 88.055 44.105 ;
    RECT 84.455 43.225 84.735 44.105 ;
    RECT 81.135 43.225 81.415 44.105 ;
    RECT 77.815 43.225 78.095 44.105 ;
    RECT 74.495 43.225 74.775 44.105 ;
    RECT 71.175 43.225 71.455 44.105 ;
    RECT 31.335 43.225 31.615 44.105 ;
    RECT 67.855 43.225 68.135 44.105 ;
    RECT 28.015 43.225 28.295 44.105 ;
    RECT 24.695 43.225 24.975 44.105 ;
    RECT 21.375 43.225 21.655 44.105 ;
    RECT 18.055 43.225 18.335 44.105 ;
    RECT 14.735 43.225 15.015 44.105 ;
    RECT 11.415 43.225 11.695 44.105 ;
    RECT 8.095 43.225 8.375 44.105 ;
    RECT 4.775 43.225 5.055 44.105 ;
    RECT 1.455 43.225 1.735 44.105 ;
    RECT 64.535 43.225 64.815 44.105 ;
    RECT 61.215 82.845 61.495 83.725 ;
    RECT 57.895 82.845 58.175 83.725 ;
    RECT 54.575 82.845 54.855 83.725 ;
    RECT 51.255 82.845 51.535 83.725 ;
    RECT 47.935 82.845 48.215 83.725 ;
    RECT 44.615 82.845 44.895 83.725 ;
    RECT 41.295 82.845 41.575 83.725 ;
    RECT 37.975 82.845 38.255 83.725 ;
    RECT 34.655 82.845 34.935 83.725 ;
    RECT 117.655 82.845 117.935 83.725 ;
    RECT 114.335 82.845 114.615 83.725 ;
    RECT 111.015 82.845 111.295 83.725 ;
    RECT 107.695 82.845 107.975 83.725 ;
    RECT 104.375 82.845 104.655 83.725 ;
    RECT 101.055 82.845 101.335 83.725 ;
    RECT 97.735 82.845 98.015 83.725 ;
    RECT 94.415 82.845 94.695 83.725 ;
    RECT 91.095 82.845 91.375 83.725 ;
    RECT 87.775 82.845 88.055 83.725 ;
    RECT 84.455 82.845 84.735 83.725 ;
    RECT 81.135 82.845 81.415 83.725 ;
    RECT 77.815 82.845 78.095 83.725 ;
    RECT 74.495 82.845 74.775 83.725 ;
    RECT 71.175 82.845 71.455 83.725 ;
    RECT 31.335 82.845 31.615 83.725 ;
    RECT 67.855 82.845 68.135 83.725 ;
    RECT 28.015 82.845 28.295 83.725 ;
    RECT 24.695 82.845 24.975 83.725 ;
    RECT 21.375 82.845 21.655 83.725 ;
    RECT 18.055 82.845 18.335 83.725 ;
    RECT 14.735 82.845 15.015 83.725 ;
    RECT 11.415 82.845 11.695 83.725 ;
    RECT 8.095 82.845 8.375 83.725 ;
    RECT 4.775 82.845 5.055 83.725 ;
    RECT 1.455 82.845 1.735 83.725 ;
    RECT 64.535 82.845 64.815 83.725 ;
    RECT 61.215 82.125 61.495 83.005 ;
    RECT 57.895 82.125 58.175 83.005 ;
    RECT 54.575 82.125 54.855 83.005 ;
    RECT 51.255 82.125 51.535 83.005 ;
    RECT 47.935 82.125 48.215 83.005 ;
    RECT 44.615 82.125 44.895 83.005 ;
    RECT 41.295 82.125 41.575 83.005 ;
    RECT 37.975 82.125 38.255 83.005 ;
    RECT 34.655 82.125 34.935 83.005 ;
    RECT 117.655 82.125 117.935 83.005 ;
    RECT 114.335 82.125 114.615 83.005 ;
    RECT 111.015 82.125 111.295 83.005 ;
    RECT 107.695 82.125 107.975 83.005 ;
    RECT 104.375 82.125 104.655 83.005 ;
    RECT 101.055 82.125 101.335 83.005 ;
    RECT 97.735 82.125 98.015 83.005 ;
    RECT 94.415 82.125 94.695 83.005 ;
    RECT 91.095 82.125 91.375 83.005 ;
    RECT 87.775 82.125 88.055 83.005 ;
    RECT 84.455 82.125 84.735 83.005 ;
    RECT 81.135 82.125 81.415 83.005 ;
    RECT 77.815 82.125 78.095 83.005 ;
    RECT 74.495 82.125 74.775 83.005 ;
    RECT 71.175 82.125 71.455 83.005 ;
    RECT 31.335 82.125 31.615 83.005 ;
    RECT 67.855 82.125 68.135 83.005 ;
    RECT 28.015 82.125 28.295 83.005 ;
    RECT 24.695 82.125 24.975 83.005 ;
    RECT 21.375 82.125 21.655 83.005 ;
    RECT 18.055 82.125 18.335 83.005 ;
    RECT 14.735 82.125 15.015 83.005 ;
    RECT 11.415 82.125 11.695 83.005 ;
    RECT 8.095 82.125 8.375 83.005 ;
    RECT 4.775 82.125 5.055 83.005 ;
    RECT 1.455 82.125 1.735 83.005 ;
    RECT 64.535 82.125 64.815 83.005 ;
    RECT 61.215 81.405 61.495 82.285 ;
    RECT 57.895 81.405 58.175 82.285 ;
    RECT 54.575 81.405 54.855 82.285 ;
    RECT 51.255 81.405 51.535 82.285 ;
    RECT 47.935 81.405 48.215 82.285 ;
    RECT 44.615 81.405 44.895 82.285 ;
    RECT 41.295 81.405 41.575 82.285 ;
    RECT 37.975 81.405 38.255 82.285 ;
    RECT 34.655 81.405 34.935 82.285 ;
    RECT 117.655 81.405 117.935 82.285 ;
    RECT 114.335 81.405 114.615 82.285 ;
    RECT 111.015 81.405 111.295 82.285 ;
    RECT 107.695 81.405 107.975 82.285 ;
    RECT 104.375 81.405 104.655 82.285 ;
    RECT 101.055 81.405 101.335 82.285 ;
    RECT 97.735 81.405 98.015 82.285 ;
    RECT 94.415 81.405 94.695 82.285 ;
    RECT 91.095 81.405 91.375 82.285 ;
    RECT 87.775 81.405 88.055 82.285 ;
    RECT 84.455 81.405 84.735 82.285 ;
    RECT 81.135 81.405 81.415 82.285 ;
    RECT 77.815 81.405 78.095 82.285 ;
    RECT 74.495 81.405 74.775 82.285 ;
    RECT 71.175 81.405 71.455 82.285 ;
    RECT 31.335 81.405 31.615 82.285 ;
    RECT 67.855 81.405 68.135 82.285 ;
    RECT 28.015 81.405 28.295 82.285 ;
    RECT 24.695 81.405 24.975 82.285 ;
    RECT 21.375 81.405 21.655 82.285 ;
    RECT 18.055 81.405 18.335 82.285 ;
    RECT 14.735 81.405 15.015 82.285 ;
    RECT 11.415 81.405 11.695 82.285 ;
    RECT 8.095 81.405 8.375 82.285 ;
    RECT 4.775 81.405 5.055 82.285 ;
    RECT 1.455 81.405 1.735 82.285 ;
    RECT 64.535 81.405 64.815 82.285 ;
    RECT 61.215 80.685 61.495 81.565 ;
    RECT 57.895 80.685 58.175 81.565 ;
    RECT 54.575 80.685 54.855 81.565 ;
    RECT 51.255 80.685 51.535 81.565 ;
    RECT 47.935 80.685 48.215 81.565 ;
    RECT 44.615 80.685 44.895 81.565 ;
    RECT 41.295 80.685 41.575 81.565 ;
    RECT 37.975 80.685 38.255 81.565 ;
    RECT 34.655 80.685 34.935 81.565 ;
    RECT 117.655 80.685 117.935 81.565 ;
    RECT 114.335 80.685 114.615 81.565 ;
    RECT 111.015 80.685 111.295 81.565 ;
    RECT 107.695 80.685 107.975 81.565 ;
    RECT 104.375 80.685 104.655 81.565 ;
    RECT 101.055 80.685 101.335 81.565 ;
    RECT 97.735 80.685 98.015 81.565 ;
    RECT 94.415 80.685 94.695 81.565 ;
    RECT 91.095 80.685 91.375 81.565 ;
    RECT 87.775 80.685 88.055 81.565 ;
    RECT 84.455 80.685 84.735 81.565 ;
    RECT 81.135 80.685 81.415 81.565 ;
    RECT 77.815 80.685 78.095 81.565 ;
    RECT 74.495 80.685 74.775 81.565 ;
    RECT 71.175 80.685 71.455 81.565 ;
    RECT 31.335 80.685 31.615 81.565 ;
    RECT 67.855 80.685 68.135 81.565 ;
    RECT 28.015 80.685 28.295 81.565 ;
    RECT 24.695 80.685 24.975 81.565 ;
    RECT 21.375 80.685 21.655 81.565 ;
    RECT 18.055 80.685 18.335 81.565 ;
    RECT 14.735 80.685 15.015 81.565 ;
    RECT 11.415 80.685 11.695 81.565 ;
    RECT 8.095 80.685 8.375 81.565 ;
    RECT 4.775 80.685 5.055 81.565 ;
    RECT 1.455 80.685 1.735 81.565 ;
    RECT 64.535 80.685 64.815 81.565 ;
    RECT 61.215 79.965 61.495 80.845 ;
    RECT 57.895 79.965 58.175 80.845 ;
    RECT 54.575 79.965 54.855 80.845 ;
    RECT 51.255 79.965 51.535 80.845 ;
    RECT 47.935 79.965 48.215 80.845 ;
    RECT 44.615 79.965 44.895 80.845 ;
    RECT 41.295 79.965 41.575 80.845 ;
    RECT 37.975 79.965 38.255 80.845 ;
    RECT 34.655 79.965 34.935 80.845 ;
    RECT 117.655 79.965 117.935 80.845 ;
    RECT 114.335 79.965 114.615 80.845 ;
    RECT 111.015 79.965 111.295 80.845 ;
    RECT 107.695 79.965 107.975 80.845 ;
    RECT 104.375 79.965 104.655 80.845 ;
    RECT 101.055 79.965 101.335 80.845 ;
    RECT 97.735 79.965 98.015 80.845 ;
    RECT 94.415 79.965 94.695 80.845 ;
    RECT 91.095 79.965 91.375 80.845 ;
    RECT 87.775 79.965 88.055 80.845 ;
    RECT 84.455 79.965 84.735 80.845 ;
    RECT 81.135 79.965 81.415 80.845 ;
    RECT 77.815 79.965 78.095 80.845 ;
    RECT 74.495 79.965 74.775 80.845 ;
    RECT 71.175 79.965 71.455 80.845 ;
    RECT 31.335 79.965 31.615 80.845 ;
    RECT 67.855 79.965 68.135 80.845 ;
    RECT 28.015 79.965 28.295 80.845 ;
    RECT 24.695 79.965 24.975 80.845 ;
    RECT 21.375 79.965 21.655 80.845 ;
    RECT 18.055 79.965 18.335 80.845 ;
    RECT 14.735 79.965 15.015 80.845 ;
    RECT 11.415 79.965 11.695 80.845 ;
    RECT 8.095 79.965 8.375 80.845 ;
    RECT 4.775 79.965 5.055 80.845 ;
    RECT 1.455 79.965 1.735 80.845 ;
    RECT 64.535 79.965 64.815 80.845 ;
    RECT 61.215 42.505 61.495 43.385 ;
    RECT 57.895 42.505 58.175 43.385 ;
    RECT 54.575 42.505 54.855 43.385 ;
    RECT 51.255 42.505 51.535 43.385 ;
    RECT 47.935 42.505 48.215 43.385 ;
    RECT 44.615 42.505 44.895 43.385 ;
    RECT 41.295 42.505 41.575 43.385 ;
    RECT 37.975 42.505 38.255 43.385 ;
    RECT 34.655 42.505 34.935 43.385 ;
    RECT 117.655 42.505 117.935 43.385 ;
    RECT 114.335 42.505 114.615 43.385 ;
    RECT 111.015 42.505 111.295 43.385 ;
    RECT 107.695 42.505 107.975 43.385 ;
    RECT 104.375 42.505 104.655 43.385 ;
    RECT 101.055 42.505 101.335 43.385 ;
    RECT 97.735 42.505 98.015 43.385 ;
    RECT 94.415 42.505 94.695 43.385 ;
    RECT 91.095 42.505 91.375 43.385 ;
    RECT 87.775 42.505 88.055 43.385 ;
    RECT 84.455 42.505 84.735 43.385 ;
    RECT 81.135 42.505 81.415 43.385 ;
    RECT 77.815 42.505 78.095 43.385 ;
    RECT 74.495 42.505 74.775 43.385 ;
    RECT 71.175 42.505 71.455 43.385 ;
    RECT 31.335 42.505 31.615 43.385 ;
    RECT 67.855 42.505 68.135 43.385 ;
    RECT 28.015 42.505 28.295 43.385 ;
    RECT 24.695 42.505 24.975 43.385 ;
    RECT 21.375 42.505 21.655 43.385 ;
    RECT 18.055 42.505 18.335 43.385 ;
    RECT 14.735 42.505 15.015 43.385 ;
    RECT 11.415 42.505 11.695 43.385 ;
    RECT 8.095 42.505 8.375 43.385 ;
    RECT 4.775 42.505 5.055 43.385 ;
    RECT 1.455 42.505 1.735 43.385 ;
    RECT 64.535 42.505 64.815 43.385 ;
    RECT 61.215 97.965 61.495 98.845 ;
    RECT 57.895 97.965 58.175 98.845 ;
    RECT 54.575 97.965 54.855 98.845 ;
    RECT 117.655 97.965 117.935 98.845 ;
    RECT 51.255 97.965 51.535 98.845 ;
    RECT 47.935 97.965 48.215 98.845 ;
    RECT 44.615 97.965 44.895 98.845 ;
    RECT 41.295 97.965 41.575 98.845 ;
    RECT 37.975 97.965 38.255 98.845 ;
    RECT 34.655 97.965 34.935 98.845 ;
    RECT 1.455 97.965 1.735 98.845 ;
    RECT 114.335 97.965 114.615 98.845 ;
    RECT 111.015 97.965 111.295 98.845 ;
    RECT 107.695 97.965 107.975 98.845 ;
    RECT 104.375 97.965 104.655 98.845 ;
    RECT 101.055 97.965 101.335 98.845 ;
    RECT 97.735 97.965 98.015 98.845 ;
    RECT 94.415 97.965 94.695 98.845 ;
    RECT 91.095 97.965 91.375 98.845 ;
    RECT 87.775 97.965 88.055 98.845 ;
    RECT 84.455 97.965 84.735 98.845 ;
    RECT 81.135 97.965 81.415 98.845 ;
    RECT 77.815 97.965 78.095 98.845 ;
    RECT 74.495 97.965 74.775 98.845 ;
    RECT 71.175 97.965 71.455 98.845 ;
    RECT 31.335 97.965 31.615 98.845 ;
    RECT 67.855 97.965 68.135 98.845 ;
    RECT 28.015 97.965 28.295 98.845 ;
    RECT 24.695 97.965 24.975 98.845 ;
    RECT 21.375 97.965 21.655 98.845 ;
    RECT 18.055 97.965 18.335 98.845 ;
    RECT 14.735 97.965 15.015 98.845 ;
    RECT 11.415 97.965 11.695 98.845 ;
    RECT 8.095 97.965 8.375 98.845 ;
    RECT 4.775 97.965 5.055 98.845 ;
    RECT 64.535 97.965 64.815 98.845 ;
    RECT 61.215 41.785 61.495 42.665 ;
    RECT 57.895 41.785 58.175 42.665 ;
    RECT 54.575 41.785 54.855 42.665 ;
    RECT 51.255 41.785 51.535 42.665 ;
    RECT 47.935 41.785 48.215 42.665 ;
    RECT 44.615 41.785 44.895 42.665 ;
    RECT 41.295 41.785 41.575 42.665 ;
    RECT 37.975 41.785 38.255 42.665 ;
    RECT 34.655 41.785 34.935 42.665 ;
    RECT 117.655 41.785 117.935 42.665 ;
    RECT 114.335 41.785 114.615 42.665 ;
    RECT 111.015 41.785 111.295 42.665 ;
    RECT 107.695 41.785 107.975 42.665 ;
    RECT 104.375 41.785 104.655 42.665 ;
    RECT 101.055 41.785 101.335 42.665 ;
    RECT 97.735 41.785 98.015 42.665 ;
    RECT 94.415 41.785 94.695 42.665 ;
    RECT 91.095 41.785 91.375 42.665 ;
    RECT 87.775 41.785 88.055 42.665 ;
    RECT 84.455 41.785 84.735 42.665 ;
    RECT 81.135 41.785 81.415 42.665 ;
    RECT 77.815 41.785 78.095 42.665 ;
    RECT 74.495 41.785 74.775 42.665 ;
    RECT 71.175 41.785 71.455 42.665 ;
    RECT 31.335 41.785 31.615 42.665 ;
    RECT 67.855 41.785 68.135 42.665 ;
    RECT 28.015 41.785 28.295 42.665 ;
    RECT 24.695 41.785 24.975 42.665 ;
    RECT 21.375 41.785 21.655 42.665 ;
    RECT 18.055 41.785 18.335 42.665 ;
    RECT 14.735 41.785 15.015 42.665 ;
    RECT 11.415 41.785 11.695 42.665 ;
    RECT 8.095 41.785 8.375 42.665 ;
    RECT 4.775 41.785 5.055 42.665 ;
    RECT 1.455 41.785 1.735 42.665 ;
    RECT 64.535 41.785 64.815 42.665 ;
    RECT 61.215 41.065 61.495 41.945 ;
    RECT 57.895 41.065 58.175 41.945 ;
    RECT 54.575 41.065 54.855 41.945 ;
    RECT 51.255 41.065 51.535 41.945 ;
    RECT 47.935 41.065 48.215 41.945 ;
    RECT 44.615 41.065 44.895 41.945 ;
    RECT 41.295 41.065 41.575 41.945 ;
    RECT 37.975 41.065 38.255 41.945 ;
    RECT 34.655 41.065 34.935 41.945 ;
    RECT 117.655 41.065 117.935 41.945 ;
    RECT 114.335 41.065 114.615 41.945 ;
    RECT 111.015 41.065 111.295 41.945 ;
    RECT 107.695 41.065 107.975 41.945 ;
    RECT 104.375 41.065 104.655 41.945 ;
    RECT 101.055 41.065 101.335 41.945 ;
    RECT 97.735 41.065 98.015 41.945 ;
    RECT 94.415 41.065 94.695 41.945 ;
    RECT 91.095 41.065 91.375 41.945 ;
    RECT 87.775 41.065 88.055 41.945 ;
    RECT 84.455 41.065 84.735 41.945 ;
    RECT 81.135 41.065 81.415 41.945 ;
    RECT 77.815 41.065 78.095 41.945 ;
    RECT 74.495 41.065 74.775 41.945 ;
    RECT 71.175 41.065 71.455 41.945 ;
    RECT 31.335 41.065 31.615 41.945 ;
    RECT 67.855 41.065 68.135 41.945 ;
    RECT 28.015 41.065 28.295 41.945 ;
    RECT 24.695 41.065 24.975 41.945 ;
    RECT 21.375 41.065 21.655 41.945 ;
    RECT 18.055 41.065 18.335 41.945 ;
    RECT 14.735 41.065 15.015 41.945 ;
    RECT 11.415 41.065 11.695 41.945 ;
    RECT 8.095 41.065 8.375 41.945 ;
    RECT 4.775 41.065 5.055 41.945 ;
    RECT 1.455 41.065 1.735 41.945 ;
    RECT 64.535 41.065 64.815 41.945 ;
    RECT 61.215 40.345 61.495 41.225 ;
    RECT 57.895 40.345 58.175 41.225 ;
    RECT 54.575 40.345 54.855 41.225 ;
    RECT 51.255 40.345 51.535 41.225 ;
    RECT 47.935 40.345 48.215 41.225 ;
    RECT 44.615 40.345 44.895 41.225 ;
    RECT 41.295 40.345 41.575 41.225 ;
    RECT 37.975 40.345 38.255 41.225 ;
    RECT 34.655 40.345 34.935 41.225 ;
    RECT 117.655 40.345 117.935 41.225 ;
    RECT 114.335 40.345 114.615 41.225 ;
    RECT 111.015 40.345 111.295 41.225 ;
    RECT 107.695 40.345 107.975 41.225 ;
    RECT 104.375 40.345 104.655 41.225 ;
    RECT 101.055 40.345 101.335 41.225 ;
    RECT 97.735 40.345 98.015 41.225 ;
    RECT 94.415 40.345 94.695 41.225 ;
    RECT 91.095 40.345 91.375 41.225 ;
    RECT 87.775 40.345 88.055 41.225 ;
    RECT 84.455 40.345 84.735 41.225 ;
    RECT 81.135 40.345 81.415 41.225 ;
    RECT 77.815 40.345 78.095 41.225 ;
    RECT 74.495 40.345 74.775 41.225 ;
    RECT 71.175 40.345 71.455 41.225 ;
    RECT 31.335 40.345 31.615 41.225 ;
    RECT 67.855 40.345 68.135 41.225 ;
    RECT 28.015 40.345 28.295 41.225 ;
    RECT 24.695 40.345 24.975 41.225 ;
    RECT 21.375 40.345 21.655 41.225 ;
    RECT 18.055 40.345 18.335 41.225 ;
    RECT 14.735 40.345 15.015 41.225 ;
    RECT 11.415 40.345 11.695 41.225 ;
    RECT 8.095 40.345 8.375 41.225 ;
    RECT 4.775 40.345 5.055 41.225 ;
    RECT 1.455 40.345 1.735 41.225 ;
    RECT 64.535 40.345 64.815 41.225 ;
    RECT 61.215 39.625 61.495 40.505 ;
    RECT 57.895 39.625 58.175 40.505 ;
    RECT 54.575 39.625 54.855 40.505 ;
    RECT 51.255 39.625 51.535 40.505 ;
    RECT 47.935 39.625 48.215 40.505 ;
    RECT 44.615 39.625 44.895 40.505 ;
    RECT 41.295 39.625 41.575 40.505 ;
    RECT 37.975 39.625 38.255 40.505 ;
    RECT 34.655 39.625 34.935 40.505 ;
    RECT 117.655 39.625 117.935 40.505 ;
    RECT 114.335 39.625 114.615 40.505 ;
    RECT 111.015 39.625 111.295 40.505 ;
    RECT 107.695 39.625 107.975 40.505 ;
    RECT 104.375 39.625 104.655 40.505 ;
    RECT 101.055 39.625 101.335 40.505 ;
    RECT 97.735 39.625 98.015 40.505 ;
    RECT 94.415 39.625 94.695 40.505 ;
    RECT 91.095 39.625 91.375 40.505 ;
    RECT 87.775 39.625 88.055 40.505 ;
    RECT 84.455 39.625 84.735 40.505 ;
    RECT 81.135 39.625 81.415 40.505 ;
    RECT 77.815 39.625 78.095 40.505 ;
    RECT 74.495 39.625 74.775 40.505 ;
    RECT 71.175 39.625 71.455 40.505 ;
    RECT 31.335 39.625 31.615 40.505 ;
    RECT 67.855 39.625 68.135 40.505 ;
    RECT 28.015 39.625 28.295 40.505 ;
    RECT 24.695 39.625 24.975 40.505 ;
    RECT 21.375 39.625 21.655 40.505 ;
    RECT 18.055 39.625 18.335 40.505 ;
    RECT 14.735 39.625 15.015 40.505 ;
    RECT 11.415 39.625 11.695 40.505 ;
    RECT 8.095 39.625 8.375 40.505 ;
    RECT 4.775 39.625 5.055 40.505 ;
    RECT 1.455 39.625 1.735 40.505 ;
    RECT 64.535 39.625 64.815 40.505 ;
    RECT 61.215 79.245 61.495 80.125 ;
    RECT 57.895 79.245 58.175 80.125 ;
    RECT 54.575 79.245 54.855 80.125 ;
    RECT 51.255 79.245 51.535 80.125 ;
    RECT 47.935 79.245 48.215 80.125 ;
    RECT 44.615 79.245 44.895 80.125 ;
    RECT 41.295 79.245 41.575 80.125 ;
    RECT 37.975 79.245 38.255 80.125 ;
    RECT 34.655 79.245 34.935 80.125 ;
    RECT 117.655 79.245 117.935 80.125 ;
    RECT 114.335 79.245 114.615 80.125 ;
    RECT 111.015 79.245 111.295 80.125 ;
    RECT 107.695 79.245 107.975 80.125 ;
    RECT 104.375 79.245 104.655 80.125 ;
    RECT 101.055 79.245 101.335 80.125 ;
    RECT 97.735 79.245 98.015 80.125 ;
    RECT 94.415 79.245 94.695 80.125 ;
    RECT 91.095 79.245 91.375 80.125 ;
    RECT 87.775 79.245 88.055 80.125 ;
    RECT 84.455 79.245 84.735 80.125 ;
    RECT 81.135 79.245 81.415 80.125 ;
    RECT 77.815 79.245 78.095 80.125 ;
    RECT 74.495 79.245 74.775 80.125 ;
    RECT 71.175 79.245 71.455 80.125 ;
    RECT 31.335 79.245 31.615 80.125 ;
    RECT 67.855 79.245 68.135 80.125 ;
    RECT 28.015 79.245 28.295 80.125 ;
    RECT 24.695 79.245 24.975 80.125 ;
    RECT 21.375 79.245 21.655 80.125 ;
    RECT 18.055 79.245 18.335 80.125 ;
    RECT 14.735 79.245 15.015 80.125 ;
    RECT 11.415 79.245 11.695 80.125 ;
    RECT 8.095 79.245 8.375 80.125 ;
    RECT 4.775 79.245 5.055 80.125 ;
    RECT 1.455 79.245 1.735 80.125 ;
    RECT 64.535 79.245 64.815 80.125 ;
    RECT 61.215 38.905 61.495 39.785 ;
    RECT 57.895 38.905 58.175 39.785 ;
    RECT 54.575 38.905 54.855 39.785 ;
    RECT 51.255 38.905 51.535 39.785 ;
    RECT 47.935 38.905 48.215 39.785 ;
    RECT 44.615 38.905 44.895 39.785 ;
    RECT 41.295 38.905 41.575 39.785 ;
    RECT 37.975 38.905 38.255 39.785 ;
    RECT 34.655 38.905 34.935 39.785 ;
    RECT 117.655 38.905 117.935 39.785 ;
    RECT 114.335 38.905 114.615 39.785 ;
    RECT 111.015 38.905 111.295 39.785 ;
    RECT 107.695 38.905 107.975 39.785 ;
    RECT 104.375 38.905 104.655 39.785 ;
    RECT 101.055 38.905 101.335 39.785 ;
    RECT 97.735 38.905 98.015 39.785 ;
    RECT 94.415 38.905 94.695 39.785 ;
    RECT 91.095 38.905 91.375 39.785 ;
    RECT 87.775 38.905 88.055 39.785 ;
    RECT 84.455 38.905 84.735 39.785 ;
    RECT 81.135 38.905 81.415 39.785 ;
    RECT 77.815 38.905 78.095 39.785 ;
    RECT 74.495 38.905 74.775 39.785 ;
    RECT 71.175 38.905 71.455 39.785 ;
    RECT 31.335 38.905 31.615 39.785 ;
    RECT 67.855 38.905 68.135 39.785 ;
    RECT 28.015 38.905 28.295 39.785 ;
    RECT 24.695 38.905 24.975 39.785 ;
    RECT 21.375 38.905 21.655 39.785 ;
    RECT 18.055 38.905 18.335 39.785 ;
    RECT 14.735 38.905 15.015 39.785 ;
    RECT 11.415 38.905 11.695 39.785 ;
    RECT 8.095 38.905 8.375 39.785 ;
    RECT 4.775 38.905 5.055 39.785 ;
    RECT 1.455 38.905 1.735 39.785 ;
    RECT 64.535 38.905 64.815 39.785 ;
    RECT 61.215 78.525 61.495 79.405 ;
    RECT 57.895 78.525 58.175 79.405 ;
    RECT 54.575 78.525 54.855 79.405 ;
    RECT 51.255 78.525 51.535 79.405 ;
    RECT 47.935 78.525 48.215 79.405 ;
    RECT 44.615 78.525 44.895 79.405 ;
    RECT 41.295 78.525 41.575 79.405 ;
    RECT 37.975 78.525 38.255 79.405 ;
    RECT 34.655 78.525 34.935 79.405 ;
    RECT 117.655 78.525 117.935 79.405 ;
    RECT 114.335 78.525 114.615 79.405 ;
    RECT 111.015 78.525 111.295 79.405 ;
    RECT 107.695 78.525 107.975 79.405 ;
    RECT 104.375 78.525 104.655 79.405 ;
    RECT 101.055 78.525 101.335 79.405 ;
    RECT 97.735 78.525 98.015 79.405 ;
    RECT 94.415 78.525 94.695 79.405 ;
    RECT 91.095 78.525 91.375 79.405 ;
    RECT 87.775 78.525 88.055 79.405 ;
    RECT 84.455 78.525 84.735 79.405 ;
    RECT 81.135 78.525 81.415 79.405 ;
    RECT 77.815 78.525 78.095 79.405 ;
    RECT 74.495 78.525 74.775 79.405 ;
    RECT 71.175 78.525 71.455 79.405 ;
    RECT 31.335 78.525 31.615 79.405 ;
    RECT 67.855 78.525 68.135 79.405 ;
    RECT 28.015 78.525 28.295 79.405 ;
    RECT 24.695 78.525 24.975 79.405 ;
    RECT 21.375 78.525 21.655 79.405 ;
    RECT 18.055 78.525 18.335 79.405 ;
    RECT 14.735 78.525 15.015 79.405 ;
    RECT 11.415 78.525 11.695 79.405 ;
    RECT 8.095 78.525 8.375 79.405 ;
    RECT 4.775 78.525 5.055 79.405 ;
    RECT 1.455 78.525 1.735 79.405 ;
    RECT 64.535 78.525 64.815 79.405 ;
    RECT 61.215 38.185 61.495 39.065 ;
    RECT 57.895 38.185 58.175 39.065 ;
    RECT 54.575 38.185 54.855 39.065 ;
    RECT 51.255 38.185 51.535 39.065 ;
    RECT 47.935 38.185 48.215 39.065 ;
    RECT 44.615 38.185 44.895 39.065 ;
    RECT 41.295 38.185 41.575 39.065 ;
    RECT 37.975 38.185 38.255 39.065 ;
    RECT 34.655 38.185 34.935 39.065 ;
    RECT 117.655 38.185 117.935 39.065 ;
    RECT 114.335 38.185 114.615 39.065 ;
    RECT 111.015 38.185 111.295 39.065 ;
    RECT 107.695 38.185 107.975 39.065 ;
    RECT 104.375 38.185 104.655 39.065 ;
    RECT 101.055 38.185 101.335 39.065 ;
    RECT 97.735 38.185 98.015 39.065 ;
    RECT 94.415 38.185 94.695 39.065 ;
    RECT 91.095 38.185 91.375 39.065 ;
    RECT 87.775 38.185 88.055 39.065 ;
    RECT 84.455 38.185 84.735 39.065 ;
    RECT 81.135 38.185 81.415 39.065 ;
    RECT 77.815 38.185 78.095 39.065 ;
    RECT 74.495 38.185 74.775 39.065 ;
    RECT 71.175 38.185 71.455 39.065 ;
    RECT 31.335 38.185 31.615 39.065 ;
    RECT 67.855 38.185 68.135 39.065 ;
    RECT 28.015 38.185 28.295 39.065 ;
    RECT 24.695 38.185 24.975 39.065 ;
    RECT 21.375 38.185 21.655 39.065 ;
    RECT 18.055 38.185 18.335 39.065 ;
    RECT 14.735 38.185 15.015 39.065 ;
    RECT 11.415 38.185 11.695 39.065 ;
    RECT 8.095 38.185 8.375 39.065 ;
    RECT 4.775 38.185 5.055 39.065 ;
    RECT 1.455 38.185 1.735 39.065 ;
    RECT 64.535 38.185 64.815 39.065 ;
    RECT 61.215 77.805 61.495 78.685 ;
    RECT 57.895 77.805 58.175 78.685 ;
    RECT 54.575 77.805 54.855 78.685 ;
    RECT 51.255 77.805 51.535 78.685 ;
    RECT 47.935 77.805 48.215 78.685 ;
    RECT 44.615 77.805 44.895 78.685 ;
    RECT 41.295 77.805 41.575 78.685 ;
    RECT 37.975 77.805 38.255 78.685 ;
    RECT 34.655 77.805 34.935 78.685 ;
    RECT 117.655 77.805 117.935 78.685 ;
    RECT 114.335 77.805 114.615 78.685 ;
    RECT 111.015 77.805 111.295 78.685 ;
    RECT 107.695 77.805 107.975 78.685 ;
    RECT 104.375 77.805 104.655 78.685 ;
    RECT 101.055 77.805 101.335 78.685 ;
    RECT 97.735 77.805 98.015 78.685 ;
    RECT 94.415 77.805 94.695 78.685 ;
    RECT 91.095 77.805 91.375 78.685 ;
    RECT 87.775 77.805 88.055 78.685 ;
    RECT 84.455 77.805 84.735 78.685 ;
    RECT 81.135 77.805 81.415 78.685 ;
    RECT 77.815 77.805 78.095 78.685 ;
    RECT 74.495 77.805 74.775 78.685 ;
    RECT 71.175 77.805 71.455 78.685 ;
    RECT 31.335 77.805 31.615 78.685 ;
    RECT 67.855 77.805 68.135 78.685 ;
    RECT 28.015 77.805 28.295 78.685 ;
    RECT 24.695 77.805 24.975 78.685 ;
    RECT 21.375 77.805 21.655 78.685 ;
    RECT 18.055 77.805 18.335 78.685 ;
    RECT 14.735 77.805 15.015 78.685 ;
    RECT 11.415 77.805 11.695 78.685 ;
    RECT 8.095 77.805 8.375 78.685 ;
    RECT 4.775 77.805 5.055 78.685 ;
    RECT 1.455 77.805 1.735 78.685 ;
    RECT 64.535 77.805 64.815 78.685 ;
    RECT 61.215 37.465 61.495 38.345 ;
    RECT 57.895 37.465 58.175 38.345 ;
    RECT 54.575 37.465 54.855 38.345 ;
    RECT 51.255 37.465 51.535 38.345 ;
    RECT 47.935 37.465 48.215 38.345 ;
    RECT 44.615 37.465 44.895 38.345 ;
    RECT 41.295 37.465 41.575 38.345 ;
    RECT 37.975 37.465 38.255 38.345 ;
    RECT 34.655 37.465 34.935 38.345 ;
    RECT 117.655 37.465 117.935 38.345 ;
    RECT 114.335 37.465 114.615 38.345 ;
    RECT 111.015 37.465 111.295 38.345 ;
    RECT 107.695 37.465 107.975 38.345 ;
    RECT 104.375 37.465 104.655 38.345 ;
    RECT 101.055 37.465 101.335 38.345 ;
    RECT 97.735 37.465 98.015 38.345 ;
    RECT 94.415 37.465 94.695 38.345 ;
    RECT 91.095 37.465 91.375 38.345 ;
    RECT 87.775 37.465 88.055 38.345 ;
    RECT 84.455 37.465 84.735 38.345 ;
    RECT 81.135 37.465 81.415 38.345 ;
    RECT 77.815 37.465 78.095 38.345 ;
    RECT 74.495 37.465 74.775 38.345 ;
    RECT 71.175 37.465 71.455 38.345 ;
    RECT 31.335 37.465 31.615 38.345 ;
    RECT 67.855 37.465 68.135 38.345 ;
    RECT 28.015 37.465 28.295 38.345 ;
    RECT 24.695 37.465 24.975 38.345 ;
    RECT 21.375 37.465 21.655 38.345 ;
    RECT 18.055 37.465 18.335 38.345 ;
    RECT 14.735 37.465 15.015 38.345 ;
    RECT 11.415 37.465 11.695 38.345 ;
    RECT 8.095 37.465 8.375 38.345 ;
    RECT 4.775 37.465 5.055 38.345 ;
    RECT 1.455 37.465 1.735 38.345 ;
    RECT 64.535 37.465 64.815 38.345 ;
    RECT 61.215 77.085 61.495 77.965 ;
    RECT 57.895 77.085 58.175 77.965 ;
    RECT 54.575 77.085 54.855 77.965 ;
    RECT 51.255 77.085 51.535 77.965 ;
    RECT 47.935 77.085 48.215 77.965 ;
    RECT 44.615 77.085 44.895 77.965 ;
    RECT 41.295 77.085 41.575 77.965 ;
    RECT 37.975 77.085 38.255 77.965 ;
    RECT 34.655 77.085 34.935 77.965 ;
    RECT 117.655 77.085 117.935 77.965 ;
    RECT 114.335 77.085 114.615 77.965 ;
    RECT 111.015 77.085 111.295 77.965 ;
    RECT 107.695 77.085 107.975 77.965 ;
    RECT 104.375 77.085 104.655 77.965 ;
    RECT 101.055 77.085 101.335 77.965 ;
    RECT 97.735 77.085 98.015 77.965 ;
    RECT 94.415 77.085 94.695 77.965 ;
    RECT 91.095 77.085 91.375 77.965 ;
    RECT 87.775 77.085 88.055 77.965 ;
    RECT 84.455 77.085 84.735 77.965 ;
    RECT 81.135 77.085 81.415 77.965 ;
    RECT 77.815 77.085 78.095 77.965 ;
    RECT 74.495 77.085 74.775 77.965 ;
    RECT 71.175 77.085 71.455 77.965 ;
    RECT 31.335 77.085 31.615 77.965 ;
    RECT 67.855 77.085 68.135 77.965 ;
    RECT 28.015 77.085 28.295 77.965 ;
    RECT 24.695 77.085 24.975 77.965 ;
    RECT 21.375 77.085 21.655 77.965 ;
    RECT 18.055 77.085 18.335 77.965 ;
    RECT 14.735 77.085 15.015 77.965 ;
    RECT 11.415 77.085 11.695 77.965 ;
    RECT 8.095 77.085 8.375 77.965 ;
    RECT 4.775 77.085 5.055 77.965 ;
    RECT 1.455 77.085 1.735 77.965 ;
    RECT 64.535 77.085 64.815 77.965 ;
    RECT 61.215 36.745 61.495 37.625 ;
    RECT 57.895 36.745 58.175 37.625 ;
    RECT 54.575 36.745 54.855 37.625 ;
    RECT 51.255 36.745 51.535 37.625 ;
    RECT 47.935 36.745 48.215 37.625 ;
    RECT 44.615 36.745 44.895 37.625 ;
    RECT 41.295 36.745 41.575 37.625 ;
    RECT 37.975 36.745 38.255 37.625 ;
    RECT 34.655 36.745 34.935 37.625 ;
    RECT 117.655 36.745 117.935 37.625 ;
    RECT 114.335 36.745 114.615 37.625 ;
    RECT 111.015 36.745 111.295 37.625 ;
    RECT 107.695 36.745 107.975 37.625 ;
    RECT 104.375 36.745 104.655 37.625 ;
    RECT 101.055 36.745 101.335 37.625 ;
    RECT 97.735 36.745 98.015 37.625 ;
    RECT 94.415 36.745 94.695 37.625 ;
    RECT 91.095 36.745 91.375 37.625 ;
    RECT 87.775 36.745 88.055 37.625 ;
    RECT 84.455 36.745 84.735 37.625 ;
    RECT 81.135 36.745 81.415 37.625 ;
    RECT 77.815 36.745 78.095 37.625 ;
    RECT 74.495 36.745 74.775 37.625 ;
    RECT 71.175 36.745 71.455 37.625 ;
    RECT 31.335 36.745 31.615 37.625 ;
    RECT 67.855 36.745 68.135 37.625 ;
    RECT 28.015 36.745 28.295 37.625 ;
    RECT 24.695 36.745 24.975 37.625 ;
    RECT 21.375 36.745 21.655 37.625 ;
    RECT 18.055 36.745 18.335 37.625 ;
    RECT 14.735 36.745 15.015 37.625 ;
    RECT 11.415 36.745 11.695 37.625 ;
    RECT 8.095 36.745 8.375 37.625 ;
    RECT 4.775 36.745 5.055 37.625 ;
    RECT 1.455 36.745 1.735 37.625 ;
    RECT 64.535 36.745 64.815 37.625 ;
    RECT 61.215 76.365 61.495 77.245 ;
    RECT 57.895 76.365 58.175 77.245 ;
    RECT 54.575 76.365 54.855 77.245 ;
    RECT 51.255 76.365 51.535 77.245 ;
    RECT 47.935 76.365 48.215 77.245 ;
    RECT 44.615 76.365 44.895 77.245 ;
    RECT 41.295 76.365 41.575 77.245 ;
    RECT 37.975 76.365 38.255 77.245 ;
    RECT 34.655 76.365 34.935 77.245 ;
    RECT 117.655 76.365 117.935 77.245 ;
    RECT 114.335 76.365 114.615 77.245 ;
    RECT 111.015 76.365 111.295 77.245 ;
    RECT 107.695 76.365 107.975 77.245 ;
    RECT 104.375 76.365 104.655 77.245 ;
    RECT 101.055 76.365 101.335 77.245 ;
    RECT 97.735 76.365 98.015 77.245 ;
    RECT 94.415 76.365 94.695 77.245 ;
    RECT 91.095 76.365 91.375 77.245 ;
    RECT 87.775 76.365 88.055 77.245 ;
    RECT 84.455 76.365 84.735 77.245 ;
    RECT 81.135 76.365 81.415 77.245 ;
    RECT 77.815 76.365 78.095 77.245 ;
    RECT 74.495 76.365 74.775 77.245 ;
    RECT 71.175 76.365 71.455 77.245 ;
    RECT 31.335 76.365 31.615 77.245 ;
    RECT 67.855 76.365 68.135 77.245 ;
    RECT 28.015 76.365 28.295 77.245 ;
    RECT 24.695 76.365 24.975 77.245 ;
    RECT 21.375 76.365 21.655 77.245 ;
    RECT 18.055 76.365 18.335 77.245 ;
    RECT 14.735 76.365 15.015 77.245 ;
    RECT 11.415 76.365 11.695 77.245 ;
    RECT 8.095 76.365 8.375 77.245 ;
    RECT 4.775 76.365 5.055 77.245 ;
    RECT 1.455 76.365 1.735 77.245 ;
    RECT 64.535 76.365 64.815 77.245 ;
    RECT 61.215 36.025 61.495 36.905 ;
    RECT 57.895 36.025 58.175 36.905 ;
    RECT 54.575 36.025 54.855 36.905 ;
    RECT 51.255 36.025 51.535 36.905 ;
    RECT 47.935 36.025 48.215 36.905 ;
    RECT 44.615 36.025 44.895 36.905 ;
    RECT 41.295 36.025 41.575 36.905 ;
    RECT 37.975 36.025 38.255 36.905 ;
    RECT 34.655 36.025 34.935 36.905 ;
    RECT 117.655 36.025 117.935 36.905 ;
    RECT 114.335 36.025 114.615 36.905 ;
    RECT 111.015 36.025 111.295 36.905 ;
    RECT 107.695 36.025 107.975 36.905 ;
    RECT 104.375 36.025 104.655 36.905 ;
    RECT 101.055 36.025 101.335 36.905 ;
    RECT 97.735 36.025 98.015 36.905 ;
    RECT 94.415 36.025 94.695 36.905 ;
    RECT 91.095 36.025 91.375 36.905 ;
    RECT 87.775 36.025 88.055 36.905 ;
    RECT 84.455 36.025 84.735 36.905 ;
    RECT 81.135 36.025 81.415 36.905 ;
    RECT 77.815 36.025 78.095 36.905 ;
    RECT 74.495 36.025 74.775 36.905 ;
    RECT 71.175 36.025 71.455 36.905 ;
    RECT 31.335 36.025 31.615 36.905 ;
    RECT 67.855 36.025 68.135 36.905 ;
    RECT 28.015 36.025 28.295 36.905 ;
    RECT 24.695 36.025 24.975 36.905 ;
    RECT 21.375 36.025 21.655 36.905 ;
    RECT 18.055 36.025 18.335 36.905 ;
    RECT 14.735 36.025 15.015 36.905 ;
    RECT 11.415 36.025 11.695 36.905 ;
    RECT 8.095 36.025 8.375 36.905 ;
    RECT 4.775 36.025 5.055 36.905 ;
    RECT 1.455 36.025 1.735 36.905 ;
    RECT 64.535 36.025 64.815 36.905 ;
    RECT 61.215 75.645 61.495 76.525 ;
    RECT 57.895 75.645 58.175 76.525 ;
    RECT 54.575 75.645 54.855 76.525 ;
    RECT 51.255 75.645 51.535 76.525 ;
    RECT 47.935 75.645 48.215 76.525 ;
    RECT 44.615 75.645 44.895 76.525 ;
    RECT 41.295 75.645 41.575 76.525 ;
    RECT 37.975 75.645 38.255 76.525 ;
    RECT 34.655 75.645 34.935 76.525 ;
    RECT 117.655 75.645 117.935 76.525 ;
    RECT 114.335 75.645 114.615 76.525 ;
    RECT 111.015 75.645 111.295 76.525 ;
    RECT 107.695 75.645 107.975 76.525 ;
    RECT 104.375 75.645 104.655 76.525 ;
    RECT 101.055 75.645 101.335 76.525 ;
    RECT 97.735 75.645 98.015 76.525 ;
    RECT 94.415 75.645 94.695 76.525 ;
    RECT 91.095 75.645 91.375 76.525 ;
    RECT 87.775 75.645 88.055 76.525 ;
    RECT 84.455 75.645 84.735 76.525 ;
    RECT 81.135 75.645 81.415 76.525 ;
    RECT 77.815 75.645 78.095 76.525 ;
    RECT 74.495 75.645 74.775 76.525 ;
    RECT 71.175 75.645 71.455 76.525 ;
    RECT 31.335 75.645 31.615 76.525 ;
    RECT 67.855 75.645 68.135 76.525 ;
    RECT 28.015 75.645 28.295 76.525 ;
    RECT 24.695 75.645 24.975 76.525 ;
    RECT 21.375 75.645 21.655 76.525 ;
    RECT 18.055 75.645 18.335 76.525 ;
    RECT 14.735 75.645 15.015 76.525 ;
    RECT 11.415 75.645 11.695 76.525 ;
    RECT 8.095 75.645 8.375 76.525 ;
    RECT 4.775 75.645 5.055 76.525 ;
    RECT 1.455 75.645 1.735 76.525 ;
    RECT 64.535 75.645 64.815 76.525 ;
    RECT 61.215 74.925 61.495 75.805 ;
    RECT 57.895 74.925 58.175 75.805 ;
    RECT 54.575 74.925 54.855 75.805 ;
    RECT 51.255 74.925 51.535 75.805 ;
    RECT 47.935 74.925 48.215 75.805 ;
    RECT 44.615 74.925 44.895 75.805 ;
    RECT 41.295 74.925 41.575 75.805 ;
    RECT 37.975 74.925 38.255 75.805 ;
    RECT 34.655 74.925 34.935 75.805 ;
    RECT 117.655 74.925 117.935 75.805 ;
    RECT 114.335 74.925 114.615 75.805 ;
    RECT 111.015 74.925 111.295 75.805 ;
    RECT 107.695 74.925 107.975 75.805 ;
    RECT 104.375 74.925 104.655 75.805 ;
    RECT 101.055 74.925 101.335 75.805 ;
    RECT 97.735 74.925 98.015 75.805 ;
    RECT 94.415 74.925 94.695 75.805 ;
    RECT 91.095 74.925 91.375 75.805 ;
    RECT 87.775 74.925 88.055 75.805 ;
    RECT 84.455 74.925 84.735 75.805 ;
    RECT 81.135 74.925 81.415 75.805 ;
    RECT 77.815 74.925 78.095 75.805 ;
    RECT 74.495 74.925 74.775 75.805 ;
    RECT 71.175 74.925 71.455 75.805 ;
    RECT 31.335 74.925 31.615 75.805 ;
    RECT 67.855 74.925 68.135 75.805 ;
    RECT 28.015 74.925 28.295 75.805 ;
    RECT 24.695 74.925 24.975 75.805 ;
    RECT 21.375 74.925 21.655 75.805 ;
    RECT 18.055 74.925 18.335 75.805 ;
    RECT 14.735 74.925 15.015 75.805 ;
    RECT 11.415 74.925 11.695 75.805 ;
    RECT 8.095 74.925 8.375 75.805 ;
    RECT 4.775 74.925 5.055 75.805 ;
    RECT 1.455 74.925 1.735 75.805 ;
    RECT 64.535 74.925 64.815 75.805 ;
    RECT 61.215 74.205 61.495 75.085 ;
    RECT 57.895 74.205 58.175 75.085 ;
    RECT 54.575 74.205 54.855 75.085 ;
    RECT 51.255 74.205 51.535 75.085 ;
    RECT 47.935 74.205 48.215 75.085 ;
    RECT 44.615 74.205 44.895 75.085 ;
    RECT 41.295 74.205 41.575 75.085 ;
    RECT 37.975 74.205 38.255 75.085 ;
    RECT 34.655 74.205 34.935 75.085 ;
    RECT 117.655 74.205 117.935 75.085 ;
    RECT 114.335 74.205 114.615 75.085 ;
    RECT 111.015 74.205 111.295 75.085 ;
    RECT 107.695 74.205 107.975 75.085 ;
    RECT 104.375 74.205 104.655 75.085 ;
    RECT 101.055 74.205 101.335 75.085 ;
    RECT 97.735 74.205 98.015 75.085 ;
    RECT 94.415 74.205 94.695 75.085 ;
    RECT 91.095 74.205 91.375 75.085 ;
    RECT 87.775 74.205 88.055 75.085 ;
    RECT 84.455 74.205 84.735 75.085 ;
    RECT 81.135 74.205 81.415 75.085 ;
    RECT 77.815 74.205 78.095 75.085 ;
    RECT 74.495 74.205 74.775 75.085 ;
    RECT 71.175 74.205 71.455 75.085 ;
    RECT 31.335 74.205 31.615 75.085 ;
    RECT 67.855 74.205 68.135 75.085 ;
    RECT 28.015 74.205 28.295 75.085 ;
    RECT 24.695 74.205 24.975 75.085 ;
    RECT 21.375 74.205 21.655 75.085 ;
    RECT 18.055 74.205 18.335 75.085 ;
    RECT 14.735 74.205 15.015 75.085 ;
    RECT 11.415 74.205 11.695 75.085 ;
    RECT 8.095 74.205 8.375 75.085 ;
    RECT 4.775 74.205 5.055 75.085 ;
    RECT 1.455 74.205 1.735 75.085 ;
    RECT 64.535 74.205 64.815 75.085 ;
    RECT 61.215 73.485 61.495 74.365 ;
    RECT 57.895 73.485 58.175 74.365 ;
    RECT 54.575 73.485 54.855 74.365 ;
    RECT 51.255 73.485 51.535 74.365 ;
    RECT 47.935 73.485 48.215 74.365 ;
    RECT 44.615 73.485 44.895 74.365 ;
    RECT 41.295 73.485 41.575 74.365 ;
    RECT 37.975 73.485 38.255 74.365 ;
    RECT 34.655 73.485 34.935 74.365 ;
    RECT 117.655 73.485 117.935 74.365 ;
    RECT 114.335 73.485 114.615 74.365 ;
    RECT 111.015 73.485 111.295 74.365 ;
    RECT 107.695 73.485 107.975 74.365 ;
    RECT 104.375 73.485 104.655 74.365 ;
    RECT 101.055 73.485 101.335 74.365 ;
    RECT 97.735 73.485 98.015 74.365 ;
    RECT 94.415 73.485 94.695 74.365 ;
    RECT 91.095 73.485 91.375 74.365 ;
    RECT 87.775 73.485 88.055 74.365 ;
    RECT 84.455 73.485 84.735 74.365 ;
    RECT 81.135 73.485 81.415 74.365 ;
    RECT 77.815 73.485 78.095 74.365 ;
    RECT 74.495 73.485 74.775 74.365 ;
    RECT 71.175 73.485 71.455 74.365 ;
    RECT 31.335 73.485 31.615 74.365 ;
    RECT 67.855 73.485 68.135 74.365 ;
    RECT 28.015 73.485 28.295 74.365 ;
    RECT 24.695 73.485 24.975 74.365 ;
    RECT 21.375 73.485 21.655 74.365 ;
    RECT 18.055 73.485 18.335 74.365 ;
    RECT 14.735 73.485 15.015 74.365 ;
    RECT 11.415 73.485 11.695 74.365 ;
    RECT 8.095 73.485 8.375 74.365 ;
    RECT 4.775 73.485 5.055 74.365 ;
    RECT 1.455 73.485 1.735 74.365 ;
    RECT 64.535 73.485 64.815 74.365 ;
    RECT 61.215 72.765 61.495 73.645 ;
    RECT 57.895 72.765 58.175 73.645 ;
    RECT 54.575 72.765 54.855 73.645 ;
    RECT 51.255 72.765 51.535 73.645 ;
    RECT 47.935 72.765 48.215 73.645 ;
    RECT 44.615 72.765 44.895 73.645 ;
    RECT 41.295 72.765 41.575 73.645 ;
    RECT 37.975 72.765 38.255 73.645 ;
    RECT 34.655 72.765 34.935 73.645 ;
    RECT 117.655 72.765 117.935 73.645 ;
    RECT 114.335 72.765 114.615 73.645 ;
    RECT 111.015 72.765 111.295 73.645 ;
    RECT 107.695 72.765 107.975 73.645 ;
    RECT 104.375 72.765 104.655 73.645 ;
    RECT 101.055 72.765 101.335 73.645 ;
    RECT 97.735 72.765 98.015 73.645 ;
    RECT 94.415 72.765 94.695 73.645 ;
    RECT 91.095 72.765 91.375 73.645 ;
    RECT 87.775 72.765 88.055 73.645 ;
    RECT 84.455 72.765 84.735 73.645 ;
    RECT 81.135 72.765 81.415 73.645 ;
    RECT 77.815 72.765 78.095 73.645 ;
    RECT 74.495 72.765 74.775 73.645 ;
    RECT 71.175 72.765 71.455 73.645 ;
    RECT 31.335 72.765 31.615 73.645 ;
    RECT 67.855 72.765 68.135 73.645 ;
    RECT 28.015 72.765 28.295 73.645 ;
    RECT 24.695 72.765 24.975 73.645 ;
    RECT 21.375 72.765 21.655 73.645 ;
    RECT 18.055 72.765 18.335 73.645 ;
    RECT 14.735 72.765 15.015 73.645 ;
    RECT 11.415 72.765 11.695 73.645 ;
    RECT 8.095 72.765 8.375 73.645 ;
    RECT 4.775 72.765 5.055 73.645 ;
    RECT 1.455 72.765 1.735 73.645 ;
    RECT 64.535 72.765 64.815 73.645 ;
    RECT 61.215 35.305 61.495 36.185 ;
    RECT 57.895 35.305 58.175 36.185 ;
    RECT 54.575 35.305 54.855 36.185 ;
    RECT 51.255 35.305 51.535 36.185 ;
    RECT 47.935 35.305 48.215 36.185 ;
    RECT 44.615 35.305 44.895 36.185 ;
    RECT 41.295 35.305 41.575 36.185 ;
    RECT 37.975 35.305 38.255 36.185 ;
    RECT 34.655 35.305 34.935 36.185 ;
    RECT 117.655 35.305 117.935 36.185 ;
    RECT 114.335 35.305 114.615 36.185 ;
    RECT 111.015 35.305 111.295 36.185 ;
    RECT 107.695 35.305 107.975 36.185 ;
    RECT 104.375 35.305 104.655 36.185 ;
    RECT 101.055 35.305 101.335 36.185 ;
    RECT 97.735 35.305 98.015 36.185 ;
    RECT 94.415 35.305 94.695 36.185 ;
    RECT 91.095 35.305 91.375 36.185 ;
    RECT 87.775 35.305 88.055 36.185 ;
    RECT 84.455 35.305 84.735 36.185 ;
    RECT 81.135 35.305 81.415 36.185 ;
    RECT 77.815 35.305 78.095 36.185 ;
    RECT 74.495 35.305 74.775 36.185 ;
    RECT 71.175 35.305 71.455 36.185 ;
    RECT 31.335 35.305 31.615 36.185 ;
    RECT 67.855 35.305 68.135 36.185 ;
    RECT 28.015 35.305 28.295 36.185 ;
    RECT 24.695 35.305 24.975 36.185 ;
    RECT 21.375 35.305 21.655 36.185 ;
    RECT 18.055 35.305 18.335 36.185 ;
    RECT 14.735 35.305 15.015 36.185 ;
    RECT 11.415 35.305 11.695 36.185 ;
    RECT 8.095 35.305 8.375 36.185 ;
    RECT 4.775 35.305 5.055 36.185 ;
    RECT 1.455 35.305 1.735 36.185 ;
    RECT 64.535 35.305 64.815 36.185 ;
    RECT 61.215 34.585 61.495 35.465 ;
    RECT 57.895 34.585 58.175 35.465 ;
    RECT 54.575 34.585 54.855 35.465 ;
    RECT 51.255 34.585 51.535 35.465 ;
    RECT 47.935 34.585 48.215 35.465 ;
    RECT 44.615 34.585 44.895 35.465 ;
    RECT 41.295 34.585 41.575 35.465 ;
    RECT 37.975 34.585 38.255 35.465 ;
    RECT 34.655 34.585 34.935 35.465 ;
    RECT 117.655 34.585 117.935 35.465 ;
    RECT 114.335 34.585 114.615 35.465 ;
    RECT 111.015 34.585 111.295 35.465 ;
    RECT 107.695 34.585 107.975 35.465 ;
    RECT 104.375 34.585 104.655 35.465 ;
    RECT 101.055 34.585 101.335 35.465 ;
    RECT 97.735 34.585 98.015 35.465 ;
    RECT 94.415 34.585 94.695 35.465 ;
    RECT 91.095 34.585 91.375 35.465 ;
    RECT 87.775 34.585 88.055 35.465 ;
    RECT 84.455 34.585 84.735 35.465 ;
    RECT 81.135 34.585 81.415 35.465 ;
    RECT 77.815 34.585 78.095 35.465 ;
    RECT 74.495 34.585 74.775 35.465 ;
    RECT 71.175 34.585 71.455 35.465 ;
    RECT 31.335 34.585 31.615 35.465 ;
    RECT 67.855 34.585 68.135 35.465 ;
    RECT 28.015 34.585 28.295 35.465 ;
    RECT 24.695 34.585 24.975 35.465 ;
    RECT 21.375 34.585 21.655 35.465 ;
    RECT 18.055 34.585 18.335 35.465 ;
    RECT 14.735 34.585 15.015 35.465 ;
    RECT 11.415 34.585 11.695 35.465 ;
    RECT 8.095 34.585 8.375 35.465 ;
    RECT 4.775 34.585 5.055 35.465 ;
    RECT 1.455 34.585 1.735 35.465 ;
    RECT 64.535 34.585 64.815 35.465 ;
    RECT 61.215 33.865 61.495 34.745 ;
    RECT 57.895 33.865 58.175 34.745 ;
    RECT 54.575 33.865 54.855 34.745 ;
    RECT 51.255 33.865 51.535 34.745 ;
    RECT 47.935 33.865 48.215 34.745 ;
    RECT 44.615 33.865 44.895 34.745 ;
    RECT 41.295 33.865 41.575 34.745 ;
    RECT 37.975 33.865 38.255 34.745 ;
    RECT 34.655 33.865 34.935 34.745 ;
    RECT 117.655 33.865 117.935 34.745 ;
    RECT 114.335 33.865 114.615 34.745 ;
    RECT 111.015 33.865 111.295 34.745 ;
    RECT 107.695 33.865 107.975 34.745 ;
    RECT 104.375 33.865 104.655 34.745 ;
    RECT 101.055 33.865 101.335 34.745 ;
    RECT 97.735 33.865 98.015 34.745 ;
    RECT 94.415 33.865 94.695 34.745 ;
    RECT 91.095 33.865 91.375 34.745 ;
    RECT 87.775 33.865 88.055 34.745 ;
    RECT 84.455 33.865 84.735 34.745 ;
    RECT 81.135 33.865 81.415 34.745 ;
    RECT 77.815 33.865 78.095 34.745 ;
    RECT 74.495 33.865 74.775 34.745 ;
    RECT 71.175 33.865 71.455 34.745 ;
    RECT 31.335 33.865 31.615 34.745 ;
    RECT 67.855 33.865 68.135 34.745 ;
    RECT 28.015 33.865 28.295 34.745 ;
    RECT 24.695 33.865 24.975 34.745 ;
    RECT 21.375 33.865 21.655 34.745 ;
    RECT 18.055 33.865 18.335 34.745 ;
    RECT 14.735 33.865 15.015 34.745 ;
    RECT 11.415 33.865 11.695 34.745 ;
    RECT 8.095 33.865 8.375 34.745 ;
    RECT 4.775 33.865 5.055 34.745 ;
    RECT 1.455 33.865 1.735 34.745 ;
    RECT 64.535 33.865 64.815 34.745 ;
    RECT 61.215 33.145 61.495 34.025 ;
    RECT 57.895 33.145 58.175 34.025 ;
    RECT 54.575 33.145 54.855 34.025 ;
    RECT 51.255 33.145 51.535 34.025 ;
    RECT 47.935 33.145 48.215 34.025 ;
    RECT 44.615 33.145 44.895 34.025 ;
    RECT 41.295 33.145 41.575 34.025 ;
    RECT 37.975 33.145 38.255 34.025 ;
    RECT 34.655 33.145 34.935 34.025 ;
    RECT 117.655 33.145 117.935 34.025 ;
    RECT 114.335 33.145 114.615 34.025 ;
    RECT 111.015 33.145 111.295 34.025 ;
    RECT 107.695 33.145 107.975 34.025 ;
    RECT 104.375 33.145 104.655 34.025 ;
    RECT 101.055 33.145 101.335 34.025 ;
    RECT 97.735 33.145 98.015 34.025 ;
    RECT 94.415 33.145 94.695 34.025 ;
    RECT 91.095 33.145 91.375 34.025 ;
    RECT 87.775 33.145 88.055 34.025 ;
    RECT 84.455 33.145 84.735 34.025 ;
    RECT 81.135 33.145 81.415 34.025 ;
    RECT 77.815 33.145 78.095 34.025 ;
    RECT 74.495 33.145 74.775 34.025 ;
    RECT 71.175 33.145 71.455 34.025 ;
    RECT 31.335 33.145 31.615 34.025 ;
    RECT 67.855 33.145 68.135 34.025 ;
    RECT 28.015 33.145 28.295 34.025 ;
    RECT 24.695 33.145 24.975 34.025 ;
    RECT 21.375 33.145 21.655 34.025 ;
    RECT 18.055 33.145 18.335 34.025 ;
    RECT 14.735 33.145 15.015 34.025 ;
    RECT 11.415 33.145 11.695 34.025 ;
    RECT 8.095 33.145 8.375 34.025 ;
    RECT 4.775 33.145 5.055 34.025 ;
    RECT 1.455 33.145 1.735 34.025 ;
    RECT 64.535 33.145 64.815 34.025 ;
    RECT 61.215 32.425 61.495 33.305 ;
    RECT 57.895 32.425 58.175 33.305 ;
    RECT 54.575 32.425 54.855 33.305 ;
    RECT 51.255 32.425 51.535 33.305 ;
    RECT 47.935 32.425 48.215 33.305 ;
    RECT 44.615 32.425 44.895 33.305 ;
    RECT 41.295 32.425 41.575 33.305 ;
    RECT 37.975 32.425 38.255 33.305 ;
    RECT 34.655 32.425 34.935 33.305 ;
    RECT 117.655 32.425 117.935 33.305 ;
    RECT 114.335 32.425 114.615 33.305 ;
    RECT 111.015 32.425 111.295 33.305 ;
    RECT 107.695 32.425 107.975 33.305 ;
    RECT 104.375 32.425 104.655 33.305 ;
    RECT 101.055 32.425 101.335 33.305 ;
    RECT 97.735 32.425 98.015 33.305 ;
    RECT 94.415 32.425 94.695 33.305 ;
    RECT 91.095 32.425 91.375 33.305 ;
    RECT 87.775 32.425 88.055 33.305 ;
    RECT 84.455 32.425 84.735 33.305 ;
    RECT 81.135 32.425 81.415 33.305 ;
    RECT 77.815 32.425 78.095 33.305 ;
    RECT 74.495 32.425 74.775 33.305 ;
    RECT 71.175 32.425 71.455 33.305 ;
    RECT 31.335 32.425 31.615 33.305 ;
    RECT 67.855 32.425 68.135 33.305 ;
    RECT 28.015 32.425 28.295 33.305 ;
    RECT 24.695 32.425 24.975 33.305 ;
    RECT 21.375 32.425 21.655 33.305 ;
    RECT 18.055 32.425 18.335 33.305 ;
    RECT 14.735 32.425 15.015 33.305 ;
    RECT 11.415 32.425 11.695 33.305 ;
    RECT 8.095 32.425 8.375 33.305 ;
    RECT 4.775 32.425 5.055 33.305 ;
    RECT 1.455 32.425 1.735 33.305 ;
    RECT 64.535 32.425 64.815 33.305 ;
    RECT 61.215 72.045 61.495 72.925 ;
    RECT 57.895 72.045 58.175 72.925 ;
    RECT 54.575 72.045 54.855 72.925 ;
    RECT 51.255 72.045 51.535 72.925 ;
    RECT 47.935 72.045 48.215 72.925 ;
    RECT 44.615 72.045 44.895 72.925 ;
    RECT 41.295 72.045 41.575 72.925 ;
    RECT 37.975 72.045 38.255 72.925 ;
    RECT 34.655 72.045 34.935 72.925 ;
    RECT 117.655 72.045 117.935 72.925 ;
    RECT 114.335 72.045 114.615 72.925 ;
    RECT 111.015 72.045 111.295 72.925 ;
    RECT 107.695 72.045 107.975 72.925 ;
    RECT 104.375 72.045 104.655 72.925 ;
    RECT 101.055 72.045 101.335 72.925 ;
    RECT 97.735 72.045 98.015 72.925 ;
    RECT 94.415 72.045 94.695 72.925 ;
    RECT 91.095 72.045 91.375 72.925 ;
    RECT 87.775 72.045 88.055 72.925 ;
    RECT 84.455 72.045 84.735 72.925 ;
    RECT 81.135 72.045 81.415 72.925 ;
    RECT 77.815 72.045 78.095 72.925 ;
    RECT 74.495 72.045 74.775 72.925 ;
    RECT 71.175 72.045 71.455 72.925 ;
    RECT 31.335 72.045 31.615 72.925 ;
    RECT 67.855 72.045 68.135 72.925 ;
    RECT 28.015 72.045 28.295 72.925 ;
    RECT 24.695 72.045 24.975 72.925 ;
    RECT 21.375 72.045 21.655 72.925 ;
    RECT 18.055 72.045 18.335 72.925 ;
    RECT 14.735 72.045 15.015 72.925 ;
    RECT 11.415 72.045 11.695 72.925 ;
    RECT 8.095 72.045 8.375 72.925 ;
    RECT 4.775 72.045 5.055 72.925 ;
    RECT 1.455 72.045 1.735 72.925 ;
    RECT 64.535 72.045 64.815 72.925 ;
    RECT 61.215 31.705 61.495 32.585 ;
    RECT 57.895 31.705 58.175 32.585 ;
    RECT 54.575 31.705 54.855 32.585 ;
    RECT 51.255 31.705 51.535 32.585 ;
    RECT 47.935 31.705 48.215 32.585 ;
    RECT 44.615 31.705 44.895 32.585 ;
    RECT 41.295 31.705 41.575 32.585 ;
    RECT 37.975 31.705 38.255 32.585 ;
    RECT 34.655 31.705 34.935 32.585 ;
    RECT 117.655 31.705 117.935 32.585 ;
    RECT 114.335 31.705 114.615 32.585 ;
    RECT 111.015 31.705 111.295 32.585 ;
    RECT 107.695 31.705 107.975 32.585 ;
    RECT 104.375 31.705 104.655 32.585 ;
    RECT 101.055 31.705 101.335 32.585 ;
    RECT 97.735 31.705 98.015 32.585 ;
    RECT 94.415 31.705 94.695 32.585 ;
    RECT 91.095 31.705 91.375 32.585 ;
    RECT 87.775 31.705 88.055 32.585 ;
    RECT 84.455 31.705 84.735 32.585 ;
    RECT 81.135 31.705 81.415 32.585 ;
    RECT 77.815 31.705 78.095 32.585 ;
    RECT 74.495 31.705 74.775 32.585 ;
    RECT 71.175 31.705 71.455 32.585 ;
    RECT 31.335 31.705 31.615 32.585 ;
    RECT 67.855 31.705 68.135 32.585 ;
    RECT 28.015 31.705 28.295 32.585 ;
    RECT 24.695 31.705 24.975 32.585 ;
    RECT 21.375 31.705 21.655 32.585 ;
    RECT 18.055 31.705 18.335 32.585 ;
    RECT 14.735 31.705 15.015 32.585 ;
    RECT 11.415 31.705 11.695 32.585 ;
    RECT 8.095 31.705 8.375 32.585 ;
    RECT 4.775 31.705 5.055 32.585 ;
    RECT 1.455 31.705 1.735 32.585 ;
    RECT 64.535 31.705 64.815 32.585 ;
    RECT 61.215 71.325 61.495 72.205 ;
    RECT 57.895 71.325 58.175 72.205 ;
    RECT 54.575 71.325 54.855 72.205 ;
    RECT 51.255 71.325 51.535 72.205 ;
    RECT 47.935 71.325 48.215 72.205 ;
    RECT 44.615 71.325 44.895 72.205 ;
    RECT 41.295 71.325 41.575 72.205 ;
    RECT 37.975 71.325 38.255 72.205 ;
    RECT 34.655 71.325 34.935 72.205 ;
    RECT 117.655 71.325 117.935 72.205 ;
    RECT 114.335 71.325 114.615 72.205 ;
    RECT 111.015 71.325 111.295 72.205 ;
    RECT 107.695 71.325 107.975 72.205 ;
    RECT 104.375 71.325 104.655 72.205 ;
    RECT 101.055 71.325 101.335 72.205 ;
    RECT 97.735 71.325 98.015 72.205 ;
    RECT 94.415 71.325 94.695 72.205 ;
    RECT 91.095 71.325 91.375 72.205 ;
    RECT 87.775 71.325 88.055 72.205 ;
    RECT 84.455 71.325 84.735 72.205 ;
    RECT 81.135 71.325 81.415 72.205 ;
    RECT 77.815 71.325 78.095 72.205 ;
    RECT 74.495 71.325 74.775 72.205 ;
    RECT 71.175 71.325 71.455 72.205 ;
    RECT 31.335 71.325 31.615 72.205 ;
    RECT 67.855 71.325 68.135 72.205 ;
    RECT 28.015 71.325 28.295 72.205 ;
    RECT 24.695 71.325 24.975 72.205 ;
    RECT 21.375 71.325 21.655 72.205 ;
    RECT 18.055 71.325 18.335 72.205 ;
    RECT 14.735 71.325 15.015 72.205 ;
    RECT 11.415 71.325 11.695 72.205 ;
    RECT 8.095 71.325 8.375 72.205 ;
    RECT 4.775 71.325 5.055 72.205 ;
    RECT 1.455 71.325 1.735 72.205 ;
    RECT 64.535 71.325 64.815 72.205 ;
    RECT 61.215 30.985 61.495 31.865 ;
    RECT 57.895 30.985 58.175 31.865 ;
    RECT 54.575 30.985 54.855 31.865 ;
    RECT 51.255 30.985 51.535 31.865 ;
    RECT 47.935 30.985 48.215 31.865 ;
    RECT 44.615 30.985 44.895 31.865 ;
    RECT 41.295 30.985 41.575 31.865 ;
    RECT 37.975 30.985 38.255 31.865 ;
    RECT 34.655 30.985 34.935 31.865 ;
    RECT 117.655 30.985 117.935 31.865 ;
    RECT 114.335 30.985 114.615 31.865 ;
    RECT 111.015 30.985 111.295 31.865 ;
    RECT 107.695 30.985 107.975 31.865 ;
    RECT 104.375 30.985 104.655 31.865 ;
    RECT 101.055 30.985 101.335 31.865 ;
    RECT 97.735 30.985 98.015 31.865 ;
    RECT 94.415 30.985 94.695 31.865 ;
    RECT 91.095 30.985 91.375 31.865 ;
    RECT 87.775 30.985 88.055 31.865 ;
    RECT 84.455 30.985 84.735 31.865 ;
    RECT 81.135 30.985 81.415 31.865 ;
    RECT 77.815 30.985 78.095 31.865 ;
    RECT 74.495 30.985 74.775 31.865 ;
    RECT 71.175 30.985 71.455 31.865 ;
    RECT 31.335 30.985 31.615 31.865 ;
    RECT 67.855 30.985 68.135 31.865 ;
    RECT 28.015 30.985 28.295 31.865 ;
    RECT 24.695 30.985 24.975 31.865 ;
    RECT 21.375 30.985 21.655 31.865 ;
    RECT 18.055 30.985 18.335 31.865 ;
    RECT 14.735 30.985 15.015 31.865 ;
    RECT 11.415 30.985 11.695 31.865 ;
    RECT 8.095 30.985 8.375 31.865 ;
    RECT 4.775 30.985 5.055 31.865 ;
    RECT 1.455 30.985 1.735 31.865 ;
    RECT 64.535 30.985 64.815 31.865 ;
    RECT 61.215 70.605 61.495 71.485 ;
    RECT 57.895 70.605 58.175 71.485 ;
    RECT 54.575 70.605 54.855 71.485 ;
    RECT 51.255 70.605 51.535 71.485 ;
    RECT 47.935 70.605 48.215 71.485 ;
    RECT 44.615 70.605 44.895 71.485 ;
    RECT 41.295 70.605 41.575 71.485 ;
    RECT 37.975 70.605 38.255 71.485 ;
    RECT 34.655 70.605 34.935 71.485 ;
    RECT 117.655 70.605 117.935 71.485 ;
    RECT 114.335 70.605 114.615 71.485 ;
    RECT 111.015 70.605 111.295 71.485 ;
    RECT 107.695 70.605 107.975 71.485 ;
    RECT 104.375 70.605 104.655 71.485 ;
    RECT 101.055 70.605 101.335 71.485 ;
    RECT 97.735 70.605 98.015 71.485 ;
    RECT 94.415 70.605 94.695 71.485 ;
    RECT 91.095 70.605 91.375 71.485 ;
    RECT 87.775 70.605 88.055 71.485 ;
    RECT 84.455 70.605 84.735 71.485 ;
    RECT 81.135 70.605 81.415 71.485 ;
    RECT 77.815 70.605 78.095 71.485 ;
    RECT 74.495 70.605 74.775 71.485 ;
    RECT 71.175 70.605 71.455 71.485 ;
    RECT 31.335 70.605 31.615 71.485 ;
    RECT 67.855 70.605 68.135 71.485 ;
    RECT 28.015 70.605 28.295 71.485 ;
    RECT 24.695 70.605 24.975 71.485 ;
    RECT 21.375 70.605 21.655 71.485 ;
    RECT 18.055 70.605 18.335 71.485 ;
    RECT 14.735 70.605 15.015 71.485 ;
    RECT 11.415 70.605 11.695 71.485 ;
    RECT 8.095 70.605 8.375 71.485 ;
    RECT 4.775 70.605 5.055 71.485 ;
    RECT 1.455 70.605 1.735 71.485 ;
    RECT 64.535 70.605 64.815 71.485 ;
    RECT 61.215 30.265 61.495 31.145 ;
    RECT 57.895 30.265 58.175 31.145 ;
    RECT 54.575 30.265 54.855 31.145 ;
    RECT 51.255 30.265 51.535 31.145 ;
    RECT 47.935 30.265 48.215 31.145 ;
    RECT 44.615 30.265 44.895 31.145 ;
    RECT 41.295 30.265 41.575 31.145 ;
    RECT 37.975 30.265 38.255 31.145 ;
    RECT 34.655 30.265 34.935 31.145 ;
    RECT 117.655 30.265 117.935 31.145 ;
    RECT 114.335 30.265 114.615 31.145 ;
    RECT 111.015 30.265 111.295 31.145 ;
    RECT 107.695 30.265 107.975 31.145 ;
    RECT 104.375 30.265 104.655 31.145 ;
    RECT 101.055 30.265 101.335 31.145 ;
    RECT 97.735 30.265 98.015 31.145 ;
    RECT 94.415 30.265 94.695 31.145 ;
    RECT 91.095 30.265 91.375 31.145 ;
    RECT 87.775 30.265 88.055 31.145 ;
    RECT 84.455 30.265 84.735 31.145 ;
    RECT 81.135 30.265 81.415 31.145 ;
    RECT 77.815 30.265 78.095 31.145 ;
    RECT 74.495 30.265 74.775 31.145 ;
    RECT 71.175 30.265 71.455 31.145 ;
    RECT 31.335 30.265 31.615 31.145 ;
    RECT 67.855 30.265 68.135 31.145 ;
    RECT 28.015 30.265 28.295 31.145 ;
    RECT 24.695 30.265 24.975 31.145 ;
    RECT 21.375 30.265 21.655 31.145 ;
    RECT 18.055 30.265 18.335 31.145 ;
    RECT 14.735 30.265 15.015 31.145 ;
    RECT 11.415 30.265 11.695 31.145 ;
    RECT 8.095 30.265 8.375 31.145 ;
    RECT 4.775 30.265 5.055 31.145 ;
    RECT 1.455 30.265 1.735 31.145 ;
    RECT 64.535 30.265 64.815 31.145 ;
    RECT 61.215 69.885 61.495 70.765 ;
    RECT 57.895 69.885 58.175 70.765 ;
    RECT 54.575 69.885 54.855 70.765 ;
    RECT 51.255 69.885 51.535 70.765 ;
    RECT 47.935 69.885 48.215 70.765 ;
    RECT 44.615 69.885 44.895 70.765 ;
    RECT 41.295 69.885 41.575 70.765 ;
    RECT 37.975 69.885 38.255 70.765 ;
    RECT 34.655 69.885 34.935 70.765 ;
    RECT 117.655 69.885 117.935 70.765 ;
    RECT 114.335 69.885 114.615 70.765 ;
    RECT 111.015 69.885 111.295 70.765 ;
    RECT 107.695 69.885 107.975 70.765 ;
    RECT 104.375 69.885 104.655 70.765 ;
    RECT 101.055 69.885 101.335 70.765 ;
    RECT 97.735 69.885 98.015 70.765 ;
    RECT 94.415 69.885 94.695 70.765 ;
    RECT 91.095 69.885 91.375 70.765 ;
    RECT 87.775 69.885 88.055 70.765 ;
    RECT 84.455 69.885 84.735 70.765 ;
    RECT 81.135 69.885 81.415 70.765 ;
    RECT 77.815 69.885 78.095 70.765 ;
    RECT 74.495 69.885 74.775 70.765 ;
    RECT 71.175 69.885 71.455 70.765 ;
    RECT 31.335 69.885 31.615 70.765 ;
    RECT 67.855 69.885 68.135 70.765 ;
    RECT 28.015 69.885 28.295 70.765 ;
    RECT 24.695 69.885 24.975 70.765 ;
    RECT 21.375 69.885 21.655 70.765 ;
    RECT 18.055 69.885 18.335 70.765 ;
    RECT 14.735 69.885 15.015 70.765 ;
    RECT 11.415 69.885 11.695 70.765 ;
    RECT 8.095 69.885 8.375 70.765 ;
    RECT 4.775 69.885 5.055 70.765 ;
    RECT 1.455 69.885 1.735 70.765 ;
    RECT 64.535 69.885 64.815 70.765 ;
    RECT 61.215 29.545 61.495 30.425 ;
    RECT 57.895 29.545 58.175 30.425 ;
    RECT 54.575 29.545 54.855 30.425 ;
    RECT 51.255 29.545 51.535 30.425 ;
    RECT 47.935 29.545 48.215 30.425 ;
    RECT 44.615 29.545 44.895 30.425 ;
    RECT 41.295 29.545 41.575 30.425 ;
    RECT 37.975 29.545 38.255 30.425 ;
    RECT 34.655 29.545 34.935 30.425 ;
    RECT 117.655 29.545 117.935 30.425 ;
    RECT 114.335 29.545 114.615 30.425 ;
    RECT 111.015 29.545 111.295 30.425 ;
    RECT 107.695 29.545 107.975 30.425 ;
    RECT 104.375 29.545 104.655 30.425 ;
    RECT 101.055 29.545 101.335 30.425 ;
    RECT 97.735 29.545 98.015 30.425 ;
    RECT 94.415 29.545 94.695 30.425 ;
    RECT 91.095 29.545 91.375 30.425 ;
    RECT 87.775 29.545 88.055 30.425 ;
    RECT 84.455 29.545 84.735 30.425 ;
    RECT 81.135 29.545 81.415 30.425 ;
    RECT 77.815 29.545 78.095 30.425 ;
    RECT 74.495 29.545 74.775 30.425 ;
    RECT 71.175 29.545 71.455 30.425 ;
    RECT 31.335 29.545 31.615 30.425 ;
    RECT 67.855 29.545 68.135 30.425 ;
    RECT 28.015 29.545 28.295 30.425 ;
    RECT 24.695 29.545 24.975 30.425 ;
    RECT 21.375 29.545 21.655 30.425 ;
    RECT 18.055 29.545 18.335 30.425 ;
    RECT 14.735 29.545 15.015 30.425 ;
    RECT 11.415 29.545 11.695 30.425 ;
    RECT 8.095 29.545 8.375 30.425 ;
    RECT 4.775 29.545 5.055 30.425 ;
    RECT 1.455 29.545 1.735 30.425 ;
    RECT 64.535 29.545 64.815 30.425 ;
    RECT 61.215 69.165 61.495 70.045 ;
    RECT 57.895 69.165 58.175 70.045 ;
    RECT 54.575 69.165 54.855 70.045 ;
    RECT 51.255 69.165 51.535 70.045 ;
    RECT 47.935 69.165 48.215 70.045 ;
    RECT 44.615 69.165 44.895 70.045 ;
    RECT 41.295 69.165 41.575 70.045 ;
    RECT 37.975 69.165 38.255 70.045 ;
    RECT 34.655 69.165 34.935 70.045 ;
    RECT 117.655 69.165 117.935 70.045 ;
    RECT 114.335 69.165 114.615 70.045 ;
    RECT 111.015 69.165 111.295 70.045 ;
    RECT 107.695 69.165 107.975 70.045 ;
    RECT 104.375 69.165 104.655 70.045 ;
    RECT 101.055 69.165 101.335 70.045 ;
    RECT 97.735 69.165 98.015 70.045 ;
    RECT 94.415 69.165 94.695 70.045 ;
    RECT 91.095 69.165 91.375 70.045 ;
    RECT 87.775 69.165 88.055 70.045 ;
    RECT 84.455 69.165 84.735 70.045 ;
    RECT 81.135 69.165 81.415 70.045 ;
    RECT 77.815 69.165 78.095 70.045 ;
    RECT 74.495 69.165 74.775 70.045 ;
    RECT 71.175 69.165 71.455 70.045 ;
    RECT 31.335 69.165 31.615 70.045 ;
    RECT 67.855 69.165 68.135 70.045 ;
    RECT 28.015 69.165 28.295 70.045 ;
    RECT 24.695 69.165 24.975 70.045 ;
    RECT 21.375 69.165 21.655 70.045 ;
    RECT 18.055 69.165 18.335 70.045 ;
    RECT 14.735 69.165 15.015 70.045 ;
    RECT 11.415 69.165 11.695 70.045 ;
    RECT 8.095 69.165 8.375 70.045 ;
    RECT 4.775 69.165 5.055 70.045 ;
    RECT 1.455 69.165 1.735 70.045 ;
    RECT 64.535 69.165 64.815 70.045 ;
    RECT 61.215 28.825 61.495 29.705 ;
    RECT 57.895 28.825 58.175 29.705 ;
    RECT 54.575 28.825 54.855 29.705 ;
    RECT 51.255 28.825 51.535 29.705 ;
    RECT 47.935 28.825 48.215 29.705 ;
    RECT 44.615 28.825 44.895 29.705 ;
    RECT 41.295 28.825 41.575 29.705 ;
    RECT 37.975 28.825 38.255 29.705 ;
    RECT 34.655 28.825 34.935 29.705 ;
    RECT 117.655 28.825 117.935 29.705 ;
    RECT 114.335 28.825 114.615 29.705 ;
    RECT 111.015 28.825 111.295 29.705 ;
    RECT 107.695 28.825 107.975 29.705 ;
    RECT 104.375 28.825 104.655 29.705 ;
    RECT 101.055 28.825 101.335 29.705 ;
    RECT 97.735 28.825 98.015 29.705 ;
    RECT 94.415 28.825 94.695 29.705 ;
    RECT 91.095 28.825 91.375 29.705 ;
    RECT 87.775 28.825 88.055 29.705 ;
    RECT 84.455 28.825 84.735 29.705 ;
    RECT 81.135 28.825 81.415 29.705 ;
    RECT 77.815 28.825 78.095 29.705 ;
    RECT 74.495 28.825 74.775 29.705 ;
    RECT 71.175 28.825 71.455 29.705 ;
    RECT 31.335 28.825 31.615 29.705 ;
    RECT 67.855 28.825 68.135 29.705 ;
    RECT 28.015 28.825 28.295 29.705 ;
    RECT 24.695 28.825 24.975 29.705 ;
    RECT 21.375 28.825 21.655 29.705 ;
    RECT 18.055 28.825 18.335 29.705 ;
    RECT 14.735 28.825 15.015 29.705 ;
    RECT 11.415 28.825 11.695 29.705 ;
    RECT 8.095 28.825 8.375 29.705 ;
    RECT 4.775 28.825 5.055 29.705 ;
    RECT 1.455 28.825 1.735 29.705 ;
    RECT 64.535 28.825 64.815 29.705 ;
    RECT 61.215 68.445 61.495 69.325 ;
    RECT 57.895 68.445 58.175 69.325 ;
    RECT 54.575 68.445 54.855 69.325 ;
    RECT 51.255 68.445 51.535 69.325 ;
    RECT 47.935 68.445 48.215 69.325 ;
    RECT 44.615 68.445 44.895 69.325 ;
    RECT 41.295 68.445 41.575 69.325 ;
    RECT 37.975 68.445 38.255 69.325 ;
    RECT 34.655 68.445 34.935 69.325 ;
    RECT 117.655 68.445 117.935 69.325 ;
    RECT 114.335 68.445 114.615 69.325 ;
    RECT 111.015 68.445 111.295 69.325 ;
    RECT 107.695 68.445 107.975 69.325 ;
    RECT 104.375 68.445 104.655 69.325 ;
    RECT 101.055 68.445 101.335 69.325 ;
    RECT 97.735 68.445 98.015 69.325 ;
    RECT 94.415 68.445 94.695 69.325 ;
    RECT 91.095 68.445 91.375 69.325 ;
    RECT 87.775 68.445 88.055 69.325 ;
    RECT 84.455 68.445 84.735 69.325 ;
    RECT 81.135 68.445 81.415 69.325 ;
    RECT 77.815 68.445 78.095 69.325 ;
    RECT 74.495 68.445 74.775 69.325 ;
    RECT 71.175 68.445 71.455 69.325 ;
    RECT 31.335 68.445 31.615 69.325 ;
    RECT 67.855 68.445 68.135 69.325 ;
    RECT 28.015 68.445 28.295 69.325 ;
    RECT 24.695 68.445 24.975 69.325 ;
    RECT 21.375 68.445 21.655 69.325 ;
    RECT 18.055 68.445 18.335 69.325 ;
    RECT 14.735 68.445 15.015 69.325 ;
    RECT 11.415 68.445 11.695 69.325 ;
    RECT 8.095 68.445 8.375 69.325 ;
    RECT 4.775 68.445 5.055 69.325 ;
    RECT 1.455 68.445 1.735 69.325 ;
    RECT 64.535 68.445 64.815 69.325 ;
    RECT 61.215 67.725 61.495 68.605 ;
    RECT 57.895 67.725 58.175 68.605 ;
    RECT 54.575 67.725 54.855 68.605 ;
    RECT 51.255 67.725 51.535 68.605 ;
    RECT 47.935 67.725 48.215 68.605 ;
    RECT 44.615 67.725 44.895 68.605 ;
    RECT 41.295 67.725 41.575 68.605 ;
    RECT 37.975 67.725 38.255 68.605 ;
    RECT 34.655 67.725 34.935 68.605 ;
    RECT 117.655 67.725 117.935 68.605 ;
    RECT 114.335 67.725 114.615 68.605 ;
    RECT 111.015 67.725 111.295 68.605 ;
    RECT 107.695 67.725 107.975 68.605 ;
    RECT 104.375 67.725 104.655 68.605 ;
    RECT 101.055 67.725 101.335 68.605 ;
    RECT 97.735 67.725 98.015 68.605 ;
    RECT 94.415 67.725 94.695 68.605 ;
    RECT 91.095 67.725 91.375 68.605 ;
    RECT 87.775 67.725 88.055 68.605 ;
    RECT 84.455 67.725 84.735 68.605 ;
    RECT 81.135 67.725 81.415 68.605 ;
    RECT 77.815 67.725 78.095 68.605 ;
    RECT 74.495 67.725 74.775 68.605 ;
    RECT 71.175 67.725 71.455 68.605 ;
    RECT 31.335 67.725 31.615 68.605 ;
    RECT 67.855 67.725 68.135 68.605 ;
    RECT 28.015 67.725 28.295 68.605 ;
    RECT 24.695 67.725 24.975 68.605 ;
    RECT 21.375 67.725 21.655 68.605 ;
    RECT 18.055 67.725 18.335 68.605 ;
    RECT 14.735 67.725 15.015 68.605 ;
    RECT 11.415 67.725 11.695 68.605 ;
    RECT 8.095 67.725 8.375 68.605 ;
    RECT 4.775 67.725 5.055 68.605 ;
    RECT 1.455 67.725 1.735 68.605 ;
    RECT 64.535 67.725 64.815 68.605 ;
    RECT 61.215 67.005 61.495 67.885 ;
    RECT 57.895 67.005 58.175 67.885 ;
    RECT 54.575 67.005 54.855 67.885 ;
    RECT 51.255 67.005 51.535 67.885 ;
    RECT 47.935 67.005 48.215 67.885 ;
    RECT 44.615 67.005 44.895 67.885 ;
    RECT 41.295 67.005 41.575 67.885 ;
    RECT 37.975 67.005 38.255 67.885 ;
    RECT 34.655 67.005 34.935 67.885 ;
    RECT 117.655 67.005 117.935 67.885 ;
    RECT 114.335 67.005 114.615 67.885 ;
    RECT 111.015 67.005 111.295 67.885 ;
    RECT 107.695 67.005 107.975 67.885 ;
    RECT 104.375 67.005 104.655 67.885 ;
    RECT 101.055 67.005 101.335 67.885 ;
    RECT 97.735 67.005 98.015 67.885 ;
    RECT 94.415 67.005 94.695 67.885 ;
    RECT 91.095 67.005 91.375 67.885 ;
    RECT 87.775 67.005 88.055 67.885 ;
    RECT 84.455 67.005 84.735 67.885 ;
    RECT 81.135 67.005 81.415 67.885 ;
    RECT 77.815 67.005 78.095 67.885 ;
    RECT 74.495 67.005 74.775 67.885 ;
    RECT 71.175 67.005 71.455 67.885 ;
    RECT 31.335 67.005 31.615 67.885 ;
    RECT 67.855 67.005 68.135 67.885 ;
    RECT 28.015 67.005 28.295 67.885 ;
    RECT 24.695 67.005 24.975 67.885 ;
    RECT 21.375 67.005 21.655 67.885 ;
    RECT 18.055 67.005 18.335 67.885 ;
    RECT 14.735 67.005 15.015 67.885 ;
    RECT 11.415 67.005 11.695 67.885 ;
    RECT 8.095 67.005 8.375 67.885 ;
    RECT 4.775 67.005 5.055 67.885 ;
    RECT 1.455 67.005 1.735 67.885 ;
    RECT 64.535 67.005 64.815 67.885 ;
    RECT 61.215 66.285 61.495 67.165 ;
    RECT 57.895 66.285 58.175 67.165 ;
    RECT 54.575 66.285 54.855 67.165 ;
    RECT 51.255 66.285 51.535 67.165 ;
    RECT 47.935 66.285 48.215 67.165 ;
    RECT 44.615 66.285 44.895 67.165 ;
    RECT 41.295 66.285 41.575 67.165 ;
    RECT 37.975 66.285 38.255 67.165 ;
    RECT 34.655 66.285 34.935 67.165 ;
    RECT 117.655 66.285 117.935 67.165 ;
    RECT 114.335 66.285 114.615 67.165 ;
    RECT 111.015 66.285 111.295 67.165 ;
    RECT 107.695 66.285 107.975 67.165 ;
    RECT 104.375 66.285 104.655 67.165 ;
    RECT 101.055 66.285 101.335 67.165 ;
    RECT 97.735 66.285 98.015 67.165 ;
    RECT 94.415 66.285 94.695 67.165 ;
    RECT 91.095 66.285 91.375 67.165 ;
    RECT 87.775 66.285 88.055 67.165 ;
    RECT 84.455 66.285 84.735 67.165 ;
    RECT 81.135 66.285 81.415 67.165 ;
    RECT 77.815 66.285 78.095 67.165 ;
    RECT 74.495 66.285 74.775 67.165 ;
    RECT 71.175 66.285 71.455 67.165 ;
    RECT 31.335 66.285 31.615 67.165 ;
    RECT 67.855 66.285 68.135 67.165 ;
    RECT 28.015 66.285 28.295 67.165 ;
    RECT 24.695 66.285 24.975 67.165 ;
    RECT 21.375 66.285 21.655 67.165 ;
    RECT 18.055 66.285 18.335 67.165 ;
    RECT 14.735 66.285 15.015 67.165 ;
    RECT 11.415 66.285 11.695 67.165 ;
    RECT 8.095 66.285 8.375 67.165 ;
    RECT 4.775 66.285 5.055 67.165 ;
    RECT 1.455 66.285 1.735 67.165 ;
    RECT 64.535 66.285 64.815 67.165 ;
    RECT 61.215 65.565 61.495 66.445 ;
    RECT 57.895 65.565 58.175 66.445 ;
    RECT 54.575 65.565 54.855 66.445 ;
    RECT 51.255 65.565 51.535 66.445 ;
    RECT 47.935 65.565 48.215 66.445 ;
    RECT 44.615 65.565 44.895 66.445 ;
    RECT 41.295 65.565 41.575 66.445 ;
    RECT 37.975 65.565 38.255 66.445 ;
    RECT 34.655 65.565 34.935 66.445 ;
    RECT 117.655 65.565 117.935 66.445 ;
    RECT 114.335 65.565 114.615 66.445 ;
    RECT 111.015 65.565 111.295 66.445 ;
    RECT 107.695 65.565 107.975 66.445 ;
    RECT 104.375 65.565 104.655 66.445 ;
    RECT 101.055 65.565 101.335 66.445 ;
    RECT 97.735 65.565 98.015 66.445 ;
    RECT 94.415 65.565 94.695 66.445 ;
    RECT 91.095 65.565 91.375 66.445 ;
    RECT 87.775 65.565 88.055 66.445 ;
    RECT 84.455 65.565 84.735 66.445 ;
    RECT 81.135 65.565 81.415 66.445 ;
    RECT 77.815 65.565 78.095 66.445 ;
    RECT 74.495 65.565 74.775 66.445 ;
    RECT 71.175 65.565 71.455 66.445 ;
    RECT 31.335 65.565 31.615 66.445 ;
    RECT 67.855 65.565 68.135 66.445 ;
    RECT 28.015 65.565 28.295 66.445 ;
    RECT 24.695 65.565 24.975 66.445 ;
    RECT 21.375 65.565 21.655 66.445 ;
    RECT 18.055 65.565 18.335 66.445 ;
    RECT 14.735 65.565 15.015 66.445 ;
    RECT 11.415 65.565 11.695 66.445 ;
    RECT 8.095 65.565 8.375 66.445 ;
    RECT 4.775 65.565 5.055 66.445 ;
    RECT 1.455 65.565 1.735 66.445 ;
    RECT 64.535 65.565 64.815 66.445 ;
    RECT 61.215 28.105 61.495 28.985 ;
    RECT 57.895 28.105 58.175 28.985 ;
    RECT 54.575 28.105 54.855 28.985 ;
    RECT 51.255 28.105 51.535 28.985 ;
    RECT 47.935 28.105 48.215 28.985 ;
    RECT 44.615 28.105 44.895 28.985 ;
    RECT 41.295 28.105 41.575 28.985 ;
    RECT 37.975 28.105 38.255 28.985 ;
    RECT 34.655 28.105 34.935 28.985 ;
    RECT 117.655 28.105 117.935 28.985 ;
    RECT 114.335 28.105 114.615 28.985 ;
    RECT 111.015 28.105 111.295 28.985 ;
    RECT 107.695 28.105 107.975 28.985 ;
    RECT 104.375 28.105 104.655 28.985 ;
    RECT 101.055 28.105 101.335 28.985 ;
    RECT 97.735 28.105 98.015 28.985 ;
    RECT 94.415 28.105 94.695 28.985 ;
    RECT 91.095 28.105 91.375 28.985 ;
    RECT 87.775 28.105 88.055 28.985 ;
    RECT 84.455 28.105 84.735 28.985 ;
    RECT 81.135 28.105 81.415 28.985 ;
    RECT 77.815 28.105 78.095 28.985 ;
    RECT 74.495 28.105 74.775 28.985 ;
    RECT 71.175 28.105 71.455 28.985 ;
    RECT 31.335 28.105 31.615 28.985 ;
    RECT 67.855 28.105 68.135 28.985 ;
    RECT 28.015 28.105 28.295 28.985 ;
    RECT 24.695 28.105 24.975 28.985 ;
    RECT 21.375 28.105 21.655 28.985 ;
    RECT 18.055 28.105 18.335 28.985 ;
    RECT 14.735 28.105 15.015 28.985 ;
    RECT 11.415 28.105 11.695 28.985 ;
    RECT 8.095 28.105 8.375 28.985 ;
    RECT 4.775 28.105 5.055 28.985 ;
    RECT 1.455 28.105 1.735 28.985 ;
    RECT 64.535 28.105 64.815 28.985 ;
    RECT 61.215 27.385 61.495 28.265 ;
    RECT 57.895 27.385 58.175 28.265 ;
    RECT 54.575 27.385 54.855 28.265 ;
    RECT 51.255 27.385 51.535 28.265 ;
    RECT 47.935 27.385 48.215 28.265 ;
    RECT 44.615 27.385 44.895 28.265 ;
    RECT 41.295 27.385 41.575 28.265 ;
    RECT 37.975 27.385 38.255 28.265 ;
    RECT 34.655 27.385 34.935 28.265 ;
    RECT 117.655 27.385 117.935 28.265 ;
    RECT 114.335 27.385 114.615 28.265 ;
    RECT 111.015 27.385 111.295 28.265 ;
    RECT 107.695 27.385 107.975 28.265 ;
    RECT 104.375 27.385 104.655 28.265 ;
    RECT 101.055 27.385 101.335 28.265 ;
    RECT 97.735 27.385 98.015 28.265 ;
    RECT 94.415 27.385 94.695 28.265 ;
    RECT 91.095 27.385 91.375 28.265 ;
    RECT 87.775 27.385 88.055 28.265 ;
    RECT 84.455 27.385 84.735 28.265 ;
    RECT 81.135 27.385 81.415 28.265 ;
    RECT 77.815 27.385 78.095 28.265 ;
    RECT 74.495 27.385 74.775 28.265 ;
    RECT 71.175 27.385 71.455 28.265 ;
    RECT 31.335 27.385 31.615 28.265 ;
    RECT 67.855 27.385 68.135 28.265 ;
    RECT 28.015 27.385 28.295 28.265 ;
    RECT 24.695 27.385 24.975 28.265 ;
    RECT 21.375 27.385 21.655 28.265 ;
    RECT 18.055 27.385 18.335 28.265 ;
    RECT 14.735 27.385 15.015 28.265 ;
    RECT 11.415 27.385 11.695 28.265 ;
    RECT 8.095 27.385 8.375 28.265 ;
    RECT 4.775 27.385 5.055 28.265 ;
    RECT 1.455 27.385 1.735 28.265 ;
    RECT 64.535 27.385 64.815 28.265 ;
    RECT 61.215 26.665 61.495 27.545 ;
    RECT 57.895 26.665 58.175 27.545 ;
    RECT 54.575 26.665 54.855 27.545 ;
    RECT 51.255 26.665 51.535 27.545 ;
    RECT 47.935 26.665 48.215 27.545 ;
    RECT 44.615 26.665 44.895 27.545 ;
    RECT 41.295 26.665 41.575 27.545 ;
    RECT 37.975 26.665 38.255 27.545 ;
    RECT 34.655 26.665 34.935 27.545 ;
    RECT 117.655 26.665 117.935 27.545 ;
    RECT 114.335 26.665 114.615 27.545 ;
    RECT 111.015 26.665 111.295 27.545 ;
    RECT 107.695 26.665 107.975 27.545 ;
    RECT 104.375 26.665 104.655 27.545 ;
    RECT 101.055 26.665 101.335 27.545 ;
    RECT 97.735 26.665 98.015 27.545 ;
    RECT 94.415 26.665 94.695 27.545 ;
    RECT 91.095 26.665 91.375 27.545 ;
    RECT 87.775 26.665 88.055 27.545 ;
    RECT 84.455 26.665 84.735 27.545 ;
    RECT 81.135 26.665 81.415 27.545 ;
    RECT 77.815 26.665 78.095 27.545 ;
    RECT 74.495 26.665 74.775 27.545 ;
    RECT 71.175 26.665 71.455 27.545 ;
    RECT 31.335 26.665 31.615 27.545 ;
    RECT 67.855 26.665 68.135 27.545 ;
    RECT 28.015 26.665 28.295 27.545 ;
    RECT 24.695 26.665 24.975 27.545 ;
    RECT 21.375 26.665 21.655 27.545 ;
    RECT 18.055 26.665 18.335 27.545 ;
    RECT 14.735 26.665 15.015 27.545 ;
    RECT 11.415 26.665 11.695 27.545 ;
    RECT 8.095 26.665 8.375 27.545 ;
    RECT 4.775 26.665 5.055 27.545 ;
    RECT 1.455 26.665 1.735 27.545 ;
    RECT 64.535 26.665 64.815 27.545 ;
    RECT 61.215 25.945 61.495 26.825 ;
    RECT 57.895 25.945 58.175 26.825 ;
    RECT 54.575 25.945 54.855 26.825 ;
    RECT 51.255 25.945 51.535 26.825 ;
    RECT 47.935 25.945 48.215 26.825 ;
    RECT 44.615 25.945 44.895 26.825 ;
    RECT 41.295 25.945 41.575 26.825 ;
    RECT 37.975 25.945 38.255 26.825 ;
    RECT 34.655 25.945 34.935 26.825 ;
    RECT 117.655 25.945 117.935 26.825 ;
    RECT 114.335 25.945 114.615 26.825 ;
    RECT 111.015 25.945 111.295 26.825 ;
    RECT 107.695 25.945 107.975 26.825 ;
    RECT 104.375 25.945 104.655 26.825 ;
    RECT 101.055 25.945 101.335 26.825 ;
    RECT 97.735 25.945 98.015 26.825 ;
    RECT 94.415 25.945 94.695 26.825 ;
    RECT 91.095 25.945 91.375 26.825 ;
    RECT 87.775 25.945 88.055 26.825 ;
    RECT 84.455 25.945 84.735 26.825 ;
    RECT 81.135 25.945 81.415 26.825 ;
    RECT 77.815 25.945 78.095 26.825 ;
    RECT 74.495 25.945 74.775 26.825 ;
    RECT 71.175 25.945 71.455 26.825 ;
    RECT 31.335 25.945 31.615 26.825 ;
    RECT 67.855 25.945 68.135 26.825 ;
    RECT 28.015 25.945 28.295 26.825 ;
    RECT 24.695 25.945 24.975 26.825 ;
    RECT 21.375 25.945 21.655 26.825 ;
    RECT 18.055 25.945 18.335 26.825 ;
    RECT 14.735 25.945 15.015 26.825 ;
    RECT 11.415 25.945 11.695 26.825 ;
    RECT 8.095 25.945 8.375 26.825 ;
    RECT 4.775 25.945 5.055 26.825 ;
    RECT 1.455 25.945 1.735 26.825 ;
    RECT 64.535 25.945 64.815 26.825 ;
    RECT 61.215 25.225 61.495 26.105 ;
    RECT 57.895 25.225 58.175 26.105 ;
    RECT 54.575 25.225 54.855 26.105 ;
    RECT 51.255 25.225 51.535 26.105 ;
    RECT 47.935 25.225 48.215 26.105 ;
    RECT 44.615 25.225 44.895 26.105 ;
    RECT 41.295 25.225 41.575 26.105 ;
    RECT 37.975 25.225 38.255 26.105 ;
    RECT 34.655 25.225 34.935 26.105 ;
    RECT 117.655 25.225 117.935 26.105 ;
    RECT 114.335 25.225 114.615 26.105 ;
    RECT 111.015 25.225 111.295 26.105 ;
    RECT 107.695 25.225 107.975 26.105 ;
    RECT 104.375 25.225 104.655 26.105 ;
    RECT 101.055 25.225 101.335 26.105 ;
    RECT 97.735 25.225 98.015 26.105 ;
    RECT 94.415 25.225 94.695 26.105 ;
    RECT 91.095 25.225 91.375 26.105 ;
    RECT 87.775 25.225 88.055 26.105 ;
    RECT 84.455 25.225 84.735 26.105 ;
    RECT 81.135 25.225 81.415 26.105 ;
    RECT 77.815 25.225 78.095 26.105 ;
    RECT 74.495 25.225 74.775 26.105 ;
    RECT 71.175 25.225 71.455 26.105 ;
    RECT 31.335 25.225 31.615 26.105 ;
    RECT 67.855 25.225 68.135 26.105 ;
    RECT 28.015 25.225 28.295 26.105 ;
    RECT 24.695 25.225 24.975 26.105 ;
    RECT 21.375 25.225 21.655 26.105 ;
    RECT 18.055 25.225 18.335 26.105 ;
    RECT 14.735 25.225 15.015 26.105 ;
    RECT 11.415 25.225 11.695 26.105 ;
    RECT 8.095 25.225 8.375 26.105 ;
    RECT 4.775 25.225 5.055 26.105 ;
    RECT 1.455 25.225 1.735 26.105 ;
    RECT 64.535 25.225 64.815 26.105 ;
    RECT 61.215 64.845 61.495 65.725 ;
    RECT 57.895 64.845 58.175 65.725 ;
    RECT 54.575 64.845 54.855 65.725 ;
    RECT 51.255 64.845 51.535 65.725 ;
    RECT 47.935 64.845 48.215 65.725 ;
    RECT 44.615 64.845 44.895 65.725 ;
    RECT 41.295 64.845 41.575 65.725 ;
    RECT 37.975 64.845 38.255 65.725 ;
    RECT 34.655 64.845 34.935 65.725 ;
    RECT 117.655 64.845 117.935 65.725 ;
    RECT 114.335 64.845 114.615 65.725 ;
    RECT 111.015 64.845 111.295 65.725 ;
    RECT 107.695 64.845 107.975 65.725 ;
    RECT 104.375 64.845 104.655 65.725 ;
    RECT 101.055 64.845 101.335 65.725 ;
    RECT 97.735 64.845 98.015 65.725 ;
    RECT 94.415 64.845 94.695 65.725 ;
    RECT 91.095 64.845 91.375 65.725 ;
    RECT 87.775 64.845 88.055 65.725 ;
    RECT 84.455 64.845 84.735 65.725 ;
    RECT 81.135 64.845 81.415 65.725 ;
    RECT 77.815 64.845 78.095 65.725 ;
    RECT 74.495 64.845 74.775 65.725 ;
    RECT 71.175 64.845 71.455 65.725 ;
    RECT 31.335 64.845 31.615 65.725 ;
    RECT 67.855 64.845 68.135 65.725 ;
    RECT 28.015 64.845 28.295 65.725 ;
    RECT 24.695 64.845 24.975 65.725 ;
    RECT 21.375 64.845 21.655 65.725 ;
    RECT 18.055 64.845 18.335 65.725 ;
    RECT 14.735 64.845 15.015 65.725 ;
    RECT 11.415 64.845 11.695 65.725 ;
    RECT 8.095 64.845 8.375 65.725 ;
    RECT 4.775 64.845 5.055 65.725 ;
    RECT 1.455 64.845 1.735 65.725 ;
    RECT 64.535 64.845 64.815 65.725 ;
    RECT 61.215 56.185 61.495 57.065 ;
    RECT 57.895 56.185 58.175 57.065 ;
    RECT 54.575 56.185 54.855 57.065 ;
    RECT 51.255 56.185 51.535 57.065 ;
    RECT 47.935 56.185 48.215 57.065 ;
    RECT 44.615 56.185 44.895 57.065 ;
    RECT 41.295 56.185 41.575 57.065 ;
    RECT 37.975 56.185 38.255 57.065 ;
    RECT 34.655 56.185 34.935 57.065 ;
    RECT 117.655 56.185 117.935 57.065 ;
    RECT 114.335 56.185 114.615 57.065 ;
    RECT 111.015 56.185 111.295 57.065 ;
    RECT 107.695 56.185 107.975 57.065 ;
    RECT 104.375 56.185 104.655 57.065 ;
    RECT 101.055 56.185 101.335 57.065 ;
    RECT 97.735 56.185 98.015 57.065 ;
    RECT 94.415 56.185 94.695 57.065 ;
    RECT 91.095 56.185 91.375 57.065 ;
    RECT 87.775 56.185 88.055 57.065 ;
    RECT 84.455 56.185 84.735 57.065 ;
    RECT 81.135 56.185 81.415 57.065 ;
    RECT 77.815 56.185 78.095 57.065 ;
    RECT 74.495 56.185 74.775 57.065 ;
    RECT 71.175 56.185 71.455 57.065 ;
    RECT 31.335 56.185 31.615 57.065 ;
    RECT 67.855 56.185 68.135 57.065 ;
    RECT 28.015 56.185 28.295 57.065 ;
    RECT 24.695 56.185 24.975 57.065 ;
    RECT 21.375 56.185 21.655 57.065 ;
    RECT 18.055 56.185 18.335 57.065 ;
    RECT 14.735 56.185 15.015 57.065 ;
    RECT 11.415 56.185 11.695 57.065 ;
    RECT 8.095 56.185 8.375 57.065 ;
    RECT 4.775 56.185 5.055 57.065 ;
    RECT 1.455 56.185 1.735 57.065 ;
    RECT 64.535 56.185 64.815 57.065 ;
    RECT 61.215 24.505 61.495 25.385 ;
    RECT 57.895 24.505 58.175 25.385 ;
    RECT 54.575 24.505 54.855 25.385 ;
    RECT 51.255 24.505 51.535 25.385 ;
    RECT 47.935 24.505 48.215 25.385 ;
    RECT 44.615 24.505 44.895 25.385 ;
    RECT 41.295 24.505 41.575 25.385 ;
    RECT 37.975 24.505 38.255 25.385 ;
    RECT 34.655 24.505 34.935 25.385 ;
    RECT 117.655 24.505 117.935 25.385 ;
    RECT 114.335 24.505 114.615 25.385 ;
    RECT 111.015 24.505 111.295 25.385 ;
    RECT 107.695 24.505 107.975 25.385 ;
    RECT 104.375 24.505 104.655 25.385 ;
    RECT 101.055 24.505 101.335 25.385 ;
    RECT 97.735 24.505 98.015 25.385 ;
    RECT 94.415 24.505 94.695 25.385 ;
    RECT 91.095 24.505 91.375 25.385 ;
    RECT 87.775 24.505 88.055 25.385 ;
    RECT 84.455 24.505 84.735 25.385 ;
    RECT 81.135 24.505 81.415 25.385 ;
    RECT 77.815 24.505 78.095 25.385 ;
    RECT 74.495 24.505 74.775 25.385 ;
    RECT 71.175 24.505 71.455 25.385 ;
    RECT 31.335 24.505 31.615 25.385 ;
    RECT 67.855 24.505 68.135 25.385 ;
    RECT 28.015 24.505 28.295 25.385 ;
    RECT 24.695 24.505 24.975 25.385 ;
    RECT 21.375 24.505 21.655 25.385 ;
    RECT 18.055 24.505 18.335 25.385 ;
    RECT 14.735 24.505 15.015 25.385 ;
    RECT 11.415 24.505 11.695 25.385 ;
    RECT 8.095 24.505 8.375 25.385 ;
    RECT 4.775 24.505 5.055 25.385 ;
    RECT 1.455 24.505 1.735 25.385 ;
    RECT 64.535 24.505 64.815 25.385 ;
    RECT 61.215 64.125 61.495 65.005 ;
    RECT 57.895 64.125 58.175 65.005 ;
    RECT 54.575 64.125 54.855 65.005 ;
    RECT 51.255 64.125 51.535 65.005 ;
    RECT 47.935 64.125 48.215 65.005 ;
    RECT 44.615 64.125 44.895 65.005 ;
    RECT 41.295 64.125 41.575 65.005 ;
    RECT 37.975 64.125 38.255 65.005 ;
    RECT 34.655 64.125 34.935 65.005 ;
    RECT 117.655 64.125 117.935 65.005 ;
    RECT 114.335 64.125 114.615 65.005 ;
    RECT 111.015 64.125 111.295 65.005 ;
    RECT 107.695 64.125 107.975 65.005 ;
    RECT 104.375 64.125 104.655 65.005 ;
    RECT 101.055 64.125 101.335 65.005 ;
    RECT 97.735 64.125 98.015 65.005 ;
    RECT 94.415 64.125 94.695 65.005 ;
    RECT 91.095 64.125 91.375 65.005 ;
    RECT 87.775 64.125 88.055 65.005 ;
    RECT 84.455 64.125 84.735 65.005 ;
    RECT 81.135 64.125 81.415 65.005 ;
    RECT 77.815 64.125 78.095 65.005 ;
    RECT 74.495 64.125 74.775 65.005 ;
    RECT 71.175 64.125 71.455 65.005 ;
    RECT 31.335 64.125 31.615 65.005 ;
    RECT 67.855 64.125 68.135 65.005 ;
    RECT 28.015 64.125 28.295 65.005 ;
    RECT 24.695 64.125 24.975 65.005 ;
    RECT 21.375 64.125 21.655 65.005 ;
    RECT 18.055 64.125 18.335 65.005 ;
    RECT 14.735 64.125 15.015 65.005 ;
    RECT 11.415 64.125 11.695 65.005 ;
    RECT 8.095 64.125 8.375 65.005 ;
    RECT 4.775 64.125 5.055 65.005 ;
    RECT 1.455 64.125 1.735 65.005 ;
    RECT 64.535 64.125 64.815 65.005 ;
    RECT 61.215 23.785 61.495 24.665 ;
    RECT 57.895 23.785 58.175 24.665 ;
    RECT 54.575 23.785 54.855 24.665 ;
    RECT 51.255 23.785 51.535 24.665 ;
    RECT 47.935 23.785 48.215 24.665 ;
    RECT 44.615 23.785 44.895 24.665 ;
    RECT 41.295 23.785 41.575 24.665 ;
    RECT 37.975 23.785 38.255 24.665 ;
    RECT 34.655 23.785 34.935 24.665 ;
    RECT 117.655 23.785 117.935 24.665 ;
    RECT 114.335 23.785 114.615 24.665 ;
    RECT 111.015 23.785 111.295 24.665 ;
    RECT 107.695 23.785 107.975 24.665 ;
    RECT 104.375 23.785 104.655 24.665 ;
    RECT 101.055 23.785 101.335 24.665 ;
    RECT 97.735 23.785 98.015 24.665 ;
    RECT 94.415 23.785 94.695 24.665 ;
    RECT 91.095 23.785 91.375 24.665 ;
    RECT 87.775 23.785 88.055 24.665 ;
    RECT 84.455 23.785 84.735 24.665 ;
    RECT 81.135 23.785 81.415 24.665 ;
    RECT 77.815 23.785 78.095 24.665 ;
    RECT 74.495 23.785 74.775 24.665 ;
    RECT 71.175 23.785 71.455 24.665 ;
    RECT 31.335 23.785 31.615 24.665 ;
    RECT 67.855 23.785 68.135 24.665 ;
    RECT 28.015 23.785 28.295 24.665 ;
    RECT 24.695 23.785 24.975 24.665 ;
    RECT 21.375 23.785 21.655 24.665 ;
    RECT 18.055 23.785 18.335 24.665 ;
    RECT 14.735 23.785 15.015 24.665 ;
    RECT 11.415 23.785 11.695 24.665 ;
    RECT 8.095 23.785 8.375 24.665 ;
    RECT 4.775 23.785 5.055 24.665 ;
    RECT 1.455 23.785 1.735 24.665 ;
    RECT 64.535 23.785 64.815 24.665 ;
    RECT 61.215 63.405 61.495 64.285 ;
    RECT 57.895 63.405 58.175 64.285 ;
    RECT 54.575 63.405 54.855 64.285 ;
    RECT 51.255 63.405 51.535 64.285 ;
    RECT 47.935 63.405 48.215 64.285 ;
    RECT 44.615 63.405 44.895 64.285 ;
    RECT 41.295 63.405 41.575 64.285 ;
    RECT 37.975 63.405 38.255 64.285 ;
    RECT 34.655 63.405 34.935 64.285 ;
    RECT 117.655 63.405 117.935 64.285 ;
    RECT 114.335 63.405 114.615 64.285 ;
    RECT 111.015 63.405 111.295 64.285 ;
    RECT 107.695 63.405 107.975 64.285 ;
    RECT 104.375 63.405 104.655 64.285 ;
    RECT 101.055 63.405 101.335 64.285 ;
    RECT 97.735 63.405 98.015 64.285 ;
    RECT 94.415 63.405 94.695 64.285 ;
    RECT 91.095 63.405 91.375 64.285 ;
    RECT 87.775 63.405 88.055 64.285 ;
    RECT 84.455 63.405 84.735 64.285 ;
    RECT 81.135 63.405 81.415 64.285 ;
    RECT 77.815 63.405 78.095 64.285 ;
    RECT 74.495 63.405 74.775 64.285 ;
    RECT 71.175 63.405 71.455 64.285 ;
    RECT 31.335 63.405 31.615 64.285 ;
    RECT 67.855 63.405 68.135 64.285 ;
    RECT 28.015 63.405 28.295 64.285 ;
    RECT 24.695 63.405 24.975 64.285 ;
    RECT 21.375 63.405 21.655 64.285 ;
    RECT 18.055 63.405 18.335 64.285 ;
    RECT 14.735 63.405 15.015 64.285 ;
    RECT 11.415 63.405 11.695 64.285 ;
    RECT 8.095 63.405 8.375 64.285 ;
    RECT 4.775 63.405 5.055 64.285 ;
    RECT 1.455 63.405 1.735 64.285 ;
    RECT 64.535 63.405 64.815 64.285 ;
    RECT 61.215 23.065 61.495 23.945 ;
    RECT 57.895 23.065 58.175 23.945 ;
    RECT 54.575 23.065 54.855 23.945 ;
    RECT 51.255 23.065 51.535 23.945 ;
    RECT 47.935 23.065 48.215 23.945 ;
    RECT 44.615 23.065 44.895 23.945 ;
    RECT 41.295 23.065 41.575 23.945 ;
    RECT 37.975 23.065 38.255 23.945 ;
    RECT 34.655 23.065 34.935 23.945 ;
    RECT 117.655 23.065 117.935 23.945 ;
    RECT 114.335 23.065 114.615 23.945 ;
    RECT 111.015 23.065 111.295 23.945 ;
    RECT 107.695 23.065 107.975 23.945 ;
    RECT 104.375 23.065 104.655 23.945 ;
    RECT 101.055 23.065 101.335 23.945 ;
    RECT 97.735 23.065 98.015 23.945 ;
    RECT 94.415 23.065 94.695 23.945 ;
    RECT 91.095 23.065 91.375 23.945 ;
    RECT 87.775 23.065 88.055 23.945 ;
    RECT 84.455 23.065 84.735 23.945 ;
    RECT 81.135 23.065 81.415 23.945 ;
    RECT 77.815 23.065 78.095 23.945 ;
    RECT 74.495 23.065 74.775 23.945 ;
    RECT 71.175 23.065 71.455 23.945 ;
    RECT 31.335 23.065 31.615 23.945 ;
    RECT 67.855 23.065 68.135 23.945 ;
    RECT 28.015 23.065 28.295 23.945 ;
    RECT 24.695 23.065 24.975 23.945 ;
    RECT 21.375 23.065 21.655 23.945 ;
    RECT 18.055 23.065 18.335 23.945 ;
    RECT 14.735 23.065 15.015 23.945 ;
    RECT 11.415 23.065 11.695 23.945 ;
    RECT 8.095 23.065 8.375 23.945 ;
    RECT 4.775 23.065 5.055 23.945 ;
    RECT 1.455 23.065 1.735 23.945 ;
    RECT 64.535 23.065 64.815 23.945 ;
    RECT 61.215 62.685 61.495 63.565 ;
    RECT 57.895 62.685 58.175 63.565 ;
    RECT 54.575 62.685 54.855 63.565 ;
    RECT 51.255 62.685 51.535 63.565 ;
    RECT 47.935 62.685 48.215 63.565 ;
    RECT 44.615 62.685 44.895 63.565 ;
    RECT 41.295 62.685 41.575 63.565 ;
    RECT 37.975 62.685 38.255 63.565 ;
    RECT 34.655 62.685 34.935 63.565 ;
    RECT 117.655 62.685 117.935 63.565 ;
    RECT 114.335 62.685 114.615 63.565 ;
    RECT 111.015 62.685 111.295 63.565 ;
    RECT 107.695 62.685 107.975 63.565 ;
    RECT 104.375 62.685 104.655 63.565 ;
    RECT 101.055 62.685 101.335 63.565 ;
    RECT 97.735 62.685 98.015 63.565 ;
    RECT 94.415 62.685 94.695 63.565 ;
    RECT 91.095 62.685 91.375 63.565 ;
    RECT 87.775 62.685 88.055 63.565 ;
    RECT 84.455 62.685 84.735 63.565 ;
    RECT 81.135 62.685 81.415 63.565 ;
    RECT 77.815 62.685 78.095 63.565 ;
    RECT 74.495 62.685 74.775 63.565 ;
    RECT 71.175 62.685 71.455 63.565 ;
    RECT 31.335 62.685 31.615 63.565 ;
    RECT 67.855 62.685 68.135 63.565 ;
    RECT 28.015 62.685 28.295 63.565 ;
    RECT 24.695 62.685 24.975 63.565 ;
    RECT 21.375 62.685 21.655 63.565 ;
    RECT 18.055 62.685 18.335 63.565 ;
    RECT 14.735 62.685 15.015 63.565 ;
    RECT 11.415 62.685 11.695 63.565 ;
    RECT 8.095 62.685 8.375 63.565 ;
    RECT 4.775 62.685 5.055 63.565 ;
    RECT 1.455 62.685 1.735 63.565 ;
    RECT 64.535 62.685 64.815 63.565 ;
    RECT 61.215 22.345 61.495 23.225 ;
    RECT 57.895 22.345 58.175 23.225 ;
    RECT 54.575 22.345 54.855 23.225 ;
    RECT 51.255 22.345 51.535 23.225 ;
    RECT 47.935 22.345 48.215 23.225 ;
    RECT 44.615 22.345 44.895 23.225 ;
    RECT 41.295 22.345 41.575 23.225 ;
    RECT 37.975 22.345 38.255 23.225 ;
    RECT 34.655 22.345 34.935 23.225 ;
    RECT 117.655 22.345 117.935 23.225 ;
    RECT 114.335 22.345 114.615 23.225 ;
    RECT 111.015 22.345 111.295 23.225 ;
    RECT 107.695 22.345 107.975 23.225 ;
    RECT 104.375 22.345 104.655 23.225 ;
    RECT 101.055 22.345 101.335 23.225 ;
    RECT 97.735 22.345 98.015 23.225 ;
    RECT 94.415 22.345 94.695 23.225 ;
    RECT 91.095 22.345 91.375 23.225 ;
    RECT 87.775 22.345 88.055 23.225 ;
    RECT 84.455 22.345 84.735 23.225 ;
    RECT 81.135 22.345 81.415 23.225 ;
    RECT 77.815 22.345 78.095 23.225 ;
    RECT 74.495 22.345 74.775 23.225 ;
    RECT 71.175 22.345 71.455 23.225 ;
    RECT 31.335 22.345 31.615 23.225 ;
    RECT 67.855 22.345 68.135 23.225 ;
    RECT 28.015 22.345 28.295 23.225 ;
    RECT 24.695 22.345 24.975 23.225 ;
    RECT 21.375 22.345 21.655 23.225 ;
    RECT 18.055 22.345 18.335 23.225 ;
    RECT 14.735 22.345 15.015 23.225 ;
    RECT 11.415 22.345 11.695 23.225 ;
    RECT 8.095 22.345 8.375 23.225 ;
    RECT 4.775 22.345 5.055 23.225 ;
    RECT 1.455 22.345 1.735 23.225 ;
    RECT 64.535 22.345 64.815 23.225 ;
    RECT 61.215 61.965 61.495 62.845 ;
    RECT 57.895 61.965 58.175 62.845 ;
    RECT 54.575 61.965 54.855 62.845 ;
    RECT 51.255 61.965 51.535 62.845 ;
    RECT 47.935 61.965 48.215 62.845 ;
    RECT 44.615 61.965 44.895 62.845 ;
    RECT 41.295 61.965 41.575 62.845 ;
    RECT 37.975 61.965 38.255 62.845 ;
    RECT 34.655 61.965 34.935 62.845 ;
    RECT 117.655 61.965 117.935 62.845 ;
    RECT 114.335 61.965 114.615 62.845 ;
    RECT 111.015 61.965 111.295 62.845 ;
    RECT 107.695 61.965 107.975 62.845 ;
    RECT 104.375 61.965 104.655 62.845 ;
    RECT 101.055 61.965 101.335 62.845 ;
    RECT 97.735 61.965 98.015 62.845 ;
    RECT 94.415 61.965 94.695 62.845 ;
    RECT 91.095 61.965 91.375 62.845 ;
    RECT 87.775 61.965 88.055 62.845 ;
    RECT 84.455 61.965 84.735 62.845 ;
    RECT 81.135 61.965 81.415 62.845 ;
    RECT 77.815 61.965 78.095 62.845 ;
    RECT 74.495 61.965 74.775 62.845 ;
    RECT 71.175 61.965 71.455 62.845 ;
    RECT 31.335 61.965 31.615 62.845 ;
    RECT 67.855 61.965 68.135 62.845 ;
    RECT 28.015 61.965 28.295 62.845 ;
    RECT 24.695 61.965 24.975 62.845 ;
    RECT 21.375 61.965 21.655 62.845 ;
    RECT 18.055 61.965 18.335 62.845 ;
    RECT 14.735 61.965 15.015 62.845 ;
    RECT 11.415 61.965 11.695 62.845 ;
    RECT 8.095 61.965 8.375 62.845 ;
    RECT 4.775 61.965 5.055 62.845 ;
    RECT 1.455 61.965 1.735 62.845 ;
    RECT 64.535 61.965 64.815 62.845 ;
    RECT 61.215 21.625 61.495 22.505 ;
    RECT 57.895 21.625 58.175 22.505 ;
    RECT 54.575 21.625 54.855 22.505 ;
    RECT 51.255 21.625 51.535 22.505 ;
    RECT 47.935 21.625 48.215 22.505 ;
    RECT 44.615 21.625 44.895 22.505 ;
    RECT 41.295 21.625 41.575 22.505 ;
    RECT 37.975 21.625 38.255 22.505 ;
    RECT 34.655 21.625 34.935 22.505 ;
    RECT 117.655 21.625 117.935 22.505 ;
    RECT 114.335 21.625 114.615 22.505 ;
    RECT 111.015 21.625 111.295 22.505 ;
    RECT 107.695 21.625 107.975 22.505 ;
    RECT 104.375 21.625 104.655 22.505 ;
    RECT 101.055 21.625 101.335 22.505 ;
    RECT 97.735 21.625 98.015 22.505 ;
    RECT 94.415 21.625 94.695 22.505 ;
    RECT 91.095 21.625 91.375 22.505 ;
    RECT 87.775 21.625 88.055 22.505 ;
    RECT 84.455 21.625 84.735 22.505 ;
    RECT 81.135 21.625 81.415 22.505 ;
    RECT 77.815 21.625 78.095 22.505 ;
    RECT 74.495 21.625 74.775 22.505 ;
    RECT 71.175 21.625 71.455 22.505 ;
    RECT 31.335 21.625 31.615 22.505 ;
    RECT 67.855 21.625 68.135 22.505 ;
    RECT 28.015 21.625 28.295 22.505 ;
    RECT 24.695 21.625 24.975 22.505 ;
    RECT 21.375 21.625 21.655 22.505 ;
    RECT 18.055 21.625 18.335 22.505 ;
    RECT 14.735 21.625 15.015 22.505 ;
    RECT 11.415 21.625 11.695 22.505 ;
    RECT 8.095 21.625 8.375 22.505 ;
    RECT 4.775 21.625 5.055 22.505 ;
    RECT 1.455 21.625 1.735 22.505 ;
    RECT 64.535 21.625 64.815 22.505 ;
    RECT 61.215 61.245 61.495 62.125 ;
    RECT 57.895 61.245 58.175 62.125 ;
    RECT 54.575 61.245 54.855 62.125 ;
    RECT 51.255 61.245 51.535 62.125 ;
    RECT 47.935 61.245 48.215 62.125 ;
    RECT 44.615 61.245 44.895 62.125 ;
    RECT 41.295 61.245 41.575 62.125 ;
    RECT 37.975 61.245 38.255 62.125 ;
    RECT 34.655 61.245 34.935 62.125 ;
    RECT 117.655 61.245 117.935 62.125 ;
    RECT 114.335 61.245 114.615 62.125 ;
    RECT 111.015 61.245 111.295 62.125 ;
    RECT 107.695 61.245 107.975 62.125 ;
    RECT 104.375 61.245 104.655 62.125 ;
    RECT 101.055 61.245 101.335 62.125 ;
    RECT 97.735 61.245 98.015 62.125 ;
    RECT 94.415 61.245 94.695 62.125 ;
    RECT 91.095 61.245 91.375 62.125 ;
    RECT 87.775 61.245 88.055 62.125 ;
    RECT 84.455 61.245 84.735 62.125 ;
    RECT 81.135 61.245 81.415 62.125 ;
    RECT 77.815 61.245 78.095 62.125 ;
    RECT 74.495 61.245 74.775 62.125 ;
    RECT 71.175 61.245 71.455 62.125 ;
    RECT 31.335 61.245 31.615 62.125 ;
    RECT 67.855 61.245 68.135 62.125 ;
    RECT 28.015 61.245 28.295 62.125 ;
    RECT 24.695 61.245 24.975 62.125 ;
    RECT 21.375 61.245 21.655 62.125 ;
    RECT 18.055 61.245 18.335 62.125 ;
    RECT 14.735 61.245 15.015 62.125 ;
    RECT 11.415 61.245 11.695 62.125 ;
    RECT 8.095 61.245 8.375 62.125 ;
    RECT 4.775 61.245 5.055 62.125 ;
    RECT 1.455 61.245 1.735 62.125 ;
    RECT 64.535 61.245 64.815 62.125 ;
    RECT 31.335 60.585 31.615 61.325 ;
    RECT 28.015 60.585 28.295 61.325 ;
    RECT 24.695 60.585 24.975 61.325 ;
    RECT 21.375 60.585 21.655 61.325 ;
    RECT 18.055 60.585 18.335 61.325 ;
    RECT 14.735 60.585 15.015 61.325 ;
    RECT 11.415 60.585 11.695 61.325 ;
    RECT 8.095 60.585 8.375 61.325 ;
    RECT 4.775 60.585 5.055 61.325 ;
    RECT 1.455 60.585 1.735 61.325 ;
    RECT 117.655 60.585 117.935 61.325 ;
    RECT 114.335 60.585 114.615 61.325 ;
    RECT 111.015 60.585 111.295 61.325 ;
    RECT 107.695 60.585 107.975 61.325 ;
    RECT 104.375 60.585 104.655 61.325 ;
    RECT 101.055 60.585 101.335 61.325 ;
    RECT 97.735 60.585 98.015 61.325 ;
    RECT 94.415 60.585 94.695 61.325 ;
    RECT 91.095 60.585 91.375 61.325 ;
    RECT 87.775 60.585 88.055 61.325 ;
    RECT 84.455 60.585 84.735 61.325 ;
    RECT 81.135 60.585 81.415 61.325 ;
    RECT 77.815 60.585 78.095 61.325 ;
    RECT 74.495 60.585 74.775 61.325 ;
    RECT 71.175 60.585 71.455 61.325 ;
    RECT 67.855 60.585 68.135 61.325 ;
    RECT 64.535 60.585 64.815 61.325 ;
    RECT 61.215 60.585 61.495 61.325 ;
    RECT 57.895 60.585 58.175 61.325 ;
    RECT 54.575 60.585 54.855 61.325 ;
    RECT 51.255 60.585 51.535 61.325 ;
    RECT 47.935 60.585 48.215 61.325 ;
    RECT 44.615 60.585 44.895 61.325 ;
    RECT 41.295 60.585 41.575 61.325 ;
    RECT 37.975 60.585 38.255 61.325 ;
    RECT 34.655 60.585 34.935 61.325 ;
    RECT 61.215 59.785 61.495 60.665 ;
    RECT 57.895 59.785 58.175 60.665 ;
    RECT 54.575 59.785 54.855 60.665 ;
    RECT 51.255 59.785 51.535 60.665 ;
    RECT 47.935 59.785 48.215 60.665 ;
    RECT 44.615 59.785 44.895 60.665 ;
    RECT 41.295 59.785 41.575 60.665 ;
    RECT 37.975 59.785 38.255 60.665 ;
    RECT 34.655 59.785 34.935 60.665 ;
    RECT 117.655 59.785 117.935 60.665 ;
    RECT 114.335 59.785 114.615 60.665 ;
    RECT 111.015 59.785 111.295 60.665 ;
    RECT 107.695 59.785 107.975 60.665 ;
    RECT 104.375 59.785 104.655 60.665 ;
    RECT 101.055 59.785 101.335 60.665 ;
    RECT 97.735 59.785 98.015 60.665 ;
    RECT 94.415 59.785 94.695 60.665 ;
    RECT 91.095 59.785 91.375 60.665 ;
    RECT 87.775 59.785 88.055 60.665 ;
    RECT 84.455 59.785 84.735 60.665 ;
    RECT 81.135 59.785 81.415 60.665 ;
    RECT 77.815 59.785 78.095 60.665 ;
    RECT 74.495 59.785 74.775 60.665 ;
    RECT 71.175 59.785 71.455 60.665 ;
    RECT 31.335 59.785 31.615 60.665 ;
    RECT 67.855 59.785 68.135 60.665 ;
    RECT 28.015 59.785 28.295 60.665 ;
    RECT 24.695 59.785 24.975 60.665 ;
    RECT 21.375 59.785 21.655 60.665 ;
    RECT 18.055 59.785 18.335 60.665 ;
    RECT 14.735 59.785 15.015 60.665 ;
    RECT 11.415 59.785 11.695 60.665 ;
    RECT 8.095 59.785 8.375 60.665 ;
    RECT 4.775 59.785 5.055 60.665 ;
    RECT 1.455 59.785 1.735 60.665 ;
    RECT 64.535 59.785 64.815 60.665 ;
    RECT 61.215 59.065 61.495 59.945 ;
    RECT 57.895 59.065 58.175 59.945 ;
    RECT 54.575 59.065 54.855 59.945 ;
    RECT 51.255 59.065 51.535 59.945 ;
    RECT 47.935 59.065 48.215 59.945 ;
    RECT 44.615 59.065 44.895 59.945 ;
    RECT 41.295 59.065 41.575 59.945 ;
    RECT 37.975 59.065 38.255 59.945 ;
    RECT 34.655 59.065 34.935 59.945 ;
    RECT 117.655 59.065 117.935 59.945 ;
    RECT 114.335 59.065 114.615 59.945 ;
    RECT 111.015 59.065 111.295 59.945 ;
    RECT 107.695 59.065 107.975 59.945 ;
    RECT 104.375 59.065 104.655 59.945 ;
    RECT 101.055 59.065 101.335 59.945 ;
    RECT 97.735 59.065 98.015 59.945 ;
    RECT 94.415 59.065 94.695 59.945 ;
    RECT 91.095 59.065 91.375 59.945 ;
    RECT 87.775 59.065 88.055 59.945 ;
    RECT 84.455 59.065 84.735 59.945 ;
    RECT 81.135 59.065 81.415 59.945 ;
    RECT 77.815 59.065 78.095 59.945 ;
    RECT 74.495 59.065 74.775 59.945 ;
    RECT 71.175 59.065 71.455 59.945 ;
    RECT 31.335 59.065 31.615 59.945 ;
    RECT 67.855 59.065 68.135 59.945 ;
    RECT 28.015 59.065 28.295 59.945 ;
    RECT 24.695 59.065 24.975 59.945 ;
    RECT 21.375 59.065 21.655 59.945 ;
    RECT 18.055 59.065 18.335 59.945 ;
    RECT 14.735 59.065 15.015 59.945 ;
    RECT 11.415 59.065 11.695 59.945 ;
    RECT 8.095 59.065 8.375 59.945 ;
    RECT 4.775 59.065 5.055 59.945 ;
    RECT 1.455 59.065 1.735 59.945 ;
    RECT 64.535 59.065 64.815 59.945 ;
    RECT 61.215 58.345 61.495 59.225 ;
    RECT 57.895 58.345 58.175 59.225 ;
    RECT 54.575 58.345 54.855 59.225 ;
    RECT 51.255 58.345 51.535 59.225 ;
    RECT 47.935 58.345 48.215 59.225 ;
    RECT 44.615 58.345 44.895 59.225 ;
    RECT 41.295 58.345 41.575 59.225 ;
    RECT 37.975 58.345 38.255 59.225 ;
    RECT 34.655 58.345 34.935 59.225 ;
    RECT 117.655 58.345 117.935 59.225 ;
    RECT 114.335 58.345 114.615 59.225 ;
    RECT 111.015 58.345 111.295 59.225 ;
    RECT 107.695 58.345 107.975 59.225 ;
    RECT 104.375 58.345 104.655 59.225 ;
    RECT 101.055 58.345 101.335 59.225 ;
    RECT 97.735 58.345 98.015 59.225 ;
    RECT 94.415 58.345 94.695 59.225 ;
    RECT 91.095 58.345 91.375 59.225 ;
    RECT 87.775 58.345 88.055 59.225 ;
    RECT 84.455 58.345 84.735 59.225 ;
    RECT 81.135 58.345 81.415 59.225 ;
    RECT 77.815 58.345 78.095 59.225 ;
    RECT 74.495 58.345 74.775 59.225 ;
    RECT 71.175 58.345 71.455 59.225 ;
    RECT 31.335 58.345 31.615 59.225 ;
    RECT 67.855 58.345 68.135 59.225 ;
    RECT 28.015 58.345 28.295 59.225 ;
    RECT 24.695 58.345 24.975 59.225 ;
    RECT 21.375 58.345 21.655 59.225 ;
    RECT 18.055 58.345 18.335 59.225 ;
    RECT 14.735 58.345 15.015 59.225 ;
    RECT 11.415 58.345 11.695 59.225 ;
    RECT 8.095 58.345 8.375 59.225 ;
    RECT 4.775 58.345 5.055 59.225 ;
    RECT 1.455 58.345 1.735 59.225 ;
    RECT 64.535 58.345 64.815 59.225 ;
    RECT 61.215 57.625 61.495 58.505 ;
    RECT 57.895 57.625 58.175 58.505 ;
    RECT 54.575 57.625 54.855 58.505 ;
    RECT 51.255 57.625 51.535 58.505 ;
    RECT 47.935 57.625 48.215 58.505 ;
    RECT 44.615 57.625 44.895 58.505 ;
    RECT 41.295 57.625 41.575 58.505 ;
    RECT 37.975 57.625 38.255 58.505 ;
    RECT 34.655 57.625 34.935 58.505 ;
    RECT 117.655 57.625 117.935 58.505 ;
    RECT 114.335 57.625 114.615 58.505 ;
    RECT 111.015 57.625 111.295 58.505 ;
    RECT 107.695 57.625 107.975 58.505 ;
    RECT 104.375 57.625 104.655 58.505 ;
    RECT 101.055 57.625 101.335 58.505 ;
    RECT 97.735 57.625 98.015 58.505 ;
    RECT 94.415 57.625 94.695 58.505 ;
    RECT 91.095 57.625 91.375 58.505 ;
    RECT 87.775 57.625 88.055 58.505 ;
    RECT 84.455 57.625 84.735 58.505 ;
    RECT 81.135 57.625 81.415 58.505 ;
    RECT 77.815 57.625 78.095 58.505 ;
    RECT 74.495 57.625 74.775 58.505 ;
    RECT 71.175 57.625 71.455 58.505 ;
    RECT 31.335 57.625 31.615 58.505 ;
    RECT 67.855 57.625 68.135 58.505 ;
    RECT 28.015 57.625 28.295 58.505 ;
    RECT 24.695 57.625 24.975 58.505 ;
    RECT 21.375 57.625 21.655 58.505 ;
    RECT 18.055 57.625 18.335 58.505 ;
    RECT 14.735 57.625 15.015 58.505 ;
    RECT 11.415 57.625 11.695 58.505 ;
    RECT 8.095 57.625 8.375 58.505 ;
    RECT 4.775 57.625 5.055 58.505 ;
    RECT 1.455 57.625 1.735 58.505 ;
    RECT 64.535 57.625 64.815 58.505 ;
    RECT 117.655 98.765 117.935 100.295 ;
    RECT 114.335 98.765 114.615 100.295 ;
    RECT 111.015 98.765 111.295 100.295 ;
    RECT 107.695 98.765 107.975 100.295 ;
    RECT 104.375 98.765 104.655 100.295 ;
    RECT 101.055 98.765 101.335 100.295 ;
    RECT 97.735 98.765 98.015 100.295 ;
    RECT 94.415 98.765 94.695 100.295 ;
    RECT 91.095 98.765 91.375 100.295 ;
    RECT 87.775 98.765 88.055 100.295 ;
    RECT 84.455 98.765 84.735 100.295 ;
    RECT 81.135 98.765 81.415 100.295 ;
    RECT 77.815 98.765 78.095 100.295 ;
    RECT 74.495 98.765 74.775 100.295 ;
    RECT 71.175 98.765 71.455 100.295 ;
    RECT 67.855 98.765 68.135 100.295 ;
    RECT 64.535 98.765 64.815 100.295 ;
    RECT 61.215 98.765 61.495 100.295 ;
    RECT 57.895 98.765 58.175 100.295 ;
    RECT 54.575 98.765 54.855 100.295 ;
    RECT 51.255 98.765 51.535 100.295 ;
    RECT 47.935 98.765 48.215 100.295 ;
    RECT 44.615 98.765 44.895 100.295 ;
    RECT 41.295 98.765 41.575 100.295 ;
    RECT 37.975 98.765 38.255 100.295 ;
    RECT 34.655 98.765 34.935 100.295 ;
    RECT 31.335 98.765 31.615 100.295 ;
    RECT 28.015 98.765 28.295 100.295 ;
    RECT 24.695 98.765 24.975 100.295 ;
    RECT 21.375 98.765 21.655 100.295 ;
    RECT 18.055 98.765 18.335 100.295 ;
    RECT 14.735 98.765 15.015 100.295 ;
    RECT 11.415 98.765 11.695 100.295 ;
    RECT 8.095 98.765 8.375 100.295 ;
    RECT 4.775 98.765 5.055 100.295 ;
    RECT 1.455 98.765 1.735 100.295 ;
    RECT 61.215 54.745 61.495 55.625 ;
    RECT 57.895 54.745 58.175 55.625 ;
    RECT 54.575 54.745 54.855 55.625 ;
    RECT 51.255 54.745 51.535 55.625 ;
    RECT 47.935 54.745 48.215 55.625 ;
    RECT 44.615 54.745 44.895 55.625 ;
    RECT 41.295 54.745 41.575 55.625 ;
    RECT 37.975 54.745 38.255 55.625 ;
    RECT 34.655 54.745 34.935 55.625 ;
    RECT 117.655 54.745 117.935 55.625 ;
    RECT 114.335 54.745 114.615 55.625 ;
    RECT 111.015 54.745 111.295 55.625 ;
    RECT 107.695 54.745 107.975 55.625 ;
    RECT 104.375 54.745 104.655 55.625 ;
    RECT 101.055 54.745 101.335 55.625 ;
    RECT 97.735 54.745 98.015 55.625 ;
    RECT 94.415 54.745 94.695 55.625 ;
    RECT 91.095 54.745 91.375 55.625 ;
    RECT 87.775 54.745 88.055 55.625 ;
    RECT 84.455 54.745 84.735 55.625 ;
    RECT 81.135 54.745 81.415 55.625 ;
    RECT 77.815 54.745 78.095 55.625 ;
    RECT 74.495 54.745 74.775 55.625 ;
    RECT 71.175 54.745 71.455 55.625 ;
    RECT 31.335 54.745 31.615 55.625 ;
    RECT 67.855 54.745 68.135 55.625 ;
    RECT 28.015 54.745 28.295 55.625 ;
    RECT 24.695 54.745 24.975 55.625 ;
    RECT 21.375 54.745 21.655 55.625 ;
    RECT 18.055 54.745 18.335 55.625 ;
    RECT 14.735 54.745 15.015 55.625 ;
    RECT 11.415 54.745 11.695 55.625 ;
    RECT 8.095 54.745 8.375 55.625 ;
    RECT 4.775 54.745 5.055 55.625 ;
    RECT 1.455 54.745 1.735 55.625 ;
    RECT 64.535 54.745 64.815 55.625 ;
    RECT 61.215 55.465 61.495 56.345 ;
    RECT 57.895 55.465 58.175 56.345 ;
    RECT 54.575 55.465 54.855 56.345 ;
    RECT 51.255 55.465 51.535 56.345 ;
    RECT 47.935 55.465 48.215 56.345 ;
    RECT 44.615 55.465 44.895 56.345 ;
    RECT 41.295 55.465 41.575 56.345 ;
    RECT 37.975 55.465 38.255 56.345 ;
    RECT 34.655 55.465 34.935 56.345 ;
    RECT 117.655 55.465 117.935 56.345 ;
    RECT 114.335 55.465 114.615 56.345 ;
    RECT 111.015 55.465 111.295 56.345 ;
    RECT 107.695 55.465 107.975 56.345 ;
    RECT 104.375 55.465 104.655 56.345 ;
    RECT 101.055 55.465 101.335 56.345 ;
    RECT 97.735 55.465 98.015 56.345 ;
    RECT 94.415 55.465 94.695 56.345 ;
    RECT 91.095 55.465 91.375 56.345 ;
    RECT 87.775 55.465 88.055 56.345 ;
    RECT 84.455 55.465 84.735 56.345 ;
    RECT 81.135 55.465 81.415 56.345 ;
    RECT 77.815 55.465 78.095 56.345 ;
    RECT 74.495 55.465 74.775 56.345 ;
    RECT 71.175 55.465 71.455 56.345 ;
    RECT 31.335 55.465 31.615 56.345 ;
    RECT 67.855 55.465 68.135 56.345 ;
    RECT 28.015 55.465 28.295 56.345 ;
    RECT 24.695 55.465 24.975 56.345 ;
    RECT 21.375 55.465 21.655 56.345 ;
    RECT 18.055 55.465 18.335 56.345 ;
    RECT 14.735 55.465 15.015 56.345 ;
    RECT 11.415 55.465 11.695 56.345 ;
    RECT 8.095 55.465 8.375 56.345 ;
    RECT 4.775 55.465 5.055 56.345 ;
    RECT 1.455 55.465 1.735 56.345 ;
    RECT 64.535 55.465 64.815 56.345 ;
    RECT 61.215 97.245 61.495 98.125 ;
    RECT 57.895 97.245 58.175 98.125 ;
    RECT 54.575 97.245 54.855 98.125 ;
    RECT 51.255 97.245 51.535 98.125 ;
    RECT 47.935 97.245 48.215 98.125 ;
    RECT 44.615 97.245 44.895 98.125 ;
    RECT 41.295 97.245 41.575 98.125 ;
    RECT 37.975 97.245 38.255 98.125 ;
    RECT 34.655 97.245 34.935 98.125 ;
    RECT 117.655 97.245 117.935 98.125 ;
    RECT 114.335 97.245 114.615 98.125 ;
    RECT 111.015 97.245 111.295 98.125 ;
    RECT 107.695 97.245 107.975 98.125 ;
    RECT 104.375 97.245 104.655 98.125 ;
    RECT 101.055 97.245 101.335 98.125 ;
    RECT 97.735 97.245 98.015 98.125 ;
    RECT 94.415 97.245 94.695 98.125 ;
    RECT 91.095 97.245 91.375 98.125 ;
    RECT 87.775 97.245 88.055 98.125 ;
    RECT 84.455 97.245 84.735 98.125 ;
    RECT 81.135 97.245 81.415 98.125 ;
    RECT 77.815 97.245 78.095 98.125 ;
    RECT 74.495 97.245 74.775 98.125 ;
    RECT 71.175 97.245 71.455 98.125 ;
    RECT 31.335 97.245 31.615 98.125 ;
    RECT 67.855 97.245 68.135 98.125 ;
    RECT 28.015 97.245 28.295 98.125 ;
    RECT 24.695 97.245 24.975 98.125 ;
    RECT 21.375 97.245 21.655 98.125 ;
    RECT 18.055 97.245 18.335 98.125 ;
    RECT 14.735 97.245 15.015 98.125 ;
    RECT 11.415 97.245 11.695 98.125 ;
    RECT 8.095 97.245 8.375 98.125 ;
    RECT 4.775 97.245 5.055 98.125 ;
    RECT 1.455 97.245 1.735 98.125 ;
    RECT 64.535 97.245 64.815 98.125 ;
    RECT 61.215 96.525 61.495 97.405 ;
    RECT 57.895 96.525 58.175 97.405 ;
    RECT 54.575 96.525 54.855 97.405 ;
    RECT 51.255 96.525 51.535 97.405 ;
    RECT 47.935 96.525 48.215 97.405 ;
    RECT 44.615 96.525 44.895 97.405 ;
    RECT 41.295 96.525 41.575 97.405 ;
    RECT 37.975 96.525 38.255 97.405 ;
    RECT 34.655 96.525 34.935 97.405 ;
    RECT 117.655 96.525 117.935 97.405 ;
    RECT 114.335 96.525 114.615 97.405 ;
    RECT 111.015 96.525 111.295 97.405 ;
    RECT 107.695 96.525 107.975 97.405 ;
    RECT 104.375 96.525 104.655 97.405 ;
    RECT 101.055 96.525 101.335 97.405 ;
    RECT 97.735 96.525 98.015 97.405 ;
    RECT 94.415 96.525 94.695 97.405 ;
    RECT 91.095 96.525 91.375 97.405 ;
    RECT 87.775 96.525 88.055 97.405 ;
    RECT 84.455 96.525 84.735 97.405 ;
    RECT 81.135 96.525 81.415 97.405 ;
    RECT 77.815 96.525 78.095 97.405 ;
    RECT 74.495 96.525 74.775 97.405 ;
    RECT 71.175 96.525 71.455 97.405 ;
    RECT 31.335 96.525 31.615 97.405 ;
    RECT 67.855 96.525 68.135 97.405 ;
    RECT 28.015 96.525 28.295 97.405 ;
    RECT 24.695 96.525 24.975 97.405 ;
    RECT 21.375 96.525 21.655 97.405 ;
    RECT 18.055 96.525 18.335 97.405 ;
    RECT 14.735 96.525 15.015 97.405 ;
    RECT 11.415 96.525 11.695 97.405 ;
    RECT 8.095 96.525 8.375 97.405 ;
    RECT 4.775 96.525 5.055 97.405 ;
    RECT 1.455 96.525 1.735 97.405 ;
    RECT 64.535 96.525 64.815 97.405 ;
    RECT 61.215 95.805 61.495 96.685 ;
    RECT 57.895 95.805 58.175 96.685 ;
    RECT 54.575 95.805 54.855 96.685 ;
    RECT 51.255 95.805 51.535 96.685 ;
    RECT 47.935 95.805 48.215 96.685 ;
    RECT 44.615 95.805 44.895 96.685 ;
    RECT 41.295 95.805 41.575 96.685 ;
    RECT 37.975 95.805 38.255 96.685 ;
    RECT 34.655 95.805 34.935 96.685 ;
    RECT 117.655 95.805 117.935 96.685 ;
    RECT 114.335 95.805 114.615 96.685 ;
    RECT 111.015 95.805 111.295 96.685 ;
    RECT 107.695 95.805 107.975 96.685 ;
    RECT 104.375 95.805 104.655 96.685 ;
    RECT 101.055 95.805 101.335 96.685 ;
    RECT 97.735 95.805 98.015 96.685 ;
    RECT 94.415 95.805 94.695 96.685 ;
    RECT 91.095 95.805 91.375 96.685 ;
    RECT 87.775 95.805 88.055 96.685 ;
    RECT 84.455 95.805 84.735 96.685 ;
    RECT 81.135 95.805 81.415 96.685 ;
    RECT 77.815 95.805 78.095 96.685 ;
    RECT 74.495 95.805 74.775 96.685 ;
    RECT 71.175 95.805 71.455 96.685 ;
    RECT 31.335 95.805 31.615 96.685 ;
    RECT 67.855 95.805 68.135 96.685 ;
    RECT 28.015 95.805 28.295 96.685 ;
    RECT 24.695 95.805 24.975 96.685 ;
    RECT 21.375 95.805 21.655 96.685 ;
    RECT 18.055 95.805 18.335 96.685 ;
    RECT 14.735 95.805 15.015 96.685 ;
    RECT 11.415 95.805 11.695 96.685 ;
    RECT 8.095 95.805 8.375 96.685 ;
    RECT 4.775 95.805 5.055 96.685 ;
    RECT 1.455 95.805 1.735 96.685 ;
    RECT 64.535 95.805 64.815 96.685 ;
    RECT 61.215 95.085 61.495 95.965 ;
    RECT 57.895 95.085 58.175 95.965 ;
    RECT 54.575 95.085 54.855 95.965 ;
    RECT 51.255 95.085 51.535 95.965 ;
    RECT 47.935 95.085 48.215 95.965 ;
    RECT 44.615 95.085 44.895 95.965 ;
    RECT 41.295 95.085 41.575 95.965 ;
    RECT 37.975 95.085 38.255 95.965 ;
    RECT 34.655 95.085 34.935 95.965 ;
    RECT 117.655 95.085 117.935 95.965 ;
    RECT 114.335 95.085 114.615 95.965 ;
    RECT 111.015 95.085 111.295 95.965 ;
    RECT 107.695 95.085 107.975 95.965 ;
    RECT 104.375 95.085 104.655 95.965 ;
    RECT 101.055 95.085 101.335 95.965 ;
    RECT 97.735 95.085 98.015 95.965 ;
    RECT 94.415 95.085 94.695 95.965 ;
    RECT 91.095 95.085 91.375 95.965 ;
    RECT 87.775 95.085 88.055 95.965 ;
    RECT 84.455 95.085 84.735 95.965 ;
    RECT 81.135 95.085 81.415 95.965 ;
    RECT 77.815 95.085 78.095 95.965 ;
    RECT 74.495 95.085 74.775 95.965 ;
    RECT 71.175 95.085 71.455 95.965 ;
    RECT 31.335 95.085 31.615 95.965 ;
    RECT 67.855 95.085 68.135 95.965 ;
    RECT 28.015 95.085 28.295 95.965 ;
    RECT 24.695 95.085 24.975 95.965 ;
    RECT 21.375 95.085 21.655 95.965 ;
    RECT 18.055 95.085 18.335 95.965 ;
    RECT 14.735 95.085 15.015 95.965 ;
    RECT 11.415 95.085 11.695 95.965 ;
    RECT 8.095 95.085 8.375 95.965 ;
    RECT 4.775 95.085 5.055 95.965 ;
    RECT 1.455 95.085 1.735 95.965 ;
    RECT 64.535 95.085 64.815 95.965 ;
    RECT 61.215 94.365 61.495 95.245 ;
    RECT 57.895 94.365 58.175 95.245 ;
    RECT 54.575 94.365 54.855 95.245 ;
    RECT 51.255 94.365 51.535 95.245 ;
    RECT 47.935 94.365 48.215 95.245 ;
    RECT 44.615 94.365 44.895 95.245 ;
    RECT 41.295 94.365 41.575 95.245 ;
    RECT 37.975 94.365 38.255 95.245 ;
    RECT 34.655 94.365 34.935 95.245 ;
    RECT 117.655 94.365 117.935 95.245 ;
    RECT 114.335 94.365 114.615 95.245 ;
    RECT 111.015 94.365 111.295 95.245 ;
    RECT 107.695 94.365 107.975 95.245 ;
    RECT 104.375 94.365 104.655 95.245 ;
    RECT 101.055 94.365 101.335 95.245 ;
    RECT 97.735 94.365 98.015 95.245 ;
    RECT 94.415 94.365 94.695 95.245 ;
    RECT 91.095 94.365 91.375 95.245 ;
    RECT 87.775 94.365 88.055 95.245 ;
    RECT 84.455 94.365 84.735 95.245 ;
    RECT 81.135 94.365 81.415 95.245 ;
    RECT 77.815 94.365 78.095 95.245 ;
    RECT 74.495 94.365 74.775 95.245 ;
    RECT 71.175 94.365 71.455 95.245 ;
    RECT 31.335 94.365 31.615 95.245 ;
    RECT 67.855 94.365 68.135 95.245 ;
    RECT 28.015 94.365 28.295 95.245 ;
    RECT 24.695 94.365 24.975 95.245 ;
    RECT 21.375 94.365 21.655 95.245 ;
    RECT 18.055 94.365 18.335 95.245 ;
    RECT 14.735 94.365 15.015 95.245 ;
    RECT 11.415 94.365 11.695 95.245 ;
    RECT 8.095 94.365 8.375 95.245 ;
    RECT 4.775 94.365 5.055 95.245 ;
    RECT 1.455 94.365 1.735 95.245 ;
    RECT 64.535 94.365 64.815 95.245 ;
    RECT 61.215 56.905 61.495 57.785 ;
    RECT 57.895 56.905 58.175 57.785 ;
    RECT 54.575 56.905 54.855 57.785 ;
    RECT 51.255 56.905 51.535 57.785 ;
    RECT 47.935 56.905 48.215 57.785 ;
    RECT 44.615 56.905 44.895 57.785 ;
    RECT 41.295 56.905 41.575 57.785 ;
    RECT 37.975 56.905 38.255 57.785 ;
    RECT 34.655 56.905 34.935 57.785 ;
    RECT 117.655 56.905 117.935 57.785 ;
    RECT 114.335 56.905 114.615 57.785 ;
    RECT 111.015 56.905 111.295 57.785 ;
    RECT 107.695 56.905 107.975 57.785 ;
    RECT 104.375 56.905 104.655 57.785 ;
    RECT 101.055 56.905 101.335 57.785 ;
    RECT 97.735 56.905 98.015 57.785 ;
    RECT 94.415 56.905 94.695 57.785 ;
    RECT 91.095 56.905 91.375 57.785 ;
    RECT 87.775 56.905 88.055 57.785 ;
    RECT 84.455 56.905 84.735 57.785 ;
    RECT 81.135 56.905 81.415 57.785 ;
    RECT 77.815 56.905 78.095 57.785 ;
    RECT 74.495 56.905 74.775 57.785 ;
    RECT 71.175 56.905 71.455 57.785 ;
    RECT 31.335 56.905 31.615 57.785 ;
    RECT 67.855 56.905 68.135 57.785 ;
    RECT 28.015 56.905 28.295 57.785 ;
    RECT 24.695 56.905 24.975 57.785 ;
    RECT 21.375 56.905 21.655 57.785 ;
    RECT 18.055 56.905 18.335 57.785 ;
    RECT 14.735 56.905 15.015 57.785 ;
    RECT 11.415 56.905 11.695 57.785 ;
    RECT 8.095 56.905 8.375 57.785 ;
    RECT 4.775 56.905 5.055 57.785 ;
    RECT 1.455 56.905 1.735 57.785 ;
    RECT 64.535 56.905 64.815 57.785 ;
    RECT 61.215 54.025 61.495 54.905 ;
    RECT 57.895 54.025 58.175 54.905 ;
    RECT 54.575 54.025 54.855 54.905 ;
    RECT 51.255 54.025 51.535 54.905 ;
    RECT 47.935 54.025 48.215 54.905 ;
    RECT 44.615 54.025 44.895 54.905 ;
    RECT 41.295 54.025 41.575 54.905 ;
    RECT 37.975 54.025 38.255 54.905 ;
    RECT 34.655 54.025 34.935 54.905 ;
    RECT 117.655 54.025 117.935 54.905 ;
    RECT 114.335 54.025 114.615 54.905 ;
    RECT 111.015 54.025 111.295 54.905 ;
    RECT 107.695 54.025 107.975 54.905 ;
    RECT 104.375 54.025 104.655 54.905 ;
    RECT 101.055 54.025 101.335 54.905 ;
    RECT 97.735 54.025 98.015 54.905 ;
    RECT 94.415 54.025 94.695 54.905 ;
    RECT 91.095 54.025 91.375 54.905 ;
    RECT 87.775 54.025 88.055 54.905 ;
    RECT 84.455 54.025 84.735 54.905 ;
    RECT 81.135 54.025 81.415 54.905 ;
    RECT 77.815 54.025 78.095 54.905 ;
    RECT 74.495 54.025 74.775 54.905 ;
    RECT 71.175 54.025 71.455 54.905 ;
    RECT 31.335 54.025 31.615 54.905 ;
    RECT 67.855 54.025 68.135 54.905 ;
    RECT 28.015 54.025 28.295 54.905 ;
    RECT 24.695 54.025 24.975 54.905 ;
    RECT 21.375 54.025 21.655 54.905 ;
    RECT 18.055 54.025 18.335 54.905 ;
    RECT 14.735 54.025 15.015 54.905 ;
    RECT 11.415 54.025 11.695 54.905 ;
    RECT 8.095 54.025 8.375 54.905 ;
    RECT 4.775 54.025 5.055 54.905 ;
    RECT 1.455 54.025 1.735 54.905 ;
    RECT 64.535 54.025 64.815 54.905 ;
    RECT 61.215 53.305 61.495 54.185 ;
    RECT 57.895 53.305 58.175 54.185 ;
    RECT 54.575 53.305 54.855 54.185 ;
    RECT 51.255 53.305 51.535 54.185 ;
    RECT 47.935 53.305 48.215 54.185 ;
    RECT 44.615 53.305 44.895 54.185 ;
    RECT 41.295 53.305 41.575 54.185 ;
    RECT 37.975 53.305 38.255 54.185 ;
    RECT 34.655 53.305 34.935 54.185 ;
    RECT 117.655 53.305 117.935 54.185 ;
    RECT 114.335 53.305 114.615 54.185 ;
    RECT 111.015 53.305 111.295 54.185 ;
    RECT 107.695 53.305 107.975 54.185 ;
    RECT 104.375 53.305 104.655 54.185 ;
    RECT 101.055 53.305 101.335 54.185 ;
    RECT 97.735 53.305 98.015 54.185 ;
    RECT 94.415 53.305 94.695 54.185 ;
    RECT 91.095 53.305 91.375 54.185 ;
    RECT 87.775 53.305 88.055 54.185 ;
    RECT 84.455 53.305 84.735 54.185 ;
    RECT 81.135 53.305 81.415 54.185 ;
    RECT 77.815 53.305 78.095 54.185 ;
    RECT 74.495 53.305 74.775 54.185 ;
    RECT 71.175 53.305 71.455 54.185 ;
    RECT 31.335 53.305 31.615 54.185 ;
    RECT 67.855 53.305 68.135 54.185 ;
    RECT 28.015 53.305 28.295 54.185 ;
    RECT 24.695 53.305 24.975 54.185 ;
    RECT 21.375 53.305 21.655 54.185 ;
    RECT 18.055 53.305 18.335 54.185 ;
    RECT 14.735 53.305 15.015 54.185 ;
    RECT 11.415 53.305 11.695 54.185 ;
    RECT 8.095 53.305 8.375 54.185 ;
    RECT 4.775 53.305 5.055 54.185 ;
    RECT 1.455 53.305 1.735 54.185 ;
    RECT 64.535 53.305 64.815 54.185 ;
    RECT 134.71 49.785 134.79 50.505 ;
    RECT 139.7 49.785 139.97 50.505 ;
    RECT 134.71 49.065 134.79 49.785 ;
    RECT 139.7 49.065 139.97 49.785 ;
    RECT 134.71 48.345 134.79 49.065 ;
    RECT 139.7 48.345 139.97 49.065 ;
    RECT 134.71 47.625 134.79 48.345 ;
    RECT 139.7 47.625 139.97 48.345 ;
    RECT 134.71 46.905 134.79 47.625 ;
    RECT 139.7 46.905 139.97 47.625 ;
    RECT 134.71 46.185 134.79 46.905 ;
    RECT 139.7 46.185 139.97 46.905 ;
    RECT 134.71 45.465 134.79 46.185 ;
    RECT 139.7 45.465 139.97 46.185 ;
    RECT 134.71 44.745 134.79 45.465 ;
    RECT 139.7 44.745 139.97 45.465 ;
    RECT 134.71 44.025 134.79 44.745 ;
    RECT 139.7 44.025 139.97 44.745 ;
    RECT 134.71 43.305 134.79 44.025 ;
    RECT 139.7 43.305 139.97 44.025 ;
    RECT 134.71 42.585 134.79 43.305 ;
    RECT 139.7 42.585 139.97 43.305 ;
    RECT 134.71 41.865 134.79 42.585 ;
    RECT 139.7 41.865 139.97 42.585 ;
    RECT 134.71 41.145 134.79 41.865 ;
    RECT 139.7 41.145 139.97 41.865 ;
    RECT 134.71 40.425 134.79 41.145 ;
    RECT 139.7 40.425 139.97 41.145 ;
    RECT 134.71 39.705 134.79 40.425 ;
    RECT 139.7 39.705 139.97 40.425 ;
    RECT 134.71 38.985 134.79 39.705 ;
    RECT 139.7 38.985 139.97 39.705 ;
    RECT 134.71 38.265 134.79 38.985 ;
    RECT 139.7 38.265 139.97 38.985 ;
    RECT 134.71 37.545 134.79 38.265 ;
    RECT 139.7 37.545 139.97 38.265 ;
    RECT 128.335 14.505 128.545 32.145 ;
    RECT 134.71 14.55 134.79 37.69 ;
    RECT 139.7 14.34 139.97 37.545 ;
    RECT 134.71 98.045 134.79 98.765 ;
    RECT 139.7 98.045 139.97 98.765 ;
    RECT 134.71 97.325 134.79 98.045 ;
    RECT 139.7 97.325 139.97 98.045 ;
    RECT 134.71 96.605 134.79 97.325 ;
    RECT 139.7 96.605 139.97 97.325 ;
    RECT 134.71 95.885 134.79 96.605 ;
    RECT 139.7 95.885 139.97 96.605 ;
    RECT 121.67 99.8 121.86 100.295 ;
    RECT 134.71 98.765 134.79 100.225 ;
    RECT 139.7 98.765 139.97 100.295 ;
    RECT 134.71 95.165 134.79 95.885 ;
    RECT 139.7 95.165 139.97 95.885 ;
    RECT 134.71 94.445 134.79 95.165 ;
    RECT 139.7 94.445 139.97 95.165 ;
    RECT 134.71 93.725 134.79 94.445 ;
    RECT 139.7 93.725 139.97 94.445 ;
    RECT 134.71 93.005 134.79 93.725 ;
    RECT 139.7 93.005 139.97 93.725 ;
    RECT 134.71 92.285 134.79 93.005 ;
    RECT 139.7 92.285 139.97 93.005 ;
    RECT 134.71 91.565 134.79 92.285 ;
    RECT 139.7 91.565 139.97 92.285 ;
    RECT 134.71 90.845 134.79 91.565 ;
    RECT 139.7 90.845 139.97 91.565 ;
    RECT 134.71 90.125 134.79 90.845 ;
    RECT 139.7 90.125 139.97 90.845 ;
    RECT 134.71 89.405 134.79 90.125 ;
    RECT 139.7 89.405 139.97 90.125 ;
    RECT 134.71 88.685 134.79 89.405 ;
    RECT 139.7 88.685 139.97 89.405 ;
    RECT 134.71 60.585 134.79 61.325 ;
    RECT 139.7 60.585 139.97 61.325 ;
    RECT 134.71 87.965 134.79 88.685 ;
    RECT 139.7 87.965 139.97 88.685 ;
    RECT 134.71 87.245 134.79 87.965 ;
    RECT 139.7 87.245 139.97 87.965 ;
    RECT 134.71 86.525 134.79 87.245 ;
    RECT 139.7 86.525 139.97 87.245 ;
    RECT 134.71 85.805 134.79 86.525 ;
    RECT 139.7 85.805 139.97 86.525 ;
    RECT 134.71 85.085 134.79 85.805 ;
    RECT 139.7 85.085 139.97 85.805 ;
    RECT 134.71 84.365 134.79 85.085 ;
    RECT 139.7 84.365 139.97 85.085 ;
    RECT 134.71 83.645 134.79 84.365 ;
    RECT 139.7 83.645 139.97 84.365 ;
    RECT 134.71 82.925 134.79 83.645 ;
    RECT 139.7 82.925 139.97 83.645 ;
    RECT 134.71 82.205 134.79 82.925 ;
    RECT 139.7 82.205 139.97 82.925 ;
    RECT 134.71 81.485 134.79 82.205 ;
    RECT 139.7 81.485 139.97 82.205 ;
    RECT 134.71 80.765 134.79 81.485 ;
    RECT 139.7 80.765 139.97 81.485 ;
    RECT 134.71 80.045 134.79 80.765 ;
    RECT 139.7 80.045 139.97 80.765 ;
    RECT 134.71 79.325 134.79 80.045 ;
    RECT 139.7 79.325 139.97 80.045 ;
    RECT 134.71 78.605 134.79 79.325 ;
    RECT 139.7 78.605 139.97 79.325 ;
    RECT 134.71 77.885 134.79 78.605 ;
    RECT 139.7 77.885 139.97 78.605 ;
    RECT 134.71 77.165 134.79 77.885 ;
    RECT 139.7 77.165 139.97 77.885 ;
    RECT 134.71 76.445 134.79 77.165 ;
    RECT 139.7 76.445 139.97 77.165 ;
    RECT 134.71 75.725 134.79 76.445 ;
    RECT 139.7 75.725 139.97 76.445 ;
    RECT 134.71 75.005 134.79 75.725 ;
    RECT 139.7 75.005 139.97 75.725 ;
    RECT 134.71 74.285 134.79 75.005 ;
    RECT 139.7 74.285 139.97 75.005 ;
    RECT 134.71 73.565 134.79 74.285 ;
    RECT 139.7 73.565 139.97 74.285 ;
    RECT 134.71 72.845 134.79 73.565 ;
    RECT 139.7 72.845 139.97 73.565 ;
    RECT 134.71 72.125 134.79 72.845 ;
    RECT 139.7 72.125 139.97 72.845 ;
    RECT 134.71 71.405 134.79 72.125 ;
    RECT 139.7 71.405 139.97 72.125 ;
    RECT 134.71 70.685 134.79 71.405 ;
    RECT 139.7 70.685 139.97 71.405 ;
    RECT 134.71 69.965 134.79 70.685 ;
    RECT 139.7 69.965 139.97 70.685 ;
    RECT 134.71 69.245 134.79 69.965 ;
    RECT 139.7 69.245 139.97 69.965 ;
    RECT 134.71 68.525 134.79 69.245 ;
    RECT 139.7 68.525 139.97 69.245 ;
    RECT 134.71 67.805 134.79 68.525 ;
    RECT 139.7 67.805 139.97 68.525 ;
    RECT 134.71 67.085 134.79 67.805 ;
    RECT 139.7 67.085 139.97 67.805 ;
    RECT 134.71 66.365 134.79 67.085 ;
    RECT 139.7 66.365 139.97 67.085 ;
    RECT 134.71 65.645 134.79 66.365 ;
    RECT 139.7 65.645 139.97 66.365 ;
    RECT 134.71 64.925 134.79 65.645 ;
    RECT 139.7 64.925 139.97 65.645 ;
    RECT 134.71 64.205 134.79 64.925 ;
    RECT 139.7 64.205 139.97 64.925 ;
    RECT 134.71 63.485 134.79 64.205 ;
    RECT 139.7 63.485 139.97 64.205 ;
    RECT 134.71 62.765 134.79 63.485 ;
    RECT 139.7 62.765 139.97 63.485 ;
    RECT 134.71 62.045 134.79 62.765 ;
    RECT 139.7 62.045 139.97 62.765 ;
    RECT 134.71 61.325 134.79 62.045 ;
    RECT 139.7 61.325 139.97 62.045 ;
    RECT 134.71 59.865 134.79 60.585 ;
    RECT 139.7 59.865 139.97 60.585 ;
    RECT 134.71 59.145 134.79 59.865 ;
    RECT 139.7 59.145 139.97 59.865 ;
    RECT 134.71 58.425 134.79 59.145 ;
    RECT 139.7 58.425 139.97 59.145 ;
    RECT 134.71 57.705 134.79 58.425 ;
    RECT 139.7 57.705 139.97 58.425 ;
    RECT 134.71 56.985 134.79 57.705 ;
    RECT 139.7 56.985 139.97 57.705 ;
    RECT 134.71 56.265 134.79 56.985 ;
    RECT 139.7 56.265 139.97 56.985 ;
    RECT 134.71 55.545 134.79 56.265 ;
    RECT 139.7 55.545 139.97 56.265 ;
    RECT 134.71 54.825 134.79 55.545 ;
    RECT 139.7 54.825 139.97 55.545 ;
    RECT 134.71 54.105 134.79 54.825 ;
    RECT 139.7 54.105 139.97 54.825 ;
    RECT 134.71 53.385 134.79 54.105 ;
    RECT 139.7 53.385 139.97 54.105 ;
    RECT 134.71 52.665 134.79 53.385 ;
    RECT 139.7 52.665 139.97 53.385 ;
    RECT 134.71 51.945 134.79 52.665 ;
    RECT 139.7 51.945 139.97 52.665 ;
    RECT 134.71 51.225 134.79 51.945 ;
    RECT 139.7 51.225 139.97 51.945 ;
    RECT 134.71 50.505 134.79 51.225 ;
    RECT 139.7 50.505 139.97 51.225 ;
    RECT 180.325 12.695 180.605 12.975 ;
    RECT 180.39 4.14 180.46 7.295 ;
    RECT 177.005 12.695 177.285 12.975 ;
    RECT 177.07 4.14 177.14 7.295 ;
    RECT 173.685 12.695 173.965 12.975 ;
    RECT 173.75 4.14 173.82 7.295 ;
    RECT 170.365 12.695 170.645 12.975 ;
    RECT 170.43 4.14 170.5 7.295 ;
    RECT 167.045 12.695 167.325 12.975 ;
    RECT 167.11 4.14 167.18 7.295 ;
    RECT 163.725 12.695 164.005 12.975 ;
    RECT 163.79 4.14 163.86 7.295 ;
    RECT 160.405 12.695 160.685 12.975 ;
    RECT 160.47 4.14 160.54 7.295 ;
    RECT 157.085 12.695 157.365 12.975 ;
    RECT 157.15 4.14 157.22 7.295 ;
    RECT 153.765 12.695 154.045 12.975 ;
    RECT 153.83 4.14 153.9 7.295 ;
    RECT 266.645 12.695 266.925 12.975 ;
    RECT 266.71 4.14 266.78 7.295 ;
    RECT 150.445 12.695 150.725 12.975 ;
    RECT 150.51 4.14 150.58 7.295 ;
    RECT 263.325 12.695 263.605 12.975 ;
    RECT 263.39 4.14 263.46 7.295 ;
    RECT 260.005 12.695 260.285 12.975 ;
    RECT 260.07 4.14 260.14 7.295 ;
    RECT 256.685 12.695 256.965 12.975 ;
    RECT 256.75 4.14 256.82 7.295 ;
    RECT 253.365 12.695 253.645 12.975 ;
    RECT 253.43 4.14 253.5 7.295 ;
    RECT 250.045 12.695 250.325 12.975 ;
    RECT 250.11 4.14 250.18 7.295 ;
    RECT 246.725 12.695 247.005 12.975 ;
    RECT 246.79 4.14 246.86 7.295 ;
    RECT 243.405 12.695 243.685 12.975 ;
    RECT 243.47 4.14 243.54 7.295 ;
    RECT 240.085 12.695 240.365 12.975 ;
    RECT 240.15 4.14 240.22 7.295 ;
    RECT 236.765 12.695 237.045 12.975 ;
    RECT 236.83 4.14 236.9 7.295 ;
    RECT 233.445 12.695 233.725 12.975 ;
    RECT 233.51 4.14 233.58 7.295 ;
    RECT 230.125 12.695 230.405 12.975 ;
    RECT 230.19 4.14 230.26 7.295 ;
    RECT 226.805 12.695 227.085 12.975 ;
    RECT 226.87 4.14 226.94 7.295 ;
    RECT 223.485 12.695 223.765 12.975 ;
    RECT 223.55 4.14 223.62 7.295 ;
    RECT 220.165 12.695 220.445 12.975 ;
    RECT 220.23 4.14 220.3 7.295 ;
    RECT 216.845 12.695 217.125 12.975 ;
    RECT 216.91 4.14 216.98 7.295 ;
    RECT 213.525 12.695 213.805 12.975 ;
    RECT 213.59 4.14 213.66 7.295 ;
    RECT 210.205 12.695 210.485 12.975 ;
    RECT 210.27 4.14 210.34 7.295 ;
    RECT 206.885 12.695 207.165 12.975 ;
    RECT 206.95 4.14 207.02 7.295 ;
    RECT 203.565 12.695 203.845 12.975 ;
    RECT 203.63 4.14 203.7 7.295 ;
    RECT 200.245 12.695 200.525 12.975 ;
    RECT 200.31 4.14 200.38 7.295 ;
    RECT 196.925 12.695 197.205 12.975 ;
    RECT 196.99 4.14 197.06 7.295 ;
    RECT 193.605 12.695 193.885 12.975 ;
    RECT 193.67 4.14 193.74 7.295 ;
    RECT 190.285 12.695 190.565 12.975 ;
    RECT 190.35 4.14 190.42 7.295 ;
    RECT 186.965 12.695 187.245 12.975 ;
    RECT 187.03 4.14 187.1 7.295 ;
    RECT 183.645 12.695 183.925 12.975 ;
    RECT 183.71 4.14 183.78 7.295 ;
    RECT 213.525 12.975 213.805 14.505 ;
    RECT 210.205 12.975 210.485 14.505 ;
    RECT 206.885 12.975 207.165 14.505 ;
    RECT 203.565 12.975 203.845 14.505 ;
    RECT 200.245 12.975 200.525 14.505 ;
    RECT 196.925 12.975 197.205 14.505 ;
    RECT 193.605 12.975 193.885 14.505 ;
    RECT 190.285 12.975 190.565 14.505 ;
    RECT 186.965 12.975 187.245 14.505 ;
    RECT 183.645 12.975 183.925 14.505 ;
    RECT 180.325 12.975 180.605 14.505 ;
    RECT 177.005 12.975 177.285 14.505 ;
    RECT 173.685 12.975 173.965 14.505 ;
    RECT 170.365 12.975 170.645 14.505 ;
    RECT 167.045 12.975 167.325 14.505 ;
    RECT 163.725 12.975 164.005 14.505 ;
    RECT 160.405 12.975 160.685 14.505 ;
    RECT 157.085 12.975 157.365 14.505 ;
    RECT 153.765 12.975 154.045 14.505 ;
    RECT 150.445 12.975 150.725 14.505 ;
    RECT 266.645 12.975 266.925 14.505 ;
    RECT 263.325 12.975 263.605 14.505 ;
    RECT 260.005 12.975 260.285 14.505 ;
    RECT 256.685 12.975 256.965 14.505 ;
    RECT 253.365 12.975 253.645 14.505 ;
    RECT 250.045 12.975 250.325 14.505 ;
    RECT 246.725 12.975 247.005 14.505 ;
    RECT 243.405 12.975 243.685 14.505 ;
    RECT 240.085 12.975 240.365 14.505 ;
    RECT 236.765 12.975 237.045 14.505 ;
    RECT 233.445 12.975 233.725 14.505 ;
    RECT 230.125 12.975 230.405 14.505 ;
    RECT 226.805 12.975 227.085 14.505 ;
    RECT 223.485 12.975 223.765 14.505 ;
    RECT 220.165 12.975 220.445 14.505 ;
    RECT 216.845 12.975 217.125 14.505 ;
    RECT 128.335 6.62 128.545 14.505 ;
    RECT 138.48 7.095 138.58 7.225 ;
    RECT 139.7 1.015 139.97 14.505 ;
    RECT 64.535 12.975 64.815 14.505 ;
    RECT 61.215 12.975 61.495 14.505 ;
    RECT 57.895 12.975 58.175 14.505 ;
    RECT 54.575 12.975 54.855 14.505 ;
    RECT 51.255 12.975 51.535 14.505 ;
    RECT 47.935 12.975 48.215 14.505 ;
    RECT 44.615 12.975 44.895 14.505 ;
    RECT 41.295 12.975 41.575 14.505 ;
    RECT 37.975 12.975 38.255 14.505 ;
    RECT 34.655 12.975 34.935 14.505 ;
    RECT 31.335 12.975 31.615 14.505 ;
    RECT 28.015 12.975 28.295 14.505 ;
    RECT 24.695 12.975 24.975 14.505 ;
    RECT 21.375 12.975 21.655 14.505 ;
    RECT 18.055 12.975 18.335 14.505 ;
    RECT 14.735 12.975 15.015 14.505 ;
    RECT 11.415 12.975 11.695 14.505 ;
    RECT 8.095 12.975 8.375 14.505 ;
    RECT 4.775 12.975 5.055 14.505 ;
    RECT 1.455 12.975 1.735 14.505 ;
    RECT 117.655 12.975 117.935 14.505 ;
    RECT 114.335 12.975 114.615 14.505 ;
    RECT 111.015 12.975 111.295 14.505 ;
    RECT 107.695 12.975 107.975 14.505 ;
    RECT 104.375 12.975 104.655 14.505 ;
    RECT 101.055 12.975 101.335 14.505 ;
    RECT 97.735 12.975 98.015 14.505 ;
    RECT 94.415 12.975 94.695 14.505 ;
    RECT 91.095 12.975 91.375 14.505 ;
    RECT 87.775 12.975 88.055 14.505 ;
    RECT 84.455 12.975 84.735 14.505 ;
    RECT 81.135 12.975 81.415 14.505 ;
    RECT 77.815 12.975 78.095 14.505 ;
    RECT 74.495 12.975 74.775 14.505 ;
    RECT 71.175 12.975 71.455 14.505 ;
    RECT 67.855 12.975 68.135 14.505 ;
    RECT 117.655 12.695 117.935 12.975 ;
    RECT 117.8 4.14 117.87 7.295 ;
    RECT 1.455 12.695 1.735 12.975 ;
    RECT 1.6 4.14 1.67 7.295 ;
    RECT 31.335 12.695 31.615 12.975 ;
    RECT 31.48 4.14 31.55 7.295 ;
    RECT 28.015 12.695 28.295 12.975 ;
    RECT 28.16 4.14 28.23 7.295 ;
    RECT 24.695 12.695 24.975 12.975 ;
    RECT 24.84 4.14 24.91 7.295 ;
    RECT 21.375 12.695 21.655 12.975 ;
    RECT 21.52 4.14 21.59 7.295 ;
    RECT 18.055 12.695 18.335 12.975 ;
    RECT 18.2 4.14 18.27 7.295 ;
    RECT 14.735 12.695 15.015 12.975 ;
    RECT 14.88 4.14 14.95 7.295 ;
    RECT 11.415 12.695 11.695 12.975 ;
    RECT 11.56 4.14 11.63 7.295 ;
    RECT 8.095 12.695 8.375 12.975 ;
    RECT 8.24 4.14 8.31 7.295 ;
    RECT 4.775 12.695 5.055 12.975 ;
    RECT 4.92 4.14 4.99 7.295 ;
    RECT 114.335 12.695 114.615 12.975 ;
    RECT 114.48 4.14 114.55 7.295 ;
    RECT 111.015 12.695 111.295 12.975 ;
    RECT 111.16 4.14 111.23 7.295 ;
    RECT 107.695 12.695 107.975 12.975 ;
    RECT 107.84 4.14 107.91 7.295 ;
    RECT 104.375 12.695 104.655 12.975 ;
    RECT 104.52 4.14 104.59 7.295 ;
    RECT 101.055 12.695 101.335 12.975 ;
    RECT 101.2 4.14 101.27 7.295 ;
    RECT 97.735 12.695 98.015 12.975 ;
    RECT 97.88 4.14 97.95 7.295 ;
    RECT 94.415 12.695 94.695 12.975 ;
    RECT 94.56 4.14 94.63 7.295 ;
    RECT 91.095 12.695 91.375 12.975 ;
    RECT 91.24 4.14 91.31 7.295 ;
    RECT 87.775 12.695 88.055 12.975 ;
    RECT 87.92 4.14 87.99 7.295 ;
    RECT 84.455 12.695 84.735 12.975 ;
    RECT 84.6 4.14 84.67 7.295 ;
    RECT 81.135 12.695 81.415 12.975 ;
    RECT 81.28 4.14 81.35 7.295 ;
    RECT 77.815 12.695 78.095 12.975 ;
    RECT 77.96 4.14 78.03 7.295 ;
    RECT 74.495 12.695 74.775 12.975 ;
    RECT 74.64 4.14 74.71 7.295 ;
    RECT 71.175 12.695 71.455 12.975 ;
    RECT 71.32 4.14 71.39 7.295 ;
    RECT 67.855 12.695 68.135 12.975 ;
    RECT 68.0 4.14 68.07 7.295 ;
    RECT 64.535 12.695 64.815 12.975 ;
    RECT 64.68 4.14 64.75 7.295 ;
    RECT 61.215 12.695 61.495 12.975 ;
    RECT 61.36 4.14 61.43 7.295 ;
    RECT 57.895 12.695 58.175 12.975 ;
    RECT 58.04 4.14 58.11 7.295 ;
    RECT 54.575 12.695 54.855 12.975 ;
    RECT 54.72 4.14 54.79 7.295 ;
    RECT 51.255 12.695 51.535 12.975 ;
    RECT 51.4 4.14 51.47 7.295 ;
    RECT 47.935 12.695 48.215 12.975 ;
    RECT 48.08 4.14 48.15 7.295 ;
    RECT 44.615 12.695 44.895 12.975 ;
    RECT 44.76 4.14 44.83 7.295 ;
    RECT 41.295 12.695 41.575 12.975 ;
    RECT 41.44 4.14 41.51 7.295 ;
    RECT 37.975 12.695 38.255 12.975 ;
    RECT 38.12 4.14 38.19 7.295 ;
    RECT 34.655 12.695 34.935 12.975 ;
    RECT 34.8 4.14 34.87 7.295 ;
    RECT 57.895 100.295 58.175 100.81 ;
    RECT 54.575 100.295 54.855 100.81 ;
    RECT 51.255 100.295 51.535 100.81 ;
    RECT 47.935 100.295 48.215 100.81 ;
    RECT 44.615 100.295 44.895 100.81 ;
    RECT 41.295 100.295 41.575 100.81 ;
    RECT 37.975 100.295 38.255 100.81 ;
    RECT 34.655 100.295 34.935 100.81 ;
    RECT 266.645 100.295 266.925 100.81 ;
    RECT 263.325 100.295 263.605 100.81 ;
    RECT 260.005 100.295 260.285 100.81 ;
    RECT 256.685 100.295 256.965 100.81 ;
    RECT 253.365 100.295 253.645 100.81 ;
    RECT 121.67 100.295 121.86 100.615 ;
    RECT 139.7 100.295 139.97 100.81 ;
    RECT 250.045 100.295 250.325 100.81 ;
    RECT 180.325 100.295 180.605 100.81 ;
    RECT 177.005 100.295 177.285 100.81 ;
    RECT 246.725 100.295 247.005 100.81 ;
    RECT 173.685 100.295 173.965 100.81 ;
    RECT 243.405 100.295 243.685 100.81 ;
    RECT 170.365 100.295 170.645 100.81 ;
    RECT 240.085 100.295 240.365 100.81 ;
    RECT 167.045 100.295 167.325 100.81 ;
    RECT 236.765 100.295 237.045 100.81 ;
    RECT 163.725 100.295 164.005 100.81 ;
    RECT 233.445 100.295 233.725 100.81 ;
    RECT 160.405 100.295 160.685 100.81 ;
    RECT 230.125 100.295 230.405 100.81 ;
    RECT 157.085 100.295 157.365 100.81 ;
    RECT 226.805 100.295 227.085 100.81 ;
    RECT 153.765 100.295 154.045 100.81 ;
    RECT 223.485 100.295 223.765 100.81 ;
    RECT 150.445 100.295 150.725 100.81 ;
    RECT 220.165 100.295 220.445 100.81 ;
    RECT 216.845 100.295 217.125 100.81 ;
    RECT 213.525 100.295 213.805 100.81 ;
    RECT 210.205 100.295 210.485 100.81 ;
    RECT 206.885 100.295 207.165 100.81 ;
    RECT 203.565 100.295 203.845 100.81 ;
    RECT 200.245 100.295 200.525 100.81 ;
    RECT 196.925 100.295 197.205 100.81 ;
    RECT 193.605 100.295 193.885 100.81 ;
    RECT 190.285 100.295 190.565 100.81 ;
    RECT 186.965 100.295 187.245 100.81 ;
    RECT 31.335 100.295 31.615 100.81 ;
    RECT 183.645 100.295 183.925 100.81 ;
    RECT 28.015 100.295 28.295 100.81 ;
    RECT 24.695 100.295 24.975 100.81 ;
    RECT 21.375 100.295 21.655 100.81 ;
    RECT 18.055 100.295 18.335 100.81 ;
    RECT 14.735 100.295 15.015 100.81 ;
    RECT 11.415 100.295 11.695 100.81 ;
    RECT 8.095 100.295 8.375 100.81 ;
    RECT 4.775 100.295 5.055 100.81 ;
    RECT 1.455 100.295 1.735 100.81 ;
    RECT 117.655 100.295 117.935 100.81 ;
    RECT 114.335 100.295 114.615 100.81 ;
    RECT 111.015 100.295 111.295 100.81 ;
    RECT 107.695 100.295 107.975 100.81 ;
    RECT 104.375 100.295 104.655 100.81 ;
    RECT 101.055 100.295 101.335 100.81 ;
    RECT 97.735 100.295 98.015 100.81 ;
    RECT 94.415 100.295 94.695 100.81 ;
    RECT 91.095 100.295 91.375 100.81 ;
    RECT 87.775 100.295 88.055 100.81 ;
    RECT 84.455 100.295 84.735 100.81 ;
    RECT 81.135 100.295 81.415 100.81 ;
    RECT 77.815 100.295 78.095 100.81 ;
    RECT 74.495 100.295 74.775 100.81 ;
    RECT 71.175 100.295 71.455 100.81 ;
    RECT 67.855 100.295 68.135 100.81 ;
    RECT 64.535 100.295 64.815 100.81 ;
    RECT 61.215 100.295 61.495 100.81 ;
    END
  END sram464x144

END LIBRARY

