# Confidential Information of ARM, Inc.
# Use subject to ARM license.
# Copyright (c) 2022 ARM, Inc.

# ACI Version r1p1

# Reifier 4.0.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;

#name: High Density Single Port Register File RVT RVT Compiler | LOGIC0040LL 40nm Process 0.299um^2 Bit Cell
#version: r1p1
#comment: This is a memory instance
#configuration:  -activity_factor 50 -back_biasing off -bits 104 -bmux off -bus_notation on -check_instname on -diodes on -drive 6 -ema on -frequency 200 -instname sram520x104 -left_bus_delim "[" -mux 4 -mvt "" -name_case upper -power_type otc -prefix "" -pwr_gnd_rename vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -retention on -right_bus_delim "]" -ser none -site_def off -top_layer m5-m10 -words 520 -write_mask off -write_thru off -corners ss_0p99v_0p99v_125c,tt_1p10v_1p10v_125c
MACRO sram520x104
  FOREIGN sram520x104 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 374.62 BY 61.255 ;
  CLASS BLOCK ;
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 187.255 0.0 187.395 0.25 ;
      LAYER M2 ;
      RECT 187.255 0.0 187.395 0.25 ;
      LAYER M1 ;
      RECT 187.255 0.0 187.395 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[6]
  PIN EMA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 189.61 0.0 189.75 0.25 ;
      LAYER M2 ;
      RECT 189.61 0.0 189.75 0.25 ;
      LAYER M3 ;
      RECT 189.61 0.0 189.75 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMA[0]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 185.65 0.0 185.79 0.25 ;
      LAYER M2 ;
      RECT 185.65 0.0 185.79 0.25 ;
      LAYER M1 ;
      RECT 185.65 0.0 185.79 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END WEN
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 190.41 0.0 190.55 0.25 ;
      LAYER M2 ;
      RECT 190.41 0.0 190.55 0.25 ;
      LAYER M3 ;
      RECT 190.41 0.0 190.55 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[9]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 185.23 0.0 185.37 0.25 ;
      LAYER M2 ;
      RECT 185.23 0.0 185.37 0.25 ;
      LAYER M1 ;
      RECT 185.23 0.0 185.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[5]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 190.69 0.0 190.83 0.25 ;
      LAYER M2 ;
      RECT 190.69 0.0 190.83 0.25 ;
      LAYER M3 ;
      RECT 190.69 0.0 190.83 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[8]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.83 0.0 181.97 0.25 ;
      LAYER M2 ;
      RECT 181.83 0.0 181.97 0.25 ;
      LAYER M1 ;
      RECT 181.83 0.0 181.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[2]
  PIN EMA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 191.26 0.0 191.4 0.25 ;
      LAYER M2 ;
      RECT 191.26 0.0 191.4 0.25 ;
      LAYER M3 ;
      RECT 191.26 0.0 191.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMA[1]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.55 0.0 181.69 0.25 ;
      LAYER M2 ;
      RECT 181.55 0.0 181.69 0.25 ;
      LAYER M1 ;
      RECT 181.55 0.0 181.69 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[3]
  PIN EMA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 191.655 0.0 191.795 0.25 ;
      LAYER M2 ;
      RECT 191.655 0.0 191.795 0.25 ;
      LAYER M3 ;
      RECT 191.655 0.0 191.795 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMA[2]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 179.54 0.0 179.68 0.25 ;
      LAYER M2 ;
      RECT 179.54 0.0 179.68 0.25 ;
      LAYER M1 ;
      RECT 179.54 0.0 179.68 0.25 ;
      LAYER M4 ;
      RECT 179.5 0.0 179.71 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CLK
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 193.805 0.0 193.945 0.25 ;
      LAYER M2 ;
      RECT 193.805 0.0 193.945 0.25 ;
      LAYER M3 ;
      RECT 193.805 0.0 193.945 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[4]
  PIN EMAW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 178.565 0.0 178.705 0.25 ;
      LAYER M2 ;
      RECT 178.565 0.0 178.705 0.25 ;
      LAYER M1 ;
      RECT 178.565 0.0 178.705 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAW[1]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 194.09 0.0 194.23 0.25 ;
      LAYER M2 ;
      RECT 194.09 0.0 194.23 0.25 ;
      LAYER M3 ;
      RECT 194.09 0.0 194.23 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[7]
  PIN EMAW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 177.75 0.0 177.89 0.25 ;
      LAYER M2 ;
      RECT 177.75 0.0 177.89 0.25 ;
      LAYER M1 ;
      RECT 177.75 0.0 177.89 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAW[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 197.485 0.0 197.625 0.25 ;
      LAYER M2 ;
      RECT 197.485 0.0 197.625 0.25 ;
      LAYER M3 ;
      RECT 197.485 0.0 197.625 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[1]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.475 0.0 174.615 0.25 ;
      LAYER M2 ;
      RECT 174.475 0.0 174.615 0.25 ;
      LAYER M1 ;
      RECT 174.475 0.0 174.615 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CEN
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 200.64 0.0 200.78 0.25 ;
      LAYER M2 ;
      RECT 200.64 0.0 200.78 0.25 ;
      LAYER M3 ;
      RECT 200.64 0.0 200.78 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END A[0]
  PIN RET1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 173.83 0.0 173.97 0.25 ;
      LAYER M2 ;
      RECT 173.83 0.0 173.97 0.25 ;
      LAYER M1 ;
      RECT 173.83 0.0 173.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END RET1N
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 201.695 0.0 201.835 0.25 ;
      LAYER M2 ;
      RECT 201.695 0.0 201.835 0.25 ;
      LAYER M3 ;
      RECT 201.695 0.0 201.835 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 172.785 0.0 172.925 0.25 ;
      LAYER M2 ;
      RECT 172.785 0.0 172.925 0.25 ;
      LAYER M1 ;
      RECT 172.785 0.0 172.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[51]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 203.325 0.0 203.465 0.25 ;
      LAYER M2 ;
      RECT 203.325 0.0 203.465 0.25 ;
      LAYER M3 ;
      RECT 203.325 0.0 203.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 171.155 0.0 171.295 0.25 ;
      LAYER M2 ;
      RECT 171.155 0.0 171.295 0.25 ;
      LAYER M1 ;
      RECT 171.155 0.0 171.295 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[51]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 205.015 0.0 205.155 0.25 ;
      LAYER M2 ;
      RECT 205.015 0.0 205.155 0.25 ;
      LAYER M3 ;
      RECT 205.015 0.0 205.155 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[53]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 169.465 0.0 169.605 0.25 ;
      LAYER M2 ;
      RECT 169.465 0.0 169.605 0.25 ;
      LAYER M1 ;
      RECT 169.465 0.0 169.605 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[50]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 206.645 0.0 206.785 0.25 ;
      LAYER M2 ;
      RECT 206.645 0.0 206.785 0.25 ;
      LAYER M3 ;
      RECT 206.645 0.0 206.785 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[53]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 167.835 0.0 167.975 0.25 ;
      LAYER M2 ;
      RECT 167.835 0.0 167.975 0.25 ;
      LAYER M1 ;
      RECT 167.835 0.0 167.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[50]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 208.335 0.0 208.475 0.25 ;
      LAYER M2 ;
      RECT 208.335 0.0 208.475 0.25 ;
      LAYER M3 ;
      RECT 208.335 0.0 208.475 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[54]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 166.145 0.0 166.285 0.25 ;
      LAYER M2 ;
      RECT 166.145 0.0 166.285 0.25 ;
      LAYER M1 ;
      RECT 166.145 0.0 166.285 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[49]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 209.965 0.0 210.105 0.25 ;
      LAYER M2 ;
      RECT 209.965 0.0 210.105 0.25 ;
      LAYER M3 ;
      RECT 209.965 0.0 210.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[54]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 164.515 0.0 164.655 0.25 ;
      LAYER M2 ;
      RECT 164.515 0.0 164.655 0.25 ;
      LAYER M1 ;
      RECT 164.515 0.0 164.655 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[49]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 211.655 0.0 211.795 0.25 ;
      LAYER M2 ;
      RECT 211.655 0.0 211.795 0.25 ;
      LAYER M3 ;
      RECT 211.655 0.0 211.795 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[55]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 162.825 0.0 162.965 0.25 ;
      LAYER M2 ;
      RECT 162.825 0.0 162.965 0.25 ;
      LAYER M1 ;
      RECT 162.825 0.0 162.965 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[48]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 213.285 0.0 213.425 0.25 ;
      LAYER M2 ;
      RECT 213.285 0.0 213.425 0.25 ;
      LAYER M3 ;
      RECT 213.285 0.0 213.425 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[55]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 161.195 0.0 161.335 0.25 ;
      LAYER M2 ;
      RECT 161.195 0.0 161.335 0.25 ;
      LAYER M1 ;
      RECT 161.195 0.0 161.335 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[48]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 214.975 0.0 215.115 0.25 ;
      LAYER M2 ;
      RECT 214.975 0.0 215.115 0.25 ;
      LAYER M3 ;
      RECT 214.975 0.0 215.115 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[56]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 159.505 0.0 159.645 0.25 ;
      LAYER M2 ;
      RECT 159.505 0.0 159.645 0.25 ;
      LAYER M1 ;
      RECT 159.505 0.0 159.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[47]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 216.605 0.0 216.745 0.25 ;
      LAYER M2 ;
      RECT 216.605 0.0 216.745 0.25 ;
      LAYER M3 ;
      RECT 216.605 0.0 216.745 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[56]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 157.875 0.0 158.015 0.25 ;
      LAYER M2 ;
      RECT 157.875 0.0 158.015 0.25 ;
      LAYER M1 ;
      RECT 157.875 0.0 158.015 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[47]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 218.295 0.0 218.435 0.25 ;
      LAYER M2 ;
      RECT 218.295 0.0 218.435 0.25 ;
      LAYER M3 ;
      RECT 218.295 0.0 218.435 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[57]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 156.185 0.0 156.325 0.25 ;
      LAYER M2 ;
      RECT 156.185 0.0 156.325 0.25 ;
      LAYER M1 ;
      RECT 156.185 0.0 156.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[46]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 219.925 0.0 220.065 0.25 ;
      LAYER M2 ;
      RECT 219.925 0.0 220.065 0.25 ;
      LAYER M3 ;
      RECT 219.925 0.0 220.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[57]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 154.555 0.0 154.695 0.25 ;
      LAYER M2 ;
      RECT 154.555 0.0 154.695 0.25 ;
      LAYER M1 ;
      RECT 154.555 0.0 154.695 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[46]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 221.615 0.0 221.755 0.25 ;
      LAYER M2 ;
      RECT 221.615 0.0 221.755 0.25 ;
      LAYER M3 ;
      RECT 221.615 0.0 221.755 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[58]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 152.865 0.0 153.005 0.25 ;
      LAYER M2 ;
      RECT 152.865 0.0 153.005 0.25 ;
      LAYER M1 ;
      RECT 152.865 0.0 153.005 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[45]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 223.245 0.0 223.385 0.25 ;
      LAYER M2 ;
      RECT 223.245 0.0 223.385 0.25 ;
      LAYER M3 ;
      RECT 223.245 0.0 223.385 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[58]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 151.235 0.0 151.375 0.25 ;
      LAYER M2 ;
      RECT 151.235 0.0 151.375 0.25 ;
      LAYER M1 ;
      RECT 151.235 0.0 151.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[45]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 224.935 0.0 225.075 0.25 ;
      LAYER M2 ;
      RECT 224.935 0.0 225.075 0.25 ;
      LAYER M3 ;
      RECT 224.935 0.0 225.075 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[59]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 149.545 0.0 149.685 0.25 ;
      LAYER M2 ;
      RECT 149.545 0.0 149.685 0.25 ;
      LAYER M1 ;
      RECT 149.545 0.0 149.685 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[44]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 226.565 0.0 226.705 0.25 ;
      LAYER M2 ;
      RECT 226.565 0.0 226.705 0.25 ;
      LAYER M3 ;
      RECT 226.565 0.0 226.705 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[59]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 147.915 0.0 148.055 0.25 ;
      LAYER M2 ;
      RECT 147.915 0.0 148.055 0.25 ;
      LAYER M1 ;
      RECT 147.915 0.0 148.055 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[44]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 228.255 0.0 228.395 0.25 ;
      LAYER M2 ;
      RECT 228.255 0.0 228.395 0.25 ;
      LAYER M3 ;
      RECT 228.255 0.0 228.395 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[60]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 146.225 0.0 146.365 0.25 ;
      LAYER M2 ;
      RECT 146.225 0.0 146.365 0.25 ;
      LAYER M1 ;
      RECT 146.225 0.0 146.365 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[43]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 229.885 0.0 230.025 0.25 ;
      LAYER M2 ;
      RECT 229.885 0.0 230.025 0.25 ;
      LAYER M3 ;
      RECT 229.885 0.0 230.025 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[60]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 144.595 0.0 144.735 0.25 ;
      LAYER M2 ;
      RECT 144.595 0.0 144.735 0.25 ;
      LAYER M1 ;
      RECT 144.595 0.0 144.735 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[43]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 231.575 0.0 231.715 0.25 ;
      LAYER M2 ;
      RECT 231.575 0.0 231.715 0.25 ;
      LAYER M3 ;
      RECT 231.575 0.0 231.715 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[61]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 142.905 0.0 143.045 0.25 ;
      LAYER M2 ;
      RECT 142.905 0.0 143.045 0.25 ;
      LAYER M1 ;
      RECT 142.905 0.0 143.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[42]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 233.205 0.0 233.345 0.25 ;
      LAYER M2 ;
      RECT 233.205 0.0 233.345 0.25 ;
      LAYER M3 ;
      RECT 233.205 0.0 233.345 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[61]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 141.275 0.0 141.415 0.25 ;
      LAYER M2 ;
      RECT 141.275 0.0 141.415 0.25 ;
      LAYER M1 ;
      RECT 141.275 0.0 141.415 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[42]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 234.895 0.0 235.035 0.25 ;
      LAYER M2 ;
      RECT 234.895 0.0 235.035 0.25 ;
      LAYER M3 ;
      RECT 234.895 0.0 235.035 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[62]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 139.585 0.0 139.725 0.25 ;
      LAYER M2 ;
      RECT 139.585 0.0 139.725 0.25 ;
      LAYER M1 ;
      RECT 139.585 0.0 139.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[41]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 236.525 0.0 236.665 0.25 ;
      LAYER M2 ;
      RECT 236.525 0.0 236.665 0.25 ;
      LAYER M3 ;
      RECT 236.525 0.0 236.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[62]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 137.955 0.0 138.095 0.25 ;
      LAYER M2 ;
      RECT 137.955 0.0 138.095 0.25 ;
      LAYER M1 ;
      RECT 137.955 0.0 138.095 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[41]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 238.215 0.0 238.355 0.25 ;
      LAYER M2 ;
      RECT 238.215 0.0 238.355 0.25 ;
      LAYER M3 ;
      RECT 238.215 0.0 238.355 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[63]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 136.265 0.0 136.405 0.25 ;
      LAYER M2 ;
      RECT 136.265 0.0 136.405 0.25 ;
      LAYER M1 ;
      RECT 136.265 0.0 136.405 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[40]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 239.845 0.0 239.985 0.25 ;
      LAYER M2 ;
      RECT 239.845 0.0 239.985 0.25 ;
      LAYER M3 ;
      RECT 239.845 0.0 239.985 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[63]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 134.635 0.0 134.775 0.25 ;
      LAYER M2 ;
      RECT 134.635 0.0 134.775 0.25 ;
      LAYER M1 ;
      RECT 134.635 0.0 134.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[40]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 241.535 0.0 241.675 0.25 ;
      LAYER M2 ;
      RECT 241.535 0.0 241.675 0.25 ;
      LAYER M3 ;
      RECT 241.535 0.0 241.675 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[64]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.945 0.0 133.085 0.25 ;
      LAYER M2 ;
      RECT 132.945 0.0 133.085 0.25 ;
      LAYER M1 ;
      RECT 132.945 0.0 133.085 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[39]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 243.165 0.0 243.305 0.25 ;
      LAYER M2 ;
      RECT 243.165 0.0 243.305 0.25 ;
      LAYER M3 ;
      RECT 243.165 0.0 243.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[64]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.315 0.0 131.455 0.25 ;
      LAYER M2 ;
      RECT 131.315 0.0 131.455 0.25 ;
      LAYER M1 ;
      RECT 131.315 0.0 131.455 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[39]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 244.855 0.0 244.995 0.25 ;
      LAYER M2 ;
      RECT 244.855 0.0 244.995 0.25 ;
      LAYER M3 ;
      RECT 244.855 0.0 244.995 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[65]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 129.625 0.0 129.765 0.25 ;
      LAYER M2 ;
      RECT 129.625 0.0 129.765 0.25 ;
      LAYER M1 ;
      RECT 129.625 0.0 129.765 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[38]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 246.485 0.0 246.625 0.25 ;
      LAYER M2 ;
      RECT 246.485 0.0 246.625 0.25 ;
      LAYER M3 ;
      RECT 246.485 0.0 246.625 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[65]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 127.995 0.0 128.135 0.25 ;
      LAYER M2 ;
      RECT 127.995 0.0 128.135 0.25 ;
      LAYER M1 ;
      RECT 127.995 0.0 128.135 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[38]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 248.175 0.0 248.315 0.25 ;
      LAYER M2 ;
      RECT 248.175 0.0 248.315 0.25 ;
      LAYER M3 ;
      RECT 248.175 0.0 248.315 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[66]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 126.305 0.0 126.445 0.25 ;
      LAYER M2 ;
      RECT 126.305 0.0 126.445 0.25 ;
      LAYER M1 ;
      RECT 126.305 0.0 126.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[37]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 249.805 0.0 249.945 0.25 ;
      LAYER M2 ;
      RECT 249.805 0.0 249.945 0.25 ;
      LAYER M3 ;
      RECT 249.805 0.0 249.945 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[66]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.675 0.0 124.815 0.25 ;
      LAYER M2 ;
      RECT 124.675 0.0 124.815 0.25 ;
      LAYER M1 ;
      RECT 124.675 0.0 124.815 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[37]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 251.495 0.0 251.635 0.25 ;
      LAYER M2 ;
      RECT 251.495 0.0 251.635 0.25 ;
      LAYER M3 ;
      RECT 251.495 0.0 251.635 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[67]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 122.985 0.0 123.125 0.25 ;
      LAYER M2 ;
      RECT 122.985 0.0 123.125 0.25 ;
      LAYER M1 ;
      RECT 122.985 0.0 123.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[36]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 253.125 0.0 253.265 0.25 ;
      LAYER M2 ;
      RECT 253.125 0.0 253.265 0.25 ;
      LAYER M3 ;
      RECT 253.125 0.0 253.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[67]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 121.355 0.0 121.495 0.25 ;
      LAYER M2 ;
      RECT 121.355 0.0 121.495 0.25 ;
      LAYER M1 ;
      RECT 121.355 0.0 121.495 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[36]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 254.815 0.0 254.955 0.25 ;
      LAYER M2 ;
      RECT 254.815 0.0 254.955 0.25 ;
      LAYER M3 ;
      RECT 254.815 0.0 254.955 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[68]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.665 0.0 119.805 0.25 ;
      LAYER M2 ;
      RECT 119.665 0.0 119.805 0.25 ;
      LAYER M1 ;
      RECT 119.665 0.0 119.805 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[35]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 256.445 0.0 256.585 0.25 ;
      LAYER M2 ;
      RECT 256.445 0.0 256.585 0.25 ;
      LAYER M3 ;
      RECT 256.445 0.0 256.585 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[68]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.035 0.0 118.175 0.25 ;
      LAYER M2 ;
      RECT 118.035 0.0 118.175 0.25 ;
      LAYER M1 ;
      RECT 118.035 0.0 118.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[35]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 258.135 0.0 258.275 0.25 ;
      LAYER M2 ;
      RECT 258.135 0.0 258.275 0.25 ;
      LAYER M3 ;
      RECT 258.135 0.0 258.275 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[69]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 116.345 0.0 116.485 0.25 ;
      LAYER M2 ;
      RECT 116.345 0.0 116.485 0.25 ;
      LAYER M1 ;
      RECT 116.345 0.0 116.485 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[34]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 259.765 0.0 259.905 0.25 ;
      LAYER M2 ;
      RECT 259.765 0.0 259.905 0.25 ;
      LAYER M3 ;
      RECT 259.765 0.0 259.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[69]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 114.715 0.0 114.855 0.25 ;
      LAYER M2 ;
      RECT 114.715 0.0 114.855 0.25 ;
      LAYER M1 ;
      RECT 114.715 0.0 114.855 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[34]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 261.455 0.0 261.595 0.25 ;
      LAYER M2 ;
      RECT 261.455 0.0 261.595 0.25 ;
      LAYER M3 ;
      RECT 261.455 0.0 261.595 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[70]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 113.025 0.0 113.165 0.25 ;
      LAYER M2 ;
      RECT 113.025 0.0 113.165 0.25 ;
      LAYER M1 ;
      RECT 113.025 0.0 113.165 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[33]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 263.085 0.0 263.225 0.25 ;
      LAYER M2 ;
      RECT 263.085 0.0 263.225 0.25 ;
      LAYER M3 ;
      RECT 263.085 0.0 263.225 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[70]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 111.395 0.0 111.535 0.25 ;
      LAYER M2 ;
      RECT 111.395 0.0 111.535 0.25 ;
      LAYER M1 ;
      RECT 111.395 0.0 111.535 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[33]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 264.775 0.0 264.915 0.25 ;
      LAYER M2 ;
      RECT 264.775 0.0 264.915 0.25 ;
      LAYER M3 ;
      RECT 264.775 0.0 264.915 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[71]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 109.705 0.0 109.845 0.25 ;
      LAYER M2 ;
      RECT 109.705 0.0 109.845 0.25 ;
      LAYER M1 ;
      RECT 109.705 0.0 109.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[32]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 266.405 0.0 266.545 0.25 ;
      LAYER M2 ;
      RECT 266.405 0.0 266.545 0.25 ;
      LAYER M3 ;
      RECT 266.405 0.0 266.545 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[71]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 108.075 0.0 108.215 0.25 ;
      LAYER M2 ;
      RECT 108.075 0.0 108.215 0.25 ;
      LAYER M1 ;
      RECT 108.075 0.0 108.215 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[32]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 268.095 0.0 268.235 0.25 ;
      LAYER M2 ;
      RECT 268.095 0.0 268.235 0.25 ;
      LAYER M3 ;
      RECT 268.095 0.0 268.235 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[72]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.385 0.0 106.525 0.25 ;
      LAYER M2 ;
      RECT 106.385 0.0 106.525 0.25 ;
      LAYER M1 ;
      RECT 106.385 0.0 106.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[31]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 269.725 0.0 269.865 0.25 ;
      LAYER M2 ;
      RECT 269.725 0.0 269.865 0.25 ;
      LAYER M3 ;
      RECT 269.725 0.0 269.865 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[72]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 104.755 0.0 104.895 0.25 ;
      LAYER M2 ;
      RECT 104.755 0.0 104.895 0.25 ;
      LAYER M1 ;
      RECT 104.755 0.0 104.895 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[31]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 271.415 0.0 271.555 0.25 ;
      LAYER M2 ;
      RECT 271.415 0.0 271.555 0.25 ;
      LAYER M3 ;
      RECT 271.415 0.0 271.555 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[73]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 103.065 0.0 103.205 0.25 ;
      LAYER M2 ;
      RECT 103.065 0.0 103.205 0.25 ;
      LAYER M1 ;
      RECT 103.065 0.0 103.205 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[30]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 273.045 0.0 273.185 0.25 ;
      LAYER M2 ;
      RECT 273.045 0.0 273.185 0.25 ;
      LAYER M3 ;
      RECT 273.045 0.0 273.185 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[73]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 101.435 0.0 101.575 0.25 ;
      LAYER M2 ;
      RECT 101.435 0.0 101.575 0.25 ;
      LAYER M1 ;
      RECT 101.435 0.0 101.575 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[30]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 274.735 0.0 274.875 0.25 ;
      LAYER M2 ;
      RECT 274.735 0.0 274.875 0.25 ;
      LAYER M3 ;
      RECT 274.735 0.0 274.875 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[74]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 99.745 0.0 99.885 0.25 ;
      LAYER M2 ;
      RECT 99.745 0.0 99.885 0.25 ;
      LAYER M1 ;
      RECT 99.745 0.0 99.885 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[29]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 276.365 0.0 276.505 0.25 ;
      LAYER M2 ;
      RECT 276.365 0.0 276.505 0.25 ;
      LAYER M3 ;
      RECT 276.365 0.0 276.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[74]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.115 0.0 98.255 0.25 ;
      LAYER M2 ;
      RECT 98.115 0.0 98.255 0.25 ;
      LAYER M1 ;
      RECT 98.115 0.0 98.255 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[29]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 278.055 0.0 278.195 0.25 ;
      LAYER M2 ;
      RECT 278.055 0.0 278.195 0.25 ;
      LAYER M3 ;
      RECT 278.055 0.0 278.195 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[75]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 96.425 0.0 96.565 0.25 ;
      LAYER M2 ;
      RECT 96.425 0.0 96.565 0.25 ;
      LAYER M1 ;
      RECT 96.425 0.0 96.565 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[28]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 279.685 0.0 279.825 0.25 ;
      LAYER M2 ;
      RECT 279.685 0.0 279.825 0.25 ;
      LAYER M3 ;
      RECT 279.685 0.0 279.825 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[75]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 94.795 0.0 94.935 0.25 ;
      LAYER M2 ;
      RECT 94.795 0.0 94.935 0.25 ;
      LAYER M1 ;
      RECT 94.795 0.0 94.935 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[28]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 281.375 0.0 281.515 0.25 ;
      LAYER M2 ;
      RECT 281.375 0.0 281.515 0.25 ;
      LAYER M3 ;
      RECT 281.375 0.0 281.515 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[76]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.105 0.0 93.245 0.25 ;
      LAYER M2 ;
      RECT 93.105 0.0 93.245 0.25 ;
      LAYER M1 ;
      RECT 93.105 0.0 93.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[27]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 283.005 0.0 283.145 0.25 ;
      LAYER M2 ;
      RECT 283.005 0.0 283.145 0.25 ;
      LAYER M3 ;
      RECT 283.005 0.0 283.145 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[76]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 91.475 0.0 91.615 0.25 ;
      LAYER M2 ;
      RECT 91.475 0.0 91.615 0.25 ;
      LAYER M1 ;
      RECT 91.475 0.0 91.615 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[27]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 284.695 0.0 284.835 0.25 ;
      LAYER M2 ;
      RECT 284.695 0.0 284.835 0.25 ;
      LAYER M3 ;
      RECT 284.695 0.0 284.835 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[77]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 89.785 0.0 89.925 0.25 ;
      LAYER M2 ;
      RECT 89.785 0.0 89.925 0.25 ;
      LAYER M1 ;
      RECT 89.785 0.0 89.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[26]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 286.325 0.0 286.465 0.25 ;
      LAYER M2 ;
      RECT 286.325 0.0 286.465 0.25 ;
      LAYER M3 ;
      RECT 286.325 0.0 286.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[77]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.155 0.0 88.295 0.25 ;
      LAYER M2 ;
      RECT 88.155 0.0 88.295 0.25 ;
      LAYER M1 ;
      RECT 88.155 0.0 88.295 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[26]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 288.015 0.0 288.155 0.25 ;
      LAYER M2 ;
      RECT 288.015 0.0 288.155 0.25 ;
      LAYER M3 ;
      RECT 288.015 0.0 288.155 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[78]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 86.465 0.0 86.605 0.25 ;
      LAYER M2 ;
      RECT 86.465 0.0 86.605 0.25 ;
      LAYER M1 ;
      RECT 86.465 0.0 86.605 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[25]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 289.645 0.0 289.785 0.25 ;
      LAYER M2 ;
      RECT 289.645 0.0 289.785 0.25 ;
      LAYER M3 ;
      RECT 289.645 0.0 289.785 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[78]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 84.835 0.0 84.975 0.25 ;
      LAYER M2 ;
      RECT 84.835 0.0 84.975 0.25 ;
      LAYER M1 ;
      RECT 84.835 0.0 84.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[25]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 291.335 0.0 291.475 0.25 ;
      LAYER M2 ;
      RECT 291.335 0.0 291.475 0.25 ;
      LAYER M3 ;
      RECT 291.335 0.0 291.475 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[79]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 83.145 0.0 83.285 0.25 ;
      LAYER M2 ;
      RECT 83.145 0.0 83.285 0.25 ;
      LAYER M1 ;
      RECT 83.145 0.0 83.285 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[24]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 292.965 0.0 293.105 0.25 ;
      LAYER M2 ;
      RECT 292.965 0.0 293.105 0.25 ;
      LAYER M3 ;
      RECT 292.965 0.0 293.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[79]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.515 0.0 81.655 0.25 ;
      LAYER M2 ;
      RECT 81.515 0.0 81.655 0.25 ;
      LAYER M1 ;
      RECT 81.515 0.0 81.655 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[24]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 294.655 0.0 294.795 0.25 ;
      LAYER M2 ;
      RECT 294.655 0.0 294.795 0.25 ;
      LAYER M3 ;
      RECT 294.655 0.0 294.795 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[80]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 79.825 0.0 79.965 0.25 ;
      LAYER M2 ;
      RECT 79.825 0.0 79.965 0.25 ;
      LAYER M1 ;
      RECT 79.825 0.0 79.965 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[23]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 296.285 0.0 296.425 0.25 ;
      LAYER M2 ;
      RECT 296.285 0.0 296.425 0.25 ;
      LAYER M3 ;
      RECT 296.285 0.0 296.425 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[80]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 78.195 0.0 78.335 0.25 ;
      LAYER M2 ;
      RECT 78.195 0.0 78.335 0.25 ;
      LAYER M1 ;
      RECT 78.195 0.0 78.335 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[23]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 297.975 0.0 298.115 0.25 ;
      LAYER M2 ;
      RECT 297.975 0.0 298.115 0.25 ;
      LAYER M3 ;
      RECT 297.975 0.0 298.115 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[81]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.505 0.0 76.645 0.25 ;
      LAYER M2 ;
      RECT 76.505 0.0 76.645 0.25 ;
      LAYER M1 ;
      RECT 76.505 0.0 76.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[22]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 299.605 0.0 299.745 0.25 ;
      LAYER M2 ;
      RECT 299.605 0.0 299.745 0.25 ;
      LAYER M3 ;
      RECT 299.605 0.0 299.745 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[81]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 74.875 0.0 75.015 0.25 ;
      LAYER M2 ;
      RECT 74.875 0.0 75.015 0.25 ;
      LAYER M1 ;
      RECT 74.875 0.0 75.015 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[22]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 301.295 0.0 301.435 0.25 ;
      LAYER M2 ;
      RECT 301.295 0.0 301.435 0.25 ;
      LAYER M3 ;
      RECT 301.295 0.0 301.435 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[82]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 73.185 0.0 73.325 0.25 ;
      LAYER M2 ;
      RECT 73.185 0.0 73.325 0.25 ;
      LAYER M1 ;
      RECT 73.185 0.0 73.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[21]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 302.925 0.0 303.065 0.25 ;
      LAYER M2 ;
      RECT 302.925 0.0 303.065 0.25 ;
      LAYER M3 ;
      RECT 302.925 0.0 303.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[82]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 71.555 0.0 71.695 0.25 ;
      LAYER M2 ;
      RECT 71.555 0.0 71.695 0.25 ;
      LAYER M1 ;
      RECT 71.555 0.0 71.695 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[21]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 304.615 0.0 304.755 0.25 ;
      LAYER M2 ;
      RECT 304.615 0.0 304.755 0.25 ;
      LAYER M3 ;
      RECT 304.615 0.0 304.755 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[83]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.865 0.0 70.005 0.25 ;
      LAYER M2 ;
      RECT 69.865 0.0 70.005 0.25 ;
      LAYER M1 ;
      RECT 69.865 0.0 70.005 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[20]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 306.245 0.0 306.385 0.25 ;
      LAYER M2 ;
      RECT 306.245 0.0 306.385 0.25 ;
      LAYER M3 ;
      RECT 306.245 0.0 306.385 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[83]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 68.235 0.0 68.375 0.25 ;
      LAYER M2 ;
      RECT 68.235 0.0 68.375 0.25 ;
      LAYER M1 ;
      RECT 68.235 0.0 68.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[20]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 307.935 0.0 308.075 0.25 ;
      LAYER M2 ;
      RECT 307.935 0.0 308.075 0.25 ;
      LAYER M3 ;
      RECT 307.935 0.0 308.075 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[84]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 66.545 0.0 66.685 0.25 ;
      LAYER M2 ;
      RECT 66.545 0.0 66.685 0.25 ;
      LAYER M1 ;
      RECT 66.545 0.0 66.685 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[19]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 309.565 0.0 309.705 0.25 ;
      LAYER M2 ;
      RECT 309.565 0.0 309.705 0.25 ;
      LAYER M3 ;
      RECT 309.565 0.0 309.705 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[84]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 64.915 0.0 65.055 0.25 ;
      LAYER M2 ;
      RECT 64.915 0.0 65.055 0.25 ;
      LAYER M1 ;
      RECT 64.915 0.0 65.055 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[19]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 311.255 0.0 311.395 0.25 ;
      LAYER M2 ;
      RECT 311.255 0.0 311.395 0.25 ;
      LAYER M3 ;
      RECT 311.255 0.0 311.395 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[85]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.225 0.0 63.365 0.25 ;
      LAYER M2 ;
      RECT 63.225 0.0 63.365 0.25 ;
      LAYER M1 ;
      RECT 63.225 0.0 63.365 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[18]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 312.885 0.0 313.025 0.25 ;
      LAYER M2 ;
      RECT 312.885 0.0 313.025 0.25 ;
      LAYER M3 ;
      RECT 312.885 0.0 313.025 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[85]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 61.595 0.0 61.735 0.25 ;
      LAYER M2 ;
      RECT 61.595 0.0 61.735 0.25 ;
      LAYER M1 ;
      RECT 61.595 0.0 61.735 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[18]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 314.575 0.0 314.715 0.25 ;
      LAYER M2 ;
      RECT 314.575 0.0 314.715 0.25 ;
      LAYER M3 ;
      RECT 314.575 0.0 314.715 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[86]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 59.905 0.0 60.045 0.25 ;
      LAYER M2 ;
      RECT 59.905 0.0 60.045 0.25 ;
      LAYER M1 ;
      RECT 59.905 0.0 60.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[17]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 316.205 0.0 316.345 0.25 ;
      LAYER M2 ;
      RECT 316.205 0.0 316.345 0.25 ;
      LAYER M3 ;
      RECT 316.205 0.0 316.345 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[86]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 58.275 0.0 58.415 0.25 ;
      LAYER M2 ;
      RECT 58.275 0.0 58.415 0.25 ;
      LAYER M1 ;
      RECT 58.275 0.0 58.415 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[17]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 317.895 0.0 318.035 0.25 ;
      LAYER M2 ;
      RECT 317.895 0.0 318.035 0.25 ;
      LAYER M3 ;
      RECT 317.895 0.0 318.035 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[87]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.585 0.0 56.725 0.25 ;
      LAYER M2 ;
      RECT 56.585 0.0 56.725 0.25 ;
      LAYER M1 ;
      RECT 56.585 0.0 56.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[16]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 319.525 0.0 319.665 0.25 ;
      LAYER M2 ;
      RECT 319.525 0.0 319.665 0.25 ;
      LAYER M3 ;
      RECT 319.525 0.0 319.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[87]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 54.955 0.0 55.095 0.25 ;
      LAYER M2 ;
      RECT 54.955 0.0 55.095 0.25 ;
      LAYER M1 ;
      RECT 54.955 0.0 55.095 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[16]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 321.215 0.0 321.355 0.25 ;
      LAYER M2 ;
      RECT 321.215 0.0 321.355 0.25 ;
      LAYER M3 ;
      RECT 321.215 0.0 321.355 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[88]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 53.265 0.0 53.405 0.25 ;
      LAYER M2 ;
      RECT 53.265 0.0 53.405 0.25 ;
      LAYER M1 ;
      RECT 53.265 0.0 53.405 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[15]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 322.845 0.0 322.985 0.25 ;
      LAYER M2 ;
      RECT 322.845 0.0 322.985 0.25 ;
      LAYER M3 ;
      RECT 322.845 0.0 322.985 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[88]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 51.635 0.0 51.775 0.25 ;
      LAYER M2 ;
      RECT 51.635 0.0 51.775 0.25 ;
      LAYER M1 ;
      RECT 51.635 0.0 51.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[15]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 324.535 0.0 324.675 0.25 ;
      LAYER M2 ;
      RECT 324.535 0.0 324.675 0.25 ;
      LAYER M3 ;
      RECT 324.535 0.0 324.675 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[89]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.945 0.0 50.085 0.25 ;
      LAYER M2 ;
      RECT 49.945 0.0 50.085 0.25 ;
      LAYER M1 ;
      RECT 49.945 0.0 50.085 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[14]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 326.165 0.0 326.305 0.25 ;
      LAYER M2 ;
      RECT 326.165 0.0 326.305 0.25 ;
      LAYER M3 ;
      RECT 326.165 0.0 326.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[89]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 48.315 0.0 48.455 0.25 ;
      LAYER M2 ;
      RECT 48.315 0.0 48.455 0.25 ;
      LAYER M1 ;
      RECT 48.315 0.0 48.455 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[14]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 327.855 0.0 327.995 0.25 ;
      LAYER M2 ;
      RECT 327.855 0.0 327.995 0.25 ;
      LAYER M3 ;
      RECT 327.855 0.0 327.995 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[90]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 46.625 0.0 46.765 0.25 ;
      LAYER M2 ;
      RECT 46.625 0.0 46.765 0.25 ;
      LAYER M1 ;
      RECT 46.625 0.0 46.765 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[13]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 329.485 0.0 329.625 0.25 ;
      LAYER M2 ;
      RECT 329.485 0.0 329.625 0.25 ;
      LAYER M3 ;
      RECT 329.485 0.0 329.625 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[90]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.995 0.0 45.135 0.25 ;
      LAYER M2 ;
      RECT 44.995 0.0 45.135 0.25 ;
      LAYER M1 ;
      RECT 44.995 0.0 45.135 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[13]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 331.175 0.0 331.315 0.25 ;
      LAYER M2 ;
      RECT 331.175 0.0 331.315 0.25 ;
      LAYER M3 ;
      RECT 331.175 0.0 331.315 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[91]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.305 0.0 43.445 0.25 ;
      LAYER M2 ;
      RECT 43.305 0.0 43.445 0.25 ;
      LAYER M1 ;
      RECT 43.305 0.0 43.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[12]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 332.805 0.0 332.945 0.25 ;
      LAYER M2 ;
      RECT 332.805 0.0 332.945 0.25 ;
      LAYER M3 ;
      RECT 332.805 0.0 332.945 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[91]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 41.675 0.0 41.815 0.25 ;
      LAYER M2 ;
      RECT 41.675 0.0 41.815 0.25 ;
      LAYER M1 ;
      RECT 41.675 0.0 41.815 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[12]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 334.495 0.0 334.635 0.25 ;
      LAYER M2 ;
      RECT 334.495 0.0 334.635 0.25 ;
      LAYER M3 ;
      RECT 334.495 0.0 334.635 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[92]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.985 0.0 40.125 0.25 ;
      LAYER M2 ;
      RECT 39.985 0.0 40.125 0.25 ;
      LAYER M1 ;
      RECT 39.985 0.0 40.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[11]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 336.125 0.0 336.265 0.25 ;
      LAYER M2 ;
      RECT 336.125 0.0 336.265 0.25 ;
      LAYER M3 ;
      RECT 336.125 0.0 336.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[92]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.355 0.0 38.495 0.25 ;
      LAYER M2 ;
      RECT 38.355 0.0 38.495 0.25 ;
      LAYER M1 ;
      RECT 38.355 0.0 38.495 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[11]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 337.815 0.0 337.955 0.25 ;
      LAYER M2 ;
      RECT 337.815 0.0 337.955 0.25 ;
      LAYER M3 ;
      RECT 337.815 0.0 337.955 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[93]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 36.665 0.0 36.805 0.25 ;
      LAYER M2 ;
      RECT 36.665 0.0 36.805 0.25 ;
      LAYER M1 ;
      RECT 36.665 0.0 36.805 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[10]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 339.445 0.0 339.585 0.25 ;
      LAYER M2 ;
      RECT 339.445 0.0 339.585 0.25 ;
      LAYER M3 ;
      RECT 339.445 0.0 339.585 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[93]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 35.035 0.0 35.175 0.25 ;
      LAYER M2 ;
      RECT 35.035 0.0 35.175 0.25 ;
      LAYER M1 ;
      RECT 35.035 0.0 35.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[10]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 341.135 0.0 341.275 0.25 ;
      LAYER M2 ;
      RECT 341.135 0.0 341.275 0.25 ;
      LAYER M3 ;
      RECT 341.135 0.0 341.275 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[94]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 33.345 0.0 33.485 0.25 ;
      LAYER M2 ;
      RECT 33.345 0.0 33.485 0.25 ;
      LAYER M1 ;
      RECT 33.345 0.0 33.485 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[9]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 342.765 0.0 342.905 0.25 ;
      LAYER M2 ;
      RECT 342.765 0.0 342.905 0.25 ;
      LAYER M3 ;
      RECT 342.765 0.0 342.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[94]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 31.715 0.0 31.855 0.25 ;
      LAYER M2 ;
      RECT 31.715 0.0 31.855 0.25 ;
      LAYER M1 ;
      RECT 31.715 0.0 31.855 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[9]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 344.455 0.0 344.595 0.25 ;
      LAYER M2 ;
      RECT 344.455 0.0 344.595 0.25 ;
      LAYER M3 ;
      RECT 344.455 0.0 344.595 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[95]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 30.025 0.0 30.165 0.25 ;
      LAYER M2 ;
      RECT 30.025 0.0 30.165 0.25 ;
      LAYER M1 ;
      RECT 30.025 0.0 30.165 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[8]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 346.085 0.0 346.225 0.25 ;
      LAYER M2 ;
      RECT 346.085 0.0 346.225 0.25 ;
      LAYER M3 ;
      RECT 346.085 0.0 346.225 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[95]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 28.395 0.0 28.535 0.25 ;
      LAYER M2 ;
      RECT 28.395 0.0 28.535 0.25 ;
      LAYER M1 ;
      RECT 28.395 0.0 28.535 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[8]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 347.775 0.0 347.915 0.25 ;
      LAYER M2 ;
      RECT 347.775 0.0 347.915 0.25 ;
      LAYER M3 ;
      RECT 347.775 0.0 347.915 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[96]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.705 0.0 26.845 0.25 ;
      LAYER M2 ;
      RECT 26.705 0.0 26.845 0.25 ;
      LAYER M1 ;
      RECT 26.705 0.0 26.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[7]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 349.405 0.0 349.545 0.25 ;
      LAYER M2 ;
      RECT 349.405 0.0 349.545 0.25 ;
      LAYER M3 ;
      RECT 349.405 0.0 349.545 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[96]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.075 0.0 25.215 0.25 ;
      LAYER M2 ;
      RECT 25.075 0.0 25.215 0.25 ;
      LAYER M1 ;
      RECT 25.075 0.0 25.215 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[7]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 351.095 0.0 351.235 0.25 ;
      LAYER M2 ;
      RECT 351.095 0.0 351.235 0.25 ;
      LAYER M3 ;
      RECT 351.095 0.0 351.235 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[97]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 23.385 0.0 23.525 0.25 ;
      LAYER M2 ;
      RECT 23.385 0.0 23.525 0.25 ;
      LAYER M1 ;
      RECT 23.385 0.0 23.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[6]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 352.725 0.0 352.865 0.25 ;
      LAYER M2 ;
      RECT 352.725 0.0 352.865 0.25 ;
      LAYER M3 ;
      RECT 352.725 0.0 352.865 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[97]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 21.755 0.0 21.895 0.25 ;
      LAYER M2 ;
      RECT 21.755 0.0 21.895 0.25 ;
      LAYER M1 ;
      RECT 21.755 0.0 21.895 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[6]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 354.415 0.0 354.555 0.25 ;
      LAYER M2 ;
      RECT 354.415 0.0 354.555 0.25 ;
      LAYER M3 ;
      RECT 354.415 0.0 354.555 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[98]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 20.065 0.0 20.205 0.25 ;
      LAYER M2 ;
      RECT 20.065 0.0 20.205 0.25 ;
      LAYER M1 ;
      RECT 20.065 0.0 20.205 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[5]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 356.045 0.0 356.185 0.25 ;
      LAYER M2 ;
      RECT 356.045 0.0 356.185 0.25 ;
      LAYER M3 ;
      RECT 356.045 0.0 356.185 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[98]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 18.435 0.0 18.575 0.25 ;
      LAYER M2 ;
      RECT 18.435 0.0 18.575 0.25 ;
      LAYER M1 ;
      RECT 18.435 0.0 18.575 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[5]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 357.735 0.0 357.875 0.25 ;
      LAYER M2 ;
      RECT 357.735 0.0 357.875 0.25 ;
      LAYER M3 ;
      RECT 357.735 0.0 357.875 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[99]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 16.745 0.0 16.885 0.25 ;
      LAYER M2 ;
      RECT 16.745 0.0 16.885 0.25 ;
      LAYER M1 ;
      RECT 16.745 0.0 16.885 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[4]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 359.365 0.0 359.505 0.25 ;
      LAYER M2 ;
      RECT 359.365 0.0 359.505 0.25 ;
      LAYER M3 ;
      RECT 359.365 0.0 359.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[99]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 15.115 0.0 15.255 0.25 ;
      LAYER M2 ;
      RECT 15.115 0.0 15.255 0.25 ;
      LAYER M1 ;
      RECT 15.115 0.0 15.255 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[4]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 361.055 0.0 361.195 0.25 ;
      LAYER M2 ;
      RECT 361.055 0.0 361.195 0.25 ;
      LAYER M3 ;
      RECT 361.055 0.0 361.195 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[100]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.425 0.0 13.565 0.25 ;
      LAYER M2 ;
      RECT 13.425 0.0 13.565 0.25 ;
      LAYER M1 ;
      RECT 13.425 0.0 13.565 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[3]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 362.685 0.0 362.825 0.25 ;
      LAYER M2 ;
      RECT 362.685 0.0 362.825 0.25 ;
      LAYER M3 ;
      RECT 362.685 0.0 362.825 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[100]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 11.795 0.0 11.935 0.25 ;
      LAYER M2 ;
      RECT 11.795 0.0 11.935 0.25 ;
      LAYER M1 ;
      RECT 11.795 0.0 11.935 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[3]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 364.375 0.0 364.515 0.25 ;
      LAYER M2 ;
      RECT 364.375 0.0 364.515 0.25 ;
      LAYER M3 ;
      RECT 364.375 0.0 364.515 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[101]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.105 0.0 10.245 0.25 ;
      LAYER M2 ;
      RECT 10.105 0.0 10.245 0.25 ;
      LAYER M1 ;
      RECT 10.105 0.0 10.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[2]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 366.005 0.0 366.145 0.25 ;
      LAYER M2 ;
      RECT 366.005 0.0 366.145 0.25 ;
      LAYER M3 ;
      RECT 366.005 0.0 366.145 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[101]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.475 0.0 8.615 0.25 ;
      LAYER M2 ;
      RECT 8.475 0.0 8.615 0.25 ;
      LAYER M1 ;
      RECT 8.475 0.0 8.615 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[2]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 367.695 0.0 367.835 0.25 ;
      LAYER M2 ;
      RECT 367.695 0.0 367.835 0.25 ;
      LAYER M3 ;
      RECT 367.695 0.0 367.835 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[102]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.785 0.0 6.925 0.25 ;
      LAYER M2 ;
      RECT 6.785 0.0 6.925 0.25 ;
      LAYER M1 ;
      RECT 6.785 0.0 6.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[1]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 369.325 0.0 369.465 0.25 ;
      LAYER M2 ;
      RECT 369.325 0.0 369.465 0.25 ;
      LAYER M3 ;
      RECT 369.325 0.0 369.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[102]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.155 0.0 5.295 0.25 ;
      LAYER M2 ;
      RECT 5.155 0.0 5.295 0.25 ;
      LAYER M1 ;
      RECT 5.155 0.0 5.295 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[1]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 371.015 0.0 371.155 0.25 ;
      LAYER M2 ;
      RECT 371.015 0.0 371.155 0.25 ;
      LAYER M3 ;
      RECT 371.015 0.0 371.155 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[103]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.465 0.0 3.605 0.25 ;
      LAYER M2 ;
      RECT 3.465 0.0 3.605 0.25 ;
      LAYER M1 ;
      RECT 3.465 0.0 3.605 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END D[0]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 372.645 0.0 372.785 0.25 ;
      LAYER M2 ;
      RECT 372.645 0.0 372.785 0.25 ;
      LAYER M3 ;
      RECT 372.645 0.0 372.785 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[103]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.835 0.0 1.975 0.25 ;
      LAYER M2 ;
      RECT 1.835 0.0 1.975 0.25 ;
      LAYER M1 ;
      RECT 1.835 0.0 1.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END Q[0]
  PIN VDDPE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.59 0.0 0.7 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 0.995 0.0 1.275 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 4.315 0.0 4.595 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.635 0.0 7.915 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.955 0.0 11.235 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 14.275 0.0 14.555 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.595 0.0 17.875 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.915 0.0 21.195 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 24.235 0.0 24.515 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.555 0.0 27.835 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.875 0.0 31.155 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 34.195 0.0 34.475 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.515 0.0 37.795 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 40.835 0.0 41.115 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.155 0.0 44.435 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.475 0.0 47.755 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.795 0.0 51.075 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 54.115 0.0 54.395 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 57.435 0.0 57.715 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 60.755 0.0 61.035 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.075 0.0 64.355 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.395 0.0 67.675 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.715 0.0 70.995 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.035 0.0 74.315 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 77.355 0.0 77.635 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 80.675 0.0 80.955 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 83.995 0.0 84.275 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.315 0.0 87.595 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.635 0.0 90.915 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 93.955 0.0 94.235 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 97.275 0.0 97.555 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.595 0.0 100.875 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.915 0.0 104.195 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 107.235 0.0 107.515 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 110.555 0.0 110.835 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 113.875 0.0 114.155 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 117.195 0.0 117.475 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.515 0.0 120.795 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.835 0.0 124.115 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 127.155 0.0 127.435 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 130.475 0.0 130.755 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 133.795 0.0 134.075 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 137.115 0.0 137.395 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 140.435 0.0 140.715 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.755 0.0 144.035 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.075 0.0 147.355 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 150.395 0.0 150.675 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 153.715 0.0 153.995 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 157.035 0.0 157.315 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 160.355 0.0 160.635 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 163.675 0.0 163.955 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 166.995 0.0 167.275 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 170.315 0.0 170.595 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 173.715 0.0 173.825 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 175.495 0.0 175.605 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.8 0.0 178.08 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 180.44 0.0 180.65 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 181.185 0.0 181.335 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 181.825 0.0 182.055 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 182.535 0.0 182.805 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 184.505 0.0 184.775 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 186.695 0.0 186.905 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 189.62 0.0 189.9 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.71 0.0 190.85 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 191.45 0.0 191.6 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 191.81 0.0 192.08 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 195.02 0.0 195.3 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.43 0.0 196.64 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 198.955 0.0 199.095 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.885 0.0 200.095 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 200.795 0.0 200.905 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 204.025 0.0 204.305 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.345 0.0 207.625 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 210.665 0.0 210.945 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.985 0.0 214.265 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 217.305 0.0 217.585 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 220.625 0.0 220.905 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 223.945 0.0 224.225 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 227.265 0.0 227.545 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 230.585 0.0 230.865 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 233.905 0.0 234.185 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 237.225 0.0 237.505 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 240.545 0.0 240.825 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 243.865 0.0 244.145 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 247.185 0.0 247.465 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 250.505 0.0 250.785 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 253.825 0.0 254.105 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 257.145 0.0 257.425 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 260.465 0.0 260.745 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 263.785 0.0 264.065 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 267.105 0.0 267.385 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 270.425 0.0 270.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 273.745 0.0 274.025 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 277.065 0.0 277.345 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 280.385 0.0 280.665 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 283.705 0.0 283.985 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 287.025 0.0 287.305 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 290.345 0.0 290.625 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 293.665 0.0 293.945 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 296.985 0.0 297.265 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 300.305 0.0 300.585 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 303.625 0.0 303.905 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 306.945 0.0 307.225 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 310.265 0.0 310.545 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 313.585 0.0 313.865 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 316.905 0.0 317.185 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 320.225 0.0 320.505 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 323.545 0.0 323.825 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 326.865 0.0 327.145 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 330.185 0.0 330.465 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 333.505 0.0 333.785 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 336.825 0.0 337.105 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 340.145 0.0 340.425 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 343.465 0.0 343.745 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 346.785 0.0 347.065 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 350.105 0.0 350.385 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 353.425 0.0 353.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 356.745 0.0 357.025 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 360.065 0.0 360.345 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 363.385 0.0 363.665 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 366.705 0.0 366.985 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 370.025 0.0 370.305 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 373.345 0.0 373.625 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 373.92 0.0 374.03 61.255 ;
      END
    END VDDPE
  PIN VDDCE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.17 0.0 0.28 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 2.405 0.0 2.685 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 5.725 0.0 6.005 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 9.045 0.0 9.325 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.365 0.0 12.645 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.685 0.0 15.965 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.005 0.0 19.285 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 22.325 0.0 22.605 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.645 0.0 25.925 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.965 0.0 29.245 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.285 0.0 32.565 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.605 0.0 35.885 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.925 0.0 39.205 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.245 0.0 42.525 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.565 0.0 45.845 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.885 0.0 49.165 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 52.205 0.0 52.485 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.525 0.0 55.805 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.845 0.0 59.125 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 62.165 0.0 62.445 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 65.485 0.0 65.765 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.805 0.0 69.085 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.125 0.0 72.405 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.445 0.0 75.725 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.765 0.0 79.045 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.085 0.0 82.365 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 85.405 0.0 85.685 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.725 0.0 89.005 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.045 0.0 92.325 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 95.365 0.0 95.645 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.685 0.0 98.965 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 102.005 0.0 102.285 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 105.325 0.0 105.605 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.645 0.0 108.925 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 111.965 0.0 112.245 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 115.285 0.0 115.565 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.605 0.0 118.885 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 121.925 0.0 122.205 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 125.245 0.0 125.525 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.565 0.0 128.845 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 131.885 0.0 132.165 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 135.205 0.0 135.485 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 138.525 0.0 138.805 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 141.845 0.0 142.125 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 145.165 0.0 145.445 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 148.485 0.0 148.765 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 151.805 0.0 152.085 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 155.125 0.0 155.405 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 158.445 0.0 158.725 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 161.765 0.0 162.045 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 165.085 0.0 165.365 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 168.405 0.0 168.685 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 171.725 0.0 172.005 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 174.135 0.0 174.245 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 176.325 0.0 176.595 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 176.855 0.0 177.125 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 178.765 0.0 179.025 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 195.63 0.0 195.84 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 197.435 0.0 197.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 198.045 0.0 198.255 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 200.375 0.0 200.485 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 202.615 0.0 202.895 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 205.935 0.0 206.215 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 209.255 0.0 209.535 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 212.575 0.0 212.855 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.895 0.0 216.175 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 219.215 0.0 219.495 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 222.535 0.0 222.815 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.855 0.0 226.135 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.175 0.0 229.455 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.495 0.0 232.775 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.815 0.0 236.095 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.135 0.0 239.415 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.455 0.0 242.735 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 245.775 0.0 246.055 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.095 0.0 249.375 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.415 0.0 252.695 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 255.735 0.0 256.015 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 259.055 0.0 259.335 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.375 0.0 262.655 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 265.695 0.0 265.975 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 269.015 0.0 269.295 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 272.335 0.0 272.615 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 275.655 0.0 275.935 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 278.975 0.0 279.255 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 282.295 0.0 282.575 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 285.615 0.0 285.895 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 288.935 0.0 289.215 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 292.255 0.0 292.535 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 295.575 0.0 295.855 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 298.895 0.0 299.175 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 302.215 0.0 302.495 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 305.535 0.0 305.815 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 308.855 0.0 309.135 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 312.175 0.0 312.455 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 315.495 0.0 315.775 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 318.815 0.0 319.095 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 322.135 0.0 322.415 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 325.455 0.0 325.735 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 328.775 0.0 329.055 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 332.095 0.0 332.375 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 335.415 0.0 335.695 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 338.735 0.0 339.015 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 342.055 0.0 342.335 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 345.375 0.0 345.655 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 348.695 0.0 348.975 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 352.015 0.0 352.295 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 355.335 0.0 355.615 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 358.655 0.0 358.935 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 361.975 0.0 362.255 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 365.295 0.0 365.575 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 368.615 0.0 368.895 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 371.935 0.0 372.215 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 374.34 0.0 374.45 61.255 ;
      END
    END VDDCE
  PIN VSSE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.38 0.0 0.49 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 1.915 0.0 2.195 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 5.235 0.0 5.515 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 8.555 0.0 8.835 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 11.875 0.0 12.155 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.195 0.0 15.475 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 18.515 0.0 18.795 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 21.835 0.0 22.115 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.155 0.0 25.435 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.475 0.0 28.755 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 31.795 0.0 32.075 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.115 0.0 35.395 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.435 0.0 38.715 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 41.755 0.0 42.035 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.075 0.0 45.355 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.395 0.0 48.675 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.715 0.0 51.995 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.035 0.0 55.315 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.355 0.0 58.635 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.675 0.0 61.955 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.995 0.0 65.275 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.315 0.0 68.595 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 71.635 0.0 71.915 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.955 0.0 75.235 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.275 0.0 78.555 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.595 0.0 81.875 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.915 0.0 85.195 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.235 0.0 88.515 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 91.555 0.0 91.835 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.875 0.0 95.155 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.195 0.0 98.475 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 101.515 0.0 101.795 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 104.835 0.0 105.115 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.155 0.0 108.435 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 111.475 0.0 111.755 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 114.795 0.0 115.075 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.115 0.0 118.395 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 121.435 0.0 121.715 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 124.755 0.0 125.035 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.075 0.0 128.355 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 131.395 0.0 131.675 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 134.715 0.0 134.995 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 138.035 0.0 138.315 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 141.355 0.0 141.635 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.675 0.0 144.955 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.995 0.0 148.275 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 151.315 0.0 151.595 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 154.635 0.0 154.915 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 157.955 0.0 158.235 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 161.275 0.0 161.555 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 164.595 0.0 164.875 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 167.915 0.0 168.195 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 171.235 0.0 171.515 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 173.925 0.0 174.035 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 174.52 0.0 174.67 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 175.16 0.0 175.37 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.34 0.0 177.62 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 178.23 0.0 178.44 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 179.85 0.0 180.12 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 183.675 0.0 183.825 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 184.895 0.0 185.005 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.425 0.0 187.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.04 0.0 190.25 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 193.975 0.0 194.125 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 194.5 0.0 194.78 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.15 0.0 196.29 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.78 0.0 197.05 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.245 0.0 199.525 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 200.585 0.0 200.695 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 203.105 0.0 203.385 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 206.425 0.0 206.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 209.745 0.0 210.025 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.065 0.0 213.345 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 216.385 0.0 216.665 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 219.705 0.0 219.985 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 223.025 0.0 223.305 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 226.345 0.0 226.625 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.665 0.0 229.945 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.985 0.0 233.265 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 236.305 0.0 236.585 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.625 0.0 239.905 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.945 0.0 243.225 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 246.265 0.0 246.545 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.585 0.0 249.865 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.905 0.0 253.185 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 256.225 0.0 256.505 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 259.545 0.0 259.825 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.865 0.0 263.145 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 266.185 0.0 266.465 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 269.505 0.0 269.785 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 272.825 0.0 273.105 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 276.145 0.0 276.425 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 279.465 0.0 279.745 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 282.785 0.0 283.065 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 286.105 0.0 286.385 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 289.425 0.0 289.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 292.745 0.0 293.025 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 296.065 0.0 296.345 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 299.385 0.0 299.665 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 302.705 0.0 302.985 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 306.025 0.0 306.305 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 309.345 0.0 309.625 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 312.665 0.0 312.945 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 315.985 0.0 316.265 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 319.305 0.0 319.585 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 322.625 0.0 322.905 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 325.945 0.0 326.225 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 329.265 0.0 329.545 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 332.585 0.0 332.865 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 335.905 0.0 336.185 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 339.225 0.0 339.505 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 342.545 0.0 342.825 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 345.865 0.0 346.145 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 349.185 0.0 349.465 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 352.505 0.0 352.785 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 355.825 0.0 356.105 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 359.145 0.0 359.425 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 362.465 0.0 362.745 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 365.785 0.0 366.065 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 369.105 0.0 369.385 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 372.425 0.0 372.705 61.255 ;
      END
    PORT
      LAYER M4 ;
      RECT 374.13 0.0 374.24 61.255 ;
      END
    END VSSE
  OBS
    #otc obstructions
    LAYER M1 DESIGNRULEWIDTH 0.07 ;
    RECT 372.925 0.0 374.62 0.32 ;
    RECT 371.295 0.0 372.505 0.32 ;
    RECT 369.605 0.0 370.875 0.32 ;
    RECT 367.975 0.0 369.185 0.32 ;
    RECT 366.285 0.0 367.555 0.32 ;
    RECT 364.655 0.0 365.865 0.32 ;
    RECT 362.965 0.0 364.235 0.32 ;
    RECT 361.335 0.0 362.545 0.32 ;
    RECT 359.645 0.0 360.915 0.32 ;
    RECT 358.015 0.0 359.225 0.32 ;
    RECT 356.325 0.0 357.595 0.32 ;
    RECT 354.695 0.0 355.905 0.32 ;
    RECT 353.005 0.0 354.275 0.32 ;
    RECT 351.375 0.0 352.585 0.32 ;
    RECT 349.685 0.0 350.955 0.32 ;
    RECT 348.055 0.0 349.265 0.32 ;
    RECT 346.365 0.0 347.635 0.32 ;
    RECT 344.735 0.0 345.945 0.32 ;
    RECT 343.045 0.0 344.315 0.32 ;
    RECT 341.415 0.0 342.625 0.32 ;
    RECT 339.725 0.0 340.995 0.32 ;
    RECT 338.095 0.0 339.305 0.32 ;
    RECT 336.405 0.0 337.675 0.32 ;
    RECT 334.775 0.0 335.985 0.32 ;
    RECT 333.085 0.0 334.355 0.32 ;
    RECT 331.455 0.0 332.665 0.32 ;
    RECT 329.765 0.0 331.035 0.32 ;
    RECT 328.135 0.0 329.345 0.32 ;
    RECT 326.445 0.0 327.715 0.32 ;
    RECT 324.815 0.0 326.025 0.32 ;
    RECT 323.125 0.0 324.395 0.32 ;
    RECT 321.495 0.0 322.705 0.32 ;
    RECT 319.805 0.0 321.075 0.32 ;
    RECT 318.175 0.0 319.385 0.32 ;
    RECT 316.485 0.0 317.755 0.32 ;
    RECT 314.855 0.0 316.065 0.32 ;
    RECT 313.165 0.0 314.435 0.32 ;
    RECT 311.535 0.0 312.745 0.32 ;
    RECT 309.845 0.0 311.115 0.32 ;
    RECT 308.215 0.0 309.425 0.32 ;
    RECT 306.525 0.0 307.795 0.32 ;
    RECT 304.895 0.0 306.105 0.32 ;
    RECT 303.205 0.0 304.475 0.32 ;
    RECT 301.575 0.0 302.785 0.32 ;
    RECT 299.885 0.0 301.155 0.32 ;
    RECT 298.255 0.0 299.465 0.32 ;
    RECT 296.565 0.0 297.835 0.32 ;
    RECT 294.935 0.0 296.145 0.32 ;
    RECT 293.245 0.0 294.515 0.32 ;
    RECT 291.615 0.0 292.825 0.32 ;
    RECT 289.925 0.0 291.195 0.32 ;
    RECT 288.295 0.0 289.505 0.32 ;
    RECT 286.605 0.0 287.875 0.32 ;
    RECT 284.975 0.0 286.185 0.32 ;
    RECT 283.285 0.0 284.555 0.32 ;
    RECT 281.655 0.0 282.865 0.32 ;
    RECT 279.965 0.0 281.235 0.32 ;
    RECT 278.335 0.0 279.545 0.32 ;
    RECT 276.645 0.0 277.915 0.32 ;
    RECT 275.015 0.0 276.225 0.32 ;
    RECT 273.325 0.0 274.595 0.32 ;
    RECT 271.695 0.0 272.905 0.32 ;
    RECT 270.005 0.0 271.275 0.32 ;
    RECT 268.375 0.0 269.585 0.32 ;
    RECT 266.685 0.0 267.955 0.32 ;
    RECT 265.055 0.0 266.265 0.32 ;
    RECT 263.365 0.0 264.635 0.32 ;
    RECT 261.735 0.0 262.945 0.32 ;
    RECT 260.045 0.0 261.315 0.32 ;
    RECT 258.415 0.0 259.625 0.32 ;
    RECT 256.725 0.0 257.995 0.32 ;
    RECT 255.095 0.0 256.305 0.32 ;
    RECT 253.405 0.0 254.675 0.32 ;
    RECT 251.775 0.0 252.985 0.32 ;
    RECT 250.085 0.0 251.355 0.32 ;
    RECT 248.455 0.0 249.665 0.32 ;
    RECT 246.765 0.0 248.035 0.32 ;
    RECT 245.135 0.0 246.345 0.32 ;
    RECT 243.445 0.0 244.715 0.32 ;
    RECT 241.815 0.0 243.025 0.32 ;
    RECT 240.125 0.0 241.395 0.32 ;
    RECT 238.495 0.0 239.705 0.32 ;
    RECT 236.805 0.0 238.075 0.32 ;
    RECT 235.175 0.0 236.385 0.32 ;
    RECT 233.485 0.0 234.755 0.32 ;
    RECT 231.855 0.0 233.065 0.32 ;
    RECT 230.165 0.0 231.435 0.32 ;
    RECT 228.535 0.0 229.745 0.32 ;
    RECT 226.845 0.0 228.115 0.32 ;
    RECT 225.215 0.0 226.425 0.32 ;
    RECT 223.525 0.0 224.795 0.32 ;
    RECT 221.895 0.0 223.105 0.32 ;
    RECT 220.205 0.0 221.475 0.32 ;
    RECT 218.575 0.0 219.785 0.32 ;
    RECT 216.885 0.0 218.155 0.32 ;
    RECT 215.255 0.0 216.465 0.32 ;
    RECT 213.565 0.0 214.835 0.32 ;
    RECT 211.935 0.0 213.145 0.32 ;
    RECT 210.245 0.0 211.515 0.32 ;
    RECT 208.615 0.0 209.825 0.32 ;
    RECT 206.925 0.0 208.195 0.32 ;
    RECT 205.295 0.0 206.505 0.32 ;
    RECT 203.605 0.0 204.875 0.32 ;
    RECT 201.975 0.0 203.185 0.32 ;
    RECT 200.92 0.0 201.555 0.32 ;
    RECT 197.765 0.0 200.5 0.32 ;
    RECT 194.37 0.0 197.345 0.32 ;
    RECT 191.935 0.0 193.665 0.32 ;
    RECT 190.97 0.0 191.12 0.32 ;
    RECT 189.89 0.0 190.27 0.32 ;
    RECT 187.535 0.0 189.47 0.32 ;
    RECT 185.93 0.0 187.115 0.32 ;
    RECT 182.11 0.0 185.09 0.32 ;
    RECT 179.82 0.0 181.41 0.32 ;
    RECT 178.845 0.0 179.4 0.32 ;
    RECT 178.03 0.0 178.425 0.32 ;
    RECT 174.755 0.0 177.61 0.32 ;
    RECT 174.11 0.0 174.335 0.32 ;
    RECT 173.065 0.0 173.69 0.32 ;
    RECT 171.435 0.0 172.645 0.32 ;
    RECT 169.745 0.0 171.015 0.32 ;
    RECT 168.115 0.0 169.325 0.32 ;
    RECT 166.425 0.0 167.695 0.32 ;
    RECT 164.795 0.0 166.005 0.32 ;
    RECT 163.105 0.0 164.375 0.32 ;
    RECT 161.475 0.0 162.685 0.32 ;
    RECT 159.785 0.0 161.055 0.32 ;
    RECT 158.155 0.0 159.365 0.32 ;
    RECT 156.465 0.0 157.735 0.32 ;
    RECT 154.835 0.0 156.045 0.32 ;
    RECT 153.145 0.0 154.415 0.32 ;
    RECT 151.515 0.0 152.725 0.32 ;
    RECT 149.825 0.0 151.095 0.32 ;
    RECT 148.195 0.0 149.405 0.32 ;
    RECT 146.505 0.0 147.775 0.32 ;
    RECT 144.875 0.0 146.085 0.32 ;
    RECT 143.185 0.0 144.455 0.32 ;
    RECT 141.555 0.0 142.765 0.32 ;
    RECT 139.865 0.0 141.135 0.32 ;
    RECT 138.235 0.0 139.445 0.32 ;
    RECT 136.545 0.0 137.815 0.32 ;
    RECT 134.915 0.0 136.125 0.32 ;
    RECT 133.225 0.0 134.495 0.32 ;
    RECT 131.595 0.0 132.805 0.32 ;
    RECT 129.905 0.0 131.175 0.32 ;
    RECT 128.275 0.0 129.485 0.32 ;
    RECT 126.585 0.0 127.855 0.32 ;
    RECT 124.955 0.0 126.165 0.32 ;
    RECT 123.265 0.0 124.535 0.32 ;
    RECT 121.635 0.0 122.845 0.32 ;
    RECT 119.945 0.0 121.215 0.32 ;
    RECT 118.315 0.0 119.525 0.32 ;
    RECT 116.625 0.0 117.895 0.32 ;
    RECT 114.995 0.0 116.205 0.32 ;
    RECT 113.305 0.0 114.575 0.32 ;
    RECT 111.675 0.0 112.885 0.32 ;
    RECT 109.985 0.0 111.255 0.32 ;
    RECT 108.355 0.0 109.565 0.32 ;
    RECT 106.665 0.0 107.935 0.32 ;
    RECT 105.035 0.0 106.245 0.32 ;
    RECT 103.345 0.0 104.615 0.32 ;
    RECT 101.715 0.0 102.925 0.32 ;
    RECT 100.025 0.0 101.295 0.32 ;
    RECT 98.395 0.0 99.605 0.32 ;
    RECT 96.705 0.0 97.975 0.32 ;
    RECT 95.075 0.0 96.285 0.32 ;
    RECT 93.385 0.0 94.655 0.32 ;
    RECT 91.755 0.0 92.965 0.32 ;
    RECT 90.065 0.0 91.335 0.32 ;
    RECT 88.435 0.0 89.645 0.32 ;
    RECT 86.745 0.0 88.015 0.32 ;
    RECT 85.115 0.0 86.325 0.32 ;
    RECT 83.425 0.0 84.695 0.32 ;
    RECT 81.795 0.0 83.005 0.32 ;
    RECT 80.105 0.0 81.375 0.32 ;
    RECT 78.475 0.0 79.685 0.32 ;
    RECT 76.785 0.0 78.055 0.32 ;
    RECT 75.155 0.0 76.365 0.32 ;
    RECT 73.465 0.0 74.735 0.32 ;
    RECT 71.835 0.0 73.045 0.32 ;
    RECT 70.145 0.0 71.415 0.32 ;
    RECT 68.515 0.0 69.725 0.32 ;
    RECT 66.825 0.0 68.095 0.32 ;
    RECT 65.195 0.0 66.405 0.32 ;
    RECT 63.505 0.0 64.775 0.32 ;
    RECT 61.875 0.0 63.085 0.32 ;
    RECT 60.185 0.0 61.455 0.32 ;
    RECT 58.555 0.0 59.765 0.32 ;
    RECT 56.865 0.0 58.135 0.32 ;
    RECT 55.235 0.0 56.445 0.32 ;
    RECT 53.545 0.0 54.815 0.32 ;
    RECT 51.915 0.0 53.125 0.32 ;
    RECT 50.225 0.0 51.495 0.32 ;
    RECT 48.595 0.0 49.805 0.32 ;
    RECT 46.905 0.0 48.175 0.32 ;
    RECT 45.275 0.0 46.485 0.32 ;
    RECT 43.585 0.0 44.855 0.32 ;
    RECT 41.955 0.0 43.165 0.32 ;
    RECT 40.265 0.0 41.535 0.32 ;
    RECT 38.635 0.0 39.845 0.32 ;
    RECT 36.945 0.0 38.215 0.32 ;
    RECT 35.315 0.0 36.525 0.32 ;
    RECT 33.625 0.0 34.895 0.32 ;
    RECT 31.995 0.0 33.205 0.32 ;
    RECT 30.305 0.0 31.575 0.32 ;
    RECT 28.675 0.0 29.885 0.32 ;
    RECT 26.985 0.0 28.255 0.32 ;
    RECT 25.355 0.0 26.565 0.32 ;
    RECT 23.665 0.0 24.935 0.32 ;
    RECT 22.035 0.0 23.245 0.32 ;
    RECT 20.345 0.0 21.615 0.32 ;
    RECT 18.715 0.0 19.925 0.32 ;
    RECT 17.025 0.0 18.295 0.32 ;
    RECT 15.395 0.0 16.605 0.32 ;
    RECT 13.705 0.0 14.975 0.32 ;
    RECT 12.075 0.0 13.285 0.32 ;
    RECT 10.385 0.0 11.655 0.32 ;
    RECT 8.755 0.0 9.965 0.32 ;
    RECT 7.065 0.0 8.335 0.32 ;
    RECT 5.435 0.0 6.645 0.32 ;
    RECT 3.745 0.0 5.015 0.32 ;
    RECT 2.115 0.0 3.325 0.32 ;
    RECT 0.0 0.0 1.695 0.32 ;
    RECT 0.0 0.32 374.62 61.255 ;
    LAYER V1 ;
    RECT 0.0 0.0 374.62 61.255 ;
    LAYER M2 DESIGNRULEWIDTH 0.07 ;
    RECT 372.925 0.0 374.62 0.32 ;
    RECT 371.295 0.0 372.505 0.32 ;
    RECT 369.605 0.0 370.875 0.32 ;
    RECT 367.975 0.0 369.185 0.32 ;
    RECT 366.285 0.0 367.555 0.32 ;
    RECT 364.655 0.0 365.865 0.32 ;
    RECT 362.965 0.0 364.235 0.32 ;
    RECT 361.335 0.0 362.545 0.32 ;
    RECT 359.645 0.0 360.915 0.32 ;
    RECT 358.015 0.0 359.225 0.32 ;
    RECT 356.325 0.0 357.595 0.32 ;
    RECT 354.695 0.0 355.905 0.32 ;
    RECT 353.005 0.0 354.275 0.32 ;
    RECT 351.375 0.0 352.585 0.32 ;
    RECT 349.685 0.0 350.955 0.32 ;
    RECT 348.055 0.0 349.265 0.32 ;
    RECT 346.365 0.0 347.635 0.32 ;
    RECT 344.735 0.0 345.945 0.32 ;
    RECT 343.045 0.0 344.315 0.32 ;
    RECT 341.415 0.0 342.625 0.32 ;
    RECT 339.725 0.0 340.995 0.32 ;
    RECT 338.095 0.0 339.305 0.32 ;
    RECT 336.405 0.0 337.675 0.32 ;
    RECT 334.775 0.0 335.985 0.32 ;
    RECT 333.085 0.0 334.355 0.32 ;
    RECT 331.455 0.0 332.665 0.32 ;
    RECT 329.765 0.0 331.035 0.32 ;
    RECT 328.135 0.0 329.345 0.32 ;
    RECT 326.445 0.0 327.715 0.32 ;
    RECT 324.815 0.0 326.025 0.32 ;
    RECT 323.125 0.0 324.395 0.32 ;
    RECT 321.495 0.0 322.705 0.32 ;
    RECT 319.805 0.0 321.075 0.32 ;
    RECT 318.175 0.0 319.385 0.32 ;
    RECT 316.485 0.0 317.755 0.32 ;
    RECT 314.855 0.0 316.065 0.32 ;
    RECT 313.165 0.0 314.435 0.32 ;
    RECT 311.535 0.0 312.745 0.32 ;
    RECT 309.845 0.0 311.115 0.32 ;
    RECT 308.215 0.0 309.425 0.32 ;
    RECT 306.525 0.0 307.795 0.32 ;
    RECT 304.895 0.0 306.105 0.32 ;
    RECT 303.205 0.0 304.475 0.32 ;
    RECT 301.575 0.0 302.785 0.32 ;
    RECT 299.885 0.0 301.155 0.32 ;
    RECT 298.255 0.0 299.465 0.32 ;
    RECT 296.565 0.0 297.835 0.32 ;
    RECT 294.935 0.0 296.145 0.32 ;
    RECT 293.245 0.0 294.515 0.32 ;
    RECT 291.615 0.0 292.825 0.32 ;
    RECT 289.925 0.0 291.195 0.32 ;
    RECT 288.295 0.0 289.505 0.32 ;
    RECT 286.605 0.0 287.875 0.32 ;
    RECT 284.975 0.0 286.185 0.32 ;
    RECT 283.285 0.0 284.555 0.32 ;
    RECT 281.655 0.0 282.865 0.32 ;
    RECT 279.965 0.0 281.235 0.32 ;
    RECT 278.335 0.0 279.545 0.32 ;
    RECT 276.645 0.0 277.915 0.32 ;
    RECT 275.015 0.0 276.225 0.32 ;
    RECT 273.325 0.0 274.595 0.32 ;
    RECT 271.695 0.0 272.905 0.32 ;
    RECT 270.005 0.0 271.275 0.32 ;
    RECT 268.375 0.0 269.585 0.32 ;
    RECT 266.685 0.0 267.955 0.32 ;
    RECT 265.055 0.0 266.265 0.32 ;
    RECT 263.365 0.0 264.635 0.32 ;
    RECT 261.735 0.0 262.945 0.32 ;
    RECT 260.045 0.0 261.315 0.32 ;
    RECT 258.415 0.0 259.625 0.32 ;
    RECT 256.725 0.0 257.995 0.32 ;
    RECT 255.095 0.0 256.305 0.32 ;
    RECT 253.405 0.0 254.675 0.32 ;
    RECT 251.775 0.0 252.985 0.32 ;
    RECT 250.085 0.0 251.355 0.32 ;
    RECT 248.455 0.0 249.665 0.32 ;
    RECT 246.765 0.0 248.035 0.32 ;
    RECT 245.135 0.0 246.345 0.32 ;
    RECT 243.445 0.0 244.715 0.32 ;
    RECT 241.815 0.0 243.025 0.32 ;
    RECT 240.125 0.0 241.395 0.32 ;
    RECT 238.495 0.0 239.705 0.32 ;
    RECT 236.805 0.0 238.075 0.32 ;
    RECT 235.175 0.0 236.385 0.32 ;
    RECT 233.485 0.0 234.755 0.32 ;
    RECT 231.855 0.0 233.065 0.32 ;
    RECT 230.165 0.0 231.435 0.32 ;
    RECT 228.535 0.0 229.745 0.32 ;
    RECT 226.845 0.0 228.115 0.32 ;
    RECT 225.215 0.0 226.425 0.32 ;
    RECT 223.525 0.0 224.795 0.32 ;
    RECT 221.895 0.0 223.105 0.32 ;
    RECT 220.205 0.0 221.475 0.32 ;
    RECT 218.575 0.0 219.785 0.32 ;
    RECT 216.885 0.0 218.155 0.32 ;
    RECT 215.255 0.0 216.465 0.32 ;
    RECT 213.565 0.0 214.835 0.32 ;
    RECT 211.935 0.0 213.145 0.32 ;
    RECT 210.245 0.0 211.515 0.32 ;
    RECT 208.615 0.0 209.825 0.32 ;
    RECT 206.925 0.0 208.195 0.32 ;
    RECT 205.295 0.0 206.505 0.32 ;
    RECT 203.605 0.0 204.875 0.32 ;
    RECT 201.975 0.0 203.185 0.32 ;
    RECT 200.92 0.0 201.555 0.32 ;
    RECT 197.765 0.0 200.5 0.32 ;
    RECT 194.37 0.0 197.345 0.32 ;
    RECT 191.935 0.0 193.665 0.32 ;
    RECT 190.97 0.0 191.12 0.32 ;
    RECT 189.89 0.0 190.27 0.32 ;
    RECT 187.535 0.0 189.47 0.32 ;
    RECT 185.93 0.0 187.115 0.32 ;
    RECT 182.11 0.0 185.09 0.32 ;
    RECT 179.82 0.0 181.41 0.32 ;
    RECT 178.845 0.0 179.4 0.32 ;
    RECT 178.03 0.0 178.425 0.32 ;
    RECT 174.755 0.0 177.61 0.32 ;
    RECT 174.11 0.0 174.335 0.32 ;
    RECT 173.065 0.0 173.69 0.32 ;
    RECT 171.435 0.0 172.645 0.32 ;
    RECT 169.745 0.0 171.015 0.32 ;
    RECT 168.115 0.0 169.325 0.32 ;
    RECT 166.425 0.0 167.695 0.32 ;
    RECT 164.795 0.0 166.005 0.32 ;
    RECT 163.105 0.0 164.375 0.32 ;
    RECT 161.475 0.0 162.685 0.32 ;
    RECT 159.785 0.0 161.055 0.32 ;
    RECT 158.155 0.0 159.365 0.32 ;
    RECT 156.465 0.0 157.735 0.32 ;
    RECT 154.835 0.0 156.045 0.32 ;
    RECT 153.145 0.0 154.415 0.32 ;
    RECT 151.515 0.0 152.725 0.32 ;
    RECT 149.825 0.0 151.095 0.32 ;
    RECT 148.195 0.0 149.405 0.32 ;
    RECT 146.505 0.0 147.775 0.32 ;
    RECT 144.875 0.0 146.085 0.32 ;
    RECT 143.185 0.0 144.455 0.32 ;
    RECT 141.555 0.0 142.765 0.32 ;
    RECT 139.865 0.0 141.135 0.32 ;
    RECT 138.235 0.0 139.445 0.32 ;
    RECT 136.545 0.0 137.815 0.32 ;
    RECT 134.915 0.0 136.125 0.32 ;
    RECT 133.225 0.0 134.495 0.32 ;
    RECT 131.595 0.0 132.805 0.32 ;
    RECT 129.905 0.0 131.175 0.32 ;
    RECT 128.275 0.0 129.485 0.32 ;
    RECT 126.585 0.0 127.855 0.32 ;
    RECT 124.955 0.0 126.165 0.32 ;
    RECT 123.265 0.0 124.535 0.32 ;
    RECT 121.635 0.0 122.845 0.32 ;
    RECT 119.945 0.0 121.215 0.32 ;
    RECT 118.315 0.0 119.525 0.32 ;
    RECT 116.625 0.0 117.895 0.32 ;
    RECT 114.995 0.0 116.205 0.32 ;
    RECT 113.305 0.0 114.575 0.32 ;
    RECT 111.675 0.0 112.885 0.32 ;
    RECT 109.985 0.0 111.255 0.32 ;
    RECT 108.355 0.0 109.565 0.32 ;
    RECT 106.665 0.0 107.935 0.32 ;
    RECT 105.035 0.0 106.245 0.32 ;
    RECT 103.345 0.0 104.615 0.32 ;
    RECT 101.715 0.0 102.925 0.32 ;
    RECT 100.025 0.0 101.295 0.32 ;
    RECT 98.395 0.0 99.605 0.32 ;
    RECT 96.705 0.0 97.975 0.32 ;
    RECT 95.075 0.0 96.285 0.32 ;
    RECT 93.385 0.0 94.655 0.32 ;
    RECT 91.755 0.0 92.965 0.32 ;
    RECT 90.065 0.0 91.335 0.32 ;
    RECT 88.435 0.0 89.645 0.32 ;
    RECT 86.745 0.0 88.015 0.32 ;
    RECT 85.115 0.0 86.325 0.32 ;
    RECT 83.425 0.0 84.695 0.32 ;
    RECT 81.795 0.0 83.005 0.32 ;
    RECT 80.105 0.0 81.375 0.32 ;
    RECT 78.475 0.0 79.685 0.32 ;
    RECT 76.785 0.0 78.055 0.32 ;
    RECT 75.155 0.0 76.365 0.32 ;
    RECT 73.465 0.0 74.735 0.32 ;
    RECT 71.835 0.0 73.045 0.32 ;
    RECT 70.145 0.0 71.415 0.32 ;
    RECT 68.515 0.0 69.725 0.32 ;
    RECT 66.825 0.0 68.095 0.32 ;
    RECT 65.195 0.0 66.405 0.32 ;
    RECT 63.505 0.0 64.775 0.32 ;
    RECT 61.875 0.0 63.085 0.32 ;
    RECT 60.185 0.0 61.455 0.32 ;
    RECT 58.555 0.0 59.765 0.32 ;
    RECT 56.865 0.0 58.135 0.32 ;
    RECT 55.235 0.0 56.445 0.32 ;
    RECT 53.545 0.0 54.815 0.32 ;
    RECT 51.915 0.0 53.125 0.32 ;
    RECT 50.225 0.0 51.495 0.32 ;
    RECT 48.595 0.0 49.805 0.32 ;
    RECT 46.905 0.0 48.175 0.32 ;
    RECT 45.275 0.0 46.485 0.32 ;
    RECT 43.585 0.0 44.855 0.32 ;
    RECT 41.955 0.0 43.165 0.32 ;
    RECT 40.265 0.0 41.535 0.32 ;
    RECT 38.635 0.0 39.845 0.32 ;
    RECT 36.945 0.0 38.215 0.32 ;
    RECT 35.315 0.0 36.525 0.32 ;
    RECT 33.625 0.0 34.895 0.32 ;
    RECT 31.995 0.0 33.205 0.32 ;
    RECT 30.305 0.0 31.575 0.32 ;
    RECT 28.675 0.0 29.885 0.32 ;
    RECT 26.985 0.0 28.255 0.32 ;
    RECT 25.355 0.0 26.565 0.32 ;
    RECT 23.665 0.0 24.935 0.32 ;
    RECT 22.035 0.0 23.245 0.32 ;
    RECT 20.345 0.0 21.615 0.32 ;
    RECT 18.715 0.0 19.925 0.32 ;
    RECT 17.025 0.0 18.295 0.32 ;
    RECT 15.395 0.0 16.605 0.32 ;
    RECT 13.705 0.0 14.975 0.32 ;
    RECT 12.075 0.0 13.285 0.32 ;
    RECT 10.385 0.0 11.655 0.32 ;
    RECT 8.755 0.0 9.965 0.32 ;
    RECT 7.065 0.0 8.335 0.32 ;
    RECT 5.435 0.0 6.645 0.32 ;
    RECT 3.745 0.0 5.015 0.32 ;
    RECT 2.115 0.0 3.325 0.32 ;
    RECT 0.0 0.0 1.695 0.32 ;
    RECT 0.0 0.32 374.62 61.255 ;
    LAYER V2 ;
    RECT 0.0 0.0 374.62 61.255 ;
    LAYER M3 DESIGNRULEWIDTH 0.07 ;
    RECT 372.925 0.0 374.62 0.32 ;
    RECT 371.295 0.0 372.505 0.32 ;
    RECT 369.605 0.0 370.875 0.32 ;
    RECT 367.975 0.0 369.185 0.32 ;
    RECT 366.285 0.0 367.555 0.32 ;
    RECT 364.655 0.0 365.865 0.32 ;
    RECT 362.965 0.0 364.235 0.32 ;
    RECT 361.335 0.0 362.545 0.32 ;
    RECT 359.645 0.0 360.915 0.32 ;
    RECT 358.015 0.0 359.225 0.32 ;
    RECT 356.325 0.0 357.595 0.32 ;
    RECT 354.695 0.0 355.905 0.32 ;
    RECT 353.005 0.0 354.275 0.32 ;
    RECT 351.375 0.0 352.585 0.32 ;
    RECT 349.685 0.0 350.955 0.32 ;
    RECT 348.055 0.0 349.265 0.32 ;
    RECT 346.365 0.0 347.635 0.32 ;
    RECT 344.735 0.0 345.945 0.32 ;
    RECT 343.045 0.0 344.315 0.32 ;
    RECT 341.415 0.0 342.625 0.32 ;
    RECT 339.725 0.0 340.995 0.32 ;
    RECT 338.095 0.0 339.305 0.32 ;
    RECT 336.405 0.0 337.675 0.32 ;
    RECT 334.775 0.0 335.985 0.32 ;
    RECT 333.085 0.0 334.355 0.32 ;
    RECT 331.455 0.0 332.665 0.32 ;
    RECT 329.765 0.0 331.035 0.32 ;
    RECT 328.135 0.0 329.345 0.32 ;
    RECT 326.445 0.0 327.715 0.32 ;
    RECT 324.815 0.0 326.025 0.32 ;
    RECT 323.125 0.0 324.395 0.32 ;
    RECT 321.495 0.0 322.705 0.32 ;
    RECT 319.805 0.0 321.075 0.32 ;
    RECT 318.175 0.0 319.385 0.32 ;
    RECT 316.485 0.0 317.755 0.32 ;
    RECT 314.855 0.0 316.065 0.32 ;
    RECT 313.165 0.0 314.435 0.32 ;
    RECT 311.535 0.0 312.745 0.32 ;
    RECT 309.845 0.0 311.115 0.32 ;
    RECT 308.215 0.0 309.425 0.32 ;
    RECT 306.525 0.0 307.795 0.32 ;
    RECT 304.895 0.0 306.105 0.32 ;
    RECT 303.205 0.0 304.475 0.32 ;
    RECT 301.575 0.0 302.785 0.32 ;
    RECT 299.885 0.0 301.155 0.32 ;
    RECT 298.255 0.0 299.465 0.32 ;
    RECT 296.565 0.0 297.835 0.32 ;
    RECT 294.935 0.0 296.145 0.32 ;
    RECT 293.245 0.0 294.515 0.32 ;
    RECT 291.615 0.0 292.825 0.32 ;
    RECT 289.925 0.0 291.195 0.32 ;
    RECT 288.295 0.0 289.505 0.32 ;
    RECT 286.605 0.0 287.875 0.32 ;
    RECT 284.975 0.0 286.185 0.32 ;
    RECT 283.285 0.0 284.555 0.32 ;
    RECT 281.655 0.0 282.865 0.32 ;
    RECT 279.965 0.0 281.235 0.32 ;
    RECT 278.335 0.0 279.545 0.32 ;
    RECT 276.645 0.0 277.915 0.32 ;
    RECT 275.015 0.0 276.225 0.32 ;
    RECT 273.325 0.0 274.595 0.32 ;
    RECT 271.695 0.0 272.905 0.32 ;
    RECT 270.005 0.0 271.275 0.32 ;
    RECT 268.375 0.0 269.585 0.32 ;
    RECT 266.685 0.0 267.955 0.32 ;
    RECT 265.055 0.0 266.265 0.32 ;
    RECT 263.365 0.0 264.635 0.32 ;
    RECT 261.735 0.0 262.945 0.32 ;
    RECT 260.045 0.0 261.315 0.32 ;
    RECT 258.415 0.0 259.625 0.32 ;
    RECT 256.725 0.0 257.995 0.32 ;
    RECT 255.095 0.0 256.305 0.32 ;
    RECT 253.405 0.0 254.675 0.32 ;
    RECT 251.775 0.0 252.985 0.32 ;
    RECT 250.085 0.0 251.355 0.32 ;
    RECT 248.455 0.0 249.665 0.32 ;
    RECT 246.765 0.0 248.035 0.32 ;
    RECT 245.135 0.0 246.345 0.32 ;
    RECT 243.445 0.0 244.715 0.32 ;
    RECT 241.815 0.0 243.025 0.32 ;
    RECT 240.125 0.0 241.395 0.32 ;
    RECT 238.495 0.0 239.705 0.32 ;
    RECT 236.805 0.0 238.075 0.32 ;
    RECT 235.175 0.0 236.385 0.32 ;
    RECT 233.485 0.0 234.755 0.32 ;
    RECT 231.855 0.0 233.065 0.32 ;
    RECT 230.165 0.0 231.435 0.32 ;
    RECT 228.535 0.0 229.745 0.32 ;
    RECT 226.845 0.0 228.115 0.32 ;
    RECT 225.215 0.0 226.425 0.32 ;
    RECT 223.525 0.0 224.795 0.32 ;
    RECT 221.895 0.0 223.105 0.32 ;
    RECT 220.205 0.0 221.475 0.32 ;
    RECT 218.575 0.0 219.785 0.32 ;
    RECT 216.885 0.0 218.155 0.32 ;
    RECT 215.255 0.0 216.465 0.32 ;
    RECT 213.565 0.0 214.835 0.32 ;
    RECT 211.935 0.0 213.145 0.32 ;
    RECT 210.245 0.0 211.515 0.32 ;
    RECT 208.615 0.0 209.825 0.32 ;
    RECT 206.925 0.0 208.195 0.32 ;
    RECT 205.295 0.0 206.505 0.32 ;
    RECT 203.605 0.0 204.875 0.32 ;
    RECT 201.975 0.0 203.185 0.32 ;
    RECT 200.92 0.0 201.555 0.32 ;
    RECT 197.765 0.0 200.5 0.32 ;
    RECT 194.37 0.0 197.345 0.32 ;
    RECT 191.935 0.0 193.665 0.32 ;
    RECT 190.97 0.0 191.12 0.32 ;
    RECT 189.89 0.0 190.27 0.32 ;
    RECT 187.535 0.0 189.47 0.32 ;
    RECT 185.93 0.0 187.115 0.32 ;
    RECT 182.11 0.0 185.09 0.32 ;
    RECT 179.82 0.0 181.41 0.32 ;
    RECT 178.845 0.0 179.4 0.32 ;
    RECT 178.03 0.0 178.425 0.32 ;
    RECT 174.755 0.0 177.61 0.32 ;
    RECT 174.11 0.0 174.335 0.32 ;
    RECT 173.065 0.0 173.69 0.32 ;
    RECT 171.435 0.0 172.645 0.32 ;
    RECT 169.745 0.0 171.015 0.32 ;
    RECT 168.115 0.0 169.325 0.32 ;
    RECT 166.425 0.0 167.695 0.32 ;
    RECT 164.795 0.0 166.005 0.32 ;
    RECT 163.105 0.0 164.375 0.32 ;
    RECT 161.475 0.0 162.685 0.32 ;
    RECT 159.785 0.0 161.055 0.32 ;
    RECT 158.155 0.0 159.365 0.32 ;
    RECT 156.465 0.0 157.735 0.32 ;
    RECT 154.835 0.0 156.045 0.32 ;
    RECT 153.145 0.0 154.415 0.32 ;
    RECT 151.515 0.0 152.725 0.32 ;
    RECT 149.825 0.0 151.095 0.32 ;
    RECT 148.195 0.0 149.405 0.32 ;
    RECT 146.505 0.0 147.775 0.32 ;
    RECT 144.875 0.0 146.085 0.32 ;
    RECT 143.185 0.0 144.455 0.32 ;
    RECT 141.555 0.0 142.765 0.32 ;
    RECT 139.865 0.0 141.135 0.32 ;
    RECT 138.235 0.0 139.445 0.32 ;
    RECT 136.545 0.0 137.815 0.32 ;
    RECT 134.915 0.0 136.125 0.32 ;
    RECT 133.225 0.0 134.495 0.32 ;
    RECT 131.595 0.0 132.805 0.32 ;
    RECT 129.905 0.0 131.175 0.32 ;
    RECT 128.275 0.0 129.485 0.32 ;
    RECT 126.585 0.0 127.855 0.32 ;
    RECT 124.955 0.0 126.165 0.32 ;
    RECT 123.265 0.0 124.535 0.32 ;
    RECT 121.635 0.0 122.845 0.32 ;
    RECT 119.945 0.0 121.215 0.32 ;
    RECT 118.315 0.0 119.525 0.32 ;
    RECT 116.625 0.0 117.895 0.32 ;
    RECT 114.995 0.0 116.205 0.32 ;
    RECT 113.305 0.0 114.575 0.32 ;
    RECT 111.675 0.0 112.885 0.32 ;
    RECT 109.985 0.0 111.255 0.32 ;
    RECT 108.355 0.0 109.565 0.32 ;
    RECT 106.665 0.0 107.935 0.32 ;
    RECT 105.035 0.0 106.245 0.32 ;
    RECT 103.345 0.0 104.615 0.32 ;
    RECT 101.715 0.0 102.925 0.32 ;
    RECT 100.025 0.0 101.295 0.32 ;
    RECT 98.395 0.0 99.605 0.32 ;
    RECT 96.705 0.0 97.975 0.32 ;
    RECT 95.075 0.0 96.285 0.32 ;
    RECT 93.385 0.0 94.655 0.32 ;
    RECT 91.755 0.0 92.965 0.32 ;
    RECT 90.065 0.0 91.335 0.32 ;
    RECT 88.435 0.0 89.645 0.32 ;
    RECT 86.745 0.0 88.015 0.32 ;
    RECT 85.115 0.0 86.325 0.32 ;
    RECT 83.425 0.0 84.695 0.32 ;
    RECT 81.795 0.0 83.005 0.32 ;
    RECT 80.105 0.0 81.375 0.32 ;
    RECT 78.475 0.0 79.685 0.32 ;
    RECT 76.785 0.0 78.055 0.32 ;
    RECT 75.155 0.0 76.365 0.32 ;
    RECT 73.465 0.0 74.735 0.32 ;
    RECT 71.835 0.0 73.045 0.32 ;
    RECT 70.145 0.0 71.415 0.32 ;
    RECT 68.515 0.0 69.725 0.32 ;
    RECT 66.825 0.0 68.095 0.32 ;
    RECT 65.195 0.0 66.405 0.32 ;
    RECT 63.505 0.0 64.775 0.32 ;
    RECT 61.875 0.0 63.085 0.32 ;
    RECT 60.185 0.0 61.455 0.32 ;
    RECT 58.555 0.0 59.765 0.32 ;
    RECT 56.865 0.0 58.135 0.32 ;
    RECT 55.235 0.0 56.445 0.32 ;
    RECT 53.545 0.0 54.815 0.32 ;
    RECT 51.915 0.0 53.125 0.32 ;
    RECT 50.225 0.0 51.495 0.32 ;
    RECT 48.595 0.0 49.805 0.32 ;
    RECT 46.905 0.0 48.175 0.32 ;
    RECT 45.275 0.0 46.485 0.32 ;
    RECT 43.585 0.0 44.855 0.32 ;
    RECT 41.955 0.0 43.165 0.32 ;
    RECT 40.265 0.0 41.535 0.32 ;
    RECT 38.635 0.0 39.845 0.32 ;
    RECT 36.945 0.0 38.215 0.32 ;
    RECT 35.315 0.0 36.525 0.32 ;
    RECT 33.625 0.0 34.895 0.32 ;
    RECT 31.995 0.0 33.205 0.32 ;
    RECT 30.305 0.0 31.575 0.32 ;
    RECT 28.675 0.0 29.885 0.32 ;
    RECT 26.985 0.0 28.255 0.32 ;
    RECT 25.355 0.0 26.565 0.32 ;
    RECT 23.665 0.0 24.935 0.32 ;
    RECT 22.035 0.0 23.245 0.32 ;
    RECT 20.345 0.0 21.615 0.32 ;
    RECT 18.715 0.0 19.925 0.32 ;
    RECT 17.025 0.0 18.295 0.32 ;
    RECT 15.395 0.0 16.605 0.32 ;
    RECT 13.705 0.0 14.975 0.32 ;
    RECT 12.075 0.0 13.285 0.32 ;
    RECT 10.385 0.0 11.655 0.32 ;
    RECT 8.755 0.0 9.965 0.32 ;
    RECT 7.065 0.0 8.335 0.32 ;
    RECT 5.435 0.0 6.645 0.32 ;
    RECT 3.745 0.0 5.015 0.32 ;
    RECT 2.115 0.0 3.325 0.32 ;
    RECT 0.0 0.0 1.695 0.32 ;
    RECT 0.0 0.32 374.62 61.255 ;
    LAYER V3 ;
    RECT 0.0 0.0 374.62 61.255 ;
    LAYER V3 ;
    RECT 59.31 0.415 59.57 0.485 ;
    RECT 58.39 0.432 58.6 0.502 ;
    RECT 55.99 0.415 56.25 0.485 ;
    RECT 55.07 0.432 55.28 0.502 ;
    RECT 52.67 0.415 52.93 0.485 ;
    RECT 51.75 0.432 51.96 0.502 ;
    RECT 49.35 0.415 49.61 0.485 ;
    RECT 48.43 0.432 48.64 0.502 ;
    RECT 331.65 0.415 331.91 0.485 ;
    RECT 332.62 0.432 332.83 0.502 ;
    RECT 46.03 0.415 46.29 0.485 ;
    RECT 45.11 0.432 45.32 0.502 ;
    RECT 328.33 0.415 328.59 0.485 ;
    RECT 329.3 0.432 329.51 0.502 ;
    RECT 42.71 0.415 42.97 0.485 ;
    RECT 41.79 0.432 42.0 0.502 ;
    RECT 325.01 0.415 325.27 0.485 ;
    RECT 325.98 0.432 326.19 0.502 ;
    RECT 39.39 0.415 39.65 0.485 ;
    RECT 38.47 0.432 38.68 0.502 ;
    RECT 321.69 0.415 321.95 0.485 ;
    RECT 322.66 0.432 322.87 0.502 ;
    RECT 36.07 0.415 36.33 0.485 ;
    RECT 35.15 0.432 35.36 0.502 ;
    RECT 318.37 0.415 318.63 0.485 ;
    RECT 319.34 0.432 319.55 0.502 ;
    RECT 315.05 0.415 315.31 0.485 ;
    RECT 316.02 0.432 316.23 0.502 ;
    RECT 311.73 0.415 311.99 0.485 ;
    RECT 312.7 0.432 312.91 0.502 ;
    RECT 308.41 0.415 308.67 0.485 ;
    RECT 309.38 0.432 309.59 0.502 ;
    RECT 305.09 0.415 305.35 0.485 ;
    RECT 306.06 0.432 306.27 0.502 ;
    RECT 175.735 0.435 175.975 0.505 ;
    RECT 176.35 0.18 177.1 0.25 ;
    RECT 179.575 0.06 179.645 0.27 ;
    RECT 180.79 0.435 181.04 0.505 ;
    RECT 183.055 0.435 183.32 0.505 ;
    RECT 184.1 0.435 184.35 0.505 ;
    RECT 191.0 0.435 191.25 0.505 ;
    RECT 193.565 0.435 193.835 0.505 ;
    RECT 198.4 0.605 198.47 0.675 ;
    RECT 198.605 0.435 198.815 0.505 ;
    RECT 301.77 0.415 302.03 0.485 ;
    RECT 302.74 0.432 302.95 0.502 ;
    RECT 232.05 0.415 232.31 0.485 ;
    RECT 233.02 0.432 233.23 0.502 ;
    RECT 228.73 0.415 228.99 0.485 ;
    RECT 229.7 0.432 229.91 0.502 ;
    RECT 298.45 0.415 298.71 0.485 ;
    RECT 299.42 0.432 299.63 0.502 ;
    RECT 225.41 0.415 225.67 0.485 ;
    RECT 226.38 0.432 226.59 0.502 ;
    RECT 295.13 0.415 295.39 0.485 ;
    RECT 296.1 0.432 296.31 0.502 ;
    RECT 222.09 0.415 222.35 0.485 ;
    RECT 223.06 0.432 223.27 0.502 ;
    RECT 291.81 0.415 292.07 0.485 ;
    RECT 292.78 0.432 292.99 0.502 ;
    RECT 218.77 0.415 219.03 0.485 ;
    RECT 219.74 0.432 219.95 0.502 ;
    RECT 288.49 0.415 288.75 0.485 ;
    RECT 289.46 0.432 289.67 0.502 ;
    RECT 215.45 0.415 215.71 0.485 ;
    RECT 216.42 0.432 216.63 0.502 ;
    RECT 285.17 0.415 285.43 0.485 ;
    RECT 286.14 0.432 286.35 0.502 ;
    RECT 212.13 0.415 212.39 0.485 ;
    RECT 213.1 0.432 213.31 0.502 ;
    RECT 281.85 0.415 282.11 0.485 ;
    RECT 282.82 0.432 283.03 0.502 ;
    RECT 208.81 0.415 209.07 0.485 ;
    RECT 209.78 0.432 209.99 0.502 ;
    RECT 278.53 0.415 278.79 0.485 ;
    RECT 279.5 0.432 279.71 0.502 ;
    RECT 172.19 0.415 172.45 0.485 ;
    RECT 171.27 0.432 171.48 0.502 ;
    RECT 205.49 0.415 205.75 0.485 ;
    RECT 206.46 0.432 206.67 0.502 ;
    RECT 275.21 0.415 275.47 0.485 ;
    RECT 276.18 0.432 276.39 0.502 ;
    RECT 168.87 0.415 169.13 0.485 ;
    RECT 167.95 0.432 168.16 0.502 ;
    RECT 202.17 0.415 202.43 0.485 ;
    RECT 203.14 0.432 203.35 0.502 ;
    RECT 271.89 0.415 272.15 0.485 ;
    RECT 272.86 0.432 273.07 0.502 ;
    RECT 268.57 0.415 268.83 0.485 ;
    RECT 269.54 0.432 269.75 0.502 ;
    RECT 165.55 0.415 165.81 0.485 ;
    RECT 164.63 0.432 164.84 0.502 ;
    RECT 162.23 0.415 162.49 0.485 ;
    RECT 161.31 0.432 161.52 0.502 ;
    RECT 265.25 0.415 265.51 0.485 ;
    RECT 266.22 0.432 266.43 0.502 ;
    RECT 158.91 0.415 159.17 0.485 ;
    RECT 157.99 0.432 158.2 0.502 ;
    RECT 261.93 0.415 262.19 0.485 ;
    RECT 262.9 0.432 263.11 0.502 ;
    RECT 155.59 0.415 155.85 0.485 ;
    RECT 154.67 0.432 154.88 0.502 ;
    RECT 258.61 0.415 258.87 0.485 ;
    RECT 259.58 0.432 259.79 0.502 ;
    RECT 152.27 0.415 152.53 0.485 ;
    RECT 151.35 0.432 151.56 0.502 ;
    RECT 255.29 0.415 255.55 0.485 ;
    RECT 256.26 0.432 256.47 0.502 ;
    RECT 148.95 0.415 149.21 0.485 ;
    RECT 148.03 0.432 148.24 0.502 ;
    RECT 251.97 0.415 252.23 0.485 ;
    RECT 252.94 0.432 253.15 0.502 ;
    RECT 145.63 0.415 145.89 0.485 ;
    RECT 144.71 0.432 144.92 0.502 ;
    RECT 248.65 0.415 248.91 0.485 ;
    RECT 249.62 0.432 249.83 0.502 ;
    RECT 142.31 0.415 142.57 0.485 ;
    RECT 141.39 0.432 141.6 0.502 ;
    RECT 245.33 0.415 245.59 0.485 ;
    RECT 246.3 0.432 246.51 0.502 ;
    RECT 138.99 0.415 139.25 0.485 ;
    RECT 138.07 0.432 138.28 0.502 ;
    RECT 242.01 0.415 242.27 0.485 ;
    RECT 242.98 0.432 243.19 0.502 ;
    RECT 135.67 0.415 135.93 0.485 ;
    RECT 134.75 0.432 134.96 0.502 ;
    RECT 238.69 0.415 238.95 0.485 ;
    RECT 239.66 0.432 239.87 0.502 ;
    RECT 32.75 0.415 33.01 0.485 ;
    RECT 31.83 0.432 32.04 0.502 ;
    RECT 235.37 0.415 235.63 0.485 ;
    RECT 236.34 0.432 236.55 0.502 ;
    RECT 29.43 0.415 29.69 0.485 ;
    RECT 28.51 0.432 28.72 0.502 ;
    RECT 26.11 0.415 26.37 0.485 ;
    RECT 25.19 0.432 25.4 0.502 ;
    RECT 22.79 0.415 23.05 0.485 ;
    RECT 21.87 0.432 22.08 0.502 ;
    RECT 19.47 0.415 19.73 0.485 ;
    RECT 18.55 0.432 18.76 0.502 ;
    RECT 16.15 0.415 16.41 0.485 ;
    RECT 15.23 0.432 15.44 0.502 ;
    RECT 12.83 0.415 13.09 0.485 ;
    RECT 11.91 0.432 12.12 0.502 ;
    RECT 9.51 0.415 9.77 0.485 ;
    RECT 8.59 0.432 8.8 0.502 ;
    RECT 6.19 0.415 6.45 0.485 ;
    RECT 5.27 0.432 5.48 0.502 ;
    RECT 2.87 0.415 3.13 0.485 ;
    RECT 1.95 0.432 2.16 0.502 ;
    RECT 132.35 0.415 132.61 0.485 ;
    RECT 131.43 0.432 131.64 0.502 ;
    RECT 129.03 0.415 129.29 0.485 ;
    RECT 128.11 0.432 128.32 0.502 ;
    RECT 125.71 0.415 125.97 0.485 ;
    RECT 124.79 0.432 125.0 0.502 ;
    RECT 122.39 0.415 122.65 0.485 ;
    RECT 121.47 0.432 121.68 0.502 ;
    RECT 119.07 0.415 119.33 0.485 ;
    RECT 118.15 0.432 118.36 0.502 ;
    RECT 115.75 0.415 116.01 0.485 ;
    RECT 114.83 0.432 115.04 0.502 ;
    RECT 112.43 0.415 112.69 0.485 ;
    RECT 111.51 0.432 111.72 0.502 ;
    RECT 109.11 0.415 109.37 0.485 ;
    RECT 108.19 0.432 108.4 0.502 ;
    RECT 105.79 0.415 106.05 0.485 ;
    RECT 104.87 0.432 105.08 0.502 ;
    RECT 102.47 0.415 102.73 0.485 ;
    RECT 101.55 0.432 101.76 0.502 ;
    RECT 371.49 0.415 371.75 0.485 ;
    RECT 372.46 0.432 372.67 0.502 ;
    RECT 368.17 0.415 368.43 0.485 ;
    RECT 369.14 0.432 369.35 0.502 ;
    RECT 99.15 0.415 99.41 0.485 ;
    RECT 98.23 0.432 98.44 0.502 ;
    RECT 95.83 0.415 96.09 0.485 ;
    RECT 94.91 0.432 95.12 0.502 ;
    RECT 92.51 0.415 92.77 0.485 ;
    RECT 91.59 0.432 91.8 0.502 ;
    RECT 89.19 0.415 89.45 0.485 ;
    RECT 88.27 0.432 88.48 0.502 ;
    RECT 85.87 0.415 86.13 0.485 ;
    RECT 84.95 0.432 85.16 0.502 ;
    RECT 364.85 0.415 365.11 0.485 ;
    RECT 365.82 0.432 366.03 0.502 ;
    RECT 82.55 0.415 82.81 0.485 ;
    RECT 81.63 0.432 81.84 0.502 ;
    RECT 361.53 0.415 361.79 0.485 ;
    RECT 362.5 0.432 362.71 0.502 ;
    RECT 79.23 0.415 79.49 0.485 ;
    RECT 78.31 0.432 78.52 0.502 ;
    RECT 358.21 0.415 358.47 0.485 ;
    RECT 359.18 0.432 359.39 0.502 ;
    RECT 75.91 0.415 76.17 0.485 ;
    RECT 74.99 0.432 75.2 0.502 ;
    RECT 354.89 0.415 355.15 0.485 ;
    RECT 355.86 0.432 356.07 0.502 ;
    RECT 72.59 0.415 72.85 0.485 ;
    RECT 71.67 0.432 71.88 0.502 ;
    RECT 351.57 0.415 351.83 0.485 ;
    RECT 352.54 0.432 352.75 0.502 ;
    RECT 69.27 0.415 69.53 0.485 ;
    RECT 68.35 0.432 68.56 0.502 ;
    RECT 348.25 0.415 348.51 0.485 ;
    RECT 349.22 0.432 349.43 0.502 ;
    RECT 344.93 0.415 345.19 0.485 ;
    RECT 345.9 0.432 346.11 0.502 ;
    RECT 341.61 0.415 341.87 0.485 ;
    RECT 342.58 0.432 342.79 0.502 ;
    RECT 338.29 0.415 338.55 0.485 ;
    RECT 339.26 0.432 339.47 0.502 ;
    RECT 334.97 0.415 335.23 0.485 ;
    RECT 335.94 0.432 336.15 0.502 ;
    RECT 65.95 0.415 66.21 0.485 ;
    RECT 65.03 0.432 65.24 0.502 ;
    RECT 62.63 0.415 62.89 0.485 ;
    RECT 61.71 0.432 61.92 0.502 ;
    RECT 303.2 33.165 303.41 33.235 ;
    RECT 303.2 33.525 303.41 33.595 ;
    RECT 303.2 33.885 303.41 33.955 ;
    RECT 302.74 33.165 302.95 33.235 ;
    RECT 302.74 33.525 302.95 33.595 ;
    RECT 302.74 33.885 302.95 33.955 ;
    RECT 372.92 33.165 373.13 33.235 ;
    RECT 372.92 33.525 373.13 33.595 ;
    RECT 372.92 33.885 373.13 33.955 ;
    RECT 372.46 33.165 372.67 33.235 ;
    RECT 372.46 33.525 372.67 33.595 ;
    RECT 372.46 33.885 372.67 33.955 ;
    RECT 369.6 33.165 369.81 33.235 ;
    RECT 369.6 33.525 369.81 33.595 ;
    RECT 369.6 33.885 369.81 33.955 ;
    RECT 369.14 33.165 369.35 33.235 ;
    RECT 369.14 33.525 369.35 33.595 ;
    RECT 369.14 33.885 369.35 33.955 ;
    RECT 200.605 33.525 200.675 33.595 ;
    RECT 299.88 33.165 300.09 33.235 ;
    RECT 299.88 33.525 300.09 33.595 ;
    RECT 299.88 33.885 300.09 33.955 ;
    RECT 299.42 33.165 299.63 33.235 ;
    RECT 299.42 33.525 299.63 33.595 ;
    RECT 299.42 33.885 299.63 33.955 ;
    RECT 296.56 33.165 296.77 33.235 ;
    RECT 296.56 33.525 296.77 33.595 ;
    RECT 296.56 33.885 296.77 33.955 ;
    RECT 296.1 33.165 296.31 33.235 ;
    RECT 296.1 33.525 296.31 33.595 ;
    RECT 296.1 33.885 296.31 33.955 ;
    RECT 293.24 33.165 293.45 33.235 ;
    RECT 293.24 33.525 293.45 33.595 ;
    RECT 293.24 33.885 293.45 33.955 ;
    RECT 292.78 33.165 292.99 33.235 ;
    RECT 292.78 33.525 292.99 33.595 ;
    RECT 292.78 33.885 292.99 33.955 ;
    RECT 289.92 33.165 290.13 33.235 ;
    RECT 289.92 33.525 290.13 33.595 ;
    RECT 289.92 33.885 290.13 33.955 ;
    RECT 289.46 33.165 289.67 33.235 ;
    RECT 289.46 33.525 289.67 33.595 ;
    RECT 289.46 33.885 289.67 33.955 ;
    RECT 286.6 33.165 286.81 33.235 ;
    RECT 286.6 33.525 286.81 33.595 ;
    RECT 286.6 33.885 286.81 33.955 ;
    RECT 286.14 33.165 286.35 33.235 ;
    RECT 286.14 33.525 286.35 33.595 ;
    RECT 286.14 33.885 286.35 33.955 ;
    RECT 283.28 33.165 283.49 33.235 ;
    RECT 283.28 33.525 283.49 33.595 ;
    RECT 283.28 33.885 283.49 33.955 ;
    RECT 282.82 33.165 283.03 33.235 ;
    RECT 282.82 33.525 283.03 33.595 ;
    RECT 282.82 33.885 283.03 33.955 ;
    RECT 279.96 33.165 280.17 33.235 ;
    RECT 279.96 33.525 280.17 33.595 ;
    RECT 279.96 33.885 280.17 33.955 ;
    RECT 279.5 33.165 279.71 33.235 ;
    RECT 279.5 33.525 279.71 33.595 ;
    RECT 279.5 33.885 279.71 33.955 ;
    RECT 276.64 33.165 276.85 33.235 ;
    RECT 276.64 33.525 276.85 33.595 ;
    RECT 276.64 33.885 276.85 33.955 ;
    RECT 276.18 33.165 276.39 33.235 ;
    RECT 276.18 33.525 276.39 33.595 ;
    RECT 276.18 33.885 276.39 33.955 ;
    RECT 273.32 33.165 273.53 33.235 ;
    RECT 273.32 33.525 273.53 33.595 ;
    RECT 273.32 33.885 273.53 33.955 ;
    RECT 272.86 33.165 273.07 33.235 ;
    RECT 272.86 33.525 273.07 33.595 ;
    RECT 272.86 33.885 273.07 33.955 ;
    RECT 270.0 33.165 270.21 33.235 ;
    RECT 270.0 33.525 270.21 33.595 ;
    RECT 270.0 33.885 270.21 33.955 ;
    RECT 269.54 33.165 269.75 33.235 ;
    RECT 269.54 33.525 269.75 33.595 ;
    RECT 269.54 33.885 269.75 33.955 ;
    RECT 233.48 33.165 233.69 33.235 ;
    RECT 233.48 33.525 233.69 33.595 ;
    RECT 233.48 33.885 233.69 33.955 ;
    RECT 233.02 33.165 233.23 33.235 ;
    RECT 233.02 33.525 233.23 33.595 ;
    RECT 233.02 33.885 233.23 33.955 ;
    RECT 230.16 33.165 230.37 33.235 ;
    RECT 230.16 33.525 230.37 33.595 ;
    RECT 230.16 33.885 230.37 33.955 ;
    RECT 229.7 33.165 229.91 33.235 ;
    RECT 229.7 33.525 229.91 33.595 ;
    RECT 229.7 33.885 229.91 33.955 ;
    RECT 366.28 33.165 366.49 33.235 ;
    RECT 366.28 33.525 366.49 33.595 ;
    RECT 366.28 33.885 366.49 33.955 ;
    RECT 365.82 33.165 366.03 33.235 ;
    RECT 365.82 33.525 366.03 33.595 ;
    RECT 365.82 33.885 366.03 33.955 ;
    RECT 226.84 33.165 227.05 33.235 ;
    RECT 226.84 33.525 227.05 33.595 ;
    RECT 226.84 33.885 227.05 33.955 ;
    RECT 226.38 33.165 226.59 33.235 ;
    RECT 226.38 33.525 226.59 33.595 ;
    RECT 226.38 33.885 226.59 33.955 ;
    RECT 362.96 33.165 363.17 33.235 ;
    RECT 362.96 33.525 363.17 33.595 ;
    RECT 362.96 33.885 363.17 33.955 ;
    RECT 362.5 33.165 362.71 33.235 ;
    RECT 362.5 33.525 362.71 33.595 ;
    RECT 362.5 33.885 362.71 33.955 ;
    RECT 223.52 33.165 223.73 33.235 ;
    RECT 223.52 33.525 223.73 33.595 ;
    RECT 223.52 33.885 223.73 33.955 ;
    RECT 223.06 33.165 223.27 33.235 ;
    RECT 223.06 33.525 223.27 33.595 ;
    RECT 223.06 33.885 223.27 33.955 ;
    RECT 359.64 33.165 359.85 33.235 ;
    RECT 359.64 33.525 359.85 33.595 ;
    RECT 359.64 33.885 359.85 33.955 ;
    RECT 359.18 33.165 359.39 33.235 ;
    RECT 359.18 33.525 359.39 33.595 ;
    RECT 359.18 33.885 359.39 33.955 ;
    RECT 220.2 33.165 220.41 33.235 ;
    RECT 220.2 33.525 220.41 33.595 ;
    RECT 220.2 33.885 220.41 33.955 ;
    RECT 219.74 33.165 219.95 33.235 ;
    RECT 219.74 33.525 219.95 33.595 ;
    RECT 219.74 33.885 219.95 33.955 ;
    RECT 356.32 33.165 356.53 33.235 ;
    RECT 356.32 33.525 356.53 33.595 ;
    RECT 356.32 33.885 356.53 33.955 ;
    RECT 355.86 33.165 356.07 33.235 ;
    RECT 355.86 33.525 356.07 33.595 ;
    RECT 355.86 33.885 356.07 33.955 ;
    RECT 353.0 33.165 353.21 33.235 ;
    RECT 353.0 33.525 353.21 33.595 ;
    RECT 353.0 33.885 353.21 33.955 ;
    RECT 352.54 33.165 352.75 33.235 ;
    RECT 352.54 33.525 352.75 33.595 ;
    RECT 352.54 33.885 352.75 33.955 ;
    RECT 216.88 33.165 217.09 33.235 ;
    RECT 216.88 33.525 217.09 33.595 ;
    RECT 216.88 33.885 217.09 33.955 ;
    RECT 216.42 33.165 216.63 33.235 ;
    RECT 216.42 33.525 216.63 33.595 ;
    RECT 216.42 33.885 216.63 33.955 ;
    RECT 349.68 33.165 349.89 33.235 ;
    RECT 349.68 33.525 349.89 33.595 ;
    RECT 349.68 33.885 349.89 33.955 ;
    RECT 349.22 33.165 349.43 33.235 ;
    RECT 349.22 33.525 349.43 33.595 ;
    RECT 349.22 33.885 349.43 33.955 ;
    RECT 213.56 33.165 213.77 33.235 ;
    RECT 213.56 33.525 213.77 33.595 ;
    RECT 213.56 33.885 213.77 33.955 ;
    RECT 213.1 33.165 213.31 33.235 ;
    RECT 213.1 33.525 213.31 33.595 ;
    RECT 213.1 33.885 213.31 33.955 ;
    RECT 346.36 33.165 346.57 33.235 ;
    RECT 346.36 33.525 346.57 33.595 ;
    RECT 346.36 33.885 346.57 33.955 ;
    RECT 345.9 33.165 346.11 33.235 ;
    RECT 345.9 33.525 346.11 33.595 ;
    RECT 345.9 33.885 346.11 33.955 ;
    RECT 210.24 33.165 210.45 33.235 ;
    RECT 210.24 33.525 210.45 33.595 ;
    RECT 210.24 33.885 210.45 33.955 ;
    RECT 209.78 33.165 209.99 33.235 ;
    RECT 209.78 33.525 209.99 33.595 ;
    RECT 209.78 33.885 209.99 33.955 ;
    RECT 343.04 33.165 343.25 33.235 ;
    RECT 343.04 33.525 343.25 33.595 ;
    RECT 343.04 33.885 343.25 33.955 ;
    RECT 342.58 33.165 342.79 33.235 ;
    RECT 342.58 33.525 342.79 33.595 ;
    RECT 342.58 33.885 342.79 33.955 ;
    RECT 206.92 33.165 207.13 33.235 ;
    RECT 206.92 33.525 207.13 33.595 ;
    RECT 206.92 33.885 207.13 33.955 ;
    RECT 206.46 33.165 206.67 33.235 ;
    RECT 206.46 33.525 206.67 33.595 ;
    RECT 206.46 33.885 206.67 33.955 ;
    RECT 339.72 33.165 339.93 33.235 ;
    RECT 339.72 33.525 339.93 33.595 ;
    RECT 339.72 33.885 339.93 33.955 ;
    RECT 339.26 33.165 339.47 33.235 ;
    RECT 339.26 33.525 339.47 33.595 ;
    RECT 339.26 33.885 339.47 33.955 ;
    RECT 203.6 33.165 203.81 33.235 ;
    RECT 203.6 33.525 203.81 33.595 ;
    RECT 203.6 33.885 203.81 33.955 ;
    RECT 203.14 33.165 203.35 33.235 ;
    RECT 203.14 33.525 203.35 33.595 ;
    RECT 203.14 33.885 203.35 33.955 ;
    RECT 336.4 33.165 336.61 33.235 ;
    RECT 336.4 33.525 336.61 33.595 ;
    RECT 336.4 33.885 336.61 33.955 ;
    RECT 335.94 33.165 336.15 33.235 ;
    RECT 335.94 33.525 336.15 33.595 ;
    RECT 335.94 33.885 336.15 33.955 ;
    RECT 266.68 33.165 266.89 33.235 ;
    RECT 266.68 33.525 266.89 33.595 ;
    RECT 266.68 33.885 266.89 33.955 ;
    RECT 266.22 33.165 266.43 33.235 ;
    RECT 266.22 33.525 266.43 33.595 ;
    RECT 266.22 33.885 266.43 33.955 ;
    RECT 263.36 33.165 263.57 33.235 ;
    RECT 263.36 33.525 263.57 33.595 ;
    RECT 263.36 33.885 263.57 33.955 ;
    RECT 262.9 33.165 263.11 33.235 ;
    RECT 262.9 33.525 263.11 33.595 ;
    RECT 262.9 33.885 263.11 33.955 ;
    RECT 260.04 33.165 260.25 33.235 ;
    RECT 260.04 33.525 260.25 33.595 ;
    RECT 260.04 33.885 260.25 33.955 ;
    RECT 259.58 33.165 259.79 33.235 ;
    RECT 259.58 33.525 259.79 33.595 ;
    RECT 259.58 33.885 259.79 33.955 ;
    RECT 256.72 33.165 256.93 33.235 ;
    RECT 256.72 33.525 256.93 33.595 ;
    RECT 256.72 33.885 256.93 33.955 ;
    RECT 256.26 33.165 256.47 33.235 ;
    RECT 256.26 33.525 256.47 33.595 ;
    RECT 256.26 33.885 256.47 33.955 ;
    RECT 253.4 33.165 253.61 33.235 ;
    RECT 253.4 33.525 253.61 33.595 ;
    RECT 253.4 33.885 253.61 33.955 ;
    RECT 252.94 33.165 253.15 33.235 ;
    RECT 252.94 33.525 253.15 33.595 ;
    RECT 252.94 33.885 253.15 33.955 ;
    RECT 250.08 33.165 250.29 33.235 ;
    RECT 250.08 33.525 250.29 33.595 ;
    RECT 250.08 33.885 250.29 33.955 ;
    RECT 249.62 33.165 249.83 33.235 ;
    RECT 249.62 33.525 249.83 33.595 ;
    RECT 249.62 33.885 249.83 33.955 ;
    RECT 246.76 33.165 246.97 33.235 ;
    RECT 246.76 33.525 246.97 33.595 ;
    RECT 246.76 33.885 246.97 33.955 ;
    RECT 246.3 33.165 246.51 33.235 ;
    RECT 246.3 33.525 246.51 33.595 ;
    RECT 246.3 33.885 246.51 33.955 ;
    RECT 243.44 33.165 243.65 33.235 ;
    RECT 243.44 33.525 243.65 33.595 ;
    RECT 243.44 33.885 243.65 33.955 ;
    RECT 242.98 33.165 243.19 33.235 ;
    RECT 242.98 33.525 243.19 33.595 ;
    RECT 242.98 33.885 243.19 33.955 ;
    RECT 240.12 33.165 240.33 33.235 ;
    RECT 240.12 33.525 240.33 33.595 ;
    RECT 240.12 33.885 240.33 33.955 ;
    RECT 239.66 33.165 239.87 33.235 ;
    RECT 239.66 33.525 239.87 33.595 ;
    RECT 239.66 33.885 239.87 33.955 ;
    RECT 236.8 33.165 237.01 33.235 ;
    RECT 236.8 33.525 237.01 33.595 ;
    RECT 236.8 33.885 237.01 33.955 ;
    RECT 236.34 33.165 236.55 33.235 ;
    RECT 236.34 33.525 236.55 33.595 ;
    RECT 236.34 33.885 236.55 33.955 ;
    RECT 374.15 33.525 374.22 33.595 ;
    RECT 333.08 33.165 333.29 33.235 ;
    RECT 333.08 33.525 333.29 33.595 ;
    RECT 333.08 33.885 333.29 33.955 ;
    RECT 332.62 33.165 332.83 33.235 ;
    RECT 332.62 33.525 332.83 33.595 ;
    RECT 332.62 33.885 332.83 33.955 ;
    RECT 329.76 33.165 329.97 33.235 ;
    RECT 329.76 33.525 329.97 33.595 ;
    RECT 329.76 33.885 329.97 33.955 ;
    RECT 329.3 33.165 329.51 33.235 ;
    RECT 329.3 33.525 329.51 33.595 ;
    RECT 329.3 33.885 329.51 33.955 ;
    RECT 326.44 33.165 326.65 33.235 ;
    RECT 326.44 33.525 326.65 33.595 ;
    RECT 326.44 33.885 326.65 33.955 ;
    RECT 325.98 33.165 326.19 33.235 ;
    RECT 325.98 33.525 326.19 33.595 ;
    RECT 325.98 33.885 326.19 33.955 ;
    RECT 323.12 33.165 323.33 33.235 ;
    RECT 323.12 33.525 323.33 33.595 ;
    RECT 323.12 33.885 323.33 33.955 ;
    RECT 322.66 33.165 322.87 33.235 ;
    RECT 322.66 33.525 322.87 33.595 ;
    RECT 322.66 33.885 322.87 33.955 ;
    RECT 319.8 33.165 320.01 33.235 ;
    RECT 319.8 33.525 320.01 33.595 ;
    RECT 319.8 33.885 320.01 33.955 ;
    RECT 319.34 33.165 319.55 33.235 ;
    RECT 319.34 33.525 319.55 33.595 ;
    RECT 319.34 33.885 319.55 33.955 ;
    RECT 316.48 33.165 316.69 33.235 ;
    RECT 316.48 33.525 316.69 33.595 ;
    RECT 316.48 33.885 316.69 33.955 ;
    RECT 316.02 33.165 316.23 33.235 ;
    RECT 316.02 33.525 316.23 33.595 ;
    RECT 316.02 33.885 316.23 33.955 ;
    RECT 313.16 33.165 313.37 33.235 ;
    RECT 313.16 33.525 313.37 33.595 ;
    RECT 313.16 33.885 313.37 33.955 ;
    RECT 312.7 33.165 312.91 33.235 ;
    RECT 312.7 33.525 312.91 33.595 ;
    RECT 312.7 33.885 312.91 33.955 ;
    RECT 309.84 33.165 310.05 33.235 ;
    RECT 309.84 33.525 310.05 33.595 ;
    RECT 309.84 33.885 310.05 33.955 ;
    RECT 309.38 33.165 309.59 33.235 ;
    RECT 309.38 33.525 309.59 33.595 ;
    RECT 309.38 33.885 309.59 33.955 ;
    RECT 306.52 33.165 306.73 33.235 ;
    RECT 306.52 33.525 306.73 33.595 ;
    RECT 306.52 33.885 306.73 33.955 ;
    RECT 306.06 33.165 306.27 33.235 ;
    RECT 306.06 33.525 306.27 33.595 ;
    RECT 306.06 33.885 306.27 33.955 ;
    RECT 303.2 18.045 303.41 18.115 ;
    RECT 303.2 18.405 303.41 18.475 ;
    RECT 303.2 18.765 303.41 18.835 ;
    RECT 302.74 18.045 302.95 18.115 ;
    RECT 302.74 18.405 302.95 18.475 ;
    RECT 302.74 18.765 302.95 18.835 ;
    RECT 372.92 18.045 373.13 18.115 ;
    RECT 372.92 18.405 373.13 18.475 ;
    RECT 372.92 18.765 373.13 18.835 ;
    RECT 372.46 18.045 372.67 18.115 ;
    RECT 372.46 18.405 372.67 18.475 ;
    RECT 372.46 18.765 372.67 18.835 ;
    RECT 369.6 18.045 369.81 18.115 ;
    RECT 369.6 18.405 369.81 18.475 ;
    RECT 369.6 18.765 369.81 18.835 ;
    RECT 369.14 18.045 369.35 18.115 ;
    RECT 369.14 18.405 369.35 18.475 ;
    RECT 369.14 18.765 369.35 18.835 ;
    RECT 200.605 18.405 200.675 18.475 ;
    RECT 299.88 18.045 300.09 18.115 ;
    RECT 299.88 18.405 300.09 18.475 ;
    RECT 299.88 18.765 300.09 18.835 ;
    RECT 299.42 18.045 299.63 18.115 ;
    RECT 299.42 18.405 299.63 18.475 ;
    RECT 299.42 18.765 299.63 18.835 ;
    RECT 296.56 18.045 296.77 18.115 ;
    RECT 296.56 18.405 296.77 18.475 ;
    RECT 296.56 18.765 296.77 18.835 ;
    RECT 296.1 18.045 296.31 18.115 ;
    RECT 296.1 18.405 296.31 18.475 ;
    RECT 296.1 18.765 296.31 18.835 ;
    RECT 293.24 18.045 293.45 18.115 ;
    RECT 293.24 18.405 293.45 18.475 ;
    RECT 293.24 18.765 293.45 18.835 ;
    RECT 292.78 18.045 292.99 18.115 ;
    RECT 292.78 18.405 292.99 18.475 ;
    RECT 292.78 18.765 292.99 18.835 ;
    RECT 289.92 18.045 290.13 18.115 ;
    RECT 289.92 18.405 290.13 18.475 ;
    RECT 289.92 18.765 290.13 18.835 ;
    RECT 289.46 18.045 289.67 18.115 ;
    RECT 289.46 18.405 289.67 18.475 ;
    RECT 289.46 18.765 289.67 18.835 ;
    RECT 286.6 18.045 286.81 18.115 ;
    RECT 286.6 18.405 286.81 18.475 ;
    RECT 286.6 18.765 286.81 18.835 ;
    RECT 286.14 18.045 286.35 18.115 ;
    RECT 286.14 18.405 286.35 18.475 ;
    RECT 286.14 18.765 286.35 18.835 ;
    RECT 283.28 18.045 283.49 18.115 ;
    RECT 283.28 18.405 283.49 18.475 ;
    RECT 283.28 18.765 283.49 18.835 ;
    RECT 282.82 18.045 283.03 18.115 ;
    RECT 282.82 18.405 283.03 18.475 ;
    RECT 282.82 18.765 283.03 18.835 ;
    RECT 279.96 18.045 280.17 18.115 ;
    RECT 279.96 18.405 280.17 18.475 ;
    RECT 279.96 18.765 280.17 18.835 ;
    RECT 279.5 18.045 279.71 18.115 ;
    RECT 279.5 18.405 279.71 18.475 ;
    RECT 279.5 18.765 279.71 18.835 ;
    RECT 276.64 18.045 276.85 18.115 ;
    RECT 276.64 18.405 276.85 18.475 ;
    RECT 276.64 18.765 276.85 18.835 ;
    RECT 276.18 18.045 276.39 18.115 ;
    RECT 276.18 18.405 276.39 18.475 ;
    RECT 276.18 18.765 276.39 18.835 ;
    RECT 273.32 18.045 273.53 18.115 ;
    RECT 273.32 18.405 273.53 18.475 ;
    RECT 273.32 18.765 273.53 18.835 ;
    RECT 272.86 18.045 273.07 18.115 ;
    RECT 272.86 18.405 273.07 18.475 ;
    RECT 272.86 18.765 273.07 18.835 ;
    RECT 270.0 18.045 270.21 18.115 ;
    RECT 270.0 18.405 270.21 18.475 ;
    RECT 270.0 18.765 270.21 18.835 ;
    RECT 269.54 18.045 269.75 18.115 ;
    RECT 269.54 18.405 269.75 18.475 ;
    RECT 269.54 18.765 269.75 18.835 ;
    RECT 233.48 18.045 233.69 18.115 ;
    RECT 233.48 18.405 233.69 18.475 ;
    RECT 233.48 18.765 233.69 18.835 ;
    RECT 233.02 18.045 233.23 18.115 ;
    RECT 233.02 18.405 233.23 18.475 ;
    RECT 233.02 18.765 233.23 18.835 ;
    RECT 230.16 18.045 230.37 18.115 ;
    RECT 230.16 18.405 230.37 18.475 ;
    RECT 230.16 18.765 230.37 18.835 ;
    RECT 229.7 18.045 229.91 18.115 ;
    RECT 229.7 18.405 229.91 18.475 ;
    RECT 229.7 18.765 229.91 18.835 ;
    RECT 366.28 18.045 366.49 18.115 ;
    RECT 366.28 18.405 366.49 18.475 ;
    RECT 366.28 18.765 366.49 18.835 ;
    RECT 365.82 18.045 366.03 18.115 ;
    RECT 365.82 18.405 366.03 18.475 ;
    RECT 365.82 18.765 366.03 18.835 ;
    RECT 226.84 18.045 227.05 18.115 ;
    RECT 226.84 18.405 227.05 18.475 ;
    RECT 226.84 18.765 227.05 18.835 ;
    RECT 226.38 18.045 226.59 18.115 ;
    RECT 226.38 18.405 226.59 18.475 ;
    RECT 226.38 18.765 226.59 18.835 ;
    RECT 362.96 18.045 363.17 18.115 ;
    RECT 362.96 18.405 363.17 18.475 ;
    RECT 362.96 18.765 363.17 18.835 ;
    RECT 362.5 18.045 362.71 18.115 ;
    RECT 362.5 18.405 362.71 18.475 ;
    RECT 362.5 18.765 362.71 18.835 ;
    RECT 223.52 18.045 223.73 18.115 ;
    RECT 223.52 18.405 223.73 18.475 ;
    RECT 223.52 18.765 223.73 18.835 ;
    RECT 223.06 18.045 223.27 18.115 ;
    RECT 223.06 18.405 223.27 18.475 ;
    RECT 223.06 18.765 223.27 18.835 ;
    RECT 359.64 18.045 359.85 18.115 ;
    RECT 359.64 18.405 359.85 18.475 ;
    RECT 359.64 18.765 359.85 18.835 ;
    RECT 359.18 18.045 359.39 18.115 ;
    RECT 359.18 18.405 359.39 18.475 ;
    RECT 359.18 18.765 359.39 18.835 ;
    RECT 220.2 18.045 220.41 18.115 ;
    RECT 220.2 18.405 220.41 18.475 ;
    RECT 220.2 18.765 220.41 18.835 ;
    RECT 219.74 18.045 219.95 18.115 ;
    RECT 219.74 18.405 219.95 18.475 ;
    RECT 219.74 18.765 219.95 18.835 ;
    RECT 356.32 18.045 356.53 18.115 ;
    RECT 356.32 18.405 356.53 18.475 ;
    RECT 356.32 18.765 356.53 18.835 ;
    RECT 355.86 18.045 356.07 18.115 ;
    RECT 355.86 18.405 356.07 18.475 ;
    RECT 355.86 18.765 356.07 18.835 ;
    RECT 353.0 18.045 353.21 18.115 ;
    RECT 353.0 18.405 353.21 18.475 ;
    RECT 353.0 18.765 353.21 18.835 ;
    RECT 352.54 18.045 352.75 18.115 ;
    RECT 352.54 18.405 352.75 18.475 ;
    RECT 352.54 18.765 352.75 18.835 ;
    RECT 216.88 18.045 217.09 18.115 ;
    RECT 216.88 18.405 217.09 18.475 ;
    RECT 216.88 18.765 217.09 18.835 ;
    RECT 216.42 18.045 216.63 18.115 ;
    RECT 216.42 18.405 216.63 18.475 ;
    RECT 216.42 18.765 216.63 18.835 ;
    RECT 349.68 18.045 349.89 18.115 ;
    RECT 349.68 18.405 349.89 18.475 ;
    RECT 349.68 18.765 349.89 18.835 ;
    RECT 349.22 18.045 349.43 18.115 ;
    RECT 349.22 18.405 349.43 18.475 ;
    RECT 349.22 18.765 349.43 18.835 ;
    RECT 213.56 18.045 213.77 18.115 ;
    RECT 213.56 18.405 213.77 18.475 ;
    RECT 213.56 18.765 213.77 18.835 ;
    RECT 213.1 18.045 213.31 18.115 ;
    RECT 213.1 18.405 213.31 18.475 ;
    RECT 213.1 18.765 213.31 18.835 ;
    RECT 346.36 18.045 346.57 18.115 ;
    RECT 346.36 18.405 346.57 18.475 ;
    RECT 346.36 18.765 346.57 18.835 ;
    RECT 345.9 18.045 346.11 18.115 ;
    RECT 345.9 18.405 346.11 18.475 ;
    RECT 345.9 18.765 346.11 18.835 ;
    RECT 210.24 18.045 210.45 18.115 ;
    RECT 210.24 18.405 210.45 18.475 ;
    RECT 210.24 18.765 210.45 18.835 ;
    RECT 209.78 18.045 209.99 18.115 ;
    RECT 209.78 18.405 209.99 18.475 ;
    RECT 209.78 18.765 209.99 18.835 ;
    RECT 343.04 18.045 343.25 18.115 ;
    RECT 343.04 18.405 343.25 18.475 ;
    RECT 343.04 18.765 343.25 18.835 ;
    RECT 342.58 18.045 342.79 18.115 ;
    RECT 342.58 18.405 342.79 18.475 ;
    RECT 342.58 18.765 342.79 18.835 ;
    RECT 206.92 18.045 207.13 18.115 ;
    RECT 206.92 18.405 207.13 18.475 ;
    RECT 206.92 18.765 207.13 18.835 ;
    RECT 206.46 18.045 206.67 18.115 ;
    RECT 206.46 18.405 206.67 18.475 ;
    RECT 206.46 18.765 206.67 18.835 ;
    RECT 339.72 18.045 339.93 18.115 ;
    RECT 339.72 18.405 339.93 18.475 ;
    RECT 339.72 18.765 339.93 18.835 ;
    RECT 339.26 18.045 339.47 18.115 ;
    RECT 339.26 18.405 339.47 18.475 ;
    RECT 339.26 18.765 339.47 18.835 ;
    RECT 203.6 18.045 203.81 18.115 ;
    RECT 203.6 18.405 203.81 18.475 ;
    RECT 203.6 18.765 203.81 18.835 ;
    RECT 203.14 18.045 203.35 18.115 ;
    RECT 203.14 18.405 203.35 18.475 ;
    RECT 203.14 18.765 203.35 18.835 ;
    RECT 336.4 18.045 336.61 18.115 ;
    RECT 336.4 18.405 336.61 18.475 ;
    RECT 336.4 18.765 336.61 18.835 ;
    RECT 335.94 18.045 336.15 18.115 ;
    RECT 335.94 18.405 336.15 18.475 ;
    RECT 335.94 18.765 336.15 18.835 ;
    RECT 266.68 18.045 266.89 18.115 ;
    RECT 266.68 18.405 266.89 18.475 ;
    RECT 266.68 18.765 266.89 18.835 ;
    RECT 266.22 18.045 266.43 18.115 ;
    RECT 266.22 18.405 266.43 18.475 ;
    RECT 266.22 18.765 266.43 18.835 ;
    RECT 263.36 18.045 263.57 18.115 ;
    RECT 263.36 18.405 263.57 18.475 ;
    RECT 263.36 18.765 263.57 18.835 ;
    RECT 262.9 18.045 263.11 18.115 ;
    RECT 262.9 18.405 263.11 18.475 ;
    RECT 262.9 18.765 263.11 18.835 ;
    RECT 260.04 18.045 260.25 18.115 ;
    RECT 260.04 18.405 260.25 18.475 ;
    RECT 260.04 18.765 260.25 18.835 ;
    RECT 259.58 18.045 259.79 18.115 ;
    RECT 259.58 18.405 259.79 18.475 ;
    RECT 259.58 18.765 259.79 18.835 ;
    RECT 256.72 18.045 256.93 18.115 ;
    RECT 256.72 18.405 256.93 18.475 ;
    RECT 256.72 18.765 256.93 18.835 ;
    RECT 256.26 18.045 256.47 18.115 ;
    RECT 256.26 18.405 256.47 18.475 ;
    RECT 256.26 18.765 256.47 18.835 ;
    RECT 253.4 18.045 253.61 18.115 ;
    RECT 253.4 18.405 253.61 18.475 ;
    RECT 253.4 18.765 253.61 18.835 ;
    RECT 252.94 18.045 253.15 18.115 ;
    RECT 252.94 18.405 253.15 18.475 ;
    RECT 252.94 18.765 253.15 18.835 ;
    RECT 250.08 18.045 250.29 18.115 ;
    RECT 250.08 18.405 250.29 18.475 ;
    RECT 250.08 18.765 250.29 18.835 ;
    RECT 249.62 18.045 249.83 18.115 ;
    RECT 249.62 18.405 249.83 18.475 ;
    RECT 249.62 18.765 249.83 18.835 ;
    RECT 246.76 18.045 246.97 18.115 ;
    RECT 246.76 18.405 246.97 18.475 ;
    RECT 246.76 18.765 246.97 18.835 ;
    RECT 246.3 18.045 246.51 18.115 ;
    RECT 246.3 18.405 246.51 18.475 ;
    RECT 246.3 18.765 246.51 18.835 ;
    RECT 243.44 18.045 243.65 18.115 ;
    RECT 243.44 18.405 243.65 18.475 ;
    RECT 243.44 18.765 243.65 18.835 ;
    RECT 242.98 18.045 243.19 18.115 ;
    RECT 242.98 18.405 243.19 18.475 ;
    RECT 242.98 18.765 243.19 18.835 ;
    RECT 240.12 18.045 240.33 18.115 ;
    RECT 240.12 18.405 240.33 18.475 ;
    RECT 240.12 18.765 240.33 18.835 ;
    RECT 239.66 18.045 239.87 18.115 ;
    RECT 239.66 18.405 239.87 18.475 ;
    RECT 239.66 18.765 239.87 18.835 ;
    RECT 236.8 18.045 237.01 18.115 ;
    RECT 236.8 18.405 237.01 18.475 ;
    RECT 236.8 18.765 237.01 18.835 ;
    RECT 236.34 18.045 236.55 18.115 ;
    RECT 236.34 18.405 236.55 18.475 ;
    RECT 236.34 18.765 236.55 18.835 ;
    RECT 374.15 18.405 374.22 18.475 ;
    RECT 333.08 18.045 333.29 18.115 ;
    RECT 333.08 18.405 333.29 18.475 ;
    RECT 333.08 18.765 333.29 18.835 ;
    RECT 332.62 18.045 332.83 18.115 ;
    RECT 332.62 18.405 332.83 18.475 ;
    RECT 332.62 18.765 332.83 18.835 ;
    RECT 329.76 18.045 329.97 18.115 ;
    RECT 329.76 18.405 329.97 18.475 ;
    RECT 329.76 18.765 329.97 18.835 ;
    RECT 329.3 18.045 329.51 18.115 ;
    RECT 329.3 18.405 329.51 18.475 ;
    RECT 329.3 18.765 329.51 18.835 ;
    RECT 326.44 18.045 326.65 18.115 ;
    RECT 326.44 18.405 326.65 18.475 ;
    RECT 326.44 18.765 326.65 18.835 ;
    RECT 325.98 18.045 326.19 18.115 ;
    RECT 325.98 18.405 326.19 18.475 ;
    RECT 325.98 18.765 326.19 18.835 ;
    RECT 323.12 18.045 323.33 18.115 ;
    RECT 323.12 18.405 323.33 18.475 ;
    RECT 323.12 18.765 323.33 18.835 ;
    RECT 322.66 18.045 322.87 18.115 ;
    RECT 322.66 18.405 322.87 18.475 ;
    RECT 322.66 18.765 322.87 18.835 ;
    RECT 319.8 18.045 320.01 18.115 ;
    RECT 319.8 18.405 320.01 18.475 ;
    RECT 319.8 18.765 320.01 18.835 ;
    RECT 319.34 18.045 319.55 18.115 ;
    RECT 319.34 18.405 319.55 18.475 ;
    RECT 319.34 18.765 319.55 18.835 ;
    RECT 316.48 18.045 316.69 18.115 ;
    RECT 316.48 18.405 316.69 18.475 ;
    RECT 316.48 18.765 316.69 18.835 ;
    RECT 316.02 18.045 316.23 18.115 ;
    RECT 316.02 18.405 316.23 18.475 ;
    RECT 316.02 18.765 316.23 18.835 ;
    RECT 313.16 18.045 313.37 18.115 ;
    RECT 313.16 18.405 313.37 18.475 ;
    RECT 313.16 18.765 313.37 18.835 ;
    RECT 312.7 18.045 312.91 18.115 ;
    RECT 312.7 18.405 312.91 18.475 ;
    RECT 312.7 18.765 312.91 18.835 ;
    RECT 309.84 18.045 310.05 18.115 ;
    RECT 309.84 18.405 310.05 18.475 ;
    RECT 309.84 18.765 310.05 18.835 ;
    RECT 309.38 18.045 309.59 18.115 ;
    RECT 309.38 18.405 309.59 18.475 ;
    RECT 309.38 18.765 309.59 18.835 ;
    RECT 306.52 18.045 306.73 18.115 ;
    RECT 306.52 18.405 306.73 18.475 ;
    RECT 306.52 18.765 306.73 18.835 ;
    RECT 306.06 18.045 306.27 18.115 ;
    RECT 306.06 18.405 306.27 18.475 ;
    RECT 306.06 18.765 306.27 18.835 ;
    RECT 303.2 17.325 303.41 17.395 ;
    RECT 303.2 17.685 303.41 17.755 ;
    RECT 303.2 18.045 303.41 18.115 ;
    RECT 302.74 17.325 302.95 17.395 ;
    RECT 302.74 17.685 302.95 17.755 ;
    RECT 302.74 18.045 302.95 18.115 ;
    RECT 372.92 17.325 373.13 17.395 ;
    RECT 372.92 17.685 373.13 17.755 ;
    RECT 372.92 18.045 373.13 18.115 ;
    RECT 372.46 17.325 372.67 17.395 ;
    RECT 372.46 17.685 372.67 17.755 ;
    RECT 372.46 18.045 372.67 18.115 ;
    RECT 369.6 17.325 369.81 17.395 ;
    RECT 369.6 17.685 369.81 17.755 ;
    RECT 369.6 18.045 369.81 18.115 ;
    RECT 369.14 17.325 369.35 17.395 ;
    RECT 369.14 17.685 369.35 17.755 ;
    RECT 369.14 18.045 369.35 18.115 ;
    RECT 200.605 17.685 200.675 17.755 ;
    RECT 299.88 17.325 300.09 17.395 ;
    RECT 299.88 17.685 300.09 17.755 ;
    RECT 299.88 18.045 300.09 18.115 ;
    RECT 299.42 17.325 299.63 17.395 ;
    RECT 299.42 17.685 299.63 17.755 ;
    RECT 299.42 18.045 299.63 18.115 ;
    RECT 296.56 17.325 296.77 17.395 ;
    RECT 296.56 17.685 296.77 17.755 ;
    RECT 296.56 18.045 296.77 18.115 ;
    RECT 296.1 17.325 296.31 17.395 ;
    RECT 296.1 17.685 296.31 17.755 ;
    RECT 296.1 18.045 296.31 18.115 ;
    RECT 293.24 17.325 293.45 17.395 ;
    RECT 293.24 17.685 293.45 17.755 ;
    RECT 293.24 18.045 293.45 18.115 ;
    RECT 292.78 17.325 292.99 17.395 ;
    RECT 292.78 17.685 292.99 17.755 ;
    RECT 292.78 18.045 292.99 18.115 ;
    RECT 289.92 17.325 290.13 17.395 ;
    RECT 289.92 17.685 290.13 17.755 ;
    RECT 289.92 18.045 290.13 18.115 ;
    RECT 289.46 17.325 289.67 17.395 ;
    RECT 289.46 17.685 289.67 17.755 ;
    RECT 289.46 18.045 289.67 18.115 ;
    RECT 286.6 17.325 286.81 17.395 ;
    RECT 286.6 17.685 286.81 17.755 ;
    RECT 286.6 18.045 286.81 18.115 ;
    RECT 286.14 17.325 286.35 17.395 ;
    RECT 286.14 17.685 286.35 17.755 ;
    RECT 286.14 18.045 286.35 18.115 ;
    RECT 283.28 17.325 283.49 17.395 ;
    RECT 283.28 17.685 283.49 17.755 ;
    RECT 283.28 18.045 283.49 18.115 ;
    RECT 282.82 17.325 283.03 17.395 ;
    RECT 282.82 17.685 283.03 17.755 ;
    RECT 282.82 18.045 283.03 18.115 ;
    RECT 279.96 17.325 280.17 17.395 ;
    RECT 279.96 17.685 280.17 17.755 ;
    RECT 279.96 18.045 280.17 18.115 ;
    RECT 279.5 17.325 279.71 17.395 ;
    RECT 279.5 17.685 279.71 17.755 ;
    RECT 279.5 18.045 279.71 18.115 ;
    RECT 276.64 17.325 276.85 17.395 ;
    RECT 276.64 17.685 276.85 17.755 ;
    RECT 276.64 18.045 276.85 18.115 ;
    RECT 276.18 17.325 276.39 17.395 ;
    RECT 276.18 17.685 276.39 17.755 ;
    RECT 276.18 18.045 276.39 18.115 ;
    RECT 273.32 17.325 273.53 17.395 ;
    RECT 273.32 17.685 273.53 17.755 ;
    RECT 273.32 18.045 273.53 18.115 ;
    RECT 272.86 17.325 273.07 17.395 ;
    RECT 272.86 17.685 273.07 17.755 ;
    RECT 272.86 18.045 273.07 18.115 ;
    RECT 270.0 17.325 270.21 17.395 ;
    RECT 270.0 17.685 270.21 17.755 ;
    RECT 270.0 18.045 270.21 18.115 ;
    RECT 269.54 17.325 269.75 17.395 ;
    RECT 269.54 17.685 269.75 17.755 ;
    RECT 269.54 18.045 269.75 18.115 ;
    RECT 233.48 17.325 233.69 17.395 ;
    RECT 233.48 17.685 233.69 17.755 ;
    RECT 233.48 18.045 233.69 18.115 ;
    RECT 233.02 17.325 233.23 17.395 ;
    RECT 233.02 17.685 233.23 17.755 ;
    RECT 233.02 18.045 233.23 18.115 ;
    RECT 230.16 17.325 230.37 17.395 ;
    RECT 230.16 17.685 230.37 17.755 ;
    RECT 230.16 18.045 230.37 18.115 ;
    RECT 229.7 17.325 229.91 17.395 ;
    RECT 229.7 17.685 229.91 17.755 ;
    RECT 229.7 18.045 229.91 18.115 ;
    RECT 366.28 17.325 366.49 17.395 ;
    RECT 366.28 17.685 366.49 17.755 ;
    RECT 366.28 18.045 366.49 18.115 ;
    RECT 365.82 17.325 366.03 17.395 ;
    RECT 365.82 17.685 366.03 17.755 ;
    RECT 365.82 18.045 366.03 18.115 ;
    RECT 226.84 17.325 227.05 17.395 ;
    RECT 226.84 17.685 227.05 17.755 ;
    RECT 226.84 18.045 227.05 18.115 ;
    RECT 226.38 17.325 226.59 17.395 ;
    RECT 226.38 17.685 226.59 17.755 ;
    RECT 226.38 18.045 226.59 18.115 ;
    RECT 362.96 17.325 363.17 17.395 ;
    RECT 362.96 17.685 363.17 17.755 ;
    RECT 362.96 18.045 363.17 18.115 ;
    RECT 362.5 17.325 362.71 17.395 ;
    RECT 362.5 17.685 362.71 17.755 ;
    RECT 362.5 18.045 362.71 18.115 ;
    RECT 223.52 17.325 223.73 17.395 ;
    RECT 223.52 17.685 223.73 17.755 ;
    RECT 223.52 18.045 223.73 18.115 ;
    RECT 223.06 17.325 223.27 17.395 ;
    RECT 223.06 17.685 223.27 17.755 ;
    RECT 223.06 18.045 223.27 18.115 ;
    RECT 359.64 17.325 359.85 17.395 ;
    RECT 359.64 17.685 359.85 17.755 ;
    RECT 359.64 18.045 359.85 18.115 ;
    RECT 359.18 17.325 359.39 17.395 ;
    RECT 359.18 17.685 359.39 17.755 ;
    RECT 359.18 18.045 359.39 18.115 ;
    RECT 220.2 17.325 220.41 17.395 ;
    RECT 220.2 17.685 220.41 17.755 ;
    RECT 220.2 18.045 220.41 18.115 ;
    RECT 219.74 17.325 219.95 17.395 ;
    RECT 219.74 17.685 219.95 17.755 ;
    RECT 219.74 18.045 219.95 18.115 ;
    RECT 356.32 17.325 356.53 17.395 ;
    RECT 356.32 17.685 356.53 17.755 ;
    RECT 356.32 18.045 356.53 18.115 ;
    RECT 355.86 17.325 356.07 17.395 ;
    RECT 355.86 17.685 356.07 17.755 ;
    RECT 355.86 18.045 356.07 18.115 ;
    RECT 353.0 17.325 353.21 17.395 ;
    RECT 353.0 17.685 353.21 17.755 ;
    RECT 353.0 18.045 353.21 18.115 ;
    RECT 352.54 17.325 352.75 17.395 ;
    RECT 352.54 17.685 352.75 17.755 ;
    RECT 352.54 18.045 352.75 18.115 ;
    RECT 216.88 17.325 217.09 17.395 ;
    RECT 216.88 17.685 217.09 17.755 ;
    RECT 216.88 18.045 217.09 18.115 ;
    RECT 216.42 17.325 216.63 17.395 ;
    RECT 216.42 17.685 216.63 17.755 ;
    RECT 216.42 18.045 216.63 18.115 ;
    RECT 349.68 17.325 349.89 17.395 ;
    RECT 349.68 17.685 349.89 17.755 ;
    RECT 349.68 18.045 349.89 18.115 ;
    RECT 349.22 17.325 349.43 17.395 ;
    RECT 349.22 17.685 349.43 17.755 ;
    RECT 349.22 18.045 349.43 18.115 ;
    RECT 213.56 17.325 213.77 17.395 ;
    RECT 213.56 17.685 213.77 17.755 ;
    RECT 213.56 18.045 213.77 18.115 ;
    RECT 213.1 17.325 213.31 17.395 ;
    RECT 213.1 17.685 213.31 17.755 ;
    RECT 213.1 18.045 213.31 18.115 ;
    RECT 346.36 17.325 346.57 17.395 ;
    RECT 346.36 17.685 346.57 17.755 ;
    RECT 346.36 18.045 346.57 18.115 ;
    RECT 345.9 17.325 346.11 17.395 ;
    RECT 345.9 17.685 346.11 17.755 ;
    RECT 345.9 18.045 346.11 18.115 ;
    RECT 210.24 17.325 210.45 17.395 ;
    RECT 210.24 17.685 210.45 17.755 ;
    RECT 210.24 18.045 210.45 18.115 ;
    RECT 209.78 17.325 209.99 17.395 ;
    RECT 209.78 17.685 209.99 17.755 ;
    RECT 209.78 18.045 209.99 18.115 ;
    RECT 343.04 17.325 343.25 17.395 ;
    RECT 343.04 17.685 343.25 17.755 ;
    RECT 343.04 18.045 343.25 18.115 ;
    RECT 342.58 17.325 342.79 17.395 ;
    RECT 342.58 17.685 342.79 17.755 ;
    RECT 342.58 18.045 342.79 18.115 ;
    RECT 206.92 17.325 207.13 17.395 ;
    RECT 206.92 17.685 207.13 17.755 ;
    RECT 206.92 18.045 207.13 18.115 ;
    RECT 206.46 17.325 206.67 17.395 ;
    RECT 206.46 17.685 206.67 17.755 ;
    RECT 206.46 18.045 206.67 18.115 ;
    RECT 339.72 17.325 339.93 17.395 ;
    RECT 339.72 17.685 339.93 17.755 ;
    RECT 339.72 18.045 339.93 18.115 ;
    RECT 339.26 17.325 339.47 17.395 ;
    RECT 339.26 17.685 339.47 17.755 ;
    RECT 339.26 18.045 339.47 18.115 ;
    RECT 203.6 17.325 203.81 17.395 ;
    RECT 203.6 17.685 203.81 17.755 ;
    RECT 203.6 18.045 203.81 18.115 ;
    RECT 203.14 17.325 203.35 17.395 ;
    RECT 203.14 17.685 203.35 17.755 ;
    RECT 203.14 18.045 203.35 18.115 ;
    RECT 336.4 17.325 336.61 17.395 ;
    RECT 336.4 17.685 336.61 17.755 ;
    RECT 336.4 18.045 336.61 18.115 ;
    RECT 335.94 17.325 336.15 17.395 ;
    RECT 335.94 17.685 336.15 17.755 ;
    RECT 335.94 18.045 336.15 18.115 ;
    RECT 266.68 17.325 266.89 17.395 ;
    RECT 266.68 17.685 266.89 17.755 ;
    RECT 266.68 18.045 266.89 18.115 ;
    RECT 266.22 17.325 266.43 17.395 ;
    RECT 266.22 17.685 266.43 17.755 ;
    RECT 266.22 18.045 266.43 18.115 ;
    RECT 263.36 17.325 263.57 17.395 ;
    RECT 263.36 17.685 263.57 17.755 ;
    RECT 263.36 18.045 263.57 18.115 ;
    RECT 262.9 17.325 263.11 17.395 ;
    RECT 262.9 17.685 263.11 17.755 ;
    RECT 262.9 18.045 263.11 18.115 ;
    RECT 260.04 17.325 260.25 17.395 ;
    RECT 260.04 17.685 260.25 17.755 ;
    RECT 260.04 18.045 260.25 18.115 ;
    RECT 259.58 17.325 259.79 17.395 ;
    RECT 259.58 17.685 259.79 17.755 ;
    RECT 259.58 18.045 259.79 18.115 ;
    RECT 256.72 17.325 256.93 17.395 ;
    RECT 256.72 17.685 256.93 17.755 ;
    RECT 256.72 18.045 256.93 18.115 ;
    RECT 256.26 17.325 256.47 17.395 ;
    RECT 256.26 17.685 256.47 17.755 ;
    RECT 256.26 18.045 256.47 18.115 ;
    RECT 253.4 17.325 253.61 17.395 ;
    RECT 253.4 17.685 253.61 17.755 ;
    RECT 253.4 18.045 253.61 18.115 ;
    RECT 252.94 17.325 253.15 17.395 ;
    RECT 252.94 17.685 253.15 17.755 ;
    RECT 252.94 18.045 253.15 18.115 ;
    RECT 250.08 17.325 250.29 17.395 ;
    RECT 250.08 17.685 250.29 17.755 ;
    RECT 250.08 18.045 250.29 18.115 ;
    RECT 249.62 17.325 249.83 17.395 ;
    RECT 249.62 17.685 249.83 17.755 ;
    RECT 249.62 18.045 249.83 18.115 ;
    RECT 246.76 17.325 246.97 17.395 ;
    RECT 246.76 17.685 246.97 17.755 ;
    RECT 246.76 18.045 246.97 18.115 ;
    RECT 246.3 17.325 246.51 17.395 ;
    RECT 246.3 17.685 246.51 17.755 ;
    RECT 246.3 18.045 246.51 18.115 ;
    RECT 243.44 17.325 243.65 17.395 ;
    RECT 243.44 17.685 243.65 17.755 ;
    RECT 243.44 18.045 243.65 18.115 ;
    RECT 242.98 17.325 243.19 17.395 ;
    RECT 242.98 17.685 243.19 17.755 ;
    RECT 242.98 18.045 243.19 18.115 ;
    RECT 240.12 17.325 240.33 17.395 ;
    RECT 240.12 17.685 240.33 17.755 ;
    RECT 240.12 18.045 240.33 18.115 ;
    RECT 239.66 17.325 239.87 17.395 ;
    RECT 239.66 17.685 239.87 17.755 ;
    RECT 239.66 18.045 239.87 18.115 ;
    RECT 236.8 17.325 237.01 17.395 ;
    RECT 236.8 17.685 237.01 17.755 ;
    RECT 236.8 18.045 237.01 18.115 ;
    RECT 236.34 17.325 236.55 17.395 ;
    RECT 236.34 17.685 236.55 17.755 ;
    RECT 236.34 18.045 236.55 18.115 ;
    RECT 374.15 17.685 374.22 17.755 ;
    RECT 333.08 17.325 333.29 17.395 ;
    RECT 333.08 17.685 333.29 17.755 ;
    RECT 333.08 18.045 333.29 18.115 ;
    RECT 332.62 17.325 332.83 17.395 ;
    RECT 332.62 17.685 332.83 17.755 ;
    RECT 332.62 18.045 332.83 18.115 ;
    RECT 329.76 17.325 329.97 17.395 ;
    RECT 329.76 17.685 329.97 17.755 ;
    RECT 329.76 18.045 329.97 18.115 ;
    RECT 329.3 17.325 329.51 17.395 ;
    RECT 329.3 17.685 329.51 17.755 ;
    RECT 329.3 18.045 329.51 18.115 ;
    RECT 326.44 17.325 326.65 17.395 ;
    RECT 326.44 17.685 326.65 17.755 ;
    RECT 326.44 18.045 326.65 18.115 ;
    RECT 325.98 17.325 326.19 17.395 ;
    RECT 325.98 17.685 326.19 17.755 ;
    RECT 325.98 18.045 326.19 18.115 ;
    RECT 323.12 17.325 323.33 17.395 ;
    RECT 323.12 17.685 323.33 17.755 ;
    RECT 323.12 18.045 323.33 18.115 ;
    RECT 322.66 17.325 322.87 17.395 ;
    RECT 322.66 17.685 322.87 17.755 ;
    RECT 322.66 18.045 322.87 18.115 ;
    RECT 319.8 17.325 320.01 17.395 ;
    RECT 319.8 17.685 320.01 17.755 ;
    RECT 319.8 18.045 320.01 18.115 ;
    RECT 319.34 17.325 319.55 17.395 ;
    RECT 319.34 17.685 319.55 17.755 ;
    RECT 319.34 18.045 319.55 18.115 ;
    RECT 316.48 17.325 316.69 17.395 ;
    RECT 316.48 17.685 316.69 17.755 ;
    RECT 316.48 18.045 316.69 18.115 ;
    RECT 316.02 17.325 316.23 17.395 ;
    RECT 316.02 17.685 316.23 17.755 ;
    RECT 316.02 18.045 316.23 18.115 ;
    RECT 313.16 17.325 313.37 17.395 ;
    RECT 313.16 17.685 313.37 17.755 ;
    RECT 313.16 18.045 313.37 18.115 ;
    RECT 312.7 17.325 312.91 17.395 ;
    RECT 312.7 17.685 312.91 17.755 ;
    RECT 312.7 18.045 312.91 18.115 ;
    RECT 309.84 17.325 310.05 17.395 ;
    RECT 309.84 17.685 310.05 17.755 ;
    RECT 309.84 18.045 310.05 18.115 ;
    RECT 309.38 17.325 309.59 17.395 ;
    RECT 309.38 17.685 309.59 17.755 ;
    RECT 309.38 18.045 309.59 18.115 ;
    RECT 306.52 17.325 306.73 17.395 ;
    RECT 306.52 17.685 306.73 17.755 ;
    RECT 306.52 18.045 306.73 18.115 ;
    RECT 306.06 17.325 306.27 17.395 ;
    RECT 306.06 17.685 306.27 17.755 ;
    RECT 306.06 18.045 306.27 18.115 ;
    RECT 303.2 16.605 303.41 16.675 ;
    RECT 303.2 16.965 303.41 17.035 ;
    RECT 303.2 17.325 303.41 17.395 ;
    RECT 302.74 16.605 302.95 16.675 ;
    RECT 302.74 16.965 302.95 17.035 ;
    RECT 302.74 17.325 302.95 17.395 ;
    RECT 372.92 16.605 373.13 16.675 ;
    RECT 372.92 16.965 373.13 17.035 ;
    RECT 372.92 17.325 373.13 17.395 ;
    RECT 372.46 16.605 372.67 16.675 ;
    RECT 372.46 16.965 372.67 17.035 ;
    RECT 372.46 17.325 372.67 17.395 ;
    RECT 369.6 16.605 369.81 16.675 ;
    RECT 369.6 16.965 369.81 17.035 ;
    RECT 369.6 17.325 369.81 17.395 ;
    RECT 369.14 16.605 369.35 16.675 ;
    RECT 369.14 16.965 369.35 17.035 ;
    RECT 369.14 17.325 369.35 17.395 ;
    RECT 200.605 16.965 200.675 17.035 ;
    RECT 299.88 16.605 300.09 16.675 ;
    RECT 299.88 16.965 300.09 17.035 ;
    RECT 299.88 17.325 300.09 17.395 ;
    RECT 299.42 16.605 299.63 16.675 ;
    RECT 299.42 16.965 299.63 17.035 ;
    RECT 299.42 17.325 299.63 17.395 ;
    RECT 296.56 16.605 296.77 16.675 ;
    RECT 296.56 16.965 296.77 17.035 ;
    RECT 296.56 17.325 296.77 17.395 ;
    RECT 296.1 16.605 296.31 16.675 ;
    RECT 296.1 16.965 296.31 17.035 ;
    RECT 296.1 17.325 296.31 17.395 ;
    RECT 293.24 16.605 293.45 16.675 ;
    RECT 293.24 16.965 293.45 17.035 ;
    RECT 293.24 17.325 293.45 17.395 ;
    RECT 292.78 16.605 292.99 16.675 ;
    RECT 292.78 16.965 292.99 17.035 ;
    RECT 292.78 17.325 292.99 17.395 ;
    RECT 289.92 16.605 290.13 16.675 ;
    RECT 289.92 16.965 290.13 17.035 ;
    RECT 289.92 17.325 290.13 17.395 ;
    RECT 289.46 16.605 289.67 16.675 ;
    RECT 289.46 16.965 289.67 17.035 ;
    RECT 289.46 17.325 289.67 17.395 ;
    RECT 286.6 16.605 286.81 16.675 ;
    RECT 286.6 16.965 286.81 17.035 ;
    RECT 286.6 17.325 286.81 17.395 ;
    RECT 286.14 16.605 286.35 16.675 ;
    RECT 286.14 16.965 286.35 17.035 ;
    RECT 286.14 17.325 286.35 17.395 ;
    RECT 283.28 16.605 283.49 16.675 ;
    RECT 283.28 16.965 283.49 17.035 ;
    RECT 283.28 17.325 283.49 17.395 ;
    RECT 282.82 16.605 283.03 16.675 ;
    RECT 282.82 16.965 283.03 17.035 ;
    RECT 282.82 17.325 283.03 17.395 ;
    RECT 279.96 16.605 280.17 16.675 ;
    RECT 279.96 16.965 280.17 17.035 ;
    RECT 279.96 17.325 280.17 17.395 ;
    RECT 279.5 16.605 279.71 16.675 ;
    RECT 279.5 16.965 279.71 17.035 ;
    RECT 279.5 17.325 279.71 17.395 ;
    RECT 276.64 16.605 276.85 16.675 ;
    RECT 276.64 16.965 276.85 17.035 ;
    RECT 276.64 17.325 276.85 17.395 ;
    RECT 276.18 16.605 276.39 16.675 ;
    RECT 276.18 16.965 276.39 17.035 ;
    RECT 276.18 17.325 276.39 17.395 ;
    RECT 273.32 16.605 273.53 16.675 ;
    RECT 273.32 16.965 273.53 17.035 ;
    RECT 273.32 17.325 273.53 17.395 ;
    RECT 272.86 16.605 273.07 16.675 ;
    RECT 272.86 16.965 273.07 17.035 ;
    RECT 272.86 17.325 273.07 17.395 ;
    RECT 270.0 16.605 270.21 16.675 ;
    RECT 270.0 16.965 270.21 17.035 ;
    RECT 270.0 17.325 270.21 17.395 ;
    RECT 269.54 16.605 269.75 16.675 ;
    RECT 269.54 16.965 269.75 17.035 ;
    RECT 269.54 17.325 269.75 17.395 ;
    RECT 233.48 16.605 233.69 16.675 ;
    RECT 233.48 16.965 233.69 17.035 ;
    RECT 233.48 17.325 233.69 17.395 ;
    RECT 233.02 16.605 233.23 16.675 ;
    RECT 233.02 16.965 233.23 17.035 ;
    RECT 233.02 17.325 233.23 17.395 ;
    RECT 230.16 16.605 230.37 16.675 ;
    RECT 230.16 16.965 230.37 17.035 ;
    RECT 230.16 17.325 230.37 17.395 ;
    RECT 229.7 16.605 229.91 16.675 ;
    RECT 229.7 16.965 229.91 17.035 ;
    RECT 229.7 17.325 229.91 17.395 ;
    RECT 366.28 16.605 366.49 16.675 ;
    RECT 366.28 16.965 366.49 17.035 ;
    RECT 366.28 17.325 366.49 17.395 ;
    RECT 365.82 16.605 366.03 16.675 ;
    RECT 365.82 16.965 366.03 17.035 ;
    RECT 365.82 17.325 366.03 17.395 ;
    RECT 226.84 16.605 227.05 16.675 ;
    RECT 226.84 16.965 227.05 17.035 ;
    RECT 226.84 17.325 227.05 17.395 ;
    RECT 226.38 16.605 226.59 16.675 ;
    RECT 226.38 16.965 226.59 17.035 ;
    RECT 226.38 17.325 226.59 17.395 ;
    RECT 362.96 16.605 363.17 16.675 ;
    RECT 362.96 16.965 363.17 17.035 ;
    RECT 362.96 17.325 363.17 17.395 ;
    RECT 362.5 16.605 362.71 16.675 ;
    RECT 362.5 16.965 362.71 17.035 ;
    RECT 362.5 17.325 362.71 17.395 ;
    RECT 223.52 16.605 223.73 16.675 ;
    RECT 223.52 16.965 223.73 17.035 ;
    RECT 223.52 17.325 223.73 17.395 ;
    RECT 223.06 16.605 223.27 16.675 ;
    RECT 223.06 16.965 223.27 17.035 ;
    RECT 223.06 17.325 223.27 17.395 ;
    RECT 359.64 16.605 359.85 16.675 ;
    RECT 359.64 16.965 359.85 17.035 ;
    RECT 359.64 17.325 359.85 17.395 ;
    RECT 359.18 16.605 359.39 16.675 ;
    RECT 359.18 16.965 359.39 17.035 ;
    RECT 359.18 17.325 359.39 17.395 ;
    RECT 220.2 16.605 220.41 16.675 ;
    RECT 220.2 16.965 220.41 17.035 ;
    RECT 220.2 17.325 220.41 17.395 ;
    RECT 219.74 16.605 219.95 16.675 ;
    RECT 219.74 16.965 219.95 17.035 ;
    RECT 219.74 17.325 219.95 17.395 ;
    RECT 356.32 16.605 356.53 16.675 ;
    RECT 356.32 16.965 356.53 17.035 ;
    RECT 356.32 17.325 356.53 17.395 ;
    RECT 355.86 16.605 356.07 16.675 ;
    RECT 355.86 16.965 356.07 17.035 ;
    RECT 355.86 17.325 356.07 17.395 ;
    RECT 353.0 16.605 353.21 16.675 ;
    RECT 353.0 16.965 353.21 17.035 ;
    RECT 353.0 17.325 353.21 17.395 ;
    RECT 352.54 16.605 352.75 16.675 ;
    RECT 352.54 16.965 352.75 17.035 ;
    RECT 352.54 17.325 352.75 17.395 ;
    RECT 216.88 16.605 217.09 16.675 ;
    RECT 216.88 16.965 217.09 17.035 ;
    RECT 216.88 17.325 217.09 17.395 ;
    RECT 216.42 16.605 216.63 16.675 ;
    RECT 216.42 16.965 216.63 17.035 ;
    RECT 216.42 17.325 216.63 17.395 ;
    RECT 349.68 16.605 349.89 16.675 ;
    RECT 349.68 16.965 349.89 17.035 ;
    RECT 349.68 17.325 349.89 17.395 ;
    RECT 349.22 16.605 349.43 16.675 ;
    RECT 349.22 16.965 349.43 17.035 ;
    RECT 349.22 17.325 349.43 17.395 ;
    RECT 213.56 16.605 213.77 16.675 ;
    RECT 213.56 16.965 213.77 17.035 ;
    RECT 213.56 17.325 213.77 17.395 ;
    RECT 213.1 16.605 213.31 16.675 ;
    RECT 213.1 16.965 213.31 17.035 ;
    RECT 213.1 17.325 213.31 17.395 ;
    RECT 346.36 16.605 346.57 16.675 ;
    RECT 346.36 16.965 346.57 17.035 ;
    RECT 346.36 17.325 346.57 17.395 ;
    RECT 345.9 16.605 346.11 16.675 ;
    RECT 345.9 16.965 346.11 17.035 ;
    RECT 345.9 17.325 346.11 17.395 ;
    RECT 210.24 16.605 210.45 16.675 ;
    RECT 210.24 16.965 210.45 17.035 ;
    RECT 210.24 17.325 210.45 17.395 ;
    RECT 209.78 16.605 209.99 16.675 ;
    RECT 209.78 16.965 209.99 17.035 ;
    RECT 209.78 17.325 209.99 17.395 ;
    RECT 343.04 16.605 343.25 16.675 ;
    RECT 343.04 16.965 343.25 17.035 ;
    RECT 343.04 17.325 343.25 17.395 ;
    RECT 342.58 16.605 342.79 16.675 ;
    RECT 342.58 16.965 342.79 17.035 ;
    RECT 342.58 17.325 342.79 17.395 ;
    RECT 206.92 16.605 207.13 16.675 ;
    RECT 206.92 16.965 207.13 17.035 ;
    RECT 206.92 17.325 207.13 17.395 ;
    RECT 206.46 16.605 206.67 16.675 ;
    RECT 206.46 16.965 206.67 17.035 ;
    RECT 206.46 17.325 206.67 17.395 ;
    RECT 339.72 16.605 339.93 16.675 ;
    RECT 339.72 16.965 339.93 17.035 ;
    RECT 339.72 17.325 339.93 17.395 ;
    RECT 339.26 16.605 339.47 16.675 ;
    RECT 339.26 16.965 339.47 17.035 ;
    RECT 339.26 17.325 339.47 17.395 ;
    RECT 203.6 16.605 203.81 16.675 ;
    RECT 203.6 16.965 203.81 17.035 ;
    RECT 203.6 17.325 203.81 17.395 ;
    RECT 203.14 16.605 203.35 16.675 ;
    RECT 203.14 16.965 203.35 17.035 ;
    RECT 203.14 17.325 203.35 17.395 ;
    RECT 336.4 16.605 336.61 16.675 ;
    RECT 336.4 16.965 336.61 17.035 ;
    RECT 336.4 17.325 336.61 17.395 ;
    RECT 335.94 16.605 336.15 16.675 ;
    RECT 335.94 16.965 336.15 17.035 ;
    RECT 335.94 17.325 336.15 17.395 ;
    RECT 266.68 16.605 266.89 16.675 ;
    RECT 266.68 16.965 266.89 17.035 ;
    RECT 266.68 17.325 266.89 17.395 ;
    RECT 266.22 16.605 266.43 16.675 ;
    RECT 266.22 16.965 266.43 17.035 ;
    RECT 266.22 17.325 266.43 17.395 ;
    RECT 263.36 16.605 263.57 16.675 ;
    RECT 263.36 16.965 263.57 17.035 ;
    RECT 263.36 17.325 263.57 17.395 ;
    RECT 262.9 16.605 263.11 16.675 ;
    RECT 262.9 16.965 263.11 17.035 ;
    RECT 262.9 17.325 263.11 17.395 ;
    RECT 260.04 16.605 260.25 16.675 ;
    RECT 260.04 16.965 260.25 17.035 ;
    RECT 260.04 17.325 260.25 17.395 ;
    RECT 259.58 16.605 259.79 16.675 ;
    RECT 259.58 16.965 259.79 17.035 ;
    RECT 259.58 17.325 259.79 17.395 ;
    RECT 256.72 16.605 256.93 16.675 ;
    RECT 256.72 16.965 256.93 17.035 ;
    RECT 256.72 17.325 256.93 17.395 ;
    RECT 256.26 16.605 256.47 16.675 ;
    RECT 256.26 16.965 256.47 17.035 ;
    RECT 256.26 17.325 256.47 17.395 ;
    RECT 253.4 16.605 253.61 16.675 ;
    RECT 253.4 16.965 253.61 17.035 ;
    RECT 253.4 17.325 253.61 17.395 ;
    RECT 252.94 16.605 253.15 16.675 ;
    RECT 252.94 16.965 253.15 17.035 ;
    RECT 252.94 17.325 253.15 17.395 ;
    RECT 250.08 16.605 250.29 16.675 ;
    RECT 250.08 16.965 250.29 17.035 ;
    RECT 250.08 17.325 250.29 17.395 ;
    RECT 249.62 16.605 249.83 16.675 ;
    RECT 249.62 16.965 249.83 17.035 ;
    RECT 249.62 17.325 249.83 17.395 ;
    RECT 246.76 16.605 246.97 16.675 ;
    RECT 246.76 16.965 246.97 17.035 ;
    RECT 246.76 17.325 246.97 17.395 ;
    RECT 246.3 16.605 246.51 16.675 ;
    RECT 246.3 16.965 246.51 17.035 ;
    RECT 246.3 17.325 246.51 17.395 ;
    RECT 243.44 16.605 243.65 16.675 ;
    RECT 243.44 16.965 243.65 17.035 ;
    RECT 243.44 17.325 243.65 17.395 ;
    RECT 242.98 16.605 243.19 16.675 ;
    RECT 242.98 16.965 243.19 17.035 ;
    RECT 242.98 17.325 243.19 17.395 ;
    RECT 240.12 16.605 240.33 16.675 ;
    RECT 240.12 16.965 240.33 17.035 ;
    RECT 240.12 17.325 240.33 17.395 ;
    RECT 239.66 16.605 239.87 16.675 ;
    RECT 239.66 16.965 239.87 17.035 ;
    RECT 239.66 17.325 239.87 17.395 ;
    RECT 236.8 16.605 237.01 16.675 ;
    RECT 236.8 16.965 237.01 17.035 ;
    RECT 236.8 17.325 237.01 17.395 ;
    RECT 236.34 16.605 236.55 16.675 ;
    RECT 236.34 16.965 236.55 17.035 ;
    RECT 236.34 17.325 236.55 17.395 ;
    RECT 374.15 16.965 374.22 17.035 ;
    RECT 333.08 16.605 333.29 16.675 ;
    RECT 333.08 16.965 333.29 17.035 ;
    RECT 333.08 17.325 333.29 17.395 ;
    RECT 332.62 16.605 332.83 16.675 ;
    RECT 332.62 16.965 332.83 17.035 ;
    RECT 332.62 17.325 332.83 17.395 ;
    RECT 329.76 16.605 329.97 16.675 ;
    RECT 329.76 16.965 329.97 17.035 ;
    RECT 329.76 17.325 329.97 17.395 ;
    RECT 329.3 16.605 329.51 16.675 ;
    RECT 329.3 16.965 329.51 17.035 ;
    RECT 329.3 17.325 329.51 17.395 ;
    RECT 326.44 16.605 326.65 16.675 ;
    RECT 326.44 16.965 326.65 17.035 ;
    RECT 326.44 17.325 326.65 17.395 ;
    RECT 325.98 16.605 326.19 16.675 ;
    RECT 325.98 16.965 326.19 17.035 ;
    RECT 325.98 17.325 326.19 17.395 ;
    RECT 323.12 16.605 323.33 16.675 ;
    RECT 323.12 16.965 323.33 17.035 ;
    RECT 323.12 17.325 323.33 17.395 ;
    RECT 322.66 16.605 322.87 16.675 ;
    RECT 322.66 16.965 322.87 17.035 ;
    RECT 322.66 17.325 322.87 17.395 ;
    RECT 319.8 16.605 320.01 16.675 ;
    RECT 319.8 16.965 320.01 17.035 ;
    RECT 319.8 17.325 320.01 17.395 ;
    RECT 319.34 16.605 319.55 16.675 ;
    RECT 319.34 16.965 319.55 17.035 ;
    RECT 319.34 17.325 319.55 17.395 ;
    RECT 316.48 16.605 316.69 16.675 ;
    RECT 316.48 16.965 316.69 17.035 ;
    RECT 316.48 17.325 316.69 17.395 ;
    RECT 316.02 16.605 316.23 16.675 ;
    RECT 316.02 16.965 316.23 17.035 ;
    RECT 316.02 17.325 316.23 17.395 ;
    RECT 313.16 16.605 313.37 16.675 ;
    RECT 313.16 16.965 313.37 17.035 ;
    RECT 313.16 17.325 313.37 17.395 ;
    RECT 312.7 16.605 312.91 16.675 ;
    RECT 312.7 16.965 312.91 17.035 ;
    RECT 312.7 17.325 312.91 17.395 ;
    RECT 309.84 16.605 310.05 16.675 ;
    RECT 309.84 16.965 310.05 17.035 ;
    RECT 309.84 17.325 310.05 17.395 ;
    RECT 309.38 16.605 309.59 16.675 ;
    RECT 309.38 16.965 309.59 17.035 ;
    RECT 309.38 17.325 309.59 17.395 ;
    RECT 306.52 16.605 306.73 16.675 ;
    RECT 306.52 16.965 306.73 17.035 ;
    RECT 306.52 17.325 306.73 17.395 ;
    RECT 306.06 16.605 306.27 16.675 ;
    RECT 306.06 16.965 306.27 17.035 ;
    RECT 306.06 17.325 306.27 17.395 ;
    RECT 303.2 32.445 303.41 32.515 ;
    RECT 303.2 32.805 303.41 32.875 ;
    RECT 303.2 33.165 303.41 33.235 ;
    RECT 302.74 32.445 302.95 32.515 ;
    RECT 302.74 32.805 302.95 32.875 ;
    RECT 302.74 33.165 302.95 33.235 ;
    RECT 372.92 32.445 373.13 32.515 ;
    RECT 372.92 32.805 373.13 32.875 ;
    RECT 372.92 33.165 373.13 33.235 ;
    RECT 372.46 32.445 372.67 32.515 ;
    RECT 372.46 32.805 372.67 32.875 ;
    RECT 372.46 33.165 372.67 33.235 ;
    RECT 369.6 32.445 369.81 32.515 ;
    RECT 369.6 32.805 369.81 32.875 ;
    RECT 369.6 33.165 369.81 33.235 ;
    RECT 369.14 32.445 369.35 32.515 ;
    RECT 369.14 32.805 369.35 32.875 ;
    RECT 369.14 33.165 369.35 33.235 ;
    RECT 200.605 32.805 200.675 32.875 ;
    RECT 299.88 32.445 300.09 32.515 ;
    RECT 299.88 32.805 300.09 32.875 ;
    RECT 299.88 33.165 300.09 33.235 ;
    RECT 299.42 32.445 299.63 32.515 ;
    RECT 299.42 32.805 299.63 32.875 ;
    RECT 299.42 33.165 299.63 33.235 ;
    RECT 296.56 32.445 296.77 32.515 ;
    RECT 296.56 32.805 296.77 32.875 ;
    RECT 296.56 33.165 296.77 33.235 ;
    RECT 296.1 32.445 296.31 32.515 ;
    RECT 296.1 32.805 296.31 32.875 ;
    RECT 296.1 33.165 296.31 33.235 ;
    RECT 293.24 32.445 293.45 32.515 ;
    RECT 293.24 32.805 293.45 32.875 ;
    RECT 293.24 33.165 293.45 33.235 ;
    RECT 292.78 32.445 292.99 32.515 ;
    RECT 292.78 32.805 292.99 32.875 ;
    RECT 292.78 33.165 292.99 33.235 ;
    RECT 289.92 32.445 290.13 32.515 ;
    RECT 289.92 32.805 290.13 32.875 ;
    RECT 289.92 33.165 290.13 33.235 ;
    RECT 289.46 32.445 289.67 32.515 ;
    RECT 289.46 32.805 289.67 32.875 ;
    RECT 289.46 33.165 289.67 33.235 ;
    RECT 286.6 32.445 286.81 32.515 ;
    RECT 286.6 32.805 286.81 32.875 ;
    RECT 286.6 33.165 286.81 33.235 ;
    RECT 286.14 32.445 286.35 32.515 ;
    RECT 286.14 32.805 286.35 32.875 ;
    RECT 286.14 33.165 286.35 33.235 ;
    RECT 283.28 32.445 283.49 32.515 ;
    RECT 283.28 32.805 283.49 32.875 ;
    RECT 283.28 33.165 283.49 33.235 ;
    RECT 282.82 32.445 283.03 32.515 ;
    RECT 282.82 32.805 283.03 32.875 ;
    RECT 282.82 33.165 283.03 33.235 ;
    RECT 279.96 32.445 280.17 32.515 ;
    RECT 279.96 32.805 280.17 32.875 ;
    RECT 279.96 33.165 280.17 33.235 ;
    RECT 279.5 32.445 279.71 32.515 ;
    RECT 279.5 32.805 279.71 32.875 ;
    RECT 279.5 33.165 279.71 33.235 ;
    RECT 276.64 32.445 276.85 32.515 ;
    RECT 276.64 32.805 276.85 32.875 ;
    RECT 276.64 33.165 276.85 33.235 ;
    RECT 276.18 32.445 276.39 32.515 ;
    RECT 276.18 32.805 276.39 32.875 ;
    RECT 276.18 33.165 276.39 33.235 ;
    RECT 273.32 32.445 273.53 32.515 ;
    RECT 273.32 32.805 273.53 32.875 ;
    RECT 273.32 33.165 273.53 33.235 ;
    RECT 272.86 32.445 273.07 32.515 ;
    RECT 272.86 32.805 273.07 32.875 ;
    RECT 272.86 33.165 273.07 33.235 ;
    RECT 270.0 32.445 270.21 32.515 ;
    RECT 270.0 32.805 270.21 32.875 ;
    RECT 270.0 33.165 270.21 33.235 ;
    RECT 269.54 32.445 269.75 32.515 ;
    RECT 269.54 32.805 269.75 32.875 ;
    RECT 269.54 33.165 269.75 33.235 ;
    RECT 233.48 32.445 233.69 32.515 ;
    RECT 233.48 32.805 233.69 32.875 ;
    RECT 233.48 33.165 233.69 33.235 ;
    RECT 233.02 32.445 233.23 32.515 ;
    RECT 233.02 32.805 233.23 32.875 ;
    RECT 233.02 33.165 233.23 33.235 ;
    RECT 230.16 32.445 230.37 32.515 ;
    RECT 230.16 32.805 230.37 32.875 ;
    RECT 230.16 33.165 230.37 33.235 ;
    RECT 229.7 32.445 229.91 32.515 ;
    RECT 229.7 32.805 229.91 32.875 ;
    RECT 229.7 33.165 229.91 33.235 ;
    RECT 366.28 32.445 366.49 32.515 ;
    RECT 366.28 32.805 366.49 32.875 ;
    RECT 366.28 33.165 366.49 33.235 ;
    RECT 365.82 32.445 366.03 32.515 ;
    RECT 365.82 32.805 366.03 32.875 ;
    RECT 365.82 33.165 366.03 33.235 ;
    RECT 226.84 32.445 227.05 32.515 ;
    RECT 226.84 32.805 227.05 32.875 ;
    RECT 226.84 33.165 227.05 33.235 ;
    RECT 226.38 32.445 226.59 32.515 ;
    RECT 226.38 32.805 226.59 32.875 ;
    RECT 226.38 33.165 226.59 33.235 ;
    RECT 362.96 32.445 363.17 32.515 ;
    RECT 362.96 32.805 363.17 32.875 ;
    RECT 362.96 33.165 363.17 33.235 ;
    RECT 362.5 32.445 362.71 32.515 ;
    RECT 362.5 32.805 362.71 32.875 ;
    RECT 362.5 33.165 362.71 33.235 ;
    RECT 223.52 32.445 223.73 32.515 ;
    RECT 223.52 32.805 223.73 32.875 ;
    RECT 223.52 33.165 223.73 33.235 ;
    RECT 223.06 32.445 223.27 32.515 ;
    RECT 223.06 32.805 223.27 32.875 ;
    RECT 223.06 33.165 223.27 33.235 ;
    RECT 359.64 32.445 359.85 32.515 ;
    RECT 359.64 32.805 359.85 32.875 ;
    RECT 359.64 33.165 359.85 33.235 ;
    RECT 359.18 32.445 359.39 32.515 ;
    RECT 359.18 32.805 359.39 32.875 ;
    RECT 359.18 33.165 359.39 33.235 ;
    RECT 220.2 32.445 220.41 32.515 ;
    RECT 220.2 32.805 220.41 32.875 ;
    RECT 220.2 33.165 220.41 33.235 ;
    RECT 219.74 32.445 219.95 32.515 ;
    RECT 219.74 32.805 219.95 32.875 ;
    RECT 219.74 33.165 219.95 33.235 ;
    RECT 356.32 32.445 356.53 32.515 ;
    RECT 356.32 32.805 356.53 32.875 ;
    RECT 356.32 33.165 356.53 33.235 ;
    RECT 355.86 32.445 356.07 32.515 ;
    RECT 355.86 32.805 356.07 32.875 ;
    RECT 355.86 33.165 356.07 33.235 ;
    RECT 353.0 32.445 353.21 32.515 ;
    RECT 353.0 32.805 353.21 32.875 ;
    RECT 353.0 33.165 353.21 33.235 ;
    RECT 352.54 32.445 352.75 32.515 ;
    RECT 352.54 32.805 352.75 32.875 ;
    RECT 352.54 33.165 352.75 33.235 ;
    RECT 216.88 32.445 217.09 32.515 ;
    RECT 216.88 32.805 217.09 32.875 ;
    RECT 216.88 33.165 217.09 33.235 ;
    RECT 216.42 32.445 216.63 32.515 ;
    RECT 216.42 32.805 216.63 32.875 ;
    RECT 216.42 33.165 216.63 33.235 ;
    RECT 349.68 32.445 349.89 32.515 ;
    RECT 349.68 32.805 349.89 32.875 ;
    RECT 349.68 33.165 349.89 33.235 ;
    RECT 349.22 32.445 349.43 32.515 ;
    RECT 349.22 32.805 349.43 32.875 ;
    RECT 349.22 33.165 349.43 33.235 ;
    RECT 213.56 32.445 213.77 32.515 ;
    RECT 213.56 32.805 213.77 32.875 ;
    RECT 213.56 33.165 213.77 33.235 ;
    RECT 213.1 32.445 213.31 32.515 ;
    RECT 213.1 32.805 213.31 32.875 ;
    RECT 213.1 33.165 213.31 33.235 ;
    RECT 346.36 32.445 346.57 32.515 ;
    RECT 346.36 32.805 346.57 32.875 ;
    RECT 346.36 33.165 346.57 33.235 ;
    RECT 345.9 32.445 346.11 32.515 ;
    RECT 345.9 32.805 346.11 32.875 ;
    RECT 345.9 33.165 346.11 33.235 ;
    RECT 210.24 32.445 210.45 32.515 ;
    RECT 210.24 32.805 210.45 32.875 ;
    RECT 210.24 33.165 210.45 33.235 ;
    RECT 209.78 32.445 209.99 32.515 ;
    RECT 209.78 32.805 209.99 32.875 ;
    RECT 209.78 33.165 209.99 33.235 ;
    RECT 343.04 32.445 343.25 32.515 ;
    RECT 343.04 32.805 343.25 32.875 ;
    RECT 343.04 33.165 343.25 33.235 ;
    RECT 342.58 32.445 342.79 32.515 ;
    RECT 342.58 32.805 342.79 32.875 ;
    RECT 342.58 33.165 342.79 33.235 ;
    RECT 206.92 32.445 207.13 32.515 ;
    RECT 206.92 32.805 207.13 32.875 ;
    RECT 206.92 33.165 207.13 33.235 ;
    RECT 206.46 32.445 206.67 32.515 ;
    RECT 206.46 32.805 206.67 32.875 ;
    RECT 206.46 33.165 206.67 33.235 ;
    RECT 339.72 32.445 339.93 32.515 ;
    RECT 339.72 32.805 339.93 32.875 ;
    RECT 339.72 33.165 339.93 33.235 ;
    RECT 339.26 32.445 339.47 32.515 ;
    RECT 339.26 32.805 339.47 32.875 ;
    RECT 339.26 33.165 339.47 33.235 ;
    RECT 203.6 32.445 203.81 32.515 ;
    RECT 203.6 32.805 203.81 32.875 ;
    RECT 203.6 33.165 203.81 33.235 ;
    RECT 203.14 32.445 203.35 32.515 ;
    RECT 203.14 32.805 203.35 32.875 ;
    RECT 203.14 33.165 203.35 33.235 ;
    RECT 336.4 32.445 336.61 32.515 ;
    RECT 336.4 32.805 336.61 32.875 ;
    RECT 336.4 33.165 336.61 33.235 ;
    RECT 335.94 32.445 336.15 32.515 ;
    RECT 335.94 32.805 336.15 32.875 ;
    RECT 335.94 33.165 336.15 33.235 ;
    RECT 266.68 32.445 266.89 32.515 ;
    RECT 266.68 32.805 266.89 32.875 ;
    RECT 266.68 33.165 266.89 33.235 ;
    RECT 266.22 32.445 266.43 32.515 ;
    RECT 266.22 32.805 266.43 32.875 ;
    RECT 266.22 33.165 266.43 33.235 ;
    RECT 263.36 32.445 263.57 32.515 ;
    RECT 263.36 32.805 263.57 32.875 ;
    RECT 263.36 33.165 263.57 33.235 ;
    RECT 262.9 32.445 263.11 32.515 ;
    RECT 262.9 32.805 263.11 32.875 ;
    RECT 262.9 33.165 263.11 33.235 ;
    RECT 260.04 32.445 260.25 32.515 ;
    RECT 260.04 32.805 260.25 32.875 ;
    RECT 260.04 33.165 260.25 33.235 ;
    RECT 259.58 32.445 259.79 32.515 ;
    RECT 259.58 32.805 259.79 32.875 ;
    RECT 259.58 33.165 259.79 33.235 ;
    RECT 256.72 32.445 256.93 32.515 ;
    RECT 256.72 32.805 256.93 32.875 ;
    RECT 256.72 33.165 256.93 33.235 ;
    RECT 256.26 32.445 256.47 32.515 ;
    RECT 256.26 32.805 256.47 32.875 ;
    RECT 256.26 33.165 256.47 33.235 ;
    RECT 253.4 32.445 253.61 32.515 ;
    RECT 253.4 32.805 253.61 32.875 ;
    RECT 253.4 33.165 253.61 33.235 ;
    RECT 252.94 32.445 253.15 32.515 ;
    RECT 252.94 32.805 253.15 32.875 ;
    RECT 252.94 33.165 253.15 33.235 ;
    RECT 250.08 32.445 250.29 32.515 ;
    RECT 250.08 32.805 250.29 32.875 ;
    RECT 250.08 33.165 250.29 33.235 ;
    RECT 249.62 32.445 249.83 32.515 ;
    RECT 249.62 32.805 249.83 32.875 ;
    RECT 249.62 33.165 249.83 33.235 ;
    RECT 246.76 32.445 246.97 32.515 ;
    RECT 246.76 32.805 246.97 32.875 ;
    RECT 246.76 33.165 246.97 33.235 ;
    RECT 246.3 32.445 246.51 32.515 ;
    RECT 246.3 32.805 246.51 32.875 ;
    RECT 246.3 33.165 246.51 33.235 ;
    RECT 243.44 32.445 243.65 32.515 ;
    RECT 243.44 32.805 243.65 32.875 ;
    RECT 243.44 33.165 243.65 33.235 ;
    RECT 242.98 32.445 243.19 32.515 ;
    RECT 242.98 32.805 243.19 32.875 ;
    RECT 242.98 33.165 243.19 33.235 ;
    RECT 240.12 32.445 240.33 32.515 ;
    RECT 240.12 32.805 240.33 32.875 ;
    RECT 240.12 33.165 240.33 33.235 ;
    RECT 239.66 32.445 239.87 32.515 ;
    RECT 239.66 32.805 239.87 32.875 ;
    RECT 239.66 33.165 239.87 33.235 ;
    RECT 236.8 32.445 237.01 32.515 ;
    RECT 236.8 32.805 237.01 32.875 ;
    RECT 236.8 33.165 237.01 33.235 ;
    RECT 236.34 32.445 236.55 32.515 ;
    RECT 236.34 32.805 236.55 32.875 ;
    RECT 236.34 33.165 236.55 33.235 ;
    RECT 374.15 32.805 374.22 32.875 ;
    RECT 333.08 32.445 333.29 32.515 ;
    RECT 333.08 32.805 333.29 32.875 ;
    RECT 333.08 33.165 333.29 33.235 ;
    RECT 332.62 32.445 332.83 32.515 ;
    RECT 332.62 32.805 332.83 32.875 ;
    RECT 332.62 33.165 332.83 33.235 ;
    RECT 329.76 32.445 329.97 32.515 ;
    RECT 329.76 32.805 329.97 32.875 ;
    RECT 329.76 33.165 329.97 33.235 ;
    RECT 329.3 32.445 329.51 32.515 ;
    RECT 329.3 32.805 329.51 32.875 ;
    RECT 329.3 33.165 329.51 33.235 ;
    RECT 326.44 32.445 326.65 32.515 ;
    RECT 326.44 32.805 326.65 32.875 ;
    RECT 326.44 33.165 326.65 33.235 ;
    RECT 325.98 32.445 326.19 32.515 ;
    RECT 325.98 32.805 326.19 32.875 ;
    RECT 325.98 33.165 326.19 33.235 ;
    RECT 323.12 32.445 323.33 32.515 ;
    RECT 323.12 32.805 323.33 32.875 ;
    RECT 323.12 33.165 323.33 33.235 ;
    RECT 322.66 32.445 322.87 32.515 ;
    RECT 322.66 32.805 322.87 32.875 ;
    RECT 322.66 33.165 322.87 33.235 ;
    RECT 319.8 32.445 320.01 32.515 ;
    RECT 319.8 32.805 320.01 32.875 ;
    RECT 319.8 33.165 320.01 33.235 ;
    RECT 319.34 32.445 319.55 32.515 ;
    RECT 319.34 32.805 319.55 32.875 ;
    RECT 319.34 33.165 319.55 33.235 ;
    RECT 316.48 32.445 316.69 32.515 ;
    RECT 316.48 32.805 316.69 32.875 ;
    RECT 316.48 33.165 316.69 33.235 ;
    RECT 316.02 32.445 316.23 32.515 ;
    RECT 316.02 32.805 316.23 32.875 ;
    RECT 316.02 33.165 316.23 33.235 ;
    RECT 313.16 32.445 313.37 32.515 ;
    RECT 313.16 32.805 313.37 32.875 ;
    RECT 313.16 33.165 313.37 33.235 ;
    RECT 312.7 32.445 312.91 32.515 ;
    RECT 312.7 32.805 312.91 32.875 ;
    RECT 312.7 33.165 312.91 33.235 ;
    RECT 309.84 32.445 310.05 32.515 ;
    RECT 309.84 32.805 310.05 32.875 ;
    RECT 309.84 33.165 310.05 33.235 ;
    RECT 309.38 32.445 309.59 32.515 ;
    RECT 309.38 32.805 309.59 32.875 ;
    RECT 309.38 33.165 309.59 33.235 ;
    RECT 306.52 32.445 306.73 32.515 ;
    RECT 306.52 32.805 306.73 32.875 ;
    RECT 306.52 33.165 306.73 33.235 ;
    RECT 306.06 32.445 306.27 32.515 ;
    RECT 306.06 32.805 306.27 32.875 ;
    RECT 306.06 33.165 306.27 33.235 ;
    RECT 303.2 15.885 303.41 15.955 ;
    RECT 303.2 16.245 303.41 16.315 ;
    RECT 303.2 16.605 303.41 16.675 ;
    RECT 302.74 15.885 302.95 15.955 ;
    RECT 302.74 16.245 302.95 16.315 ;
    RECT 302.74 16.605 302.95 16.675 ;
    RECT 372.92 15.885 373.13 15.955 ;
    RECT 372.92 16.245 373.13 16.315 ;
    RECT 372.92 16.605 373.13 16.675 ;
    RECT 372.46 15.885 372.67 15.955 ;
    RECT 372.46 16.245 372.67 16.315 ;
    RECT 372.46 16.605 372.67 16.675 ;
    RECT 369.6 15.885 369.81 15.955 ;
    RECT 369.6 16.245 369.81 16.315 ;
    RECT 369.6 16.605 369.81 16.675 ;
    RECT 369.14 15.885 369.35 15.955 ;
    RECT 369.14 16.245 369.35 16.315 ;
    RECT 369.14 16.605 369.35 16.675 ;
    RECT 200.605 16.245 200.675 16.315 ;
    RECT 299.88 15.885 300.09 15.955 ;
    RECT 299.88 16.245 300.09 16.315 ;
    RECT 299.88 16.605 300.09 16.675 ;
    RECT 299.42 15.885 299.63 15.955 ;
    RECT 299.42 16.245 299.63 16.315 ;
    RECT 299.42 16.605 299.63 16.675 ;
    RECT 296.56 15.885 296.77 15.955 ;
    RECT 296.56 16.245 296.77 16.315 ;
    RECT 296.56 16.605 296.77 16.675 ;
    RECT 296.1 15.885 296.31 15.955 ;
    RECT 296.1 16.245 296.31 16.315 ;
    RECT 296.1 16.605 296.31 16.675 ;
    RECT 293.24 15.885 293.45 15.955 ;
    RECT 293.24 16.245 293.45 16.315 ;
    RECT 293.24 16.605 293.45 16.675 ;
    RECT 292.78 15.885 292.99 15.955 ;
    RECT 292.78 16.245 292.99 16.315 ;
    RECT 292.78 16.605 292.99 16.675 ;
    RECT 289.92 15.885 290.13 15.955 ;
    RECT 289.92 16.245 290.13 16.315 ;
    RECT 289.92 16.605 290.13 16.675 ;
    RECT 289.46 15.885 289.67 15.955 ;
    RECT 289.46 16.245 289.67 16.315 ;
    RECT 289.46 16.605 289.67 16.675 ;
    RECT 286.6 15.885 286.81 15.955 ;
    RECT 286.6 16.245 286.81 16.315 ;
    RECT 286.6 16.605 286.81 16.675 ;
    RECT 286.14 15.885 286.35 15.955 ;
    RECT 286.14 16.245 286.35 16.315 ;
    RECT 286.14 16.605 286.35 16.675 ;
    RECT 283.28 15.885 283.49 15.955 ;
    RECT 283.28 16.245 283.49 16.315 ;
    RECT 283.28 16.605 283.49 16.675 ;
    RECT 282.82 15.885 283.03 15.955 ;
    RECT 282.82 16.245 283.03 16.315 ;
    RECT 282.82 16.605 283.03 16.675 ;
    RECT 279.96 15.885 280.17 15.955 ;
    RECT 279.96 16.245 280.17 16.315 ;
    RECT 279.96 16.605 280.17 16.675 ;
    RECT 279.5 15.885 279.71 15.955 ;
    RECT 279.5 16.245 279.71 16.315 ;
    RECT 279.5 16.605 279.71 16.675 ;
    RECT 276.64 15.885 276.85 15.955 ;
    RECT 276.64 16.245 276.85 16.315 ;
    RECT 276.64 16.605 276.85 16.675 ;
    RECT 276.18 15.885 276.39 15.955 ;
    RECT 276.18 16.245 276.39 16.315 ;
    RECT 276.18 16.605 276.39 16.675 ;
    RECT 273.32 15.885 273.53 15.955 ;
    RECT 273.32 16.245 273.53 16.315 ;
    RECT 273.32 16.605 273.53 16.675 ;
    RECT 272.86 15.885 273.07 15.955 ;
    RECT 272.86 16.245 273.07 16.315 ;
    RECT 272.86 16.605 273.07 16.675 ;
    RECT 270.0 15.885 270.21 15.955 ;
    RECT 270.0 16.245 270.21 16.315 ;
    RECT 270.0 16.605 270.21 16.675 ;
    RECT 269.54 15.885 269.75 15.955 ;
    RECT 269.54 16.245 269.75 16.315 ;
    RECT 269.54 16.605 269.75 16.675 ;
    RECT 233.48 15.885 233.69 15.955 ;
    RECT 233.48 16.245 233.69 16.315 ;
    RECT 233.48 16.605 233.69 16.675 ;
    RECT 233.02 15.885 233.23 15.955 ;
    RECT 233.02 16.245 233.23 16.315 ;
    RECT 233.02 16.605 233.23 16.675 ;
    RECT 230.16 15.885 230.37 15.955 ;
    RECT 230.16 16.245 230.37 16.315 ;
    RECT 230.16 16.605 230.37 16.675 ;
    RECT 229.7 15.885 229.91 15.955 ;
    RECT 229.7 16.245 229.91 16.315 ;
    RECT 229.7 16.605 229.91 16.675 ;
    RECT 366.28 15.885 366.49 15.955 ;
    RECT 366.28 16.245 366.49 16.315 ;
    RECT 366.28 16.605 366.49 16.675 ;
    RECT 365.82 15.885 366.03 15.955 ;
    RECT 365.82 16.245 366.03 16.315 ;
    RECT 365.82 16.605 366.03 16.675 ;
    RECT 226.84 15.885 227.05 15.955 ;
    RECT 226.84 16.245 227.05 16.315 ;
    RECT 226.84 16.605 227.05 16.675 ;
    RECT 226.38 15.885 226.59 15.955 ;
    RECT 226.38 16.245 226.59 16.315 ;
    RECT 226.38 16.605 226.59 16.675 ;
    RECT 362.96 15.885 363.17 15.955 ;
    RECT 362.96 16.245 363.17 16.315 ;
    RECT 362.96 16.605 363.17 16.675 ;
    RECT 362.5 15.885 362.71 15.955 ;
    RECT 362.5 16.245 362.71 16.315 ;
    RECT 362.5 16.605 362.71 16.675 ;
    RECT 223.52 15.885 223.73 15.955 ;
    RECT 223.52 16.245 223.73 16.315 ;
    RECT 223.52 16.605 223.73 16.675 ;
    RECT 223.06 15.885 223.27 15.955 ;
    RECT 223.06 16.245 223.27 16.315 ;
    RECT 223.06 16.605 223.27 16.675 ;
    RECT 359.64 15.885 359.85 15.955 ;
    RECT 359.64 16.245 359.85 16.315 ;
    RECT 359.64 16.605 359.85 16.675 ;
    RECT 359.18 15.885 359.39 15.955 ;
    RECT 359.18 16.245 359.39 16.315 ;
    RECT 359.18 16.605 359.39 16.675 ;
    RECT 220.2 15.885 220.41 15.955 ;
    RECT 220.2 16.245 220.41 16.315 ;
    RECT 220.2 16.605 220.41 16.675 ;
    RECT 219.74 15.885 219.95 15.955 ;
    RECT 219.74 16.245 219.95 16.315 ;
    RECT 219.74 16.605 219.95 16.675 ;
    RECT 356.32 15.885 356.53 15.955 ;
    RECT 356.32 16.245 356.53 16.315 ;
    RECT 356.32 16.605 356.53 16.675 ;
    RECT 355.86 15.885 356.07 15.955 ;
    RECT 355.86 16.245 356.07 16.315 ;
    RECT 355.86 16.605 356.07 16.675 ;
    RECT 353.0 15.885 353.21 15.955 ;
    RECT 353.0 16.245 353.21 16.315 ;
    RECT 353.0 16.605 353.21 16.675 ;
    RECT 352.54 15.885 352.75 15.955 ;
    RECT 352.54 16.245 352.75 16.315 ;
    RECT 352.54 16.605 352.75 16.675 ;
    RECT 216.88 15.885 217.09 15.955 ;
    RECT 216.88 16.245 217.09 16.315 ;
    RECT 216.88 16.605 217.09 16.675 ;
    RECT 216.42 15.885 216.63 15.955 ;
    RECT 216.42 16.245 216.63 16.315 ;
    RECT 216.42 16.605 216.63 16.675 ;
    RECT 349.68 15.885 349.89 15.955 ;
    RECT 349.68 16.245 349.89 16.315 ;
    RECT 349.68 16.605 349.89 16.675 ;
    RECT 349.22 15.885 349.43 15.955 ;
    RECT 349.22 16.245 349.43 16.315 ;
    RECT 349.22 16.605 349.43 16.675 ;
    RECT 213.56 15.885 213.77 15.955 ;
    RECT 213.56 16.245 213.77 16.315 ;
    RECT 213.56 16.605 213.77 16.675 ;
    RECT 213.1 15.885 213.31 15.955 ;
    RECT 213.1 16.245 213.31 16.315 ;
    RECT 213.1 16.605 213.31 16.675 ;
    RECT 346.36 15.885 346.57 15.955 ;
    RECT 346.36 16.245 346.57 16.315 ;
    RECT 346.36 16.605 346.57 16.675 ;
    RECT 345.9 15.885 346.11 15.955 ;
    RECT 345.9 16.245 346.11 16.315 ;
    RECT 345.9 16.605 346.11 16.675 ;
    RECT 210.24 15.885 210.45 15.955 ;
    RECT 210.24 16.245 210.45 16.315 ;
    RECT 210.24 16.605 210.45 16.675 ;
    RECT 209.78 15.885 209.99 15.955 ;
    RECT 209.78 16.245 209.99 16.315 ;
    RECT 209.78 16.605 209.99 16.675 ;
    RECT 343.04 15.885 343.25 15.955 ;
    RECT 343.04 16.245 343.25 16.315 ;
    RECT 343.04 16.605 343.25 16.675 ;
    RECT 342.58 15.885 342.79 15.955 ;
    RECT 342.58 16.245 342.79 16.315 ;
    RECT 342.58 16.605 342.79 16.675 ;
    RECT 206.92 15.885 207.13 15.955 ;
    RECT 206.92 16.245 207.13 16.315 ;
    RECT 206.92 16.605 207.13 16.675 ;
    RECT 206.46 15.885 206.67 15.955 ;
    RECT 206.46 16.245 206.67 16.315 ;
    RECT 206.46 16.605 206.67 16.675 ;
    RECT 339.72 15.885 339.93 15.955 ;
    RECT 339.72 16.245 339.93 16.315 ;
    RECT 339.72 16.605 339.93 16.675 ;
    RECT 339.26 15.885 339.47 15.955 ;
    RECT 339.26 16.245 339.47 16.315 ;
    RECT 339.26 16.605 339.47 16.675 ;
    RECT 203.6 15.885 203.81 15.955 ;
    RECT 203.6 16.245 203.81 16.315 ;
    RECT 203.6 16.605 203.81 16.675 ;
    RECT 203.14 15.885 203.35 15.955 ;
    RECT 203.14 16.245 203.35 16.315 ;
    RECT 203.14 16.605 203.35 16.675 ;
    RECT 336.4 15.885 336.61 15.955 ;
    RECT 336.4 16.245 336.61 16.315 ;
    RECT 336.4 16.605 336.61 16.675 ;
    RECT 335.94 15.885 336.15 15.955 ;
    RECT 335.94 16.245 336.15 16.315 ;
    RECT 335.94 16.605 336.15 16.675 ;
    RECT 266.68 15.885 266.89 15.955 ;
    RECT 266.68 16.245 266.89 16.315 ;
    RECT 266.68 16.605 266.89 16.675 ;
    RECT 266.22 15.885 266.43 15.955 ;
    RECT 266.22 16.245 266.43 16.315 ;
    RECT 266.22 16.605 266.43 16.675 ;
    RECT 263.36 15.885 263.57 15.955 ;
    RECT 263.36 16.245 263.57 16.315 ;
    RECT 263.36 16.605 263.57 16.675 ;
    RECT 262.9 15.885 263.11 15.955 ;
    RECT 262.9 16.245 263.11 16.315 ;
    RECT 262.9 16.605 263.11 16.675 ;
    RECT 260.04 15.885 260.25 15.955 ;
    RECT 260.04 16.245 260.25 16.315 ;
    RECT 260.04 16.605 260.25 16.675 ;
    RECT 259.58 15.885 259.79 15.955 ;
    RECT 259.58 16.245 259.79 16.315 ;
    RECT 259.58 16.605 259.79 16.675 ;
    RECT 256.72 15.885 256.93 15.955 ;
    RECT 256.72 16.245 256.93 16.315 ;
    RECT 256.72 16.605 256.93 16.675 ;
    RECT 256.26 15.885 256.47 15.955 ;
    RECT 256.26 16.245 256.47 16.315 ;
    RECT 256.26 16.605 256.47 16.675 ;
    RECT 253.4 15.885 253.61 15.955 ;
    RECT 253.4 16.245 253.61 16.315 ;
    RECT 253.4 16.605 253.61 16.675 ;
    RECT 252.94 15.885 253.15 15.955 ;
    RECT 252.94 16.245 253.15 16.315 ;
    RECT 252.94 16.605 253.15 16.675 ;
    RECT 250.08 15.885 250.29 15.955 ;
    RECT 250.08 16.245 250.29 16.315 ;
    RECT 250.08 16.605 250.29 16.675 ;
    RECT 249.62 15.885 249.83 15.955 ;
    RECT 249.62 16.245 249.83 16.315 ;
    RECT 249.62 16.605 249.83 16.675 ;
    RECT 246.76 15.885 246.97 15.955 ;
    RECT 246.76 16.245 246.97 16.315 ;
    RECT 246.76 16.605 246.97 16.675 ;
    RECT 246.3 15.885 246.51 15.955 ;
    RECT 246.3 16.245 246.51 16.315 ;
    RECT 246.3 16.605 246.51 16.675 ;
    RECT 243.44 15.885 243.65 15.955 ;
    RECT 243.44 16.245 243.65 16.315 ;
    RECT 243.44 16.605 243.65 16.675 ;
    RECT 242.98 15.885 243.19 15.955 ;
    RECT 242.98 16.245 243.19 16.315 ;
    RECT 242.98 16.605 243.19 16.675 ;
    RECT 240.12 15.885 240.33 15.955 ;
    RECT 240.12 16.245 240.33 16.315 ;
    RECT 240.12 16.605 240.33 16.675 ;
    RECT 239.66 15.885 239.87 15.955 ;
    RECT 239.66 16.245 239.87 16.315 ;
    RECT 239.66 16.605 239.87 16.675 ;
    RECT 236.8 15.885 237.01 15.955 ;
    RECT 236.8 16.245 237.01 16.315 ;
    RECT 236.8 16.605 237.01 16.675 ;
    RECT 236.34 15.885 236.55 15.955 ;
    RECT 236.34 16.245 236.55 16.315 ;
    RECT 236.34 16.605 236.55 16.675 ;
    RECT 374.15 16.245 374.22 16.315 ;
    RECT 333.08 15.885 333.29 15.955 ;
    RECT 333.08 16.245 333.29 16.315 ;
    RECT 333.08 16.605 333.29 16.675 ;
    RECT 332.62 15.885 332.83 15.955 ;
    RECT 332.62 16.245 332.83 16.315 ;
    RECT 332.62 16.605 332.83 16.675 ;
    RECT 329.76 15.885 329.97 15.955 ;
    RECT 329.76 16.245 329.97 16.315 ;
    RECT 329.76 16.605 329.97 16.675 ;
    RECT 329.3 15.885 329.51 15.955 ;
    RECT 329.3 16.245 329.51 16.315 ;
    RECT 329.3 16.605 329.51 16.675 ;
    RECT 326.44 15.885 326.65 15.955 ;
    RECT 326.44 16.245 326.65 16.315 ;
    RECT 326.44 16.605 326.65 16.675 ;
    RECT 325.98 15.885 326.19 15.955 ;
    RECT 325.98 16.245 326.19 16.315 ;
    RECT 325.98 16.605 326.19 16.675 ;
    RECT 323.12 15.885 323.33 15.955 ;
    RECT 323.12 16.245 323.33 16.315 ;
    RECT 323.12 16.605 323.33 16.675 ;
    RECT 322.66 15.885 322.87 15.955 ;
    RECT 322.66 16.245 322.87 16.315 ;
    RECT 322.66 16.605 322.87 16.675 ;
    RECT 319.8 15.885 320.01 15.955 ;
    RECT 319.8 16.245 320.01 16.315 ;
    RECT 319.8 16.605 320.01 16.675 ;
    RECT 319.34 15.885 319.55 15.955 ;
    RECT 319.34 16.245 319.55 16.315 ;
    RECT 319.34 16.605 319.55 16.675 ;
    RECT 316.48 15.885 316.69 15.955 ;
    RECT 316.48 16.245 316.69 16.315 ;
    RECT 316.48 16.605 316.69 16.675 ;
    RECT 316.02 15.885 316.23 15.955 ;
    RECT 316.02 16.245 316.23 16.315 ;
    RECT 316.02 16.605 316.23 16.675 ;
    RECT 313.16 15.885 313.37 15.955 ;
    RECT 313.16 16.245 313.37 16.315 ;
    RECT 313.16 16.605 313.37 16.675 ;
    RECT 312.7 15.885 312.91 15.955 ;
    RECT 312.7 16.245 312.91 16.315 ;
    RECT 312.7 16.605 312.91 16.675 ;
    RECT 309.84 15.885 310.05 15.955 ;
    RECT 309.84 16.245 310.05 16.315 ;
    RECT 309.84 16.605 310.05 16.675 ;
    RECT 309.38 15.885 309.59 15.955 ;
    RECT 309.38 16.245 309.59 16.315 ;
    RECT 309.38 16.605 309.59 16.675 ;
    RECT 306.52 15.885 306.73 15.955 ;
    RECT 306.52 16.245 306.73 16.315 ;
    RECT 306.52 16.605 306.73 16.675 ;
    RECT 306.06 15.885 306.27 15.955 ;
    RECT 306.06 16.245 306.27 16.315 ;
    RECT 306.06 16.605 306.27 16.675 ;
    RECT 303.2 31.725 303.41 31.795 ;
    RECT 303.2 32.085 303.41 32.155 ;
    RECT 303.2 32.445 303.41 32.515 ;
    RECT 302.74 31.725 302.95 31.795 ;
    RECT 302.74 32.085 302.95 32.155 ;
    RECT 302.74 32.445 302.95 32.515 ;
    RECT 372.92 31.725 373.13 31.795 ;
    RECT 372.92 32.085 373.13 32.155 ;
    RECT 372.92 32.445 373.13 32.515 ;
    RECT 372.46 31.725 372.67 31.795 ;
    RECT 372.46 32.085 372.67 32.155 ;
    RECT 372.46 32.445 372.67 32.515 ;
    RECT 369.6 31.725 369.81 31.795 ;
    RECT 369.6 32.085 369.81 32.155 ;
    RECT 369.6 32.445 369.81 32.515 ;
    RECT 369.14 31.725 369.35 31.795 ;
    RECT 369.14 32.085 369.35 32.155 ;
    RECT 369.14 32.445 369.35 32.515 ;
    RECT 200.605 32.085 200.675 32.155 ;
    RECT 299.88 31.725 300.09 31.795 ;
    RECT 299.88 32.085 300.09 32.155 ;
    RECT 299.88 32.445 300.09 32.515 ;
    RECT 299.42 31.725 299.63 31.795 ;
    RECT 299.42 32.085 299.63 32.155 ;
    RECT 299.42 32.445 299.63 32.515 ;
    RECT 296.56 31.725 296.77 31.795 ;
    RECT 296.56 32.085 296.77 32.155 ;
    RECT 296.56 32.445 296.77 32.515 ;
    RECT 296.1 31.725 296.31 31.795 ;
    RECT 296.1 32.085 296.31 32.155 ;
    RECT 296.1 32.445 296.31 32.515 ;
    RECT 293.24 31.725 293.45 31.795 ;
    RECT 293.24 32.085 293.45 32.155 ;
    RECT 293.24 32.445 293.45 32.515 ;
    RECT 292.78 31.725 292.99 31.795 ;
    RECT 292.78 32.085 292.99 32.155 ;
    RECT 292.78 32.445 292.99 32.515 ;
    RECT 289.92 31.725 290.13 31.795 ;
    RECT 289.92 32.085 290.13 32.155 ;
    RECT 289.92 32.445 290.13 32.515 ;
    RECT 289.46 31.725 289.67 31.795 ;
    RECT 289.46 32.085 289.67 32.155 ;
    RECT 289.46 32.445 289.67 32.515 ;
    RECT 286.6 31.725 286.81 31.795 ;
    RECT 286.6 32.085 286.81 32.155 ;
    RECT 286.6 32.445 286.81 32.515 ;
    RECT 286.14 31.725 286.35 31.795 ;
    RECT 286.14 32.085 286.35 32.155 ;
    RECT 286.14 32.445 286.35 32.515 ;
    RECT 283.28 31.725 283.49 31.795 ;
    RECT 283.28 32.085 283.49 32.155 ;
    RECT 283.28 32.445 283.49 32.515 ;
    RECT 282.82 31.725 283.03 31.795 ;
    RECT 282.82 32.085 283.03 32.155 ;
    RECT 282.82 32.445 283.03 32.515 ;
    RECT 279.96 31.725 280.17 31.795 ;
    RECT 279.96 32.085 280.17 32.155 ;
    RECT 279.96 32.445 280.17 32.515 ;
    RECT 279.5 31.725 279.71 31.795 ;
    RECT 279.5 32.085 279.71 32.155 ;
    RECT 279.5 32.445 279.71 32.515 ;
    RECT 276.64 31.725 276.85 31.795 ;
    RECT 276.64 32.085 276.85 32.155 ;
    RECT 276.64 32.445 276.85 32.515 ;
    RECT 276.18 31.725 276.39 31.795 ;
    RECT 276.18 32.085 276.39 32.155 ;
    RECT 276.18 32.445 276.39 32.515 ;
    RECT 273.32 31.725 273.53 31.795 ;
    RECT 273.32 32.085 273.53 32.155 ;
    RECT 273.32 32.445 273.53 32.515 ;
    RECT 272.86 31.725 273.07 31.795 ;
    RECT 272.86 32.085 273.07 32.155 ;
    RECT 272.86 32.445 273.07 32.515 ;
    RECT 270.0 31.725 270.21 31.795 ;
    RECT 270.0 32.085 270.21 32.155 ;
    RECT 270.0 32.445 270.21 32.515 ;
    RECT 269.54 31.725 269.75 31.795 ;
    RECT 269.54 32.085 269.75 32.155 ;
    RECT 269.54 32.445 269.75 32.515 ;
    RECT 233.48 31.725 233.69 31.795 ;
    RECT 233.48 32.085 233.69 32.155 ;
    RECT 233.48 32.445 233.69 32.515 ;
    RECT 233.02 31.725 233.23 31.795 ;
    RECT 233.02 32.085 233.23 32.155 ;
    RECT 233.02 32.445 233.23 32.515 ;
    RECT 230.16 31.725 230.37 31.795 ;
    RECT 230.16 32.085 230.37 32.155 ;
    RECT 230.16 32.445 230.37 32.515 ;
    RECT 229.7 31.725 229.91 31.795 ;
    RECT 229.7 32.085 229.91 32.155 ;
    RECT 229.7 32.445 229.91 32.515 ;
    RECT 366.28 31.725 366.49 31.795 ;
    RECT 366.28 32.085 366.49 32.155 ;
    RECT 366.28 32.445 366.49 32.515 ;
    RECT 365.82 31.725 366.03 31.795 ;
    RECT 365.82 32.085 366.03 32.155 ;
    RECT 365.82 32.445 366.03 32.515 ;
    RECT 226.84 31.725 227.05 31.795 ;
    RECT 226.84 32.085 227.05 32.155 ;
    RECT 226.84 32.445 227.05 32.515 ;
    RECT 226.38 31.725 226.59 31.795 ;
    RECT 226.38 32.085 226.59 32.155 ;
    RECT 226.38 32.445 226.59 32.515 ;
    RECT 362.96 31.725 363.17 31.795 ;
    RECT 362.96 32.085 363.17 32.155 ;
    RECT 362.96 32.445 363.17 32.515 ;
    RECT 362.5 31.725 362.71 31.795 ;
    RECT 362.5 32.085 362.71 32.155 ;
    RECT 362.5 32.445 362.71 32.515 ;
    RECT 223.52 31.725 223.73 31.795 ;
    RECT 223.52 32.085 223.73 32.155 ;
    RECT 223.52 32.445 223.73 32.515 ;
    RECT 223.06 31.725 223.27 31.795 ;
    RECT 223.06 32.085 223.27 32.155 ;
    RECT 223.06 32.445 223.27 32.515 ;
    RECT 359.64 31.725 359.85 31.795 ;
    RECT 359.64 32.085 359.85 32.155 ;
    RECT 359.64 32.445 359.85 32.515 ;
    RECT 359.18 31.725 359.39 31.795 ;
    RECT 359.18 32.085 359.39 32.155 ;
    RECT 359.18 32.445 359.39 32.515 ;
    RECT 220.2 31.725 220.41 31.795 ;
    RECT 220.2 32.085 220.41 32.155 ;
    RECT 220.2 32.445 220.41 32.515 ;
    RECT 219.74 31.725 219.95 31.795 ;
    RECT 219.74 32.085 219.95 32.155 ;
    RECT 219.74 32.445 219.95 32.515 ;
    RECT 356.32 31.725 356.53 31.795 ;
    RECT 356.32 32.085 356.53 32.155 ;
    RECT 356.32 32.445 356.53 32.515 ;
    RECT 355.86 31.725 356.07 31.795 ;
    RECT 355.86 32.085 356.07 32.155 ;
    RECT 355.86 32.445 356.07 32.515 ;
    RECT 353.0 31.725 353.21 31.795 ;
    RECT 353.0 32.085 353.21 32.155 ;
    RECT 353.0 32.445 353.21 32.515 ;
    RECT 352.54 31.725 352.75 31.795 ;
    RECT 352.54 32.085 352.75 32.155 ;
    RECT 352.54 32.445 352.75 32.515 ;
    RECT 216.88 31.725 217.09 31.795 ;
    RECT 216.88 32.085 217.09 32.155 ;
    RECT 216.88 32.445 217.09 32.515 ;
    RECT 216.42 31.725 216.63 31.795 ;
    RECT 216.42 32.085 216.63 32.155 ;
    RECT 216.42 32.445 216.63 32.515 ;
    RECT 349.68 31.725 349.89 31.795 ;
    RECT 349.68 32.085 349.89 32.155 ;
    RECT 349.68 32.445 349.89 32.515 ;
    RECT 349.22 31.725 349.43 31.795 ;
    RECT 349.22 32.085 349.43 32.155 ;
    RECT 349.22 32.445 349.43 32.515 ;
    RECT 213.56 31.725 213.77 31.795 ;
    RECT 213.56 32.085 213.77 32.155 ;
    RECT 213.56 32.445 213.77 32.515 ;
    RECT 213.1 31.725 213.31 31.795 ;
    RECT 213.1 32.085 213.31 32.155 ;
    RECT 213.1 32.445 213.31 32.515 ;
    RECT 346.36 31.725 346.57 31.795 ;
    RECT 346.36 32.085 346.57 32.155 ;
    RECT 346.36 32.445 346.57 32.515 ;
    RECT 345.9 31.725 346.11 31.795 ;
    RECT 345.9 32.085 346.11 32.155 ;
    RECT 345.9 32.445 346.11 32.515 ;
    RECT 210.24 31.725 210.45 31.795 ;
    RECT 210.24 32.085 210.45 32.155 ;
    RECT 210.24 32.445 210.45 32.515 ;
    RECT 209.78 31.725 209.99 31.795 ;
    RECT 209.78 32.085 209.99 32.155 ;
    RECT 209.78 32.445 209.99 32.515 ;
    RECT 343.04 31.725 343.25 31.795 ;
    RECT 343.04 32.085 343.25 32.155 ;
    RECT 343.04 32.445 343.25 32.515 ;
    RECT 342.58 31.725 342.79 31.795 ;
    RECT 342.58 32.085 342.79 32.155 ;
    RECT 342.58 32.445 342.79 32.515 ;
    RECT 206.92 31.725 207.13 31.795 ;
    RECT 206.92 32.085 207.13 32.155 ;
    RECT 206.92 32.445 207.13 32.515 ;
    RECT 206.46 31.725 206.67 31.795 ;
    RECT 206.46 32.085 206.67 32.155 ;
    RECT 206.46 32.445 206.67 32.515 ;
    RECT 339.72 31.725 339.93 31.795 ;
    RECT 339.72 32.085 339.93 32.155 ;
    RECT 339.72 32.445 339.93 32.515 ;
    RECT 339.26 31.725 339.47 31.795 ;
    RECT 339.26 32.085 339.47 32.155 ;
    RECT 339.26 32.445 339.47 32.515 ;
    RECT 203.6 31.725 203.81 31.795 ;
    RECT 203.6 32.085 203.81 32.155 ;
    RECT 203.6 32.445 203.81 32.515 ;
    RECT 203.14 31.725 203.35 31.795 ;
    RECT 203.14 32.085 203.35 32.155 ;
    RECT 203.14 32.445 203.35 32.515 ;
    RECT 336.4 31.725 336.61 31.795 ;
    RECT 336.4 32.085 336.61 32.155 ;
    RECT 336.4 32.445 336.61 32.515 ;
    RECT 335.94 31.725 336.15 31.795 ;
    RECT 335.94 32.085 336.15 32.155 ;
    RECT 335.94 32.445 336.15 32.515 ;
    RECT 266.68 31.725 266.89 31.795 ;
    RECT 266.68 32.085 266.89 32.155 ;
    RECT 266.68 32.445 266.89 32.515 ;
    RECT 266.22 31.725 266.43 31.795 ;
    RECT 266.22 32.085 266.43 32.155 ;
    RECT 266.22 32.445 266.43 32.515 ;
    RECT 263.36 31.725 263.57 31.795 ;
    RECT 263.36 32.085 263.57 32.155 ;
    RECT 263.36 32.445 263.57 32.515 ;
    RECT 262.9 31.725 263.11 31.795 ;
    RECT 262.9 32.085 263.11 32.155 ;
    RECT 262.9 32.445 263.11 32.515 ;
    RECT 260.04 31.725 260.25 31.795 ;
    RECT 260.04 32.085 260.25 32.155 ;
    RECT 260.04 32.445 260.25 32.515 ;
    RECT 259.58 31.725 259.79 31.795 ;
    RECT 259.58 32.085 259.79 32.155 ;
    RECT 259.58 32.445 259.79 32.515 ;
    RECT 256.72 31.725 256.93 31.795 ;
    RECT 256.72 32.085 256.93 32.155 ;
    RECT 256.72 32.445 256.93 32.515 ;
    RECT 256.26 31.725 256.47 31.795 ;
    RECT 256.26 32.085 256.47 32.155 ;
    RECT 256.26 32.445 256.47 32.515 ;
    RECT 253.4 31.725 253.61 31.795 ;
    RECT 253.4 32.085 253.61 32.155 ;
    RECT 253.4 32.445 253.61 32.515 ;
    RECT 252.94 31.725 253.15 31.795 ;
    RECT 252.94 32.085 253.15 32.155 ;
    RECT 252.94 32.445 253.15 32.515 ;
    RECT 250.08 31.725 250.29 31.795 ;
    RECT 250.08 32.085 250.29 32.155 ;
    RECT 250.08 32.445 250.29 32.515 ;
    RECT 249.62 31.725 249.83 31.795 ;
    RECT 249.62 32.085 249.83 32.155 ;
    RECT 249.62 32.445 249.83 32.515 ;
    RECT 246.76 31.725 246.97 31.795 ;
    RECT 246.76 32.085 246.97 32.155 ;
    RECT 246.76 32.445 246.97 32.515 ;
    RECT 246.3 31.725 246.51 31.795 ;
    RECT 246.3 32.085 246.51 32.155 ;
    RECT 246.3 32.445 246.51 32.515 ;
    RECT 243.44 31.725 243.65 31.795 ;
    RECT 243.44 32.085 243.65 32.155 ;
    RECT 243.44 32.445 243.65 32.515 ;
    RECT 242.98 31.725 243.19 31.795 ;
    RECT 242.98 32.085 243.19 32.155 ;
    RECT 242.98 32.445 243.19 32.515 ;
    RECT 240.12 31.725 240.33 31.795 ;
    RECT 240.12 32.085 240.33 32.155 ;
    RECT 240.12 32.445 240.33 32.515 ;
    RECT 239.66 31.725 239.87 31.795 ;
    RECT 239.66 32.085 239.87 32.155 ;
    RECT 239.66 32.445 239.87 32.515 ;
    RECT 236.8 31.725 237.01 31.795 ;
    RECT 236.8 32.085 237.01 32.155 ;
    RECT 236.8 32.445 237.01 32.515 ;
    RECT 236.34 31.725 236.55 31.795 ;
    RECT 236.34 32.085 236.55 32.155 ;
    RECT 236.34 32.445 236.55 32.515 ;
    RECT 374.15 32.085 374.22 32.155 ;
    RECT 333.08 31.725 333.29 31.795 ;
    RECT 333.08 32.085 333.29 32.155 ;
    RECT 333.08 32.445 333.29 32.515 ;
    RECT 332.62 31.725 332.83 31.795 ;
    RECT 332.62 32.085 332.83 32.155 ;
    RECT 332.62 32.445 332.83 32.515 ;
    RECT 329.76 31.725 329.97 31.795 ;
    RECT 329.76 32.085 329.97 32.155 ;
    RECT 329.76 32.445 329.97 32.515 ;
    RECT 329.3 31.725 329.51 31.795 ;
    RECT 329.3 32.085 329.51 32.155 ;
    RECT 329.3 32.445 329.51 32.515 ;
    RECT 326.44 31.725 326.65 31.795 ;
    RECT 326.44 32.085 326.65 32.155 ;
    RECT 326.44 32.445 326.65 32.515 ;
    RECT 325.98 31.725 326.19 31.795 ;
    RECT 325.98 32.085 326.19 32.155 ;
    RECT 325.98 32.445 326.19 32.515 ;
    RECT 323.12 31.725 323.33 31.795 ;
    RECT 323.12 32.085 323.33 32.155 ;
    RECT 323.12 32.445 323.33 32.515 ;
    RECT 322.66 31.725 322.87 31.795 ;
    RECT 322.66 32.085 322.87 32.155 ;
    RECT 322.66 32.445 322.87 32.515 ;
    RECT 319.8 31.725 320.01 31.795 ;
    RECT 319.8 32.085 320.01 32.155 ;
    RECT 319.8 32.445 320.01 32.515 ;
    RECT 319.34 31.725 319.55 31.795 ;
    RECT 319.34 32.085 319.55 32.155 ;
    RECT 319.34 32.445 319.55 32.515 ;
    RECT 316.48 31.725 316.69 31.795 ;
    RECT 316.48 32.085 316.69 32.155 ;
    RECT 316.48 32.445 316.69 32.515 ;
    RECT 316.02 31.725 316.23 31.795 ;
    RECT 316.02 32.085 316.23 32.155 ;
    RECT 316.02 32.445 316.23 32.515 ;
    RECT 313.16 31.725 313.37 31.795 ;
    RECT 313.16 32.085 313.37 32.155 ;
    RECT 313.16 32.445 313.37 32.515 ;
    RECT 312.7 31.725 312.91 31.795 ;
    RECT 312.7 32.085 312.91 32.155 ;
    RECT 312.7 32.445 312.91 32.515 ;
    RECT 309.84 31.725 310.05 31.795 ;
    RECT 309.84 32.085 310.05 32.155 ;
    RECT 309.84 32.445 310.05 32.515 ;
    RECT 309.38 31.725 309.59 31.795 ;
    RECT 309.38 32.085 309.59 32.155 ;
    RECT 309.38 32.445 309.59 32.515 ;
    RECT 306.52 31.725 306.73 31.795 ;
    RECT 306.52 32.085 306.73 32.155 ;
    RECT 306.52 32.445 306.73 32.515 ;
    RECT 306.06 31.725 306.27 31.795 ;
    RECT 306.06 32.085 306.27 32.155 ;
    RECT 306.06 32.445 306.27 32.515 ;
    RECT 303.2 15.165 303.41 15.235 ;
    RECT 303.2 15.525 303.41 15.595 ;
    RECT 303.2 15.885 303.41 15.955 ;
    RECT 302.74 15.165 302.95 15.235 ;
    RECT 302.74 15.525 302.95 15.595 ;
    RECT 302.74 15.885 302.95 15.955 ;
    RECT 372.92 15.165 373.13 15.235 ;
    RECT 372.92 15.525 373.13 15.595 ;
    RECT 372.92 15.885 373.13 15.955 ;
    RECT 372.46 15.165 372.67 15.235 ;
    RECT 372.46 15.525 372.67 15.595 ;
    RECT 372.46 15.885 372.67 15.955 ;
    RECT 369.6 15.165 369.81 15.235 ;
    RECT 369.6 15.525 369.81 15.595 ;
    RECT 369.6 15.885 369.81 15.955 ;
    RECT 369.14 15.165 369.35 15.235 ;
    RECT 369.14 15.525 369.35 15.595 ;
    RECT 369.14 15.885 369.35 15.955 ;
    RECT 200.605 15.525 200.675 15.595 ;
    RECT 299.88 15.165 300.09 15.235 ;
    RECT 299.88 15.525 300.09 15.595 ;
    RECT 299.88 15.885 300.09 15.955 ;
    RECT 299.42 15.165 299.63 15.235 ;
    RECT 299.42 15.525 299.63 15.595 ;
    RECT 299.42 15.885 299.63 15.955 ;
    RECT 296.56 15.165 296.77 15.235 ;
    RECT 296.56 15.525 296.77 15.595 ;
    RECT 296.56 15.885 296.77 15.955 ;
    RECT 296.1 15.165 296.31 15.235 ;
    RECT 296.1 15.525 296.31 15.595 ;
    RECT 296.1 15.885 296.31 15.955 ;
    RECT 293.24 15.165 293.45 15.235 ;
    RECT 293.24 15.525 293.45 15.595 ;
    RECT 293.24 15.885 293.45 15.955 ;
    RECT 292.78 15.165 292.99 15.235 ;
    RECT 292.78 15.525 292.99 15.595 ;
    RECT 292.78 15.885 292.99 15.955 ;
    RECT 289.92 15.165 290.13 15.235 ;
    RECT 289.92 15.525 290.13 15.595 ;
    RECT 289.92 15.885 290.13 15.955 ;
    RECT 289.46 15.165 289.67 15.235 ;
    RECT 289.46 15.525 289.67 15.595 ;
    RECT 289.46 15.885 289.67 15.955 ;
    RECT 286.6 15.165 286.81 15.235 ;
    RECT 286.6 15.525 286.81 15.595 ;
    RECT 286.6 15.885 286.81 15.955 ;
    RECT 286.14 15.165 286.35 15.235 ;
    RECT 286.14 15.525 286.35 15.595 ;
    RECT 286.14 15.885 286.35 15.955 ;
    RECT 283.28 15.165 283.49 15.235 ;
    RECT 283.28 15.525 283.49 15.595 ;
    RECT 283.28 15.885 283.49 15.955 ;
    RECT 282.82 15.165 283.03 15.235 ;
    RECT 282.82 15.525 283.03 15.595 ;
    RECT 282.82 15.885 283.03 15.955 ;
    RECT 279.96 15.165 280.17 15.235 ;
    RECT 279.96 15.525 280.17 15.595 ;
    RECT 279.96 15.885 280.17 15.955 ;
    RECT 279.5 15.165 279.71 15.235 ;
    RECT 279.5 15.525 279.71 15.595 ;
    RECT 279.5 15.885 279.71 15.955 ;
    RECT 276.64 15.165 276.85 15.235 ;
    RECT 276.64 15.525 276.85 15.595 ;
    RECT 276.64 15.885 276.85 15.955 ;
    RECT 276.18 15.165 276.39 15.235 ;
    RECT 276.18 15.525 276.39 15.595 ;
    RECT 276.18 15.885 276.39 15.955 ;
    RECT 273.32 15.165 273.53 15.235 ;
    RECT 273.32 15.525 273.53 15.595 ;
    RECT 273.32 15.885 273.53 15.955 ;
    RECT 272.86 15.165 273.07 15.235 ;
    RECT 272.86 15.525 273.07 15.595 ;
    RECT 272.86 15.885 273.07 15.955 ;
    RECT 270.0 15.165 270.21 15.235 ;
    RECT 270.0 15.525 270.21 15.595 ;
    RECT 270.0 15.885 270.21 15.955 ;
    RECT 269.54 15.165 269.75 15.235 ;
    RECT 269.54 15.525 269.75 15.595 ;
    RECT 269.54 15.885 269.75 15.955 ;
    RECT 233.48 15.165 233.69 15.235 ;
    RECT 233.48 15.525 233.69 15.595 ;
    RECT 233.48 15.885 233.69 15.955 ;
    RECT 233.02 15.165 233.23 15.235 ;
    RECT 233.02 15.525 233.23 15.595 ;
    RECT 233.02 15.885 233.23 15.955 ;
    RECT 230.16 15.165 230.37 15.235 ;
    RECT 230.16 15.525 230.37 15.595 ;
    RECT 230.16 15.885 230.37 15.955 ;
    RECT 229.7 15.165 229.91 15.235 ;
    RECT 229.7 15.525 229.91 15.595 ;
    RECT 229.7 15.885 229.91 15.955 ;
    RECT 366.28 15.165 366.49 15.235 ;
    RECT 366.28 15.525 366.49 15.595 ;
    RECT 366.28 15.885 366.49 15.955 ;
    RECT 365.82 15.165 366.03 15.235 ;
    RECT 365.82 15.525 366.03 15.595 ;
    RECT 365.82 15.885 366.03 15.955 ;
    RECT 226.84 15.165 227.05 15.235 ;
    RECT 226.84 15.525 227.05 15.595 ;
    RECT 226.84 15.885 227.05 15.955 ;
    RECT 226.38 15.165 226.59 15.235 ;
    RECT 226.38 15.525 226.59 15.595 ;
    RECT 226.38 15.885 226.59 15.955 ;
    RECT 362.96 15.165 363.17 15.235 ;
    RECT 362.96 15.525 363.17 15.595 ;
    RECT 362.96 15.885 363.17 15.955 ;
    RECT 362.5 15.165 362.71 15.235 ;
    RECT 362.5 15.525 362.71 15.595 ;
    RECT 362.5 15.885 362.71 15.955 ;
    RECT 223.52 15.165 223.73 15.235 ;
    RECT 223.52 15.525 223.73 15.595 ;
    RECT 223.52 15.885 223.73 15.955 ;
    RECT 223.06 15.165 223.27 15.235 ;
    RECT 223.06 15.525 223.27 15.595 ;
    RECT 223.06 15.885 223.27 15.955 ;
    RECT 359.64 15.165 359.85 15.235 ;
    RECT 359.64 15.525 359.85 15.595 ;
    RECT 359.64 15.885 359.85 15.955 ;
    RECT 359.18 15.165 359.39 15.235 ;
    RECT 359.18 15.525 359.39 15.595 ;
    RECT 359.18 15.885 359.39 15.955 ;
    RECT 220.2 15.165 220.41 15.235 ;
    RECT 220.2 15.525 220.41 15.595 ;
    RECT 220.2 15.885 220.41 15.955 ;
    RECT 219.74 15.165 219.95 15.235 ;
    RECT 219.74 15.525 219.95 15.595 ;
    RECT 219.74 15.885 219.95 15.955 ;
    RECT 356.32 15.165 356.53 15.235 ;
    RECT 356.32 15.525 356.53 15.595 ;
    RECT 356.32 15.885 356.53 15.955 ;
    RECT 355.86 15.165 356.07 15.235 ;
    RECT 355.86 15.525 356.07 15.595 ;
    RECT 355.86 15.885 356.07 15.955 ;
    RECT 353.0 15.165 353.21 15.235 ;
    RECT 353.0 15.525 353.21 15.595 ;
    RECT 353.0 15.885 353.21 15.955 ;
    RECT 352.54 15.165 352.75 15.235 ;
    RECT 352.54 15.525 352.75 15.595 ;
    RECT 352.54 15.885 352.75 15.955 ;
    RECT 216.88 15.165 217.09 15.235 ;
    RECT 216.88 15.525 217.09 15.595 ;
    RECT 216.88 15.885 217.09 15.955 ;
    RECT 216.42 15.165 216.63 15.235 ;
    RECT 216.42 15.525 216.63 15.595 ;
    RECT 216.42 15.885 216.63 15.955 ;
    RECT 349.68 15.165 349.89 15.235 ;
    RECT 349.68 15.525 349.89 15.595 ;
    RECT 349.68 15.885 349.89 15.955 ;
    RECT 349.22 15.165 349.43 15.235 ;
    RECT 349.22 15.525 349.43 15.595 ;
    RECT 349.22 15.885 349.43 15.955 ;
    RECT 213.56 15.165 213.77 15.235 ;
    RECT 213.56 15.525 213.77 15.595 ;
    RECT 213.56 15.885 213.77 15.955 ;
    RECT 213.1 15.165 213.31 15.235 ;
    RECT 213.1 15.525 213.31 15.595 ;
    RECT 213.1 15.885 213.31 15.955 ;
    RECT 346.36 15.165 346.57 15.235 ;
    RECT 346.36 15.525 346.57 15.595 ;
    RECT 346.36 15.885 346.57 15.955 ;
    RECT 345.9 15.165 346.11 15.235 ;
    RECT 345.9 15.525 346.11 15.595 ;
    RECT 345.9 15.885 346.11 15.955 ;
    RECT 210.24 15.165 210.45 15.235 ;
    RECT 210.24 15.525 210.45 15.595 ;
    RECT 210.24 15.885 210.45 15.955 ;
    RECT 209.78 15.165 209.99 15.235 ;
    RECT 209.78 15.525 209.99 15.595 ;
    RECT 209.78 15.885 209.99 15.955 ;
    RECT 343.04 15.165 343.25 15.235 ;
    RECT 343.04 15.525 343.25 15.595 ;
    RECT 343.04 15.885 343.25 15.955 ;
    RECT 342.58 15.165 342.79 15.235 ;
    RECT 342.58 15.525 342.79 15.595 ;
    RECT 342.58 15.885 342.79 15.955 ;
    RECT 206.92 15.165 207.13 15.235 ;
    RECT 206.92 15.525 207.13 15.595 ;
    RECT 206.92 15.885 207.13 15.955 ;
    RECT 206.46 15.165 206.67 15.235 ;
    RECT 206.46 15.525 206.67 15.595 ;
    RECT 206.46 15.885 206.67 15.955 ;
    RECT 339.72 15.165 339.93 15.235 ;
    RECT 339.72 15.525 339.93 15.595 ;
    RECT 339.72 15.885 339.93 15.955 ;
    RECT 339.26 15.165 339.47 15.235 ;
    RECT 339.26 15.525 339.47 15.595 ;
    RECT 339.26 15.885 339.47 15.955 ;
    RECT 203.6 15.165 203.81 15.235 ;
    RECT 203.6 15.525 203.81 15.595 ;
    RECT 203.6 15.885 203.81 15.955 ;
    RECT 203.14 15.165 203.35 15.235 ;
    RECT 203.14 15.525 203.35 15.595 ;
    RECT 203.14 15.885 203.35 15.955 ;
    RECT 336.4 15.165 336.61 15.235 ;
    RECT 336.4 15.525 336.61 15.595 ;
    RECT 336.4 15.885 336.61 15.955 ;
    RECT 335.94 15.165 336.15 15.235 ;
    RECT 335.94 15.525 336.15 15.595 ;
    RECT 335.94 15.885 336.15 15.955 ;
    RECT 266.68 15.165 266.89 15.235 ;
    RECT 266.68 15.525 266.89 15.595 ;
    RECT 266.68 15.885 266.89 15.955 ;
    RECT 266.22 15.165 266.43 15.235 ;
    RECT 266.22 15.525 266.43 15.595 ;
    RECT 266.22 15.885 266.43 15.955 ;
    RECT 263.36 15.165 263.57 15.235 ;
    RECT 263.36 15.525 263.57 15.595 ;
    RECT 263.36 15.885 263.57 15.955 ;
    RECT 262.9 15.165 263.11 15.235 ;
    RECT 262.9 15.525 263.11 15.595 ;
    RECT 262.9 15.885 263.11 15.955 ;
    RECT 260.04 15.165 260.25 15.235 ;
    RECT 260.04 15.525 260.25 15.595 ;
    RECT 260.04 15.885 260.25 15.955 ;
    RECT 259.58 15.165 259.79 15.235 ;
    RECT 259.58 15.525 259.79 15.595 ;
    RECT 259.58 15.885 259.79 15.955 ;
    RECT 256.72 15.165 256.93 15.235 ;
    RECT 256.72 15.525 256.93 15.595 ;
    RECT 256.72 15.885 256.93 15.955 ;
    RECT 256.26 15.165 256.47 15.235 ;
    RECT 256.26 15.525 256.47 15.595 ;
    RECT 256.26 15.885 256.47 15.955 ;
    RECT 253.4 15.165 253.61 15.235 ;
    RECT 253.4 15.525 253.61 15.595 ;
    RECT 253.4 15.885 253.61 15.955 ;
    RECT 252.94 15.165 253.15 15.235 ;
    RECT 252.94 15.525 253.15 15.595 ;
    RECT 252.94 15.885 253.15 15.955 ;
    RECT 250.08 15.165 250.29 15.235 ;
    RECT 250.08 15.525 250.29 15.595 ;
    RECT 250.08 15.885 250.29 15.955 ;
    RECT 249.62 15.165 249.83 15.235 ;
    RECT 249.62 15.525 249.83 15.595 ;
    RECT 249.62 15.885 249.83 15.955 ;
    RECT 246.76 15.165 246.97 15.235 ;
    RECT 246.76 15.525 246.97 15.595 ;
    RECT 246.76 15.885 246.97 15.955 ;
    RECT 246.3 15.165 246.51 15.235 ;
    RECT 246.3 15.525 246.51 15.595 ;
    RECT 246.3 15.885 246.51 15.955 ;
    RECT 243.44 15.165 243.65 15.235 ;
    RECT 243.44 15.525 243.65 15.595 ;
    RECT 243.44 15.885 243.65 15.955 ;
    RECT 242.98 15.165 243.19 15.235 ;
    RECT 242.98 15.525 243.19 15.595 ;
    RECT 242.98 15.885 243.19 15.955 ;
    RECT 240.12 15.165 240.33 15.235 ;
    RECT 240.12 15.525 240.33 15.595 ;
    RECT 240.12 15.885 240.33 15.955 ;
    RECT 239.66 15.165 239.87 15.235 ;
    RECT 239.66 15.525 239.87 15.595 ;
    RECT 239.66 15.885 239.87 15.955 ;
    RECT 236.8 15.165 237.01 15.235 ;
    RECT 236.8 15.525 237.01 15.595 ;
    RECT 236.8 15.885 237.01 15.955 ;
    RECT 236.34 15.165 236.55 15.235 ;
    RECT 236.34 15.525 236.55 15.595 ;
    RECT 236.34 15.885 236.55 15.955 ;
    RECT 374.15 15.525 374.22 15.595 ;
    RECT 333.08 15.165 333.29 15.235 ;
    RECT 333.08 15.525 333.29 15.595 ;
    RECT 333.08 15.885 333.29 15.955 ;
    RECT 332.62 15.165 332.83 15.235 ;
    RECT 332.62 15.525 332.83 15.595 ;
    RECT 332.62 15.885 332.83 15.955 ;
    RECT 329.76 15.165 329.97 15.235 ;
    RECT 329.76 15.525 329.97 15.595 ;
    RECT 329.76 15.885 329.97 15.955 ;
    RECT 329.3 15.165 329.51 15.235 ;
    RECT 329.3 15.525 329.51 15.595 ;
    RECT 329.3 15.885 329.51 15.955 ;
    RECT 326.44 15.165 326.65 15.235 ;
    RECT 326.44 15.525 326.65 15.595 ;
    RECT 326.44 15.885 326.65 15.955 ;
    RECT 325.98 15.165 326.19 15.235 ;
    RECT 325.98 15.525 326.19 15.595 ;
    RECT 325.98 15.885 326.19 15.955 ;
    RECT 323.12 15.165 323.33 15.235 ;
    RECT 323.12 15.525 323.33 15.595 ;
    RECT 323.12 15.885 323.33 15.955 ;
    RECT 322.66 15.165 322.87 15.235 ;
    RECT 322.66 15.525 322.87 15.595 ;
    RECT 322.66 15.885 322.87 15.955 ;
    RECT 319.8 15.165 320.01 15.235 ;
    RECT 319.8 15.525 320.01 15.595 ;
    RECT 319.8 15.885 320.01 15.955 ;
    RECT 319.34 15.165 319.55 15.235 ;
    RECT 319.34 15.525 319.55 15.595 ;
    RECT 319.34 15.885 319.55 15.955 ;
    RECT 316.48 15.165 316.69 15.235 ;
    RECT 316.48 15.525 316.69 15.595 ;
    RECT 316.48 15.885 316.69 15.955 ;
    RECT 316.02 15.165 316.23 15.235 ;
    RECT 316.02 15.525 316.23 15.595 ;
    RECT 316.02 15.885 316.23 15.955 ;
    RECT 313.16 15.165 313.37 15.235 ;
    RECT 313.16 15.525 313.37 15.595 ;
    RECT 313.16 15.885 313.37 15.955 ;
    RECT 312.7 15.165 312.91 15.235 ;
    RECT 312.7 15.525 312.91 15.595 ;
    RECT 312.7 15.885 312.91 15.955 ;
    RECT 309.84 15.165 310.05 15.235 ;
    RECT 309.84 15.525 310.05 15.595 ;
    RECT 309.84 15.885 310.05 15.955 ;
    RECT 309.38 15.165 309.59 15.235 ;
    RECT 309.38 15.525 309.59 15.595 ;
    RECT 309.38 15.885 309.59 15.955 ;
    RECT 306.52 15.165 306.73 15.235 ;
    RECT 306.52 15.525 306.73 15.595 ;
    RECT 306.52 15.885 306.73 15.955 ;
    RECT 306.06 15.165 306.27 15.235 ;
    RECT 306.06 15.525 306.27 15.595 ;
    RECT 306.06 15.885 306.27 15.955 ;
    RECT 303.2 31.005 303.41 31.075 ;
    RECT 303.2 31.365 303.41 31.435 ;
    RECT 303.2 31.725 303.41 31.795 ;
    RECT 302.74 31.005 302.95 31.075 ;
    RECT 302.74 31.365 302.95 31.435 ;
    RECT 302.74 31.725 302.95 31.795 ;
    RECT 372.92 31.005 373.13 31.075 ;
    RECT 372.92 31.365 373.13 31.435 ;
    RECT 372.92 31.725 373.13 31.795 ;
    RECT 372.46 31.005 372.67 31.075 ;
    RECT 372.46 31.365 372.67 31.435 ;
    RECT 372.46 31.725 372.67 31.795 ;
    RECT 369.6 31.005 369.81 31.075 ;
    RECT 369.6 31.365 369.81 31.435 ;
    RECT 369.6 31.725 369.81 31.795 ;
    RECT 369.14 31.005 369.35 31.075 ;
    RECT 369.14 31.365 369.35 31.435 ;
    RECT 369.14 31.725 369.35 31.795 ;
    RECT 200.605 31.365 200.675 31.435 ;
    RECT 299.88 31.005 300.09 31.075 ;
    RECT 299.88 31.365 300.09 31.435 ;
    RECT 299.88 31.725 300.09 31.795 ;
    RECT 299.42 31.005 299.63 31.075 ;
    RECT 299.42 31.365 299.63 31.435 ;
    RECT 299.42 31.725 299.63 31.795 ;
    RECT 296.56 31.005 296.77 31.075 ;
    RECT 296.56 31.365 296.77 31.435 ;
    RECT 296.56 31.725 296.77 31.795 ;
    RECT 296.1 31.005 296.31 31.075 ;
    RECT 296.1 31.365 296.31 31.435 ;
    RECT 296.1 31.725 296.31 31.795 ;
    RECT 293.24 31.005 293.45 31.075 ;
    RECT 293.24 31.365 293.45 31.435 ;
    RECT 293.24 31.725 293.45 31.795 ;
    RECT 292.78 31.005 292.99 31.075 ;
    RECT 292.78 31.365 292.99 31.435 ;
    RECT 292.78 31.725 292.99 31.795 ;
    RECT 289.92 31.005 290.13 31.075 ;
    RECT 289.92 31.365 290.13 31.435 ;
    RECT 289.92 31.725 290.13 31.795 ;
    RECT 289.46 31.005 289.67 31.075 ;
    RECT 289.46 31.365 289.67 31.435 ;
    RECT 289.46 31.725 289.67 31.795 ;
    RECT 286.6 31.005 286.81 31.075 ;
    RECT 286.6 31.365 286.81 31.435 ;
    RECT 286.6 31.725 286.81 31.795 ;
    RECT 286.14 31.005 286.35 31.075 ;
    RECT 286.14 31.365 286.35 31.435 ;
    RECT 286.14 31.725 286.35 31.795 ;
    RECT 283.28 31.005 283.49 31.075 ;
    RECT 283.28 31.365 283.49 31.435 ;
    RECT 283.28 31.725 283.49 31.795 ;
    RECT 282.82 31.005 283.03 31.075 ;
    RECT 282.82 31.365 283.03 31.435 ;
    RECT 282.82 31.725 283.03 31.795 ;
    RECT 279.96 31.005 280.17 31.075 ;
    RECT 279.96 31.365 280.17 31.435 ;
    RECT 279.96 31.725 280.17 31.795 ;
    RECT 279.5 31.005 279.71 31.075 ;
    RECT 279.5 31.365 279.71 31.435 ;
    RECT 279.5 31.725 279.71 31.795 ;
    RECT 276.64 31.005 276.85 31.075 ;
    RECT 276.64 31.365 276.85 31.435 ;
    RECT 276.64 31.725 276.85 31.795 ;
    RECT 276.18 31.005 276.39 31.075 ;
    RECT 276.18 31.365 276.39 31.435 ;
    RECT 276.18 31.725 276.39 31.795 ;
    RECT 273.32 31.005 273.53 31.075 ;
    RECT 273.32 31.365 273.53 31.435 ;
    RECT 273.32 31.725 273.53 31.795 ;
    RECT 272.86 31.005 273.07 31.075 ;
    RECT 272.86 31.365 273.07 31.435 ;
    RECT 272.86 31.725 273.07 31.795 ;
    RECT 270.0 31.005 270.21 31.075 ;
    RECT 270.0 31.365 270.21 31.435 ;
    RECT 270.0 31.725 270.21 31.795 ;
    RECT 269.54 31.005 269.75 31.075 ;
    RECT 269.54 31.365 269.75 31.435 ;
    RECT 269.54 31.725 269.75 31.795 ;
    RECT 233.48 31.005 233.69 31.075 ;
    RECT 233.48 31.365 233.69 31.435 ;
    RECT 233.48 31.725 233.69 31.795 ;
    RECT 233.02 31.005 233.23 31.075 ;
    RECT 233.02 31.365 233.23 31.435 ;
    RECT 233.02 31.725 233.23 31.795 ;
    RECT 230.16 31.005 230.37 31.075 ;
    RECT 230.16 31.365 230.37 31.435 ;
    RECT 230.16 31.725 230.37 31.795 ;
    RECT 229.7 31.005 229.91 31.075 ;
    RECT 229.7 31.365 229.91 31.435 ;
    RECT 229.7 31.725 229.91 31.795 ;
    RECT 366.28 31.005 366.49 31.075 ;
    RECT 366.28 31.365 366.49 31.435 ;
    RECT 366.28 31.725 366.49 31.795 ;
    RECT 365.82 31.005 366.03 31.075 ;
    RECT 365.82 31.365 366.03 31.435 ;
    RECT 365.82 31.725 366.03 31.795 ;
    RECT 226.84 31.005 227.05 31.075 ;
    RECT 226.84 31.365 227.05 31.435 ;
    RECT 226.84 31.725 227.05 31.795 ;
    RECT 226.38 31.005 226.59 31.075 ;
    RECT 226.38 31.365 226.59 31.435 ;
    RECT 226.38 31.725 226.59 31.795 ;
    RECT 362.96 31.005 363.17 31.075 ;
    RECT 362.96 31.365 363.17 31.435 ;
    RECT 362.96 31.725 363.17 31.795 ;
    RECT 362.5 31.005 362.71 31.075 ;
    RECT 362.5 31.365 362.71 31.435 ;
    RECT 362.5 31.725 362.71 31.795 ;
    RECT 223.52 31.005 223.73 31.075 ;
    RECT 223.52 31.365 223.73 31.435 ;
    RECT 223.52 31.725 223.73 31.795 ;
    RECT 223.06 31.005 223.27 31.075 ;
    RECT 223.06 31.365 223.27 31.435 ;
    RECT 223.06 31.725 223.27 31.795 ;
    RECT 359.64 31.005 359.85 31.075 ;
    RECT 359.64 31.365 359.85 31.435 ;
    RECT 359.64 31.725 359.85 31.795 ;
    RECT 359.18 31.005 359.39 31.075 ;
    RECT 359.18 31.365 359.39 31.435 ;
    RECT 359.18 31.725 359.39 31.795 ;
    RECT 220.2 31.005 220.41 31.075 ;
    RECT 220.2 31.365 220.41 31.435 ;
    RECT 220.2 31.725 220.41 31.795 ;
    RECT 219.74 31.005 219.95 31.075 ;
    RECT 219.74 31.365 219.95 31.435 ;
    RECT 219.74 31.725 219.95 31.795 ;
    RECT 356.32 31.005 356.53 31.075 ;
    RECT 356.32 31.365 356.53 31.435 ;
    RECT 356.32 31.725 356.53 31.795 ;
    RECT 355.86 31.005 356.07 31.075 ;
    RECT 355.86 31.365 356.07 31.435 ;
    RECT 355.86 31.725 356.07 31.795 ;
    RECT 353.0 31.005 353.21 31.075 ;
    RECT 353.0 31.365 353.21 31.435 ;
    RECT 353.0 31.725 353.21 31.795 ;
    RECT 352.54 31.005 352.75 31.075 ;
    RECT 352.54 31.365 352.75 31.435 ;
    RECT 352.54 31.725 352.75 31.795 ;
    RECT 216.88 31.005 217.09 31.075 ;
    RECT 216.88 31.365 217.09 31.435 ;
    RECT 216.88 31.725 217.09 31.795 ;
    RECT 216.42 31.005 216.63 31.075 ;
    RECT 216.42 31.365 216.63 31.435 ;
    RECT 216.42 31.725 216.63 31.795 ;
    RECT 349.68 31.005 349.89 31.075 ;
    RECT 349.68 31.365 349.89 31.435 ;
    RECT 349.68 31.725 349.89 31.795 ;
    RECT 349.22 31.005 349.43 31.075 ;
    RECT 349.22 31.365 349.43 31.435 ;
    RECT 349.22 31.725 349.43 31.795 ;
    RECT 213.56 31.005 213.77 31.075 ;
    RECT 213.56 31.365 213.77 31.435 ;
    RECT 213.56 31.725 213.77 31.795 ;
    RECT 213.1 31.005 213.31 31.075 ;
    RECT 213.1 31.365 213.31 31.435 ;
    RECT 213.1 31.725 213.31 31.795 ;
    RECT 346.36 31.005 346.57 31.075 ;
    RECT 346.36 31.365 346.57 31.435 ;
    RECT 346.36 31.725 346.57 31.795 ;
    RECT 345.9 31.005 346.11 31.075 ;
    RECT 345.9 31.365 346.11 31.435 ;
    RECT 345.9 31.725 346.11 31.795 ;
    RECT 210.24 31.005 210.45 31.075 ;
    RECT 210.24 31.365 210.45 31.435 ;
    RECT 210.24 31.725 210.45 31.795 ;
    RECT 209.78 31.005 209.99 31.075 ;
    RECT 209.78 31.365 209.99 31.435 ;
    RECT 209.78 31.725 209.99 31.795 ;
    RECT 343.04 31.005 343.25 31.075 ;
    RECT 343.04 31.365 343.25 31.435 ;
    RECT 343.04 31.725 343.25 31.795 ;
    RECT 342.58 31.005 342.79 31.075 ;
    RECT 342.58 31.365 342.79 31.435 ;
    RECT 342.58 31.725 342.79 31.795 ;
    RECT 206.92 31.005 207.13 31.075 ;
    RECT 206.92 31.365 207.13 31.435 ;
    RECT 206.92 31.725 207.13 31.795 ;
    RECT 206.46 31.005 206.67 31.075 ;
    RECT 206.46 31.365 206.67 31.435 ;
    RECT 206.46 31.725 206.67 31.795 ;
    RECT 339.72 31.005 339.93 31.075 ;
    RECT 339.72 31.365 339.93 31.435 ;
    RECT 339.72 31.725 339.93 31.795 ;
    RECT 339.26 31.005 339.47 31.075 ;
    RECT 339.26 31.365 339.47 31.435 ;
    RECT 339.26 31.725 339.47 31.795 ;
    RECT 203.6 31.005 203.81 31.075 ;
    RECT 203.6 31.365 203.81 31.435 ;
    RECT 203.6 31.725 203.81 31.795 ;
    RECT 203.14 31.005 203.35 31.075 ;
    RECT 203.14 31.365 203.35 31.435 ;
    RECT 203.14 31.725 203.35 31.795 ;
    RECT 336.4 31.005 336.61 31.075 ;
    RECT 336.4 31.365 336.61 31.435 ;
    RECT 336.4 31.725 336.61 31.795 ;
    RECT 335.94 31.005 336.15 31.075 ;
    RECT 335.94 31.365 336.15 31.435 ;
    RECT 335.94 31.725 336.15 31.795 ;
    RECT 266.68 31.005 266.89 31.075 ;
    RECT 266.68 31.365 266.89 31.435 ;
    RECT 266.68 31.725 266.89 31.795 ;
    RECT 266.22 31.005 266.43 31.075 ;
    RECT 266.22 31.365 266.43 31.435 ;
    RECT 266.22 31.725 266.43 31.795 ;
    RECT 263.36 31.005 263.57 31.075 ;
    RECT 263.36 31.365 263.57 31.435 ;
    RECT 263.36 31.725 263.57 31.795 ;
    RECT 262.9 31.005 263.11 31.075 ;
    RECT 262.9 31.365 263.11 31.435 ;
    RECT 262.9 31.725 263.11 31.795 ;
    RECT 260.04 31.005 260.25 31.075 ;
    RECT 260.04 31.365 260.25 31.435 ;
    RECT 260.04 31.725 260.25 31.795 ;
    RECT 259.58 31.005 259.79 31.075 ;
    RECT 259.58 31.365 259.79 31.435 ;
    RECT 259.58 31.725 259.79 31.795 ;
    RECT 256.72 31.005 256.93 31.075 ;
    RECT 256.72 31.365 256.93 31.435 ;
    RECT 256.72 31.725 256.93 31.795 ;
    RECT 256.26 31.005 256.47 31.075 ;
    RECT 256.26 31.365 256.47 31.435 ;
    RECT 256.26 31.725 256.47 31.795 ;
    RECT 253.4 31.005 253.61 31.075 ;
    RECT 253.4 31.365 253.61 31.435 ;
    RECT 253.4 31.725 253.61 31.795 ;
    RECT 252.94 31.005 253.15 31.075 ;
    RECT 252.94 31.365 253.15 31.435 ;
    RECT 252.94 31.725 253.15 31.795 ;
    RECT 250.08 31.005 250.29 31.075 ;
    RECT 250.08 31.365 250.29 31.435 ;
    RECT 250.08 31.725 250.29 31.795 ;
    RECT 249.62 31.005 249.83 31.075 ;
    RECT 249.62 31.365 249.83 31.435 ;
    RECT 249.62 31.725 249.83 31.795 ;
    RECT 246.76 31.005 246.97 31.075 ;
    RECT 246.76 31.365 246.97 31.435 ;
    RECT 246.76 31.725 246.97 31.795 ;
    RECT 246.3 31.005 246.51 31.075 ;
    RECT 246.3 31.365 246.51 31.435 ;
    RECT 246.3 31.725 246.51 31.795 ;
    RECT 243.44 31.005 243.65 31.075 ;
    RECT 243.44 31.365 243.65 31.435 ;
    RECT 243.44 31.725 243.65 31.795 ;
    RECT 242.98 31.005 243.19 31.075 ;
    RECT 242.98 31.365 243.19 31.435 ;
    RECT 242.98 31.725 243.19 31.795 ;
    RECT 240.12 31.005 240.33 31.075 ;
    RECT 240.12 31.365 240.33 31.435 ;
    RECT 240.12 31.725 240.33 31.795 ;
    RECT 239.66 31.005 239.87 31.075 ;
    RECT 239.66 31.365 239.87 31.435 ;
    RECT 239.66 31.725 239.87 31.795 ;
    RECT 236.8 31.005 237.01 31.075 ;
    RECT 236.8 31.365 237.01 31.435 ;
    RECT 236.8 31.725 237.01 31.795 ;
    RECT 236.34 31.005 236.55 31.075 ;
    RECT 236.34 31.365 236.55 31.435 ;
    RECT 236.34 31.725 236.55 31.795 ;
    RECT 374.15 31.365 374.22 31.435 ;
    RECT 333.08 31.005 333.29 31.075 ;
    RECT 333.08 31.365 333.29 31.435 ;
    RECT 333.08 31.725 333.29 31.795 ;
    RECT 332.62 31.005 332.83 31.075 ;
    RECT 332.62 31.365 332.83 31.435 ;
    RECT 332.62 31.725 332.83 31.795 ;
    RECT 329.76 31.005 329.97 31.075 ;
    RECT 329.76 31.365 329.97 31.435 ;
    RECT 329.76 31.725 329.97 31.795 ;
    RECT 329.3 31.005 329.51 31.075 ;
    RECT 329.3 31.365 329.51 31.435 ;
    RECT 329.3 31.725 329.51 31.795 ;
    RECT 326.44 31.005 326.65 31.075 ;
    RECT 326.44 31.365 326.65 31.435 ;
    RECT 326.44 31.725 326.65 31.795 ;
    RECT 325.98 31.005 326.19 31.075 ;
    RECT 325.98 31.365 326.19 31.435 ;
    RECT 325.98 31.725 326.19 31.795 ;
    RECT 323.12 31.005 323.33 31.075 ;
    RECT 323.12 31.365 323.33 31.435 ;
    RECT 323.12 31.725 323.33 31.795 ;
    RECT 322.66 31.005 322.87 31.075 ;
    RECT 322.66 31.365 322.87 31.435 ;
    RECT 322.66 31.725 322.87 31.795 ;
    RECT 319.8 31.005 320.01 31.075 ;
    RECT 319.8 31.365 320.01 31.435 ;
    RECT 319.8 31.725 320.01 31.795 ;
    RECT 319.34 31.005 319.55 31.075 ;
    RECT 319.34 31.365 319.55 31.435 ;
    RECT 319.34 31.725 319.55 31.795 ;
    RECT 316.48 31.005 316.69 31.075 ;
    RECT 316.48 31.365 316.69 31.435 ;
    RECT 316.48 31.725 316.69 31.795 ;
    RECT 316.02 31.005 316.23 31.075 ;
    RECT 316.02 31.365 316.23 31.435 ;
    RECT 316.02 31.725 316.23 31.795 ;
    RECT 313.16 31.005 313.37 31.075 ;
    RECT 313.16 31.365 313.37 31.435 ;
    RECT 313.16 31.725 313.37 31.795 ;
    RECT 312.7 31.005 312.91 31.075 ;
    RECT 312.7 31.365 312.91 31.435 ;
    RECT 312.7 31.725 312.91 31.795 ;
    RECT 309.84 31.005 310.05 31.075 ;
    RECT 309.84 31.365 310.05 31.435 ;
    RECT 309.84 31.725 310.05 31.795 ;
    RECT 309.38 31.005 309.59 31.075 ;
    RECT 309.38 31.365 309.59 31.435 ;
    RECT 309.38 31.725 309.59 31.795 ;
    RECT 306.52 31.005 306.73 31.075 ;
    RECT 306.52 31.365 306.73 31.435 ;
    RECT 306.52 31.725 306.73 31.795 ;
    RECT 306.06 31.005 306.27 31.075 ;
    RECT 306.06 31.365 306.27 31.435 ;
    RECT 306.06 31.725 306.27 31.795 ;
    RECT 303.2 14.445 303.41 14.515 ;
    RECT 303.2 14.805 303.41 14.875 ;
    RECT 303.2 15.165 303.41 15.235 ;
    RECT 302.74 14.445 302.95 14.515 ;
    RECT 302.74 14.805 302.95 14.875 ;
    RECT 302.74 15.165 302.95 15.235 ;
    RECT 372.92 14.445 373.13 14.515 ;
    RECT 372.92 14.805 373.13 14.875 ;
    RECT 372.92 15.165 373.13 15.235 ;
    RECT 372.46 14.445 372.67 14.515 ;
    RECT 372.46 14.805 372.67 14.875 ;
    RECT 372.46 15.165 372.67 15.235 ;
    RECT 369.6 14.445 369.81 14.515 ;
    RECT 369.6 14.805 369.81 14.875 ;
    RECT 369.6 15.165 369.81 15.235 ;
    RECT 369.14 14.445 369.35 14.515 ;
    RECT 369.14 14.805 369.35 14.875 ;
    RECT 369.14 15.165 369.35 15.235 ;
    RECT 200.605 14.805 200.675 14.875 ;
    RECT 299.88 14.445 300.09 14.515 ;
    RECT 299.88 14.805 300.09 14.875 ;
    RECT 299.88 15.165 300.09 15.235 ;
    RECT 299.42 14.445 299.63 14.515 ;
    RECT 299.42 14.805 299.63 14.875 ;
    RECT 299.42 15.165 299.63 15.235 ;
    RECT 296.56 14.445 296.77 14.515 ;
    RECT 296.56 14.805 296.77 14.875 ;
    RECT 296.56 15.165 296.77 15.235 ;
    RECT 296.1 14.445 296.31 14.515 ;
    RECT 296.1 14.805 296.31 14.875 ;
    RECT 296.1 15.165 296.31 15.235 ;
    RECT 293.24 14.445 293.45 14.515 ;
    RECT 293.24 14.805 293.45 14.875 ;
    RECT 293.24 15.165 293.45 15.235 ;
    RECT 292.78 14.445 292.99 14.515 ;
    RECT 292.78 14.805 292.99 14.875 ;
    RECT 292.78 15.165 292.99 15.235 ;
    RECT 289.92 14.445 290.13 14.515 ;
    RECT 289.92 14.805 290.13 14.875 ;
    RECT 289.92 15.165 290.13 15.235 ;
    RECT 289.46 14.445 289.67 14.515 ;
    RECT 289.46 14.805 289.67 14.875 ;
    RECT 289.46 15.165 289.67 15.235 ;
    RECT 286.6 14.445 286.81 14.515 ;
    RECT 286.6 14.805 286.81 14.875 ;
    RECT 286.6 15.165 286.81 15.235 ;
    RECT 286.14 14.445 286.35 14.515 ;
    RECT 286.14 14.805 286.35 14.875 ;
    RECT 286.14 15.165 286.35 15.235 ;
    RECT 283.28 14.445 283.49 14.515 ;
    RECT 283.28 14.805 283.49 14.875 ;
    RECT 283.28 15.165 283.49 15.235 ;
    RECT 282.82 14.445 283.03 14.515 ;
    RECT 282.82 14.805 283.03 14.875 ;
    RECT 282.82 15.165 283.03 15.235 ;
    RECT 279.96 14.445 280.17 14.515 ;
    RECT 279.96 14.805 280.17 14.875 ;
    RECT 279.96 15.165 280.17 15.235 ;
    RECT 279.5 14.445 279.71 14.515 ;
    RECT 279.5 14.805 279.71 14.875 ;
    RECT 279.5 15.165 279.71 15.235 ;
    RECT 276.64 14.445 276.85 14.515 ;
    RECT 276.64 14.805 276.85 14.875 ;
    RECT 276.64 15.165 276.85 15.235 ;
    RECT 276.18 14.445 276.39 14.515 ;
    RECT 276.18 14.805 276.39 14.875 ;
    RECT 276.18 15.165 276.39 15.235 ;
    RECT 273.32 14.445 273.53 14.515 ;
    RECT 273.32 14.805 273.53 14.875 ;
    RECT 273.32 15.165 273.53 15.235 ;
    RECT 272.86 14.445 273.07 14.515 ;
    RECT 272.86 14.805 273.07 14.875 ;
    RECT 272.86 15.165 273.07 15.235 ;
    RECT 270.0 14.445 270.21 14.515 ;
    RECT 270.0 14.805 270.21 14.875 ;
    RECT 270.0 15.165 270.21 15.235 ;
    RECT 269.54 14.445 269.75 14.515 ;
    RECT 269.54 14.805 269.75 14.875 ;
    RECT 269.54 15.165 269.75 15.235 ;
    RECT 233.48 14.445 233.69 14.515 ;
    RECT 233.48 14.805 233.69 14.875 ;
    RECT 233.48 15.165 233.69 15.235 ;
    RECT 233.02 14.445 233.23 14.515 ;
    RECT 233.02 14.805 233.23 14.875 ;
    RECT 233.02 15.165 233.23 15.235 ;
    RECT 230.16 14.445 230.37 14.515 ;
    RECT 230.16 14.805 230.37 14.875 ;
    RECT 230.16 15.165 230.37 15.235 ;
    RECT 229.7 14.445 229.91 14.515 ;
    RECT 229.7 14.805 229.91 14.875 ;
    RECT 229.7 15.165 229.91 15.235 ;
    RECT 366.28 14.445 366.49 14.515 ;
    RECT 366.28 14.805 366.49 14.875 ;
    RECT 366.28 15.165 366.49 15.235 ;
    RECT 365.82 14.445 366.03 14.515 ;
    RECT 365.82 14.805 366.03 14.875 ;
    RECT 365.82 15.165 366.03 15.235 ;
    RECT 226.84 14.445 227.05 14.515 ;
    RECT 226.84 14.805 227.05 14.875 ;
    RECT 226.84 15.165 227.05 15.235 ;
    RECT 226.38 14.445 226.59 14.515 ;
    RECT 226.38 14.805 226.59 14.875 ;
    RECT 226.38 15.165 226.59 15.235 ;
    RECT 362.96 14.445 363.17 14.515 ;
    RECT 362.96 14.805 363.17 14.875 ;
    RECT 362.96 15.165 363.17 15.235 ;
    RECT 362.5 14.445 362.71 14.515 ;
    RECT 362.5 14.805 362.71 14.875 ;
    RECT 362.5 15.165 362.71 15.235 ;
    RECT 223.52 14.445 223.73 14.515 ;
    RECT 223.52 14.805 223.73 14.875 ;
    RECT 223.52 15.165 223.73 15.235 ;
    RECT 223.06 14.445 223.27 14.515 ;
    RECT 223.06 14.805 223.27 14.875 ;
    RECT 223.06 15.165 223.27 15.235 ;
    RECT 359.64 14.445 359.85 14.515 ;
    RECT 359.64 14.805 359.85 14.875 ;
    RECT 359.64 15.165 359.85 15.235 ;
    RECT 359.18 14.445 359.39 14.515 ;
    RECT 359.18 14.805 359.39 14.875 ;
    RECT 359.18 15.165 359.39 15.235 ;
    RECT 220.2 14.445 220.41 14.515 ;
    RECT 220.2 14.805 220.41 14.875 ;
    RECT 220.2 15.165 220.41 15.235 ;
    RECT 219.74 14.445 219.95 14.515 ;
    RECT 219.74 14.805 219.95 14.875 ;
    RECT 219.74 15.165 219.95 15.235 ;
    RECT 356.32 14.445 356.53 14.515 ;
    RECT 356.32 14.805 356.53 14.875 ;
    RECT 356.32 15.165 356.53 15.235 ;
    RECT 355.86 14.445 356.07 14.515 ;
    RECT 355.86 14.805 356.07 14.875 ;
    RECT 355.86 15.165 356.07 15.235 ;
    RECT 353.0 14.445 353.21 14.515 ;
    RECT 353.0 14.805 353.21 14.875 ;
    RECT 353.0 15.165 353.21 15.235 ;
    RECT 352.54 14.445 352.75 14.515 ;
    RECT 352.54 14.805 352.75 14.875 ;
    RECT 352.54 15.165 352.75 15.235 ;
    RECT 216.88 14.445 217.09 14.515 ;
    RECT 216.88 14.805 217.09 14.875 ;
    RECT 216.88 15.165 217.09 15.235 ;
    RECT 216.42 14.445 216.63 14.515 ;
    RECT 216.42 14.805 216.63 14.875 ;
    RECT 216.42 15.165 216.63 15.235 ;
    RECT 349.68 14.445 349.89 14.515 ;
    RECT 349.68 14.805 349.89 14.875 ;
    RECT 349.68 15.165 349.89 15.235 ;
    RECT 349.22 14.445 349.43 14.515 ;
    RECT 349.22 14.805 349.43 14.875 ;
    RECT 349.22 15.165 349.43 15.235 ;
    RECT 213.56 14.445 213.77 14.515 ;
    RECT 213.56 14.805 213.77 14.875 ;
    RECT 213.56 15.165 213.77 15.235 ;
    RECT 213.1 14.445 213.31 14.515 ;
    RECT 213.1 14.805 213.31 14.875 ;
    RECT 213.1 15.165 213.31 15.235 ;
    RECT 346.36 14.445 346.57 14.515 ;
    RECT 346.36 14.805 346.57 14.875 ;
    RECT 346.36 15.165 346.57 15.235 ;
    RECT 345.9 14.445 346.11 14.515 ;
    RECT 345.9 14.805 346.11 14.875 ;
    RECT 345.9 15.165 346.11 15.235 ;
    RECT 210.24 14.445 210.45 14.515 ;
    RECT 210.24 14.805 210.45 14.875 ;
    RECT 210.24 15.165 210.45 15.235 ;
    RECT 209.78 14.445 209.99 14.515 ;
    RECT 209.78 14.805 209.99 14.875 ;
    RECT 209.78 15.165 209.99 15.235 ;
    RECT 343.04 14.445 343.25 14.515 ;
    RECT 343.04 14.805 343.25 14.875 ;
    RECT 343.04 15.165 343.25 15.235 ;
    RECT 342.58 14.445 342.79 14.515 ;
    RECT 342.58 14.805 342.79 14.875 ;
    RECT 342.58 15.165 342.79 15.235 ;
    RECT 206.92 14.445 207.13 14.515 ;
    RECT 206.92 14.805 207.13 14.875 ;
    RECT 206.92 15.165 207.13 15.235 ;
    RECT 206.46 14.445 206.67 14.515 ;
    RECT 206.46 14.805 206.67 14.875 ;
    RECT 206.46 15.165 206.67 15.235 ;
    RECT 339.72 14.445 339.93 14.515 ;
    RECT 339.72 14.805 339.93 14.875 ;
    RECT 339.72 15.165 339.93 15.235 ;
    RECT 339.26 14.445 339.47 14.515 ;
    RECT 339.26 14.805 339.47 14.875 ;
    RECT 339.26 15.165 339.47 15.235 ;
    RECT 203.6 14.445 203.81 14.515 ;
    RECT 203.6 14.805 203.81 14.875 ;
    RECT 203.6 15.165 203.81 15.235 ;
    RECT 203.14 14.445 203.35 14.515 ;
    RECT 203.14 14.805 203.35 14.875 ;
    RECT 203.14 15.165 203.35 15.235 ;
    RECT 336.4 14.445 336.61 14.515 ;
    RECT 336.4 14.805 336.61 14.875 ;
    RECT 336.4 15.165 336.61 15.235 ;
    RECT 335.94 14.445 336.15 14.515 ;
    RECT 335.94 14.805 336.15 14.875 ;
    RECT 335.94 15.165 336.15 15.235 ;
    RECT 266.68 14.445 266.89 14.515 ;
    RECT 266.68 14.805 266.89 14.875 ;
    RECT 266.68 15.165 266.89 15.235 ;
    RECT 266.22 14.445 266.43 14.515 ;
    RECT 266.22 14.805 266.43 14.875 ;
    RECT 266.22 15.165 266.43 15.235 ;
    RECT 263.36 14.445 263.57 14.515 ;
    RECT 263.36 14.805 263.57 14.875 ;
    RECT 263.36 15.165 263.57 15.235 ;
    RECT 262.9 14.445 263.11 14.515 ;
    RECT 262.9 14.805 263.11 14.875 ;
    RECT 262.9 15.165 263.11 15.235 ;
    RECT 260.04 14.445 260.25 14.515 ;
    RECT 260.04 14.805 260.25 14.875 ;
    RECT 260.04 15.165 260.25 15.235 ;
    RECT 259.58 14.445 259.79 14.515 ;
    RECT 259.58 14.805 259.79 14.875 ;
    RECT 259.58 15.165 259.79 15.235 ;
    RECT 256.72 14.445 256.93 14.515 ;
    RECT 256.72 14.805 256.93 14.875 ;
    RECT 256.72 15.165 256.93 15.235 ;
    RECT 256.26 14.445 256.47 14.515 ;
    RECT 256.26 14.805 256.47 14.875 ;
    RECT 256.26 15.165 256.47 15.235 ;
    RECT 253.4 14.445 253.61 14.515 ;
    RECT 253.4 14.805 253.61 14.875 ;
    RECT 253.4 15.165 253.61 15.235 ;
    RECT 252.94 14.445 253.15 14.515 ;
    RECT 252.94 14.805 253.15 14.875 ;
    RECT 252.94 15.165 253.15 15.235 ;
    RECT 250.08 14.445 250.29 14.515 ;
    RECT 250.08 14.805 250.29 14.875 ;
    RECT 250.08 15.165 250.29 15.235 ;
    RECT 249.62 14.445 249.83 14.515 ;
    RECT 249.62 14.805 249.83 14.875 ;
    RECT 249.62 15.165 249.83 15.235 ;
    RECT 246.76 14.445 246.97 14.515 ;
    RECT 246.76 14.805 246.97 14.875 ;
    RECT 246.76 15.165 246.97 15.235 ;
    RECT 246.3 14.445 246.51 14.515 ;
    RECT 246.3 14.805 246.51 14.875 ;
    RECT 246.3 15.165 246.51 15.235 ;
    RECT 243.44 14.445 243.65 14.515 ;
    RECT 243.44 14.805 243.65 14.875 ;
    RECT 243.44 15.165 243.65 15.235 ;
    RECT 242.98 14.445 243.19 14.515 ;
    RECT 242.98 14.805 243.19 14.875 ;
    RECT 242.98 15.165 243.19 15.235 ;
    RECT 240.12 14.445 240.33 14.515 ;
    RECT 240.12 14.805 240.33 14.875 ;
    RECT 240.12 15.165 240.33 15.235 ;
    RECT 239.66 14.445 239.87 14.515 ;
    RECT 239.66 14.805 239.87 14.875 ;
    RECT 239.66 15.165 239.87 15.235 ;
    RECT 236.8 14.445 237.01 14.515 ;
    RECT 236.8 14.805 237.01 14.875 ;
    RECT 236.8 15.165 237.01 15.235 ;
    RECT 236.34 14.445 236.55 14.515 ;
    RECT 236.34 14.805 236.55 14.875 ;
    RECT 236.34 15.165 236.55 15.235 ;
    RECT 374.15 14.805 374.22 14.875 ;
    RECT 333.08 14.445 333.29 14.515 ;
    RECT 333.08 14.805 333.29 14.875 ;
    RECT 333.08 15.165 333.29 15.235 ;
    RECT 332.62 14.445 332.83 14.515 ;
    RECT 332.62 14.805 332.83 14.875 ;
    RECT 332.62 15.165 332.83 15.235 ;
    RECT 329.76 14.445 329.97 14.515 ;
    RECT 329.76 14.805 329.97 14.875 ;
    RECT 329.76 15.165 329.97 15.235 ;
    RECT 329.3 14.445 329.51 14.515 ;
    RECT 329.3 14.805 329.51 14.875 ;
    RECT 329.3 15.165 329.51 15.235 ;
    RECT 326.44 14.445 326.65 14.515 ;
    RECT 326.44 14.805 326.65 14.875 ;
    RECT 326.44 15.165 326.65 15.235 ;
    RECT 325.98 14.445 326.19 14.515 ;
    RECT 325.98 14.805 326.19 14.875 ;
    RECT 325.98 15.165 326.19 15.235 ;
    RECT 323.12 14.445 323.33 14.515 ;
    RECT 323.12 14.805 323.33 14.875 ;
    RECT 323.12 15.165 323.33 15.235 ;
    RECT 322.66 14.445 322.87 14.515 ;
    RECT 322.66 14.805 322.87 14.875 ;
    RECT 322.66 15.165 322.87 15.235 ;
    RECT 319.8 14.445 320.01 14.515 ;
    RECT 319.8 14.805 320.01 14.875 ;
    RECT 319.8 15.165 320.01 15.235 ;
    RECT 319.34 14.445 319.55 14.515 ;
    RECT 319.34 14.805 319.55 14.875 ;
    RECT 319.34 15.165 319.55 15.235 ;
    RECT 316.48 14.445 316.69 14.515 ;
    RECT 316.48 14.805 316.69 14.875 ;
    RECT 316.48 15.165 316.69 15.235 ;
    RECT 316.02 14.445 316.23 14.515 ;
    RECT 316.02 14.805 316.23 14.875 ;
    RECT 316.02 15.165 316.23 15.235 ;
    RECT 313.16 14.445 313.37 14.515 ;
    RECT 313.16 14.805 313.37 14.875 ;
    RECT 313.16 15.165 313.37 15.235 ;
    RECT 312.7 14.445 312.91 14.515 ;
    RECT 312.7 14.805 312.91 14.875 ;
    RECT 312.7 15.165 312.91 15.235 ;
    RECT 309.84 14.445 310.05 14.515 ;
    RECT 309.84 14.805 310.05 14.875 ;
    RECT 309.84 15.165 310.05 15.235 ;
    RECT 309.38 14.445 309.59 14.515 ;
    RECT 309.38 14.805 309.59 14.875 ;
    RECT 309.38 15.165 309.59 15.235 ;
    RECT 306.52 14.445 306.73 14.515 ;
    RECT 306.52 14.805 306.73 14.875 ;
    RECT 306.52 15.165 306.73 15.235 ;
    RECT 306.06 14.445 306.27 14.515 ;
    RECT 306.06 14.805 306.27 14.875 ;
    RECT 306.06 15.165 306.27 15.235 ;
    RECT 303.2 30.285 303.41 30.355 ;
    RECT 303.2 30.645 303.41 30.715 ;
    RECT 303.2 31.005 303.41 31.075 ;
    RECT 302.74 30.285 302.95 30.355 ;
    RECT 302.74 30.645 302.95 30.715 ;
    RECT 302.74 31.005 302.95 31.075 ;
    RECT 372.92 30.285 373.13 30.355 ;
    RECT 372.92 30.645 373.13 30.715 ;
    RECT 372.92 31.005 373.13 31.075 ;
    RECT 372.46 30.285 372.67 30.355 ;
    RECT 372.46 30.645 372.67 30.715 ;
    RECT 372.46 31.005 372.67 31.075 ;
    RECT 369.6 30.285 369.81 30.355 ;
    RECT 369.6 30.645 369.81 30.715 ;
    RECT 369.6 31.005 369.81 31.075 ;
    RECT 369.14 30.285 369.35 30.355 ;
    RECT 369.14 30.645 369.35 30.715 ;
    RECT 369.14 31.005 369.35 31.075 ;
    RECT 200.605 30.645 200.675 30.715 ;
    RECT 299.88 30.285 300.09 30.355 ;
    RECT 299.88 30.645 300.09 30.715 ;
    RECT 299.88 31.005 300.09 31.075 ;
    RECT 299.42 30.285 299.63 30.355 ;
    RECT 299.42 30.645 299.63 30.715 ;
    RECT 299.42 31.005 299.63 31.075 ;
    RECT 296.56 30.285 296.77 30.355 ;
    RECT 296.56 30.645 296.77 30.715 ;
    RECT 296.56 31.005 296.77 31.075 ;
    RECT 296.1 30.285 296.31 30.355 ;
    RECT 296.1 30.645 296.31 30.715 ;
    RECT 296.1 31.005 296.31 31.075 ;
    RECT 293.24 30.285 293.45 30.355 ;
    RECT 293.24 30.645 293.45 30.715 ;
    RECT 293.24 31.005 293.45 31.075 ;
    RECT 292.78 30.285 292.99 30.355 ;
    RECT 292.78 30.645 292.99 30.715 ;
    RECT 292.78 31.005 292.99 31.075 ;
    RECT 289.92 30.285 290.13 30.355 ;
    RECT 289.92 30.645 290.13 30.715 ;
    RECT 289.92 31.005 290.13 31.075 ;
    RECT 289.46 30.285 289.67 30.355 ;
    RECT 289.46 30.645 289.67 30.715 ;
    RECT 289.46 31.005 289.67 31.075 ;
    RECT 286.6 30.285 286.81 30.355 ;
    RECT 286.6 30.645 286.81 30.715 ;
    RECT 286.6 31.005 286.81 31.075 ;
    RECT 286.14 30.285 286.35 30.355 ;
    RECT 286.14 30.645 286.35 30.715 ;
    RECT 286.14 31.005 286.35 31.075 ;
    RECT 283.28 30.285 283.49 30.355 ;
    RECT 283.28 30.645 283.49 30.715 ;
    RECT 283.28 31.005 283.49 31.075 ;
    RECT 282.82 30.285 283.03 30.355 ;
    RECT 282.82 30.645 283.03 30.715 ;
    RECT 282.82 31.005 283.03 31.075 ;
    RECT 279.96 30.285 280.17 30.355 ;
    RECT 279.96 30.645 280.17 30.715 ;
    RECT 279.96 31.005 280.17 31.075 ;
    RECT 279.5 30.285 279.71 30.355 ;
    RECT 279.5 30.645 279.71 30.715 ;
    RECT 279.5 31.005 279.71 31.075 ;
    RECT 276.64 30.285 276.85 30.355 ;
    RECT 276.64 30.645 276.85 30.715 ;
    RECT 276.64 31.005 276.85 31.075 ;
    RECT 276.18 30.285 276.39 30.355 ;
    RECT 276.18 30.645 276.39 30.715 ;
    RECT 276.18 31.005 276.39 31.075 ;
    RECT 273.32 30.285 273.53 30.355 ;
    RECT 273.32 30.645 273.53 30.715 ;
    RECT 273.32 31.005 273.53 31.075 ;
    RECT 272.86 30.285 273.07 30.355 ;
    RECT 272.86 30.645 273.07 30.715 ;
    RECT 272.86 31.005 273.07 31.075 ;
    RECT 270.0 30.285 270.21 30.355 ;
    RECT 270.0 30.645 270.21 30.715 ;
    RECT 270.0 31.005 270.21 31.075 ;
    RECT 269.54 30.285 269.75 30.355 ;
    RECT 269.54 30.645 269.75 30.715 ;
    RECT 269.54 31.005 269.75 31.075 ;
    RECT 233.48 30.285 233.69 30.355 ;
    RECT 233.48 30.645 233.69 30.715 ;
    RECT 233.48 31.005 233.69 31.075 ;
    RECT 233.02 30.285 233.23 30.355 ;
    RECT 233.02 30.645 233.23 30.715 ;
    RECT 233.02 31.005 233.23 31.075 ;
    RECT 230.16 30.285 230.37 30.355 ;
    RECT 230.16 30.645 230.37 30.715 ;
    RECT 230.16 31.005 230.37 31.075 ;
    RECT 229.7 30.285 229.91 30.355 ;
    RECT 229.7 30.645 229.91 30.715 ;
    RECT 229.7 31.005 229.91 31.075 ;
    RECT 366.28 30.285 366.49 30.355 ;
    RECT 366.28 30.645 366.49 30.715 ;
    RECT 366.28 31.005 366.49 31.075 ;
    RECT 365.82 30.285 366.03 30.355 ;
    RECT 365.82 30.645 366.03 30.715 ;
    RECT 365.82 31.005 366.03 31.075 ;
    RECT 226.84 30.285 227.05 30.355 ;
    RECT 226.84 30.645 227.05 30.715 ;
    RECT 226.84 31.005 227.05 31.075 ;
    RECT 226.38 30.285 226.59 30.355 ;
    RECT 226.38 30.645 226.59 30.715 ;
    RECT 226.38 31.005 226.59 31.075 ;
    RECT 362.96 30.285 363.17 30.355 ;
    RECT 362.96 30.645 363.17 30.715 ;
    RECT 362.96 31.005 363.17 31.075 ;
    RECT 362.5 30.285 362.71 30.355 ;
    RECT 362.5 30.645 362.71 30.715 ;
    RECT 362.5 31.005 362.71 31.075 ;
    RECT 223.52 30.285 223.73 30.355 ;
    RECT 223.52 30.645 223.73 30.715 ;
    RECT 223.52 31.005 223.73 31.075 ;
    RECT 223.06 30.285 223.27 30.355 ;
    RECT 223.06 30.645 223.27 30.715 ;
    RECT 223.06 31.005 223.27 31.075 ;
    RECT 359.64 30.285 359.85 30.355 ;
    RECT 359.64 30.645 359.85 30.715 ;
    RECT 359.64 31.005 359.85 31.075 ;
    RECT 359.18 30.285 359.39 30.355 ;
    RECT 359.18 30.645 359.39 30.715 ;
    RECT 359.18 31.005 359.39 31.075 ;
    RECT 220.2 30.285 220.41 30.355 ;
    RECT 220.2 30.645 220.41 30.715 ;
    RECT 220.2 31.005 220.41 31.075 ;
    RECT 219.74 30.285 219.95 30.355 ;
    RECT 219.74 30.645 219.95 30.715 ;
    RECT 219.74 31.005 219.95 31.075 ;
    RECT 356.32 30.285 356.53 30.355 ;
    RECT 356.32 30.645 356.53 30.715 ;
    RECT 356.32 31.005 356.53 31.075 ;
    RECT 355.86 30.285 356.07 30.355 ;
    RECT 355.86 30.645 356.07 30.715 ;
    RECT 355.86 31.005 356.07 31.075 ;
    RECT 353.0 30.285 353.21 30.355 ;
    RECT 353.0 30.645 353.21 30.715 ;
    RECT 353.0 31.005 353.21 31.075 ;
    RECT 352.54 30.285 352.75 30.355 ;
    RECT 352.54 30.645 352.75 30.715 ;
    RECT 352.54 31.005 352.75 31.075 ;
    RECT 216.88 30.285 217.09 30.355 ;
    RECT 216.88 30.645 217.09 30.715 ;
    RECT 216.88 31.005 217.09 31.075 ;
    RECT 216.42 30.285 216.63 30.355 ;
    RECT 216.42 30.645 216.63 30.715 ;
    RECT 216.42 31.005 216.63 31.075 ;
    RECT 349.68 30.285 349.89 30.355 ;
    RECT 349.68 30.645 349.89 30.715 ;
    RECT 349.68 31.005 349.89 31.075 ;
    RECT 349.22 30.285 349.43 30.355 ;
    RECT 349.22 30.645 349.43 30.715 ;
    RECT 349.22 31.005 349.43 31.075 ;
    RECT 213.56 30.285 213.77 30.355 ;
    RECT 213.56 30.645 213.77 30.715 ;
    RECT 213.56 31.005 213.77 31.075 ;
    RECT 213.1 30.285 213.31 30.355 ;
    RECT 213.1 30.645 213.31 30.715 ;
    RECT 213.1 31.005 213.31 31.075 ;
    RECT 346.36 30.285 346.57 30.355 ;
    RECT 346.36 30.645 346.57 30.715 ;
    RECT 346.36 31.005 346.57 31.075 ;
    RECT 345.9 30.285 346.11 30.355 ;
    RECT 345.9 30.645 346.11 30.715 ;
    RECT 345.9 31.005 346.11 31.075 ;
    RECT 210.24 30.285 210.45 30.355 ;
    RECT 210.24 30.645 210.45 30.715 ;
    RECT 210.24 31.005 210.45 31.075 ;
    RECT 209.78 30.285 209.99 30.355 ;
    RECT 209.78 30.645 209.99 30.715 ;
    RECT 209.78 31.005 209.99 31.075 ;
    RECT 343.04 30.285 343.25 30.355 ;
    RECT 343.04 30.645 343.25 30.715 ;
    RECT 343.04 31.005 343.25 31.075 ;
    RECT 342.58 30.285 342.79 30.355 ;
    RECT 342.58 30.645 342.79 30.715 ;
    RECT 342.58 31.005 342.79 31.075 ;
    RECT 206.92 30.285 207.13 30.355 ;
    RECT 206.92 30.645 207.13 30.715 ;
    RECT 206.92 31.005 207.13 31.075 ;
    RECT 206.46 30.285 206.67 30.355 ;
    RECT 206.46 30.645 206.67 30.715 ;
    RECT 206.46 31.005 206.67 31.075 ;
    RECT 339.72 30.285 339.93 30.355 ;
    RECT 339.72 30.645 339.93 30.715 ;
    RECT 339.72 31.005 339.93 31.075 ;
    RECT 339.26 30.285 339.47 30.355 ;
    RECT 339.26 30.645 339.47 30.715 ;
    RECT 339.26 31.005 339.47 31.075 ;
    RECT 203.6 30.285 203.81 30.355 ;
    RECT 203.6 30.645 203.81 30.715 ;
    RECT 203.6 31.005 203.81 31.075 ;
    RECT 203.14 30.285 203.35 30.355 ;
    RECT 203.14 30.645 203.35 30.715 ;
    RECT 203.14 31.005 203.35 31.075 ;
    RECT 336.4 30.285 336.61 30.355 ;
    RECT 336.4 30.645 336.61 30.715 ;
    RECT 336.4 31.005 336.61 31.075 ;
    RECT 335.94 30.285 336.15 30.355 ;
    RECT 335.94 30.645 336.15 30.715 ;
    RECT 335.94 31.005 336.15 31.075 ;
    RECT 266.68 30.285 266.89 30.355 ;
    RECT 266.68 30.645 266.89 30.715 ;
    RECT 266.68 31.005 266.89 31.075 ;
    RECT 266.22 30.285 266.43 30.355 ;
    RECT 266.22 30.645 266.43 30.715 ;
    RECT 266.22 31.005 266.43 31.075 ;
    RECT 263.36 30.285 263.57 30.355 ;
    RECT 263.36 30.645 263.57 30.715 ;
    RECT 263.36 31.005 263.57 31.075 ;
    RECT 262.9 30.285 263.11 30.355 ;
    RECT 262.9 30.645 263.11 30.715 ;
    RECT 262.9 31.005 263.11 31.075 ;
    RECT 260.04 30.285 260.25 30.355 ;
    RECT 260.04 30.645 260.25 30.715 ;
    RECT 260.04 31.005 260.25 31.075 ;
    RECT 259.58 30.285 259.79 30.355 ;
    RECT 259.58 30.645 259.79 30.715 ;
    RECT 259.58 31.005 259.79 31.075 ;
    RECT 256.72 30.285 256.93 30.355 ;
    RECT 256.72 30.645 256.93 30.715 ;
    RECT 256.72 31.005 256.93 31.075 ;
    RECT 256.26 30.285 256.47 30.355 ;
    RECT 256.26 30.645 256.47 30.715 ;
    RECT 256.26 31.005 256.47 31.075 ;
    RECT 253.4 30.285 253.61 30.355 ;
    RECT 253.4 30.645 253.61 30.715 ;
    RECT 253.4 31.005 253.61 31.075 ;
    RECT 252.94 30.285 253.15 30.355 ;
    RECT 252.94 30.645 253.15 30.715 ;
    RECT 252.94 31.005 253.15 31.075 ;
    RECT 250.08 30.285 250.29 30.355 ;
    RECT 250.08 30.645 250.29 30.715 ;
    RECT 250.08 31.005 250.29 31.075 ;
    RECT 249.62 30.285 249.83 30.355 ;
    RECT 249.62 30.645 249.83 30.715 ;
    RECT 249.62 31.005 249.83 31.075 ;
    RECT 246.76 30.285 246.97 30.355 ;
    RECT 246.76 30.645 246.97 30.715 ;
    RECT 246.76 31.005 246.97 31.075 ;
    RECT 246.3 30.285 246.51 30.355 ;
    RECT 246.3 30.645 246.51 30.715 ;
    RECT 246.3 31.005 246.51 31.075 ;
    RECT 243.44 30.285 243.65 30.355 ;
    RECT 243.44 30.645 243.65 30.715 ;
    RECT 243.44 31.005 243.65 31.075 ;
    RECT 242.98 30.285 243.19 30.355 ;
    RECT 242.98 30.645 243.19 30.715 ;
    RECT 242.98 31.005 243.19 31.075 ;
    RECT 240.12 30.285 240.33 30.355 ;
    RECT 240.12 30.645 240.33 30.715 ;
    RECT 240.12 31.005 240.33 31.075 ;
    RECT 239.66 30.285 239.87 30.355 ;
    RECT 239.66 30.645 239.87 30.715 ;
    RECT 239.66 31.005 239.87 31.075 ;
    RECT 236.8 30.285 237.01 30.355 ;
    RECT 236.8 30.645 237.01 30.715 ;
    RECT 236.8 31.005 237.01 31.075 ;
    RECT 236.34 30.285 236.55 30.355 ;
    RECT 236.34 30.645 236.55 30.715 ;
    RECT 236.34 31.005 236.55 31.075 ;
    RECT 374.15 30.645 374.22 30.715 ;
    RECT 333.08 30.285 333.29 30.355 ;
    RECT 333.08 30.645 333.29 30.715 ;
    RECT 333.08 31.005 333.29 31.075 ;
    RECT 332.62 30.285 332.83 30.355 ;
    RECT 332.62 30.645 332.83 30.715 ;
    RECT 332.62 31.005 332.83 31.075 ;
    RECT 329.76 30.285 329.97 30.355 ;
    RECT 329.76 30.645 329.97 30.715 ;
    RECT 329.76 31.005 329.97 31.075 ;
    RECT 329.3 30.285 329.51 30.355 ;
    RECT 329.3 30.645 329.51 30.715 ;
    RECT 329.3 31.005 329.51 31.075 ;
    RECT 326.44 30.285 326.65 30.355 ;
    RECT 326.44 30.645 326.65 30.715 ;
    RECT 326.44 31.005 326.65 31.075 ;
    RECT 325.98 30.285 326.19 30.355 ;
    RECT 325.98 30.645 326.19 30.715 ;
    RECT 325.98 31.005 326.19 31.075 ;
    RECT 323.12 30.285 323.33 30.355 ;
    RECT 323.12 30.645 323.33 30.715 ;
    RECT 323.12 31.005 323.33 31.075 ;
    RECT 322.66 30.285 322.87 30.355 ;
    RECT 322.66 30.645 322.87 30.715 ;
    RECT 322.66 31.005 322.87 31.075 ;
    RECT 319.8 30.285 320.01 30.355 ;
    RECT 319.8 30.645 320.01 30.715 ;
    RECT 319.8 31.005 320.01 31.075 ;
    RECT 319.34 30.285 319.55 30.355 ;
    RECT 319.34 30.645 319.55 30.715 ;
    RECT 319.34 31.005 319.55 31.075 ;
    RECT 316.48 30.285 316.69 30.355 ;
    RECT 316.48 30.645 316.69 30.715 ;
    RECT 316.48 31.005 316.69 31.075 ;
    RECT 316.02 30.285 316.23 30.355 ;
    RECT 316.02 30.645 316.23 30.715 ;
    RECT 316.02 31.005 316.23 31.075 ;
    RECT 313.16 30.285 313.37 30.355 ;
    RECT 313.16 30.645 313.37 30.715 ;
    RECT 313.16 31.005 313.37 31.075 ;
    RECT 312.7 30.285 312.91 30.355 ;
    RECT 312.7 30.645 312.91 30.715 ;
    RECT 312.7 31.005 312.91 31.075 ;
    RECT 309.84 30.285 310.05 30.355 ;
    RECT 309.84 30.645 310.05 30.715 ;
    RECT 309.84 31.005 310.05 31.075 ;
    RECT 309.38 30.285 309.59 30.355 ;
    RECT 309.38 30.645 309.59 30.715 ;
    RECT 309.38 31.005 309.59 31.075 ;
    RECT 306.52 30.285 306.73 30.355 ;
    RECT 306.52 30.645 306.73 30.715 ;
    RECT 306.52 31.005 306.73 31.075 ;
    RECT 306.06 30.285 306.27 30.355 ;
    RECT 306.06 30.645 306.27 30.715 ;
    RECT 306.06 31.005 306.27 31.075 ;
    RECT 303.2 13.725 303.41 13.795 ;
    RECT 303.2 14.085 303.41 14.155 ;
    RECT 303.2 14.445 303.41 14.515 ;
    RECT 302.74 13.725 302.95 13.795 ;
    RECT 302.74 14.085 302.95 14.155 ;
    RECT 302.74 14.445 302.95 14.515 ;
    RECT 372.92 13.725 373.13 13.795 ;
    RECT 372.92 14.085 373.13 14.155 ;
    RECT 372.92 14.445 373.13 14.515 ;
    RECT 372.46 13.725 372.67 13.795 ;
    RECT 372.46 14.085 372.67 14.155 ;
    RECT 372.46 14.445 372.67 14.515 ;
    RECT 369.6 13.725 369.81 13.795 ;
    RECT 369.6 14.085 369.81 14.155 ;
    RECT 369.6 14.445 369.81 14.515 ;
    RECT 369.14 13.725 369.35 13.795 ;
    RECT 369.14 14.085 369.35 14.155 ;
    RECT 369.14 14.445 369.35 14.515 ;
    RECT 200.605 14.085 200.675 14.155 ;
    RECT 299.88 13.725 300.09 13.795 ;
    RECT 299.88 14.085 300.09 14.155 ;
    RECT 299.88 14.445 300.09 14.515 ;
    RECT 299.42 13.725 299.63 13.795 ;
    RECT 299.42 14.085 299.63 14.155 ;
    RECT 299.42 14.445 299.63 14.515 ;
    RECT 296.56 13.725 296.77 13.795 ;
    RECT 296.56 14.085 296.77 14.155 ;
    RECT 296.56 14.445 296.77 14.515 ;
    RECT 296.1 13.725 296.31 13.795 ;
    RECT 296.1 14.085 296.31 14.155 ;
    RECT 296.1 14.445 296.31 14.515 ;
    RECT 293.24 13.725 293.45 13.795 ;
    RECT 293.24 14.085 293.45 14.155 ;
    RECT 293.24 14.445 293.45 14.515 ;
    RECT 292.78 13.725 292.99 13.795 ;
    RECT 292.78 14.085 292.99 14.155 ;
    RECT 292.78 14.445 292.99 14.515 ;
    RECT 289.92 13.725 290.13 13.795 ;
    RECT 289.92 14.085 290.13 14.155 ;
    RECT 289.92 14.445 290.13 14.515 ;
    RECT 289.46 13.725 289.67 13.795 ;
    RECT 289.46 14.085 289.67 14.155 ;
    RECT 289.46 14.445 289.67 14.515 ;
    RECT 286.6 13.725 286.81 13.795 ;
    RECT 286.6 14.085 286.81 14.155 ;
    RECT 286.6 14.445 286.81 14.515 ;
    RECT 286.14 13.725 286.35 13.795 ;
    RECT 286.14 14.085 286.35 14.155 ;
    RECT 286.14 14.445 286.35 14.515 ;
    RECT 283.28 13.725 283.49 13.795 ;
    RECT 283.28 14.085 283.49 14.155 ;
    RECT 283.28 14.445 283.49 14.515 ;
    RECT 282.82 13.725 283.03 13.795 ;
    RECT 282.82 14.085 283.03 14.155 ;
    RECT 282.82 14.445 283.03 14.515 ;
    RECT 279.96 13.725 280.17 13.795 ;
    RECT 279.96 14.085 280.17 14.155 ;
    RECT 279.96 14.445 280.17 14.515 ;
    RECT 279.5 13.725 279.71 13.795 ;
    RECT 279.5 14.085 279.71 14.155 ;
    RECT 279.5 14.445 279.71 14.515 ;
    RECT 276.64 13.725 276.85 13.795 ;
    RECT 276.64 14.085 276.85 14.155 ;
    RECT 276.64 14.445 276.85 14.515 ;
    RECT 276.18 13.725 276.39 13.795 ;
    RECT 276.18 14.085 276.39 14.155 ;
    RECT 276.18 14.445 276.39 14.515 ;
    RECT 273.32 13.725 273.53 13.795 ;
    RECT 273.32 14.085 273.53 14.155 ;
    RECT 273.32 14.445 273.53 14.515 ;
    RECT 272.86 13.725 273.07 13.795 ;
    RECT 272.86 14.085 273.07 14.155 ;
    RECT 272.86 14.445 273.07 14.515 ;
    RECT 270.0 13.725 270.21 13.795 ;
    RECT 270.0 14.085 270.21 14.155 ;
    RECT 270.0 14.445 270.21 14.515 ;
    RECT 269.54 13.725 269.75 13.795 ;
    RECT 269.54 14.085 269.75 14.155 ;
    RECT 269.54 14.445 269.75 14.515 ;
    RECT 233.48 13.725 233.69 13.795 ;
    RECT 233.48 14.085 233.69 14.155 ;
    RECT 233.48 14.445 233.69 14.515 ;
    RECT 233.02 13.725 233.23 13.795 ;
    RECT 233.02 14.085 233.23 14.155 ;
    RECT 233.02 14.445 233.23 14.515 ;
    RECT 230.16 13.725 230.37 13.795 ;
    RECT 230.16 14.085 230.37 14.155 ;
    RECT 230.16 14.445 230.37 14.515 ;
    RECT 229.7 13.725 229.91 13.795 ;
    RECT 229.7 14.085 229.91 14.155 ;
    RECT 229.7 14.445 229.91 14.515 ;
    RECT 366.28 13.725 366.49 13.795 ;
    RECT 366.28 14.085 366.49 14.155 ;
    RECT 366.28 14.445 366.49 14.515 ;
    RECT 365.82 13.725 366.03 13.795 ;
    RECT 365.82 14.085 366.03 14.155 ;
    RECT 365.82 14.445 366.03 14.515 ;
    RECT 226.84 13.725 227.05 13.795 ;
    RECT 226.84 14.085 227.05 14.155 ;
    RECT 226.84 14.445 227.05 14.515 ;
    RECT 226.38 13.725 226.59 13.795 ;
    RECT 226.38 14.085 226.59 14.155 ;
    RECT 226.38 14.445 226.59 14.515 ;
    RECT 362.96 13.725 363.17 13.795 ;
    RECT 362.96 14.085 363.17 14.155 ;
    RECT 362.96 14.445 363.17 14.515 ;
    RECT 362.5 13.725 362.71 13.795 ;
    RECT 362.5 14.085 362.71 14.155 ;
    RECT 362.5 14.445 362.71 14.515 ;
    RECT 223.52 13.725 223.73 13.795 ;
    RECT 223.52 14.085 223.73 14.155 ;
    RECT 223.52 14.445 223.73 14.515 ;
    RECT 223.06 13.725 223.27 13.795 ;
    RECT 223.06 14.085 223.27 14.155 ;
    RECT 223.06 14.445 223.27 14.515 ;
    RECT 359.64 13.725 359.85 13.795 ;
    RECT 359.64 14.085 359.85 14.155 ;
    RECT 359.64 14.445 359.85 14.515 ;
    RECT 359.18 13.725 359.39 13.795 ;
    RECT 359.18 14.085 359.39 14.155 ;
    RECT 359.18 14.445 359.39 14.515 ;
    RECT 220.2 13.725 220.41 13.795 ;
    RECT 220.2 14.085 220.41 14.155 ;
    RECT 220.2 14.445 220.41 14.515 ;
    RECT 219.74 13.725 219.95 13.795 ;
    RECT 219.74 14.085 219.95 14.155 ;
    RECT 219.74 14.445 219.95 14.515 ;
    RECT 356.32 13.725 356.53 13.795 ;
    RECT 356.32 14.085 356.53 14.155 ;
    RECT 356.32 14.445 356.53 14.515 ;
    RECT 355.86 13.725 356.07 13.795 ;
    RECT 355.86 14.085 356.07 14.155 ;
    RECT 355.86 14.445 356.07 14.515 ;
    RECT 353.0 13.725 353.21 13.795 ;
    RECT 353.0 14.085 353.21 14.155 ;
    RECT 353.0 14.445 353.21 14.515 ;
    RECT 352.54 13.725 352.75 13.795 ;
    RECT 352.54 14.085 352.75 14.155 ;
    RECT 352.54 14.445 352.75 14.515 ;
    RECT 216.88 13.725 217.09 13.795 ;
    RECT 216.88 14.085 217.09 14.155 ;
    RECT 216.88 14.445 217.09 14.515 ;
    RECT 216.42 13.725 216.63 13.795 ;
    RECT 216.42 14.085 216.63 14.155 ;
    RECT 216.42 14.445 216.63 14.515 ;
    RECT 349.68 13.725 349.89 13.795 ;
    RECT 349.68 14.085 349.89 14.155 ;
    RECT 349.68 14.445 349.89 14.515 ;
    RECT 349.22 13.725 349.43 13.795 ;
    RECT 349.22 14.085 349.43 14.155 ;
    RECT 349.22 14.445 349.43 14.515 ;
    RECT 213.56 13.725 213.77 13.795 ;
    RECT 213.56 14.085 213.77 14.155 ;
    RECT 213.56 14.445 213.77 14.515 ;
    RECT 213.1 13.725 213.31 13.795 ;
    RECT 213.1 14.085 213.31 14.155 ;
    RECT 213.1 14.445 213.31 14.515 ;
    RECT 346.36 13.725 346.57 13.795 ;
    RECT 346.36 14.085 346.57 14.155 ;
    RECT 346.36 14.445 346.57 14.515 ;
    RECT 345.9 13.725 346.11 13.795 ;
    RECT 345.9 14.085 346.11 14.155 ;
    RECT 345.9 14.445 346.11 14.515 ;
    RECT 210.24 13.725 210.45 13.795 ;
    RECT 210.24 14.085 210.45 14.155 ;
    RECT 210.24 14.445 210.45 14.515 ;
    RECT 209.78 13.725 209.99 13.795 ;
    RECT 209.78 14.085 209.99 14.155 ;
    RECT 209.78 14.445 209.99 14.515 ;
    RECT 343.04 13.725 343.25 13.795 ;
    RECT 343.04 14.085 343.25 14.155 ;
    RECT 343.04 14.445 343.25 14.515 ;
    RECT 342.58 13.725 342.79 13.795 ;
    RECT 342.58 14.085 342.79 14.155 ;
    RECT 342.58 14.445 342.79 14.515 ;
    RECT 206.92 13.725 207.13 13.795 ;
    RECT 206.92 14.085 207.13 14.155 ;
    RECT 206.92 14.445 207.13 14.515 ;
    RECT 206.46 13.725 206.67 13.795 ;
    RECT 206.46 14.085 206.67 14.155 ;
    RECT 206.46 14.445 206.67 14.515 ;
    RECT 339.72 13.725 339.93 13.795 ;
    RECT 339.72 14.085 339.93 14.155 ;
    RECT 339.72 14.445 339.93 14.515 ;
    RECT 339.26 13.725 339.47 13.795 ;
    RECT 339.26 14.085 339.47 14.155 ;
    RECT 339.26 14.445 339.47 14.515 ;
    RECT 203.6 13.725 203.81 13.795 ;
    RECT 203.6 14.085 203.81 14.155 ;
    RECT 203.6 14.445 203.81 14.515 ;
    RECT 203.14 13.725 203.35 13.795 ;
    RECT 203.14 14.085 203.35 14.155 ;
    RECT 203.14 14.445 203.35 14.515 ;
    RECT 336.4 13.725 336.61 13.795 ;
    RECT 336.4 14.085 336.61 14.155 ;
    RECT 336.4 14.445 336.61 14.515 ;
    RECT 335.94 13.725 336.15 13.795 ;
    RECT 335.94 14.085 336.15 14.155 ;
    RECT 335.94 14.445 336.15 14.515 ;
    RECT 266.68 13.725 266.89 13.795 ;
    RECT 266.68 14.085 266.89 14.155 ;
    RECT 266.68 14.445 266.89 14.515 ;
    RECT 266.22 13.725 266.43 13.795 ;
    RECT 266.22 14.085 266.43 14.155 ;
    RECT 266.22 14.445 266.43 14.515 ;
    RECT 263.36 13.725 263.57 13.795 ;
    RECT 263.36 14.085 263.57 14.155 ;
    RECT 263.36 14.445 263.57 14.515 ;
    RECT 262.9 13.725 263.11 13.795 ;
    RECT 262.9 14.085 263.11 14.155 ;
    RECT 262.9 14.445 263.11 14.515 ;
    RECT 260.04 13.725 260.25 13.795 ;
    RECT 260.04 14.085 260.25 14.155 ;
    RECT 260.04 14.445 260.25 14.515 ;
    RECT 259.58 13.725 259.79 13.795 ;
    RECT 259.58 14.085 259.79 14.155 ;
    RECT 259.58 14.445 259.79 14.515 ;
    RECT 256.72 13.725 256.93 13.795 ;
    RECT 256.72 14.085 256.93 14.155 ;
    RECT 256.72 14.445 256.93 14.515 ;
    RECT 256.26 13.725 256.47 13.795 ;
    RECT 256.26 14.085 256.47 14.155 ;
    RECT 256.26 14.445 256.47 14.515 ;
    RECT 253.4 13.725 253.61 13.795 ;
    RECT 253.4 14.085 253.61 14.155 ;
    RECT 253.4 14.445 253.61 14.515 ;
    RECT 252.94 13.725 253.15 13.795 ;
    RECT 252.94 14.085 253.15 14.155 ;
    RECT 252.94 14.445 253.15 14.515 ;
    RECT 250.08 13.725 250.29 13.795 ;
    RECT 250.08 14.085 250.29 14.155 ;
    RECT 250.08 14.445 250.29 14.515 ;
    RECT 249.62 13.725 249.83 13.795 ;
    RECT 249.62 14.085 249.83 14.155 ;
    RECT 249.62 14.445 249.83 14.515 ;
    RECT 246.76 13.725 246.97 13.795 ;
    RECT 246.76 14.085 246.97 14.155 ;
    RECT 246.76 14.445 246.97 14.515 ;
    RECT 246.3 13.725 246.51 13.795 ;
    RECT 246.3 14.085 246.51 14.155 ;
    RECT 246.3 14.445 246.51 14.515 ;
    RECT 243.44 13.725 243.65 13.795 ;
    RECT 243.44 14.085 243.65 14.155 ;
    RECT 243.44 14.445 243.65 14.515 ;
    RECT 242.98 13.725 243.19 13.795 ;
    RECT 242.98 14.085 243.19 14.155 ;
    RECT 242.98 14.445 243.19 14.515 ;
    RECT 240.12 13.725 240.33 13.795 ;
    RECT 240.12 14.085 240.33 14.155 ;
    RECT 240.12 14.445 240.33 14.515 ;
    RECT 239.66 13.725 239.87 13.795 ;
    RECT 239.66 14.085 239.87 14.155 ;
    RECT 239.66 14.445 239.87 14.515 ;
    RECT 236.8 13.725 237.01 13.795 ;
    RECT 236.8 14.085 237.01 14.155 ;
    RECT 236.8 14.445 237.01 14.515 ;
    RECT 236.34 13.725 236.55 13.795 ;
    RECT 236.34 14.085 236.55 14.155 ;
    RECT 236.34 14.445 236.55 14.515 ;
    RECT 374.15 14.085 374.22 14.155 ;
    RECT 333.08 13.725 333.29 13.795 ;
    RECT 333.08 14.085 333.29 14.155 ;
    RECT 333.08 14.445 333.29 14.515 ;
    RECT 332.62 13.725 332.83 13.795 ;
    RECT 332.62 14.085 332.83 14.155 ;
    RECT 332.62 14.445 332.83 14.515 ;
    RECT 329.76 13.725 329.97 13.795 ;
    RECT 329.76 14.085 329.97 14.155 ;
    RECT 329.76 14.445 329.97 14.515 ;
    RECT 329.3 13.725 329.51 13.795 ;
    RECT 329.3 14.085 329.51 14.155 ;
    RECT 329.3 14.445 329.51 14.515 ;
    RECT 326.44 13.725 326.65 13.795 ;
    RECT 326.44 14.085 326.65 14.155 ;
    RECT 326.44 14.445 326.65 14.515 ;
    RECT 325.98 13.725 326.19 13.795 ;
    RECT 325.98 14.085 326.19 14.155 ;
    RECT 325.98 14.445 326.19 14.515 ;
    RECT 323.12 13.725 323.33 13.795 ;
    RECT 323.12 14.085 323.33 14.155 ;
    RECT 323.12 14.445 323.33 14.515 ;
    RECT 322.66 13.725 322.87 13.795 ;
    RECT 322.66 14.085 322.87 14.155 ;
    RECT 322.66 14.445 322.87 14.515 ;
    RECT 319.8 13.725 320.01 13.795 ;
    RECT 319.8 14.085 320.01 14.155 ;
    RECT 319.8 14.445 320.01 14.515 ;
    RECT 319.34 13.725 319.55 13.795 ;
    RECT 319.34 14.085 319.55 14.155 ;
    RECT 319.34 14.445 319.55 14.515 ;
    RECT 316.48 13.725 316.69 13.795 ;
    RECT 316.48 14.085 316.69 14.155 ;
    RECT 316.48 14.445 316.69 14.515 ;
    RECT 316.02 13.725 316.23 13.795 ;
    RECT 316.02 14.085 316.23 14.155 ;
    RECT 316.02 14.445 316.23 14.515 ;
    RECT 313.16 13.725 313.37 13.795 ;
    RECT 313.16 14.085 313.37 14.155 ;
    RECT 313.16 14.445 313.37 14.515 ;
    RECT 312.7 13.725 312.91 13.795 ;
    RECT 312.7 14.085 312.91 14.155 ;
    RECT 312.7 14.445 312.91 14.515 ;
    RECT 309.84 13.725 310.05 13.795 ;
    RECT 309.84 14.085 310.05 14.155 ;
    RECT 309.84 14.445 310.05 14.515 ;
    RECT 309.38 13.725 309.59 13.795 ;
    RECT 309.38 14.085 309.59 14.155 ;
    RECT 309.38 14.445 309.59 14.515 ;
    RECT 306.52 13.725 306.73 13.795 ;
    RECT 306.52 14.085 306.73 14.155 ;
    RECT 306.52 14.445 306.73 14.515 ;
    RECT 306.06 13.725 306.27 13.795 ;
    RECT 306.06 14.085 306.27 14.155 ;
    RECT 306.06 14.445 306.27 14.515 ;
    RECT 303.2 29.565 303.41 29.635 ;
    RECT 303.2 29.925 303.41 29.995 ;
    RECT 303.2 30.285 303.41 30.355 ;
    RECT 302.74 29.565 302.95 29.635 ;
    RECT 302.74 29.925 302.95 29.995 ;
    RECT 302.74 30.285 302.95 30.355 ;
    RECT 372.92 29.565 373.13 29.635 ;
    RECT 372.92 29.925 373.13 29.995 ;
    RECT 372.92 30.285 373.13 30.355 ;
    RECT 372.46 29.565 372.67 29.635 ;
    RECT 372.46 29.925 372.67 29.995 ;
    RECT 372.46 30.285 372.67 30.355 ;
    RECT 369.6 29.565 369.81 29.635 ;
    RECT 369.6 29.925 369.81 29.995 ;
    RECT 369.6 30.285 369.81 30.355 ;
    RECT 369.14 29.565 369.35 29.635 ;
    RECT 369.14 29.925 369.35 29.995 ;
    RECT 369.14 30.285 369.35 30.355 ;
    RECT 200.605 29.925 200.675 29.995 ;
    RECT 299.88 29.565 300.09 29.635 ;
    RECT 299.88 29.925 300.09 29.995 ;
    RECT 299.88 30.285 300.09 30.355 ;
    RECT 299.42 29.565 299.63 29.635 ;
    RECT 299.42 29.925 299.63 29.995 ;
    RECT 299.42 30.285 299.63 30.355 ;
    RECT 296.56 29.565 296.77 29.635 ;
    RECT 296.56 29.925 296.77 29.995 ;
    RECT 296.56 30.285 296.77 30.355 ;
    RECT 296.1 29.565 296.31 29.635 ;
    RECT 296.1 29.925 296.31 29.995 ;
    RECT 296.1 30.285 296.31 30.355 ;
    RECT 293.24 29.565 293.45 29.635 ;
    RECT 293.24 29.925 293.45 29.995 ;
    RECT 293.24 30.285 293.45 30.355 ;
    RECT 292.78 29.565 292.99 29.635 ;
    RECT 292.78 29.925 292.99 29.995 ;
    RECT 292.78 30.285 292.99 30.355 ;
    RECT 289.92 29.565 290.13 29.635 ;
    RECT 289.92 29.925 290.13 29.995 ;
    RECT 289.92 30.285 290.13 30.355 ;
    RECT 289.46 29.565 289.67 29.635 ;
    RECT 289.46 29.925 289.67 29.995 ;
    RECT 289.46 30.285 289.67 30.355 ;
    RECT 286.6 29.565 286.81 29.635 ;
    RECT 286.6 29.925 286.81 29.995 ;
    RECT 286.6 30.285 286.81 30.355 ;
    RECT 286.14 29.565 286.35 29.635 ;
    RECT 286.14 29.925 286.35 29.995 ;
    RECT 286.14 30.285 286.35 30.355 ;
    RECT 283.28 29.565 283.49 29.635 ;
    RECT 283.28 29.925 283.49 29.995 ;
    RECT 283.28 30.285 283.49 30.355 ;
    RECT 282.82 29.565 283.03 29.635 ;
    RECT 282.82 29.925 283.03 29.995 ;
    RECT 282.82 30.285 283.03 30.355 ;
    RECT 279.96 29.565 280.17 29.635 ;
    RECT 279.96 29.925 280.17 29.995 ;
    RECT 279.96 30.285 280.17 30.355 ;
    RECT 279.5 29.565 279.71 29.635 ;
    RECT 279.5 29.925 279.71 29.995 ;
    RECT 279.5 30.285 279.71 30.355 ;
    RECT 276.64 29.565 276.85 29.635 ;
    RECT 276.64 29.925 276.85 29.995 ;
    RECT 276.64 30.285 276.85 30.355 ;
    RECT 276.18 29.565 276.39 29.635 ;
    RECT 276.18 29.925 276.39 29.995 ;
    RECT 276.18 30.285 276.39 30.355 ;
    RECT 273.32 29.565 273.53 29.635 ;
    RECT 273.32 29.925 273.53 29.995 ;
    RECT 273.32 30.285 273.53 30.355 ;
    RECT 272.86 29.565 273.07 29.635 ;
    RECT 272.86 29.925 273.07 29.995 ;
    RECT 272.86 30.285 273.07 30.355 ;
    RECT 270.0 29.565 270.21 29.635 ;
    RECT 270.0 29.925 270.21 29.995 ;
    RECT 270.0 30.285 270.21 30.355 ;
    RECT 269.54 29.565 269.75 29.635 ;
    RECT 269.54 29.925 269.75 29.995 ;
    RECT 269.54 30.285 269.75 30.355 ;
    RECT 233.48 29.565 233.69 29.635 ;
    RECT 233.48 29.925 233.69 29.995 ;
    RECT 233.48 30.285 233.69 30.355 ;
    RECT 233.02 29.565 233.23 29.635 ;
    RECT 233.02 29.925 233.23 29.995 ;
    RECT 233.02 30.285 233.23 30.355 ;
    RECT 230.16 29.565 230.37 29.635 ;
    RECT 230.16 29.925 230.37 29.995 ;
    RECT 230.16 30.285 230.37 30.355 ;
    RECT 229.7 29.565 229.91 29.635 ;
    RECT 229.7 29.925 229.91 29.995 ;
    RECT 229.7 30.285 229.91 30.355 ;
    RECT 366.28 29.565 366.49 29.635 ;
    RECT 366.28 29.925 366.49 29.995 ;
    RECT 366.28 30.285 366.49 30.355 ;
    RECT 365.82 29.565 366.03 29.635 ;
    RECT 365.82 29.925 366.03 29.995 ;
    RECT 365.82 30.285 366.03 30.355 ;
    RECT 226.84 29.565 227.05 29.635 ;
    RECT 226.84 29.925 227.05 29.995 ;
    RECT 226.84 30.285 227.05 30.355 ;
    RECT 226.38 29.565 226.59 29.635 ;
    RECT 226.38 29.925 226.59 29.995 ;
    RECT 226.38 30.285 226.59 30.355 ;
    RECT 362.96 29.565 363.17 29.635 ;
    RECT 362.96 29.925 363.17 29.995 ;
    RECT 362.96 30.285 363.17 30.355 ;
    RECT 362.5 29.565 362.71 29.635 ;
    RECT 362.5 29.925 362.71 29.995 ;
    RECT 362.5 30.285 362.71 30.355 ;
    RECT 223.52 29.565 223.73 29.635 ;
    RECT 223.52 29.925 223.73 29.995 ;
    RECT 223.52 30.285 223.73 30.355 ;
    RECT 223.06 29.565 223.27 29.635 ;
    RECT 223.06 29.925 223.27 29.995 ;
    RECT 223.06 30.285 223.27 30.355 ;
    RECT 359.64 29.565 359.85 29.635 ;
    RECT 359.64 29.925 359.85 29.995 ;
    RECT 359.64 30.285 359.85 30.355 ;
    RECT 359.18 29.565 359.39 29.635 ;
    RECT 359.18 29.925 359.39 29.995 ;
    RECT 359.18 30.285 359.39 30.355 ;
    RECT 220.2 29.565 220.41 29.635 ;
    RECT 220.2 29.925 220.41 29.995 ;
    RECT 220.2 30.285 220.41 30.355 ;
    RECT 219.74 29.565 219.95 29.635 ;
    RECT 219.74 29.925 219.95 29.995 ;
    RECT 219.74 30.285 219.95 30.355 ;
    RECT 356.32 29.565 356.53 29.635 ;
    RECT 356.32 29.925 356.53 29.995 ;
    RECT 356.32 30.285 356.53 30.355 ;
    RECT 355.86 29.565 356.07 29.635 ;
    RECT 355.86 29.925 356.07 29.995 ;
    RECT 355.86 30.285 356.07 30.355 ;
    RECT 353.0 29.565 353.21 29.635 ;
    RECT 353.0 29.925 353.21 29.995 ;
    RECT 353.0 30.285 353.21 30.355 ;
    RECT 352.54 29.565 352.75 29.635 ;
    RECT 352.54 29.925 352.75 29.995 ;
    RECT 352.54 30.285 352.75 30.355 ;
    RECT 216.88 29.565 217.09 29.635 ;
    RECT 216.88 29.925 217.09 29.995 ;
    RECT 216.88 30.285 217.09 30.355 ;
    RECT 216.42 29.565 216.63 29.635 ;
    RECT 216.42 29.925 216.63 29.995 ;
    RECT 216.42 30.285 216.63 30.355 ;
    RECT 349.68 29.565 349.89 29.635 ;
    RECT 349.68 29.925 349.89 29.995 ;
    RECT 349.68 30.285 349.89 30.355 ;
    RECT 349.22 29.565 349.43 29.635 ;
    RECT 349.22 29.925 349.43 29.995 ;
    RECT 349.22 30.285 349.43 30.355 ;
    RECT 213.56 29.565 213.77 29.635 ;
    RECT 213.56 29.925 213.77 29.995 ;
    RECT 213.56 30.285 213.77 30.355 ;
    RECT 213.1 29.565 213.31 29.635 ;
    RECT 213.1 29.925 213.31 29.995 ;
    RECT 213.1 30.285 213.31 30.355 ;
    RECT 346.36 29.565 346.57 29.635 ;
    RECT 346.36 29.925 346.57 29.995 ;
    RECT 346.36 30.285 346.57 30.355 ;
    RECT 345.9 29.565 346.11 29.635 ;
    RECT 345.9 29.925 346.11 29.995 ;
    RECT 345.9 30.285 346.11 30.355 ;
    RECT 210.24 29.565 210.45 29.635 ;
    RECT 210.24 29.925 210.45 29.995 ;
    RECT 210.24 30.285 210.45 30.355 ;
    RECT 209.78 29.565 209.99 29.635 ;
    RECT 209.78 29.925 209.99 29.995 ;
    RECT 209.78 30.285 209.99 30.355 ;
    RECT 343.04 29.565 343.25 29.635 ;
    RECT 343.04 29.925 343.25 29.995 ;
    RECT 343.04 30.285 343.25 30.355 ;
    RECT 342.58 29.565 342.79 29.635 ;
    RECT 342.58 29.925 342.79 29.995 ;
    RECT 342.58 30.285 342.79 30.355 ;
    RECT 206.92 29.565 207.13 29.635 ;
    RECT 206.92 29.925 207.13 29.995 ;
    RECT 206.92 30.285 207.13 30.355 ;
    RECT 206.46 29.565 206.67 29.635 ;
    RECT 206.46 29.925 206.67 29.995 ;
    RECT 206.46 30.285 206.67 30.355 ;
    RECT 339.72 29.565 339.93 29.635 ;
    RECT 339.72 29.925 339.93 29.995 ;
    RECT 339.72 30.285 339.93 30.355 ;
    RECT 339.26 29.565 339.47 29.635 ;
    RECT 339.26 29.925 339.47 29.995 ;
    RECT 339.26 30.285 339.47 30.355 ;
    RECT 203.6 29.565 203.81 29.635 ;
    RECT 203.6 29.925 203.81 29.995 ;
    RECT 203.6 30.285 203.81 30.355 ;
    RECT 203.14 29.565 203.35 29.635 ;
    RECT 203.14 29.925 203.35 29.995 ;
    RECT 203.14 30.285 203.35 30.355 ;
    RECT 336.4 29.565 336.61 29.635 ;
    RECT 336.4 29.925 336.61 29.995 ;
    RECT 336.4 30.285 336.61 30.355 ;
    RECT 335.94 29.565 336.15 29.635 ;
    RECT 335.94 29.925 336.15 29.995 ;
    RECT 335.94 30.285 336.15 30.355 ;
    RECT 266.68 29.565 266.89 29.635 ;
    RECT 266.68 29.925 266.89 29.995 ;
    RECT 266.68 30.285 266.89 30.355 ;
    RECT 266.22 29.565 266.43 29.635 ;
    RECT 266.22 29.925 266.43 29.995 ;
    RECT 266.22 30.285 266.43 30.355 ;
    RECT 263.36 29.565 263.57 29.635 ;
    RECT 263.36 29.925 263.57 29.995 ;
    RECT 263.36 30.285 263.57 30.355 ;
    RECT 262.9 29.565 263.11 29.635 ;
    RECT 262.9 29.925 263.11 29.995 ;
    RECT 262.9 30.285 263.11 30.355 ;
    RECT 260.04 29.565 260.25 29.635 ;
    RECT 260.04 29.925 260.25 29.995 ;
    RECT 260.04 30.285 260.25 30.355 ;
    RECT 259.58 29.565 259.79 29.635 ;
    RECT 259.58 29.925 259.79 29.995 ;
    RECT 259.58 30.285 259.79 30.355 ;
    RECT 256.72 29.565 256.93 29.635 ;
    RECT 256.72 29.925 256.93 29.995 ;
    RECT 256.72 30.285 256.93 30.355 ;
    RECT 256.26 29.565 256.47 29.635 ;
    RECT 256.26 29.925 256.47 29.995 ;
    RECT 256.26 30.285 256.47 30.355 ;
    RECT 253.4 29.565 253.61 29.635 ;
    RECT 253.4 29.925 253.61 29.995 ;
    RECT 253.4 30.285 253.61 30.355 ;
    RECT 252.94 29.565 253.15 29.635 ;
    RECT 252.94 29.925 253.15 29.995 ;
    RECT 252.94 30.285 253.15 30.355 ;
    RECT 250.08 29.565 250.29 29.635 ;
    RECT 250.08 29.925 250.29 29.995 ;
    RECT 250.08 30.285 250.29 30.355 ;
    RECT 249.62 29.565 249.83 29.635 ;
    RECT 249.62 29.925 249.83 29.995 ;
    RECT 249.62 30.285 249.83 30.355 ;
    RECT 246.76 29.565 246.97 29.635 ;
    RECT 246.76 29.925 246.97 29.995 ;
    RECT 246.76 30.285 246.97 30.355 ;
    RECT 246.3 29.565 246.51 29.635 ;
    RECT 246.3 29.925 246.51 29.995 ;
    RECT 246.3 30.285 246.51 30.355 ;
    RECT 243.44 29.565 243.65 29.635 ;
    RECT 243.44 29.925 243.65 29.995 ;
    RECT 243.44 30.285 243.65 30.355 ;
    RECT 242.98 29.565 243.19 29.635 ;
    RECT 242.98 29.925 243.19 29.995 ;
    RECT 242.98 30.285 243.19 30.355 ;
    RECT 240.12 29.565 240.33 29.635 ;
    RECT 240.12 29.925 240.33 29.995 ;
    RECT 240.12 30.285 240.33 30.355 ;
    RECT 239.66 29.565 239.87 29.635 ;
    RECT 239.66 29.925 239.87 29.995 ;
    RECT 239.66 30.285 239.87 30.355 ;
    RECT 236.8 29.565 237.01 29.635 ;
    RECT 236.8 29.925 237.01 29.995 ;
    RECT 236.8 30.285 237.01 30.355 ;
    RECT 236.34 29.565 236.55 29.635 ;
    RECT 236.34 29.925 236.55 29.995 ;
    RECT 236.34 30.285 236.55 30.355 ;
    RECT 374.15 29.925 374.22 29.995 ;
    RECT 333.08 29.565 333.29 29.635 ;
    RECT 333.08 29.925 333.29 29.995 ;
    RECT 333.08 30.285 333.29 30.355 ;
    RECT 332.62 29.565 332.83 29.635 ;
    RECT 332.62 29.925 332.83 29.995 ;
    RECT 332.62 30.285 332.83 30.355 ;
    RECT 329.76 29.565 329.97 29.635 ;
    RECT 329.76 29.925 329.97 29.995 ;
    RECT 329.76 30.285 329.97 30.355 ;
    RECT 329.3 29.565 329.51 29.635 ;
    RECT 329.3 29.925 329.51 29.995 ;
    RECT 329.3 30.285 329.51 30.355 ;
    RECT 326.44 29.565 326.65 29.635 ;
    RECT 326.44 29.925 326.65 29.995 ;
    RECT 326.44 30.285 326.65 30.355 ;
    RECT 325.98 29.565 326.19 29.635 ;
    RECT 325.98 29.925 326.19 29.995 ;
    RECT 325.98 30.285 326.19 30.355 ;
    RECT 323.12 29.565 323.33 29.635 ;
    RECT 323.12 29.925 323.33 29.995 ;
    RECT 323.12 30.285 323.33 30.355 ;
    RECT 322.66 29.565 322.87 29.635 ;
    RECT 322.66 29.925 322.87 29.995 ;
    RECT 322.66 30.285 322.87 30.355 ;
    RECT 319.8 29.565 320.01 29.635 ;
    RECT 319.8 29.925 320.01 29.995 ;
    RECT 319.8 30.285 320.01 30.355 ;
    RECT 319.34 29.565 319.55 29.635 ;
    RECT 319.34 29.925 319.55 29.995 ;
    RECT 319.34 30.285 319.55 30.355 ;
    RECT 316.48 29.565 316.69 29.635 ;
    RECT 316.48 29.925 316.69 29.995 ;
    RECT 316.48 30.285 316.69 30.355 ;
    RECT 316.02 29.565 316.23 29.635 ;
    RECT 316.02 29.925 316.23 29.995 ;
    RECT 316.02 30.285 316.23 30.355 ;
    RECT 313.16 29.565 313.37 29.635 ;
    RECT 313.16 29.925 313.37 29.995 ;
    RECT 313.16 30.285 313.37 30.355 ;
    RECT 312.7 29.565 312.91 29.635 ;
    RECT 312.7 29.925 312.91 29.995 ;
    RECT 312.7 30.285 312.91 30.355 ;
    RECT 309.84 29.565 310.05 29.635 ;
    RECT 309.84 29.925 310.05 29.995 ;
    RECT 309.84 30.285 310.05 30.355 ;
    RECT 309.38 29.565 309.59 29.635 ;
    RECT 309.38 29.925 309.59 29.995 ;
    RECT 309.38 30.285 309.59 30.355 ;
    RECT 306.52 29.565 306.73 29.635 ;
    RECT 306.52 29.925 306.73 29.995 ;
    RECT 306.52 30.285 306.73 30.355 ;
    RECT 306.06 29.565 306.27 29.635 ;
    RECT 306.06 29.925 306.27 29.995 ;
    RECT 306.06 30.285 306.27 30.355 ;
    RECT 303.2 13.005 303.41 13.075 ;
    RECT 303.2 13.365 303.41 13.435 ;
    RECT 303.2 13.725 303.41 13.795 ;
    RECT 302.74 13.005 302.95 13.075 ;
    RECT 302.74 13.365 302.95 13.435 ;
    RECT 302.74 13.725 302.95 13.795 ;
    RECT 372.92 13.005 373.13 13.075 ;
    RECT 372.92 13.365 373.13 13.435 ;
    RECT 372.92 13.725 373.13 13.795 ;
    RECT 372.46 13.005 372.67 13.075 ;
    RECT 372.46 13.365 372.67 13.435 ;
    RECT 372.46 13.725 372.67 13.795 ;
    RECT 369.6 13.005 369.81 13.075 ;
    RECT 369.6 13.365 369.81 13.435 ;
    RECT 369.6 13.725 369.81 13.795 ;
    RECT 369.14 13.005 369.35 13.075 ;
    RECT 369.14 13.365 369.35 13.435 ;
    RECT 369.14 13.725 369.35 13.795 ;
    RECT 200.605 13.365 200.675 13.435 ;
    RECT 299.88 13.005 300.09 13.075 ;
    RECT 299.88 13.365 300.09 13.435 ;
    RECT 299.88 13.725 300.09 13.795 ;
    RECT 299.42 13.005 299.63 13.075 ;
    RECT 299.42 13.365 299.63 13.435 ;
    RECT 299.42 13.725 299.63 13.795 ;
    RECT 296.56 13.005 296.77 13.075 ;
    RECT 296.56 13.365 296.77 13.435 ;
    RECT 296.56 13.725 296.77 13.795 ;
    RECT 296.1 13.005 296.31 13.075 ;
    RECT 296.1 13.365 296.31 13.435 ;
    RECT 296.1 13.725 296.31 13.795 ;
    RECT 293.24 13.005 293.45 13.075 ;
    RECT 293.24 13.365 293.45 13.435 ;
    RECT 293.24 13.725 293.45 13.795 ;
    RECT 292.78 13.005 292.99 13.075 ;
    RECT 292.78 13.365 292.99 13.435 ;
    RECT 292.78 13.725 292.99 13.795 ;
    RECT 289.92 13.005 290.13 13.075 ;
    RECT 289.92 13.365 290.13 13.435 ;
    RECT 289.92 13.725 290.13 13.795 ;
    RECT 289.46 13.005 289.67 13.075 ;
    RECT 289.46 13.365 289.67 13.435 ;
    RECT 289.46 13.725 289.67 13.795 ;
    RECT 286.6 13.005 286.81 13.075 ;
    RECT 286.6 13.365 286.81 13.435 ;
    RECT 286.6 13.725 286.81 13.795 ;
    RECT 286.14 13.005 286.35 13.075 ;
    RECT 286.14 13.365 286.35 13.435 ;
    RECT 286.14 13.725 286.35 13.795 ;
    RECT 283.28 13.005 283.49 13.075 ;
    RECT 283.28 13.365 283.49 13.435 ;
    RECT 283.28 13.725 283.49 13.795 ;
    RECT 282.82 13.005 283.03 13.075 ;
    RECT 282.82 13.365 283.03 13.435 ;
    RECT 282.82 13.725 283.03 13.795 ;
    RECT 279.96 13.005 280.17 13.075 ;
    RECT 279.96 13.365 280.17 13.435 ;
    RECT 279.96 13.725 280.17 13.795 ;
    RECT 279.5 13.005 279.71 13.075 ;
    RECT 279.5 13.365 279.71 13.435 ;
    RECT 279.5 13.725 279.71 13.795 ;
    RECT 276.64 13.005 276.85 13.075 ;
    RECT 276.64 13.365 276.85 13.435 ;
    RECT 276.64 13.725 276.85 13.795 ;
    RECT 276.18 13.005 276.39 13.075 ;
    RECT 276.18 13.365 276.39 13.435 ;
    RECT 276.18 13.725 276.39 13.795 ;
    RECT 273.32 13.005 273.53 13.075 ;
    RECT 273.32 13.365 273.53 13.435 ;
    RECT 273.32 13.725 273.53 13.795 ;
    RECT 272.86 13.005 273.07 13.075 ;
    RECT 272.86 13.365 273.07 13.435 ;
    RECT 272.86 13.725 273.07 13.795 ;
    RECT 270.0 13.005 270.21 13.075 ;
    RECT 270.0 13.365 270.21 13.435 ;
    RECT 270.0 13.725 270.21 13.795 ;
    RECT 269.54 13.005 269.75 13.075 ;
    RECT 269.54 13.365 269.75 13.435 ;
    RECT 269.54 13.725 269.75 13.795 ;
    RECT 233.48 13.005 233.69 13.075 ;
    RECT 233.48 13.365 233.69 13.435 ;
    RECT 233.48 13.725 233.69 13.795 ;
    RECT 233.02 13.005 233.23 13.075 ;
    RECT 233.02 13.365 233.23 13.435 ;
    RECT 233.02 13.725 233.23 13.795 ;
    RECT 230.16 13.005 230.37 13.075 ;
    RECT 230.16 13.365 230.37 13.435 ;
    RECT 230.16 13.725 230.37 13.795 ;
    RECT 229.7 13.005 229.91 13.075 ;
    RECT 229.7 13.365 229.91 13.435 ;
    RECT 229.7 13.725 229.91 13.795 ;
    RECT 366.28 13.005 366.49 13.075 ;
    RECT 366.28 13.365 366.49 13.435 ;
    RECT 366.28 13.725 366.49 13.795 ;
    RECT 365.82 13.005 366.03 13.075 ;
    RECT 365.82 13.365 366.03 13.435 ;
    RECT 365.82 13.725 366.03 13.795 ;
    RECT 226.84 13.005 227.05 13.075 ;
    RECT 226.84 13.365 227.05 13.435 ;
    RECT 226.84 13.725 227.05 13.795 ;
    RECT 226.38 13.005 226.59 13.075 ;
    RECT 226.38 13.365 226.59 13.435 ;
    RECT 226.38 13.725 226.59 13.795 ;
    RECT 362.96 13.005 363.17 13.075 ;
    RECT 362.96 13.365 363.17 13.435 ;
    RECT 362.96 13.725 363.17 13.795 ;
    RECT 362.5 13.005 362.71 13.075 ;
    RECT 362.5 13.365 362.71 13.435 ;
    RECT 362.5 13.725 362.71 13.795 ;
    RECT 223.52 13.005 223.73 13.075 ;
    RECT 223.52 13.365 223.73 13.435 ;
    RECT 223.52 13.725 223.73 13.795 ;
    RECT 223.06 13.005 223.27 13.075 ;
    RECT 223.06 13.365 223.27 13.435 ;
    RECT 223.06 13.725 223.27 13.795 ;
    RECT 359.64 13.005 359.85 13.075 ;
    RECT 359.64 13.365 359.85 13.435 ;
    RECT 359.64 13.725 359.85 13.795 ;
    RECT 359.18 13.005 359.39 13.075 ;
    RECT 359.18 13.365 359.39 13.435 ;
    RECT 359.18 13.725 359.39 13.795 ;
    RECT 220.2 13.005 220.41 13.075 ;
    RECT 220.2 13.365 220.41 13.435 ;
    RECT 220.2 13.725 220.41 13.795 ;
    RECT 219.74 13.005 219.95 13.075 ;
    RECT 219.74 13.365 219.95 13.435 ;
    RECT 219.74 13.725 219.95 13.795 ;
    RECT 356.32 13.005 356.53 13.075 ;
    RECT 356.32 13.365 356.53 13.435 ;
    RECT 356.32 13.725 356.53 13.795 ;
    RECT 355.86 13.005 356.07 13.075 ;
    RECT 355.86 13.365 356.07 13.435 ;
    RECT 355.86 13.725 356.07 13.795 ;
    RECT 353.0 13.005 353.21 13.075 ;
    RECT 353.0 13.365 353.21 13.435 ;
    RECT 353.0 13.725 353.21 13.795 ;
    RECT 352.54 13.005 352.75 13.075 ;
    RECT 352.54 13.365 352.75 13.435 ;
    RECT 352.54 13.725 352.75 13.795 ;
    RECT 216.88 13.005 217.09 13.075 ;
    RECT 216.88 13.365 217.09 13.435 ;
    RECT 216.88 13.725 217.09 13.795 ;
    RECT 216.42 13.005 216.63 13.075 ;
    RECT 216.42 13.365 216.63 13.435 ;
    RECT 216.42 13.725 216.63 13.795 ;
    RECT 349.68 13.005 349.89 13.075 ;
    RECT 349.68 13.365 349.89 13.435 ;
    RECT 349.68 13.725 349.89 13.795 ;
    RECT 349.22 13.005 349.43 13.075 ;
    RECT 349.22 13.365 349.43 13.435 ;
    RECT 349.22 13.725 349.43 13.795 ;
    RECT 213.56 13.005 213.77 13.075 ;
    RECT 213.56 13.365 213.77 13.435 ;
    RECT 213.56 13.725 213.77 13.795 ;
    RECT 213.1 13.005 213.31 13.075 ;
    RECT 213.1 13.365 213.31 13.435 ;
    RECT 213.1 13.725 213.31 13.795 ;
    RECT 346.36 13.005 346.57 13.075 ;
    RECT 346.36 13.365 346.57 13.435 ;
    RECT 346.36 13.725 346.57 13.795 ;
    RECT 345.9 13.005 346.11 13.075 ;
    RECT 345.9 13.365 346.11 13.435 ;
    RECT 345.9 13.725 346.11 13.795 ;
    RECT 210.24 13.005 210.45 13.075 ;
    RECT 210.24 13.365 210.45 13.435 ;
    RECT 210.24 13.725 210.45 13.795 ;
    RECT 209.78 13.005 209.99 13.075 ;
    RECT 209.78 13.365 209.99 13.435 ;
    RECT 209.78 13.725 209.99 13.795 ;
    RECT 343.04 13.005 343.25 13.075 ;
    RECT 343.04 13.365 343.25 13.435 ;
    RECT 343.04 13.725 343.25 13.795 ;
    RECT 342.58 13.005 342.79 13.075 ;
    RECT 342.58 13.365 342.79 13.435 ;
    RECT 342.58 13.725 342.79 13.795 ;
    RECT 206.92 13.005 207.13 13.075 ;
    RECT 206.92 13.365 207.13 13.435 ;
    RECT 206.92 13.725 207.13 13.795 ;
    RECT 206.46 13.005 206.67 13.075 ;
    RECT 206.46 13.365 206.67 13.435 ;
    RECT 206.46 13.725 206.67 13.795 ;
    RECT 339.72 13.005 339.93 13.075 ;
    RECT 339.72 13.365 339.93 13.435 ;
    RECT 339.72 13.725 339.93 13.795 ;
    RECT 339.26 13.005 339.47 13.075 ;
    RECT 339.26 13.365 339.47 13.435 ;
    RECT 339.26 13.725 339.47 13.795 ;
    RECT 203.6 13.005 203.81 13.075 ;
    RECT 203.6 13.365 203.81 13.435 ;
    RECT 203.6 13.725 203.81 13.795 ;
    RECT 203.14 13.005 203.35 13.075 ;
    RECT 203.14 13.365 203.35 13.435 ;
    RECT 203.14 13.725 203.35 13.795 ;
    RECT 336.4 13.005 336.61 13.075 ;
    RECT 336.4 13.365 336.61 13.435 ;
    RECT 336.4 13.725 336.61 13.795 ;
    RECT 335.94 13.005 336.15 13.075 ;
    RECT 335.94 13.365 336.15 13.435 ;
    RECT 335.94 13.725 336.15 13.795 ;
    RECT 266.68 13.005 266.89 13.075 ;
    RECT 266.68 13.365 266.89 13.435 ;
    RECT 266.68 13.725 266.89 13.795 ;
    RECT 266.22 13.005 266.43 13.075 ;
    RECT 266.22 13.365 266.43 13.435 ;
    RECT 266.22 13.725 266.43 13.795 ;
    RECT 263.36 13.005 263.57 13.075 ;
    RECT 263.36 13.365 263.57 13.435 ;
    RECT 263.36 13.725 263.57 13.795 ;
    RECT 262.9 13.005 263.11 13.075 ;
    RECT 262.9 13.365 263.11 13.435 ;
    RECT 262.9 13.725 263.11 13.795 ;
    RECT 260.04 13.005 260.25 13.075 ;
    RECT 260.04 13.365 260.25 13.435 ;
    RECT 260.04 13.725 260.25 13.795 ;
    RECT 259.58 13.005 259.79 13.075 ;
    RECT 259.58 13.365 259.79 13.435 ;
    RECT 259.58 13.725 259.79 13.795 ;
    RECT 256.72 13.005 256.93 13.075 ;
    RECT 256.72 13.365 256.93 13.435 ;
    RECT 256.72 13.725 256.93 13.795 ;
    RECT 256.26 13.005 256.47 13.075 ;
    RECT 256.26 13.365 256.47 13.435 ;
    RECT 256.26 13.725 256.47 13.795 ;
    RECT 253.4 13.005 253.61 13.075 ;
    RECT 253.4 13.365 253.61 13.435 ;
    RECT 253.4 13.725 253.61 13.795 ;
    RECT 252.94 13.005 253.15 13.075 ;
    RECT 252.94 13.365 253.15 13.435 ;
    RECT 252.94 13.725 253.15 13.795 ;
    RECT 250.08 13.005 250.29 13.075 ;
    RECT 250.08 13.365 250.29 13.435 ;
    RECT 250.08 13.725 250.29 13.795 ;
    RECT 249.62 13.005 249.83 13.075 ;
    RECT 249.62 13.365 249.83 13.435 ;
    RECT 249.62 13.725 249.83 13.795 ;
    RECT 246.76 13.005 246.97 13.075 ;
    RECT 246.76 13.365 246.97 13.435 ;
    RECT 246.76 13.725 246.97 13.795 ;
    RECT 246.3 13.005 246.51 13.075 ;
    RECT 246.3 13.365 246.51 13.435 ;
    RECT 246.3 13.725 246.51 13.795 ;
    RECT 243.44 13.005 243.65 13.075 ;
    RECT 243.44 13.365 243.65 13.435 ;
    RECT 243.44 13.725 243.65 13.795 ;
    RECT 242.98 13.005 243.19 13.075 ;
    RECT 242.98 13.365 243.19 13.435 ;
    RECT 242.98 13.725 243.19 13.795 ;
    RECT 240.12 13.005 240.33 13.075 ;
    RECT 240.12 13.365 240.33 13.435 ;
    RECT 240.12 13.725 240.33 13.795 ;
    RECT 239.66 13.005 239.87 13.075 ;
    RECT 239.66 13.365 239.87 13.435 ;
    RECT 239.66 13.725 239.87 13.795 ;
    RECT 236.8 13.005 237.01 13.075 ;
    RECT 236.8 13.365 237.01 13.435 ;
    RECT 236.8 13.725 237.01 13.795 ;
    RECT 236.34 13.005 236.55 13.075 ;
    RECT 236.34 13.365 236.55 13.435 ;
    RECT 236.34 13.725 236.55 13.795 ;
    RECT 374.15 13.365 374.22 13.435 ;
    RECT 333.08 13.005 333.29 13.075 ;
    RECT 333.08 13.365 333.29 13.435 ;
    RECT 333.08 13.725 333.29 13.795 ;
    RECT 332.62 13.005 332.83 13.075 ;
    RECT 332.62 13.365 332.83 13.435 ;
    RECT 332.62 13.725 332.83 13.795 ;
    RECT 329.76 13.005 329.97 13.075 ;
    RECT 329.76 13.365 329.97 13.435 ;
    RECT 329.76 13.725 329.97 13.795 ;
    RECT 329.3 13.005 329.51 13.075 ;
    RECT 329.3 13.365 329.51 13.435 ;
    RECT 329.3 13.725 329.51 13.795 ;
    RECT 326.44 13.005 326.65 13.075 ;
    RECT 326.44 13.365 326.65 13.435 ;
    RECT 326.44 13.725 326.65 13.795 ;
    RECT 325.98 13.005 326.19 13.075 ;
    RECT 325.98 13.365 326.19 13.435 ;
    RECT 325.98 13.725 326.19 13.795 ;
    RECT 323.12 13.005 323.33 13.075 ;
    RECT 323.12 13.365 323.33 13.435 ;
    RECT 323.12 13.725 323.33 13.795 ;
    RECT 322.66 13.005 322.87 13.075 ;
    RECT 322.66 13.365 322.87 13.435 ;
    RECT 322.66 13.725 322.87 13.795 ;
    RECT 319.8 13.005 320.01 13.075 ;
    RECT 319.8 13.365 320.01 13.435 ;
    RECT 319.8 13.725 320.01 13.795 ;
    RECT 319.34 13.005 319.55 13.075 ;
    RECT 319.34 13.365 319.55 13.435 ;
    RECT 319.34 13.725 319.55 13.795 ;
    RECT 316.48 13.005 316.69 13.075 ;
    RECT 316.48 13.365 316.69 13.435 ;
    RECT 316.48 13.725 316.69 13.795 ;
    RECT 316.02 13.005 316.23 13.075 ;
    RECT 316.02 13.365 316.23 13.435 ;
    RECT 316.02 13.725 316.23 13.795 ;
    RECT 313.16 13.005 313.37 13.075 ;
    RECT 313.16 13.365 313.37 13.435 ;
    RECT 313.16 13.725 313.37 13.795 ;
    RECT 312.7 13.005 312.91 13.075 ;
    RECT 312.7 13.365 312.91 13.435 ;
    RECT 312.7 13.725 312.91 13.795 ;
    RECT 309.84 13.005 310.05 13.075 ;
    RECT 309.84 13.365 310.05 13.435 ;
    RECT 309.84 13.725 310.05 13.795 ;
    RECT 309.38 13.005 309.59 13.075 ;
    RECT 309.38 13.365 309.59 13.435 ;
    RECT 309.38 13.725 309.59 13.795 ;
    RECT 306.52 13.005 306.73 13.075 ;
    RECT 306.52 13.365 306.73 13.435 ;
    RECT 306.52 13.725 306.73 13.795 ;
    RECT 306.06 13.005 306.27 13.075 ;
    RECT 306.06 13.365 306.27 13.435 ;
    RECT 306.06 13.725 306.27 13.795 ;
    RECT 303.2 28.845 303.41 28.915 ;
    RECT 303.2 29.205 303.41 29.275 ;
    RECT 303.2 29.565 303.41 29.635 ;
    RECT 302.74 28.845 302.95 28.915 ;
    RECT 302.74 29.205 302.95 29.275 ;
    RECT 302.74 29.565 302.95 29.635 ;
    RECT 372.92 28.845 373.13 28.915 ;
    RECT 372.92 29.205 373.13 29.275 ;
    RECT 372.92 29.565 373.13 29.635 ;
    RECT 372.46 28.845 372.67 28.915 ;
    RECT 372.46 29.205 372.67 29.275 ;
    RECT 372.46 29.565 372.67 29.635 ;
    RECT 369.6 28.845 369.81 28.915 ;
    RECT 369.6 29.205 369.81 29.275 ;
    RECT 369.6 29.565 369.81 29.635 ;
    RECT 369.14 28.845 369.35 28.915 ;
    RECT 369.14 29.205 369.35 29.275 ;
    RECT 369.14 29.565 369.35 29.635 ;
    RECT 200.605 29.205 200.675 29.275 ;
    RECT 299.88 28.845 300.09 28.915 ;
    RECT 299.88 29.205 300.09 29.275 ;
    RECT 299.88 29.565 300.09 29.635 ;
    RECT 299.42 28.845 299.63 28.915 ;
    RECT 299.42 29.205 299.63 29.275 ;
    RECT 299.42 29.565 299.63 29.635 ;
    RECT 296.56 28.845 296.77 28.915 ;
    RECT 296.56 29.205 296.77 29.275 ;
    RECT 296.56 29.565 296.77 29.635 ;
    RECT 296.1 28.845 296.31 28.915 ;
    RECT 296.1 29.205 296.31 29.275 ;
    RECT 296.1 29.565 296.31 29.635 ;
    RECT 293.24 28.845 293.45 28.915 ;
    RECT 293.24 29.205 293.45 29.275 ;
    RECT 293.24 29.565 293.45 29.635 ;
    RECT 292.78 28.845 292.99 28.915 ;
    RECT 292.78 29.205 292.99 29.275 ;
    RECT 292.78 29.565 292.99 29.635 ;
    RECT 289.92 28.845 290.13 28.915 ;
    RECT 289.92 29.205 290.13 29.275 ;
    RECT 289.92 29.565 290.13 29.635 ;
    RECT 289.46 28.845 289.67 28.915 ;
    RECT 289.46 29.205 289.67 29.275 ;
    RECT 289.46 29.565 289.67 29.635 ;
    RECT 286.6 28.845 286.81 28.915 ;
    RECT 286.6 29.205 286.81 29.275 ;
    RECT 286.6 29.565 286.81 29.635 ;
    RECT 286.14 28.845 286.35 28.915 ;
    RECT 286.14 29.205 286.35 29.275 ;
    RECT 286.14 29.565 286.35 29.635 ;
    RECT 283.28 28.845 283.49 28.915 ;
    RECT 283.28 29.205 283.49 29.275 ;
    RECT 283.28 29.565 283.49 29.635 ;
    RECT 282.82 28.845 283.03 28.915 ;
    RECT 282.82 29.205 283.03 29.275 ;
    RECT 282.82 29.565 283.03 29.635 ;
    RECT 279.96 28.845 280.17 28.915 ;
    RECT 279.96 29.205 280.17 29.275 ;
    RECT 279.96 29.565 280.17 29.635 ;
    RECT 279.5 28.845 279.71 28.915 ;
    RECT 279.5 29.205 279.71 29.275 ;
    RECT 279.5 29.565 279.71 29.635 ;
    RECT 276.64 28.845 276.85 28.915 ;
    RECT 276.64 29.205 276.85 29.275 ;
    RECT 276.64 29.565 276.85 29.635 ;
    RECT 276.18 28.845 276.39 28.915 ;
    RECT 276.18 29.205 276.39 29.275 ;
    RECT 276.18 29.565 276.39 29.635 ;
    RECT 273.32 28.845 273.53 28.915 ;
    RECT 273.32 29.205 273.53 29.275 ;
    RECT 273.32 29.565 273.53 29.635 ;
    RECT 272.86 28.845 273.07 28.915 ;
    RECT 272.86 29.205 273.07 29.275 ;
    RECT 272.86 29.565 273.07 29.635 ;
    RECT 270.0 28.845 270.21 28.915 ;
    RECT 270.0 29.205 270.21 29.275 ;
    RECT 270.0 29.565 270.21 29.635 ;
    RECT 269.54 28.845 269.75 28.915 ;
    RECT 269.54 29.205 269.75 29.275 ;
    RECT 269.54 29.565 269.75 29.635 ;
    RECT 233.48 28.845 233.69 28.915 ;
    RECT 233.48 29.205 233.69 29.275 ;
    RECT 233.48 29.565 233.69 29.635 ;
    RECT 233.02 28.845 233.23 28.915 ;
    RECT 233.02 29.205 233.23 29.275 ;
    RECT 233.02 29.565 233.23 29.635 ;
    RECT 230.16 28.845 230.37 28.915 ;
    RECT 230.16 29.205 230.37 29.275 ;
    RECT 230.16 29.565 230.37 29.635 ;
    RECT 229.7 28.845 229.91 28.915 ;
    RECT 229.7 29.205 229.91 29.275 ;
    RECT 229.7 29.565 229.91 29.635 ;
    RECT 366.28 28.845 366.49 28.915 ;
    RECT 366.28 29.205 366.49 29.275 ;
    RECT 366.28 29.565 366.49 29.635 ;
    RECT 365.82 28.845 366.03 28.915 ;
    RECT 365.82 29.205 366.03 29.275 ;
    RECT 365.82 29.565 366.03 29.635 ;
    RECT 226.84 28.845 227.05 28.915 ;
    RECT 226.84 29.205 227.05 29.275 ;
    RECT 226.84 29.565 227.05 29.635 ;
    RECT 226.38 28.845 226.59 28.915 ;
    RECT 226.38 29.205 226.59 29.275 ;
    RECT 226.38 29.565 226.59 29.635 ;
    RECT 362.96 28.845 363.17 28.915 ;
    RECT 362.96 29.205 363.17 29.275 ;
    RECT 362.96 29.565 363.17 29.635 ;
    RECT 362.5 28.845 362.71 28.915 ;
    RECT 362.5 29.205 362.71 29.275 ;
    RECT 362.5 29.565 362.71 29.635 ;
    RECT 223.52 28.845 223.73 28.915 ;
    RECT 223.52 29.205 223.73 29.275 ;
    RECT 223.52 29.565 223.73 29.635 ;
    RECT 223.06 28.845 223.27 28.915 ;
    RECT 223.06 29.205 223.27 29.275 ;
    RECT 223.06 29.565 223.27 29.635 ;
    RECT 359.64 28.845 359.85 28.915 ;
    RECT 359.64 29.205 359.85 29.275 ;
    RECT 359.64 29.565 359.85 29.635 ;
    RECT 359.18 28.845 359.39 28.915 ;
    RECT 359.18 29.205 359.39 29.275 ;
    RECT 359.18 29.565 359.39 29.635 ;
    RECT 220.2 28.845 220.41 28.915 ;
    RECT 220.2 29.205 220.41 29.275 ;
    RECT 220.2 29.565 220.41 29.635 ;
    RECT 219.74 28.845 219.95 28.915 ;
    RECT 219.74 29.205 219.95 29.275 ;
    RECT 219.74 29.565 219.95 29.635 ;
    RECT 356.32 28.845 356.53 28.915 ;
    RECT 356.32 29.205 356.53 29.275 ;
    RECT 356.32 29.565 356.53 29.635 ;
    RECT 355.86 28.845 356.07 28.915 ;
    RECT 355.86 29.205 356.07 29.275 ;
    RECT 355.86 29.565 356.07 29.635 ;
    RECT 353.0 28.845 353.21 28.915 ;
    RECT 353.0 29.205 353.21 29.275 ;
    RECT 353.0 29.565 353.21 29.635 ;
    RECT 352.54 28.845 352.75 28.915 ;
    RECT 352.54 29.205 352.75 29.275 ;
    RECT 352.54 29.565 352.75 29.635 ;
    RECT 216.88 28.845 217.09 28.915 ;
    RECT 216.88 29.205 217.09 29.275 ;
    RECT 216.88 29.565 217.09 29.635 ;
    RECT 216.42 28.845 216.63 28.915 ;
    RECT 216.42 29.205 216.63 29.275 ;
    RECT 216.42 29.565 216.63 29.635 ;
    RECT 349.68 28.845 349.89 28.915 ;
    RECT 349.68 29.205 349.89 29.275 ;
    RECT 349.68 29.565 349.89 29.635 ;
    RECT 349.22 28.845 349.43 28.915 ;
    RECT 349.22 29.205 349.43 29.275 ;
    RECT 349.22 29.565 349.43 29.635 ;
    RECT 213.56 28.845 213.77 28.915 ;
    RECT 213.56 29.205 213.77 29.275 ;
    RECT 213.56 29.565 213.77 29.635 ;
    RECT 213.1 28.845 213.31 28.915 ;
    RECT 213.1 29.205 213.31 29.275 ;
    RECT 213.1 29.565 213.31 29.635 ;
    RECT 346.36 28.845 346.57 28.915 ;
    RECT 346.36 29.205 346.57 29.275 ;
    RECT 346.36 29.565 346.57 29.635 ;
    RECT 345.9 28.845 346.11 28.915 ;
    RECT 345.9 29.205 346.11 29.275 ;
    RECT 345.9 29.565 346.11 29.635 ;
    RECT 210.24 28.845 210.45 28.915 ;
    RECT 210.24 29.205 210.45 29.275 ;
    RECT 210.24 29.565 210.45 29.635 ;
    RECT 209.78 28.845 209.99 28.915 ;
    RECT 209.78 29.205 209.99 29.275 ;
    RECT 209.78 29.565 209.99 29.635 ;
    RECT 343.04 28.845 343.25 28.915 ;
    RECT 343.04 29.205 343.25 29.275 ;
    RECT 343.04 29.565 343.25 29.635 ;
    RECT 342.58 28.845 342.79 28.915 ;
    RECT 342.58 29.205 342.79 29.275 ;
    RECT 342.58 29.565 342.79 29.635 ;
    RECT 206.92 28.845 207.13 28.915 ;
    RECT 206.92 29.205 207.13 29.275 ;
    RECT 206.92 29.565 207.13 29.635 ;
    RECT 206.46 28.845 206.67 28.915 ;
    RECT 206.46 29.205 206.67 29.275 ;
    RECT 206.46 29.565 206.67 29.635 ;
    RECT 339.72 28.845 339.93 28.915 ;
    RECT 339.72 29.205 339.93 29.275 ;
    RECT 339.72 29.565 339.93 29.635 ;
    RECT 339.26 28.845 339.47 28.915 ;
    RECT 339.26 29.205 339.47 29.275 ;
    RECT 339.26 29.565 339.47 29.635 ;
    RECT 203.6 28.845 203.81 28.915 ;
    RECT 203.6 29.205 203.81 29.275 ;
    RECT 203.6 29.565 203.81 29.635 ;
    RECT 203.14 28.845 203.35 28.915 ;
    RECT 203.14 29.205 203.35 29.275 ;
    RECT 203.14 29.565 203.35 29.635 ;
    RECT 336.4 28.845 336.61 28.915 ;
    RECT 336.4 29.205 336.61 29.275 ;
    RECT 336.4 29.565 336.61 29.635 ;
    RECT 335.94 28.845 336.15 28.915 ;
    RECT 335.94 29.205 336.15 29.275 ;
    RECT 335.94 29.565 336.15 29.635 ;
    RECT 266.68 28.845 266.89 28.915 ;
    RECT 266.68 29.205 266.89 29.275 ;
    RECT 266.68 29.565 266.89 29.635 ;
    RECT 266.22 28.845 266.43 28.915 ;
    RECT 266.22 29.205 266.43 29.275 ;
    RECT 266.22 29.565 266.43 29.635 ;
    RECT 263.36 28.845 263.57 28.915 ;
    RECT 263.36 29.205 263.57 29.275 ;
    RECT 263.36 29.565 263.57 29.635 ;
    RECT 262.9 28.845 263.11 28.915 ;
    RECT 262.9 29.205 263.11 29.275 ;
    RECT 262.9 29.565 263.11 29.635 ;
    RECT 260.04 28.845 260.25 28.915 ;
    RECT 260.04 29.205 260.25 29.275 ;
    RECT 260.04 29.565 260.25 29.635 ;
    RECT 259.58 28.845 259.79 28.915 ;
    RECT 259.58 29.205 259.79 29.275 ;
    RECT 259.58 29.565 259.79 29.635 ;
    RECT 256.72 28.845 256.93 28.915 ;
    RECT 256.72 29.205 256.93 29.275 ;
    RECT 256.72 29.565 256.93 29.635 ;
    RECT 256.26 28.845 256.47 28.915 ;
    RECT 256.26 29.205 256.47 29.275 ;
    RECT 256.26 29.565 256.47 29.635 ;
    RECT 253.4 28.845 253.61 28.915 ;
    RECT 253.4 29.205 253.61 29.275 ;
    RECT 253.4 29.565 253.61 29.635 ;
    RECT 252.94 28.845 253.15 28.915 ;
    RECT 252.94 29.205 253.15 29.275 ;
    RECT 252.94 29.565 253.15 29.635 ;
    RECT 250.08 28.845 250.29 28.915 ;
    RECT 250.08 29.205 250.29 29.275 ;
    RECT 250.08 29.565 250.29 29.635 ;
    RECT 249.62 28.845 249.83 28.915 ;
    RECT 249.62 29.205 249.83 29.275 ;
    RECT 249.62 29.565 249.83 29.635 ;
    RECT 246.76 28.845 246.97 28.915 ;
    RECT 246.76 29.205 246.97 29.275 ;
    RECT 246.76 29.565 246.97 29.635 ;
    RECT 246.3 28.845 246.51 28.915 ;
    RECT 246.3 29.205 246.51 29.275 ;
    RECT 246.3 29.565 246.51 29.635 ;
    RECT 243.44 28.845 243.65 28.915 ;
    RECT 243.44 29.205 243.65 29.275 ;
    RECT 243.44 29.565 243.65 29.635 ;
    RECT 242.98 28.845 243.19 28.915 ;
    RECT 242.98 29.205 243.19 29.275 ;
    RECT 242.98 29.565 243.19 29.635 ;
    RECT 240.12 28.845 240.33 28.915 ;
    RECT 240.12 29.205 240.33 29.275 ;
    RECT 240.12 29.565 240.33 29.635 ;
    RECT 239.66 28.845 239.87 28.915 ;
    RECT 239.66 29.205 239.87 29.275 ;
    RECT 239.66 29.565 239.87 29.635 ;
    RECT 236.8 28.845 237.01 28.915 ;
    RECT 236.8 29.205 237.01 29.275 ;
    RECT 236.8 29.565 237.01 29.635 ;
    RECT 236.34 28.845 236.55 28.915 ;
    RECT 236.34 29.205 236.55 29.275 ;
    RECT 236.34 29.565 236.55 29.635 ;
    RECT 374.15 29.205 374.22 29.275 ;
    RECT 333.08 28.845 333.29 28.915 ;
    RECT 333.08 29.205 333.29 29.275 ;
    RECT 333.08 29.565 333.29 29.635 ;
    RECT 332.62 28.845 332.83 28.915 ;
    RECT 332.62 29.205 332.83 29.275 ;
    RECT 332.62 29.565 332.83 29.635 ;
    RECT 329.76 28.845 329.97 28.915 ;
    RECT 329.76 29.205 329.97 29.275 ;
    RECT 329.76 29.565 329.97 29.635 ;
    RECT 329.3 28.845 329.51 28.915 ;
    RECT 329.3 29.205 329.51 29.275 ;
    RECT 329.3 29.565 329.51 29.635 ;
    RECT 326.44 28.845 326.65 28.915 ;
    RECT 326.44 29.205 326.65 29.275 ;
    RECT 326.44 29.565 326.65 29.635 ;
    RECT 325.98 28.845 326.19 28.915 ;
    RECT 325.98 29.205 326.19 29.275 ;
    RECT 325.98 29.565 326.19 29.635 ;
    RECT 323.12 28.845 323.33 28.915 ;
    RECT 323.12 29.205 323.33 29.275 ;
    RECT 323.12 29.565 323.33 29.635 ;
    RECT 322.66 28.845 322.87 28.915 ;
    RECT 322.66 29.205 322.87 29.275 ;
    RECT 322.66 29.565 322.87 29.635 ;
    RECT 319.8 28.845 320.01 28.915 ;
    RECT 319.8 29.205 320.01 29.275 ;
    RECT 319.8 29.565 320.01 29.635 ;
    RECT 319.34 28.845 319.55 28.915 ;
    RECT 319.34 29.205 319.55 29.275 ;
    RECT 319.34 29.565 319.55 29.635 ;
    RECT 316.48 28.845 316.69 28.915 ;
    RECT 316.48 29.205 316.69 29.275 ;
    RECT 316.48 29.565 316.69 29.635 ;
    RECT 316.02 28.845 316.23 28.915 ;
    RECT 316.02 29.205 316.23 29.275 ;
    RECT 316.02 29.565 316.23 29.635 ;
    RECT 313.16 28.845 313.37 28.915 ;
    RECT 313.16 29.205 313.37 29.275 ;
    RECT 313.16 29.565 313.37 29.635 ;
    RECT 312.7 28.845 312.91 28.915 ;
    RECT 312.7 29.205 312.91 29.275 ;
    RECT 312.7 29.565 312.91 29.635 ;
    RECT 309.84 28.845 310.05 28.915 ;
    RECT 309.84 29.205 310.05 29.275 ;
    RECT 309.84 29.565 310.05 29.635 ;
    RECT 309.38 28.845 309.59 28.915 ;
    RECT 309.38 29.205 309.59 29.275 ;
    RECT 309.38 29.565 309.59 29.635 ;
    RECT 306.52 28.845 306.73 28.915 ;
    RECT 306.52 29.205 306.73 29.275 ;
    RECT 306.52 29.565 306.73 29.635 ;
    RECT 306.06 28.845 306.27 28.915 ;
    RECT 306.06 29.205 306.27 29.275 ;
    RECT 306.06 29.565 306.27 29.635 ;
    RECT 303.2 12.285 303.41 12.355 ;
    RECT 303.2 12.645 303.41 12.715 ;
    RECT 303.2 13.005 303.41 13.075 ;
    RECT 302.74 12.285 302.95 12.355 ;
    RECT 302.74 12.645 302.95 12.715 ;
    RECT 302.74 13.005 302.95 13.075 ;
    RECT 372.92 12.285 373.13 12.355 ;
    RECT 372.92 12.645 373.13 12.715 ;
    RECT 372.92 13.005 373.13 13.075 ;
    RECT 372.46 12.285 372.67 12.355 ;
    RECT 372.46 12.645 372.67 12.715 ;
    RECT 372.46 13.005 372.67 13.075 ;
    RECT 369.6 12.285 369.81 12.355 ;
    RECT 369.6 12.645 369.81 12.715 ;
    RECT 369.6 13.005 369.81 13.075 ;
    RECT 369.14 12.285 369.35 12.355 ;
    RECT 369.14 12.645 369.35 12.715 ;
    RECT 369.14 13.005 369.35 13.075 ;
    RECT 200.605 12.645 200.675 12.715 ;
    RECT 299.88 12.285 300.09 12.355 ;
    RECT 299.88 12.645 300.09 12.715 ;
    RECT 299.88 13.005 300.09 13.075 ;
    RECT 299.42 12.285 299.63 12.355 ;
    RECT 299.42 12.645 299.63 12.715 ;
    RECT 299.42 13.005 299.63 13.075 ;
    RECT 296.56 12.285 296.77 12.355 ;
    RECT 296.56 12.645 296.77 12.715 ;
    RECT 296.56 13.005 296.77 13.075 ;
    RECT 296.1 12.285 296.31 12.355 ;
    RECT 296.1 12.645 296.31 12.715 ;
    RECT 296.1 13.005 296.31 13.075 ;
    RECT 293.24 12.285 293.45 12.355 ;
    RECT 293.24 12.645 293.45 12.715 ;
    RECT 293.24 13.005 293.45 13.075 ;
    RECT 292.78 12.285 292.99 12.355 ;
    RECT 292.78 12.645 292.99 12.715 ;
    RECT 292.78 13.005 292.99 13.075 ;
    RECT 289.92 12.285 290.13 12.355 ;
    RECT 289.92 12.645 290.13 12.715 ;
    RECT 289.92 13.005 290.13 13.075 ;
    RECT 289.46 12.285 289.67 12.355 ;
    RECT 289.46 12.645 289.67 12.715 ;
    RECT 289.46 13.005 289.67 13.075 ;
    RECT 286.6 12.285 286.81 12.355 ;
    RECT 286.6 12.645 286.81 12.715 ;
    RECT 286.6 13.005 286.81 13.075 ;
    RECT 286.14 12.285 286.35 12.355 ;
    RECT 286.14 12.645 286.35 12.715 ;
    RECT 286.14 13.005 286.35 13.075 ;
    RECT 283.28 12.285 283.49 12.355 ;
    RECT 283.28 12.645 283.49 12.715 ;
    RECT 283.28 13.005 283.49 13.075 ;
    RECT 282.82 12.285 283.03 12.355 ;
    RECT 282.82 12.645 283.03 12.715 ;
    RECT 282.82 13.005 283.03 13.075 ;
    RECT 279.96 12.285 280.17 12.355 ;
    RECT 279.96 12.645 280.17 12.715 ;
    RECT 279.96 13.005 280.17 13.075 ;
    RECT 279.5 12.285 279.71 12.355 ;
    RECT 279.5 12.645 279.71 12.715 ;
    RECT 279.5 13.005 279.71 13.075 ;
    RECT 276.64 12.285 276.85 12.355 ;
    RECT 276.64 12.645 276.85 12.715 ;
    RECT 276.64 13.005 276.85 13.075 ;
    RECT 276.18 12.285 276.39 12.355 ;
    RECT 276.18 12.645 276.39 12.715 ;
    RECT 276.18 13.005 276.39 13.075 ;
    RECT 273.32 12.285 273.53 12.355 ;
    RECT 273.32 12.645 273.53 12.715 ;
    RECT 273.32 13.005 273.53 13.075 ;
    RECT 272.86 12.285 273.07 12.355 ;
    RECT 272.86 12.645 273.07 12.715 ;
    RECT 272.86 13.005 273.07 13.075 ;
    RECT 270.0 12.285 270.21 12.355 ;
    RECT 270.0 12.645 270.21 12.715 ;
    RECT 270.0 13.005 270.21 13.075 ;
    RECT 269.54 12.285 269.75 12.355 ;
    RECT 269.54 12.645 269.75 12.715 ;
    RECT 269.54 13.005 269.75 13.075 ;
    RECT 233.48 12.285 233.69 12.355 ;
    RECT 233.48 12.645 233.69 12.715 ;
    RECT 233.48 13.005 233.69 13.075 ;
    RECT 233.02 12.285 233.23 12.355 ;
    RECT 233.02 12.645 233.23 12.715 ;
    RECT 233.02 13.005 233.23 13.075 ;
    RECT 230.16 12.285 230.37 12.355 ;
    RECT 230.16 12.645 230.37 12.715 ;
    RECT 230.16 13.005 230.37 13.075 ;
    RECT 229.7 12.285 229.91 12.355 ;
    RECT 229.7 12.645 229.91 12.715 ;
    RECT 229.7 13.005 229.91 13.075 ;
    RECT 366.28 12.285 366.49 12.355 ;
    RECT 366.28 12.645 366.49 12.715 ;
    RECT 366.28 13.005 366.49 13.075 ;
    RECT 365.82 12.285 366.03 12.355 ;
    RECT 365.82 12.645 366.03 12.715 ;
    RECT 365.82 13.005 366.03 13.075 ;
    RECT 226.84 12.285 227.05 12.355 ;
    RECT 226.84 12.645 227.05 12.715 ;
    RECT 226.84 13.005 227.05 13.075 ;
    RECT 226.38 12.285 226.59 12.355 ;
    RECT 226.38 12.645 226.59 12.715 ;
    RECT 226.38 13.005 226.59 13.075 ;
    RECT 362.96 12.285 363.17 12.355 ;
    RECT 362.96 12.645 363.17 12.715 ;
    RECT 362.96 13.005 363.17 13.075 ;
    RECT 362.5 12.285 362.71 12.355 ;
    RECT 362.5 12.645 362.71 12.715 ;
    RECT 362.5 13.005 362.71 13.075 ;
    RECT 223.52 12.285 223.73 12.355 ;
    RECT 223.52 12.645 223.73 12.715 ;
    RECT 223.52 13.005 223.73 13.075 ;
    RECT 223.06 12.285 223.27 12.355 ;
    RECT 223.06 12.645 223.27 12.715 ;
    RECT 223.06 13.005 223.27 13.075 ;
    RECT 359.64 12.285 359.85 12.355 ;
    RECT 359.64 12.645 359.85 12.715 ;
    RECT 359.64 13.005 359.85 13.075 ;
    RECT 359.18 12.285 359.39 12.355 ;
    RECT 359.18 12.645 359.39 12.715 ;
    RECT 359.18 13.005 359.39 13.075 ;
    RECT 220.2 12.285 220.41 12.355 ;
    RECT 220.2 12.645 220.41 12.715 ;
    RECT 220.2 13.005 220.41 13.075 ;
    RECT 219.74 12.285 219.95 12.355 ;
    RECT 219.74 12.645 219.95 12.715 ;
    RECT 219.74 13.005 219.95 13.075 ;
    RECT 356.32 12.285 356.53 12.355 ;
    RECT 356.32 12.645 356.53 12.715 ;
    RECT 356.32 13.005 356.53 13.075 ;
    RECT 355.86 12.285 356.07 12.355 ;
    RECT 355.86 12.645 356.07 12.715 ;
    RECT 355.86 13.005 356.07 13.075 ;
    RECT 353.0 12.285 353.21 12.355 ;
    RECT 353.0 12.645 353.21 12.715 ;
    RECT 353.0 13.005 353.21 13.075 ;
    RECT 352.54 12.285 352.75 12.355 ;
    RECT 352.54 12.645 352.75 12.715 ;
    RECT 352.54 13.005 352.75 13.075 ;
    RECT 216.88 12.285 217.09 12.355 ;
    RECT 216.88 12.645 217.09 12.715 ;
    RECT 216.88 13.005 217.09 13.075 ;
    RECT 216.42 12.285 216.63 12.355 ;
    RECT 216.42 12.645 216.63 12.715 ;
    RECT 216.42 13.005 216.63 13.075 ;
    RECT 349.68 12.285 349.89 12.355 ;
    RECT 349.68 12.645 349.89 12.715 ;
    RECT 349.68 13.005 349.89 13.075 ;
    RECT 349.22 12.285 349.43 12.355 ;
    RECT 349.22 12.645 349.43 12.715 ;
    RECT 349.22 13.005 349.43 13.075 ;
    RECT 213.56 12.285 213.77 12.355 ;
    RECT 213.56 12.645 213.77 12.715 ;
    RECT 213.56 13.005 213.77 13.075 ;
    RECT 213.1 12.285 213.31 12.355 ;
    RECT 213.1 12.645 213.31 12.715 ;
    RECT 213.1 13.005 213.31 13.075 ;
    RECT 346.36 12.285 346.57 12.355 ;
    RECT 346.36 12.645 346.57 12.715 ;
    RECT 346.36 13.005 346.57 13.075 ;
    RECT 345.9 12.285 346.11 12.355 ;
    RECT 345.9 12.645 346.11 12.715 ;
    RECT 345.9 13.005 346.11 13.075 ;
    RECT 210.24 12.285 210.45 12.355 ;
    RECT 210.24 12.645 210.45 12.715 ;
    RECT 210.24 13.005 210.45 13.075 ;
    RECT 209.78 12.285 209.99 12.355 ;
    RECT 209.78 12.645 209.99 12.715 ;
    RECT 209.78 13.005 209.99 13.075 ;
    RECT 343.04 12.285 343.25 12.355 ;
    RECT 343.04 12.645 343.25 12.715 ;
    RECT 343.04 13.005 343.25 13.075 ;
    RECT 342.58 12.285 342.79 12.355 ;
    RECT 342.58 12.645 342.79 12.715 ;
    RECT 342.58 13.005 342.79 13.075 ;
    RECT 206.92 12.285 207.13 12.355 ;
    RECT 206.92 12.645 207.13 12.715 ;
    RECT 206.92 13.005 207.13 13.075 ;
    RECT 206.46 12.285 206.67 12.355 ;
    RECT 206.46 12.645 206.67 12.715 ;
    RECT 206.46 13.005 206.67 13.075 ;
    RECT 339.72 12.285 339.93 12.355 ;
    RECT 339.72 12.645 339.93 12.715 ;
    RECT 339.72 13.005 339.93 13.075 ;
    RECT 339.26 12.285 339.47 12.355 ;
    RECT 339.26 12.645 339.47 12.715 ;
    RECT 339.26 13.005 339.47 13.075 ;
    RECT 203.6 12.285 203.81 12.355 ;
    RECT 203.6 12.645 203.81 12.715 ;
    RECT 203.6 13.005 203.81 13.075 ;
    RECT 203.14 12.285 203.35 12.355 ;
    RECT 203.14 12.645 203.35 12.715 ;
    RECT 203.14 13.005 203.35 13.075 ;
    RECT 336.4 12.285 336.61 12.355 ;
    RECT 336.4 12.645 336.61 12.715 ;
    RECT 336.4 13.005 336.61 13.075 ;
    RECT 335.94 12.285 336.15 12.355 ;
    RECT 335.94 12.645 336.15 12.715 ;
    RECT 335.94 13.005 336.15 13.075 ;
    RECT 266.68 12.285 266.89 12.355 ;
    RECT 266.68 12.645 266.89 12.715 ;
    RECT 266.68 13.005 266.89 13.075 ;
    RECT 266.22 12.285 266.43 12.355 ;
    RECT 266.22 12.645 266.43 12.715 ;
    RECT 266.22 13.005 266.43 13.075 ;
    RECT 263.36 12.285 263.57 12.355 ;
    RECT 263.36 12.645 263.57 12.715 ;
    RECT 263.36 13.005 263.57 13.075 ;
    RECT 262.9 12.285 263.11 12.355 ;
    RECT 262.9 12.645 263.11 12.715 ;
    RECT 262.9 13.005 263.11 13.075 ;
    RECT 260.04 12.285 260.25 12.355 ;
    RECT 260.04 12.645 260.25 12.715 ;
    RECT 260.04 13.005 260.25 13.075 ;
    RECT 259.58 12.285 259.79 12.355 ;
    RECT 259.58 12.645 259.79 12.715 ;
    RECT 259.58 13.005 259.79 13.075 ;
    RECT 256.72 12.285 256.93 12.355 ;
    RECT 256.72 12.645 256.93 12.715 ;
    RECT 256.72 13.005 256.93 13.075 ;
    RECT 256.26 12.285 256.47 12.355 ;
    RECT 256.26 12.645 256.47 12.715 ;
    RECT 256.26 13.005 256.47 13.075 ;
    RECT 253.4 12.285 253.61 12.355 ;
    RECT 253.4 12.645 253.61 12.715 ;
    RECT 253.4 13.005 253.61 13.075 ;
    RECT 252.94 12.285 253.15 12.355 ;
    RECT 252.94 12.645 253.15 12.715 ;
    RECT 252.94 13.005 253.15 13.075 ;
    RECT 250.08 12.285 250.29 12.355 ;
    RECT 250.08 12.645 250.29 12.715 ;
    RECT 250.08 13.005 250.29 13.075 ;
    RECT 249.62 12.285 249.83 12.355 ;
    RECT 249.62 12.645 249.83 12.715 ;
    RECT 249.62 13.005 249.83 13.075 ;
    RECT 246.76 12.285 246.97 12.355 ;
    RECT 246.76 12.645 246.97 12.715 ;
    RECT 246.76 13.005 246.97 13.075 ;
    RECT 246.3 12.285 246.51 12.355 ;
    RECT 246.3 12.645 246.51 12.715 ;
    RECT 246.3 13.005 246.51 13.075 ;
    RECT 243.44 12.285 243.65 12.355 ;
    RECT 243.44 12.645 243.65 12.715 ;
    RECT 243.44 13.005 243.65 13.075 ;
    RECT 242.98 12.285 243.19 12.355 ;
    RECT 242.98 12.645 243.19 12.715 ;
    RECT 242.98 13.005 243.19 13.075 ;
    RECT 240.12 12.285 240.33 12.355 ;
    RECT 240.12 12.645 240.33 12.715 ;
    RECT 240.12 13.005 240.33 13.075 ;
    RECT 239.66 12.285 239.87 12.355 ;
    RECT 239.66 12.645 239.87 12.715 ;
    RECT 239.66 13.005 239.87 13.075 ;
    RECT 236.8 12.285 237.01 12.355 ;
    RECT 236.8 12.645 237.01 12.715 ;
    RECT 236.8 13.005 237.01 13.075 ;
    RECT 236.34 12.285 236.55 12.355 ;
    RECT 236.34 12.645 236.55 12.715 ;
    RECT 236.34 13.005 236.55 13.075 ;
    RECT 374.15 12.645 374.22 12.715 ;
    RECT 333.08 12.285 333.29 12.355 ;
    RECT 333.08 12.645 333.29 12.715 ;
    RECT 333.08 13.005 333.29 13.075 ;
    RECT 332.62 12.285 332.83 12.355 ;
    RECT 332.62 12.645 332.83 12.715 ;
    RECT 332.62 13.005 332.83 13.075 ;
    RECT 329.76 12.285 329.97 12.355 ;
    RECT 329.76 12.645 329.97 12.715 ;
    RECT 329.76 13.005 329.97 13.075 ;
    RECT 329.3 12.285 329.51 12.355 ;
    RECT 329.3 12.645 329.51 12.715 ;
    RECT 329.3 13.005 329.51 13.075 ;
    RECT 326.44 12.285 326.65 12.355 ;
    RECT 326.44 12.645 326.65 12.715 ;
    RECT 326.44 13.005 326.65 13.075 ;
    RECT 325.98 12.285 326.19 12.355 ;
    RECT 325.98 12.645 326.19 12.715 ;
    RECT 325.98 13.005 326.19 13.075 ;
    RECT 323.12 12.285 323.33 12.355 ;
    RECT 323.12 12.645 323.33 12.715 ;
    RECT 323.12 13.005 323.33 13.075 ;
    RECT 322.66 12.285 322.87 12.355 ;
    RECT 322.66 12.645 322.87 12.715 ;
    RECT 322.66 13.005 322.87 13.075 ;
    RECT 319.8 12.285 320.01 12.355 ;
    RECT 319.8 12.645 320.01 12.715 ;
    RECT 319.8 13.005 320.01 13.075 ;
    RECT 319.34 12.285 319.55 12.355 ;
    RECT 319.34 12.645 319.55 12.715 ;
    RECT 319.34 13.005 319.55 13.075 ;
    RECT 316.48 12.285 316.69 12.355 ;
    RECT 316.48 12.645 316.69 12.715 ;
    RECT 316.48 13.005 316.69 13.075 ;
    RECT 316.02 12.285 316.23 12.355 ;
    RECT 316.02 12.645 316.23 12.715 ;
    RECT 316.02 13.005 316.23 13.075 ;
    RECT 313.16 12.285 313.37 12.355 ;
    RECT 313.16 12.645 313.37 12.715 ;
    RECT 313.16 13.005 313.37 13.075 ;
    RECT 312.7 12.285 312.91 12.355 ;
    RECT 312.7 12.645 312.91 12.715 ;
    RECT 312.7 13.005 312.91 13.075 ;
    RECT 309.84 12.285 310.05 12.355 ;
    RECT 309.84 12.645 310.05 12.715 ;
    RECT 309.84 13.005 310.05 13.075 ;
    RECT 309.38 12.285 309.59 12.355 ;
    RECT 309.38 12.645 309.59 12.715 ;
    RECT 309.38 13.005 309.59 13.075 ;
    RECT 306.52 12.285 306.73 12.355 ;
    RECT 306.52 12.645 306.73 12.715 ;
    RECT 306.52 13.005 306.73 13.075 ;
    RECT 306.06 12.285 306.27 12.355 ;
    RECT 306.06 12.645 306.27 12.715 ;
    RECT 306.06 13.005 306.27 13.075 ;
    RECT 303.2 28.125 303.41 28.195 ;
    RECT 303.2 28.485 303.41 28.555 ;
    RECT 303.2 28.845 303.41 28.915 ;
    RECT 302.74 28.125 302.95 28.195 ;
    RECT 302.74 28.485 302.95 28.555 ;
    RECT 302.74 28.845 302.95 28.915 ;
    RECT 372.92 28.125 373.13 28.195 ;
    RECT 372.92 28.485 373.13 28.555 ;
    RECT 372.92 28.845 373.13 28.915 ;
    RECT 372.46 28.125 372.67 28.195 ;
    RECT 372.46 28.485 372.67 28.555 ;
    RECT 372.46 28.845 372.67 28.915 ;
    RECT 369.6 28.125 369.81 28.195 ;
    RECT 369.6 28.485 369.81 28.555 ;
    RECT 369.6 28.845 369.81 28.915 ;
    RECT 369.14 28.125 369.35 28.195 ;
    RECT 369.14 28.485 369.35 28.555 ;
    RECT 369.14 28.845 369.35 28.915 ;
    RECT 200.605 28.485 200.675 28.555 ;
    RECT 299.88 28.125 300.09 28.195 ;
    RECT 299.88 28.485 300.09 28.555 ;
    RECT 299.88 28.845 300.09 28.915 ;
    RECT 299.42 28.125 299.63 28.195 ;
    RECT 299.42 28.485 299.63 28.555 ;
    RECT 299.42 28.845 299.63 28.915 ;
    RECT 296.56 28.125 296.77 28.195 ;
    RECT 296.56 28.485 296.77 28.555 ;
    RECT 296.56 28.845 296.77 28.915 ;
    RECT 296.1 28.125 296.31 28.195 ;
    RECT 296.1 28.485 296.31 28.555 ;
    RECT 296.1 28.845 296.31 28.915 ;
    RECT 293.24 28.125 293.45 28.195 ;
    RECT 293.24 28.485 293.45 28.555 ;
    RECT 293.24 28.845 293.45 28.915 ;
    RECT 292.78 28.125 292.99 28.195 ;
    RECT 292.78 28.485 292.99 28.555 ;
    RECT 292.78 28.845 292.99 28.915 ;
    RECT 289.92 28.125 290.13 28.195 ;
    RECT 289.92 28.485 290.13 28.555 ;
    RECT 289.92 28.845 290.13 28.915 ;
    RECT 289.46 28.125 289.67 28.195 ;
    RECT 289.46 28.485 289.67 28.555 ;
    RECT 289.46 28.845 289.67 28.915 ;
    RECT 286.6 28.125 286.81 28.195 ;
    RECT 286.6 28.485 286.81 28.555 ;
    RECT 286.6 28.845 286.81 28.915 ;
    RECT 286.14 28.125 286.35 28.195 ;
    RECT 286.14 28.485 286.35 28.555 ;
    RECT 286.14 28.845 286.35 28.915 ;
    RECT 283.28 28.125 283.49 28.195 ;
    RECT 283.28 28.485 283.49 28.555 ;
    RECT 283.28 28.845 283.49 28.915 ;
    RECT 282.82 28.125 283.03 28.195 ;
    RECT 282.82 28.485 283.03 28.555 ;
    RECT 282.82 28.845 283.03 28.915 ;
    RECT 279.96 28.125 280.17 28.195 ;
    RECT 279.96 28.485 280.17 28.555 ;
    RECT 279.96 28.845 280.17 28.915 ;
    RECT 279.5 28.125 279.71 28.195 ;
    RECT 279.5 28.485 279.71 28.555 ;
    RECT 279.5 28.845 279.71 28.915 ;
    RECT 276.64 28.125 276.85 28.195 ;
    RECT 276.64 28.485 276.85 28.555 ;
    RECT 276.64 28.845 276.85 28.915 ;
    RECT 276.18 28.125 276.39 28.195 ;
    RECT 276.18 28.485 276.39 28.555 ;
    RECT 276.18 28.845 276.39 28.915 ;
    RECT 273.32 28.125 273.53 28.195 ;
    RECT 273.32 28.485 273.53 28.555 ;
    RECT 273.32 28.845 273.53 28.915 ;
    RECT 272.86 28.125 273.07 28.195 ;
    RECT 272.86 28.485 273.07 28.555 ;
    RECT 272.86 28.845 273.07 28.915 ;
    RECT 270.0 28.125 270.21 28.195 ;
    RECT 270.0 28.485 270.21 28.555 ;
    RECT 270.0 28.845 270.21 28.915 ;
    RECT 269.54 28.125 269.75 28.195 ;
    RECT 269.54 28.485 269.75 28.555 ;
    RECT 269.54 28.845 269.75 28.915 ;
    RECT 233.48 28.125 233.69 28.195 ;
    RECT 233.48 28.485 233.69 28.555 ;
    RECT 233.48 28.845 233.69 28.915 ;
    RECT 233.02 28.125 233.23 28.195 ;
    RECT 233.02 28.485 233.23 28.555 ;
    RECT 233.02 28.845 233.23 28.915 ;
    RECT 230.16 28.125 230.37 28.195 ;
    RECT 230.16 28.485 230.37 28.555 ;
    RECT 230.16 28.845 230.37 28.915 ;
    RECT 229.7 28.125 229.91 28.195 ;
    RECT 229.7 28.485 229.91 28.555 ;
    RECT 229.7 28.845 229.91 28.915 ;
    RECT 366.28 28.125 366.49 28.195 ;
    RECT 366.28 28.485 366.49 28.555 ;
    RECT 366.28 28.845 366.49 28.915 ;
    RECT 365.82 28.125 366.03 28.195 ;
    RECT 365.82 28.485 366.03 28.555 ;
    RECT 365.82 28.845 366.03 28.915 ;
    RECT 226.84 28.125 227.05 28.195 ;
    RECT 226.84 28.485 227.05 28.555 ;
    RECT 226.84 28.845 227.05 28.915 ;
    RECT 226.38 28.125 226.59 28.195 ;
    RECT 226.38 28.485 226.59 28.555 ;
    RECT 226.38 28.845 226.59 28.915 ;
    RECT 362.96 28.125 363.17 28.195 ;
    RECT 362.96 28.485 363.17 28.555 ;
    RECT 362.96 28.845 363.17 28.915 ;
    RECT 362.5 28.125 362.71 28.195 ;
    RECT 362.5 28.485 362.71 28.555 ;
    RECT 362.5 28.845 362.71 28.915 ;
    RECT 223.52 28.125 223.73 28.195 ;
    RECT 223.52 28.485 223.73 28.555 ;
    RECT 223.52 28.845 223.73 28.915 ;
    RECT 223.06 28.125 223.27 28.195 ;
    RECT 223.06 28.485 223.27 28.555 ;
    RECT 223.06 28.845 223.27 28.915 ;
    RECT 359.64 28.125 359.85 28.195 ;
    RECT 359.64 28.485 359.85 28.555 ;
    RECT 359.64 28.845 359.85 28.915 ;
    RECT 359.18 28.125 359.39 28.195 ;
    RECT 359.18 28.485 359.39 28.555 ;
    RECT 359.18 28.845 359.39 28.915 ;
    RECT 220.2 28.125 220.41 28.195 ;
    RECT 220.2 28.485 220.41 28.555 ;
    RECT 220.2 28.845 220.41 28.915 ;
    RECT 219.74 28.125 219.95 28.195 ;
    RECT 219.74 28.485 219.95 28.555 ;
    RECT 219.74 28.845 219.95 28.915 ;
    RECT 356.32 28.125 356.53 28.195 ;
    RECT 356.32 28.485 356.53 28.555 ;
    RECT 356.32 28.845 356.53 28.915 ;
    RECT 355.86 28.125 356.07 28.195 ;
    RECT 355.86 28.485 356.07 28.555 ;
    RECT 355.86 28.845 356.07 28.915 ;
    RECT 353.0 28.125 353.21 28.195 ;
    RECT 353.0 28.485 353.21 28.555 ;
    RECT 353.0 28.845 353.21 28.915 ;
    RECT 352.54 28.125 352.75 28.195 ;
    RECT 352.54 28.485 352.75 28.555 ;
    RECT 352.54 28.845 352.75 28.915 ;
    RECT 216.88 28.125 217.09 28.195 ;
    RECT 216.88 28.485 217.09 28.555 ;
    RECT 216.88 28.845 217.09 28.915 ;
    RECT 216.42 28.125 216.63 28.195 ;
    RECT 216.42 28.485 216.63 28.555 ;
    RECT 216.42 28.845 216.63 28.915 ;
    RECT 349.68 28.125 349.89 28.195 ;
    RECT 349.68 28.485 349.89 28.555 ;
    RECT 349.68 28.845 349.89 28.915 ;
    RECT 349.22 28.125 349.43 28.195 ;
    RECT 349.22 28.485 349.43 28.555 ;
    RECT 349.22 28.845 349.43 28.915 ;
    RECT 213.56 28.125 213.77 28.195 ;
    RECT 213.56 28.485 213.77 28.555 ;
    RECT 213.56 28.845 213.77 28.915 ;
    RECT 213.1 28.125 213.31 28.195 ;
    RECT 213.1 28.485 213.31 28.555 ;
    RECT 213.1 28.845 213.31 28.915 ;
    RECT 346.36 28.125 346.57 28.195 ;
    RECT 346.36 28.485 346.57 28.555 ;
    RECT 346.36 28.845 346.57 28.915 ;
    RECT 345.9 28.125 346.11 28.195 ;
    RECT 345.9 28.485 346.11 28.555 ;
    RECT 345.9 28.845 346.11 28.915 ;
    RECT 210.24 28.125 210.45 28.195 ;
    RECT 210.24 28.485 210.45 28.555 ;
    RECT 210.24 28.845 210.45 28.915 ;
    RECT 209.78 28.125 209.99 28.195 ;
    RECT 209.78 28.485 209.99 28.555 ;
    RECT 209.78 28.845 209.99 28.915 ;
    RECT 343.04 28.125 343.25 28.195 ;
    RECT 343.04 28.485 343.25 28.555 ;
    RECT 343.04 28.845 343.25 28.915 ;
    RECT 342.58 28.125 342.79 28.195 ;
    RECT 342.58 28.485 342.79 28.555 ;
    RECT 342.58 28.845 342.79 28.915 ;
    RECT 206.92 28.125 207.13 28.195 ;
    RECT 206.92 28.485 207.13 28.555 ;
    RECT 206.92 28.845 207.13 28.915 ;
    RECT 206.46 28.125 206.67 28.195 ;
    RECT 206.46 28.485 206.67 28.555 ;
    RECT 206.46 28.845 206.67 28.915 ;
    RECT 339.72 28.125 339.93 28.195 ;
    RECT 339.72 28.485 339.93 28.555 ;
    RECT 339.72 28.845 339.93 28.915 ;
    RECT 339.26 28.125 339.47 28.195 ;
    RECT 339.26 28.485 339.47 28.555 ;
    RECT 339.26 28.845 339.47 28.915 ;
    RECT 203.6 28.125 203.81 28.195 ;
    RECT 203.6 28.485 203.81 28.555 ;
    RECT 203.6 28.845 203.81 28.915 ;
    RECT 203.14 28.125 203.35 28.195 ;
    RECT 203.14 28.485 203.35 28.555 ;
    RECT 203.14 28.845 203.35 28.915 ;
    RECT 336.4 28.125 336.61 28.195 ;
    RECT 336.4 28.485 336.61 28.555 ;
    RECT 336.4 28.845 336.61 28.915 ;
    RECT 335.94 28.125 336.15 28.195 ;
    RECT 335.94 28.485 336.15 28.555 ;
    RECT 335.94 28.845 336.15 28.915 ;
    RECT 266.68 28.125 266.89 28.195 ;
    RECT 266.68 28.485 266.89 28.555 ;
    RECT 266.68 28.845 266.89 28.915 ;
    RECT 266.22 28.125 266.43 28.195 ;
    RECT 266.22 28.485 266.43 28.555 ;
    RECT 266.22 28.845 266.43 28.915 ;
    RECT 263.36 28.125 263.57 28.195 ;
    RECT 263.36 28.485 263.57 28.555 ;
    RECT 263.36 28.845 263.57 28.915 ;
    RECT 262.9 28.125 263.11 28.195 ;
    RECT 262.9 28.485 263.11 28.555 ;
    RECT 262.9 28.845 263.11 28.915 ;
    RECT 260.04 28.125 260.25 28.195 ;
    RECT 260.04 28.485 260.25 28.555 ;
    RECT 260.04 28.845 260.25 28.915 ;
    RECT 259.58 28.125 259.79 28.195 ;
    RECT 259.58 28.485 259.79 28.555 ;
    RECT 259.58 28.845 259.79 28.915 ;
    RECT 256.72 28.125 256.93 28.195 ;
    RECT 256.72 28.485 256.93 28.555 ;
    RECT 256.72 28.845 256.93 28.915 ;
    RECT 256.26 28.125 256.47 28.195 ;
    RECT 256.26 28.485 256.47 28.555 ;
    RECT 256.26 28.845 256.47 28.915 ;
    RECT 253.4 28.125 253.61 28.195 ;
    RECT 253.4 28.485 253.61 28.555 ;
    RECT 253.4 28.845 253.61 28.915 ;
    RECT 252.94 28.125 253.15 28.195 ;
    RECT 252.94 28.485 253.15 28.555 ;
    RECT 252.94 28.845 253.15 28.915 ;
    RECT 250.08 28.125 250.29 28.195 ;
    RECT 250.08 28.485 250.29 28.555 ;
    RECT 250.08 28.845 250.29 28.915 ;
    RECT 249.62 28.125 249.83 28.195 ;
    RECT 249.62 28.485 249.83 28.555 ;
    RECT 249.62 28.845 249.83 28.915 ;
    RECT 246.76 28.125 246.97 28.195 ;
    RECT 246.76 28.485 246.97 28.555 ;
    RECT 246.76 28.845 246.97 28.915 ;
    RECT 246.3 28.125 246.51 28.195 ;
    RECT 246.3 28.485 246.51 28.555 ;
    RECT 246.3 28.845 246.51 28.915 ;
    RECT 243.44 28.125 243.65 28.195 ;
    RECT 243.44 28.485 243.65 28.555 ;
    RECT 243.44 28.845 243.65 28.915 ;
    RECT 242.98 28.125 243.19 28.195 ;
    RECT 242.98 28.485 243.19 28.555 ;
    RECT 242.98 28.845 243.19 28.915 ;
    RECT 240.12 28.125 240.33 28.195 ;
    RECT 240.12 28.485 240.33 28.555 ;
    RECT 240.12 28.845 240.33 28.915 ;
    RECT 239.66 28.125 239.87 28.195 ;
    RECT 239.66 28.485 239.87 28.555 ;
    RECT 239.66 28.845 239.87 28.915 ;
    RECT 236.8 28.125 237.01 28.195 ;
    RECT 236.8 28.485 237.01 28.555 ;
    RECT 236.8 28.845 237.01 28.915 ;
    RECT 236.34 28.125 236.55 28.195 ;
    RECT 236.34 28.485 236.55 28.555 ;
    RECT 236.34 28.845 236.55 28.915 ;
    RECT 374.15 28.485 374.22 28.555 ;
    RECT 333.08 28.125 333.29 28.195 ;
    RECT 333.08 28.485 333.29 28.555 ;
    RECT 333.08 28.845 333.29 28.915 ;
    RECT 332.62 28.125 332.83 28.195 ;
    RECT 332.62 28.485 332.83 28.555 ;
    RECT 332.62 28.845 332.83 28.915 ;
    RECT 329.76 28.125 329.97 28.195 ;
    RECT 329.76 28.485 329.97 28.555 ;
    RECT 329.76 28.845 329.97 28.915 ;
    RECT 329.3 28.125 329.51 28.195 ;
    RECT 329.3 28.485 329.51 28.555 ;
    RECT 329.3 28.845 329.51 28.915 ;
    RECT 326.44 28.125 326.65 28.195 ;
    RECT 326.44 28.485 326.65 28.555 ;
    RECT 326.44 28.845 326.65 28.915 ;
    RECT 325.98 28.125 326.19 28.195 ;
    RECT 325.98 28.485 326.19 28.555 ;
    RECT 325.98 28.845 326.19 28.915 ;
    RECT 323.12 28.125 323.33 28.195 ;
    RECT 323.12 28.485 323.33 28.555 ;
    RECT 323.12 28.845 323.33 28.915 ;
    RECT 322.66 28.125 322.87 28.195 ;
    RECT 322.66 28.485 322.87 28.555 ;
    RECT 322.66 28.845 322.87 28.915 ;
    RECT 319.8 28.125 320.01 28.195 ;
    RECT 319.8 28.485 320.01 28.555 ;
    RECT 319.8 28.845 320.01 28.915 ;
    RECT 319.34 28.125 319.55 28.195 ;
    RECT 319.34 28.485 319.55 28.555 ;
    RECT 319.34 28.845 319.55 28.915 ;
    RECT 316.48 28.125 316.69 28.195 ;
    RECT 316.48 28.485 316.69 28.555 ;
    RECT 316.48 28.845 316.69 28.915 ;
    RECT 316.02 28.125 316.23 28.195 ;
    RECT 316.02 28.485 316.23 28.555 ;
    RECT 316.02 28.845 316.23 28.915 ;
    RECT 313.16 28.125 313.37 28.195 ;
    RECT 313.16 28.485 313.37 28.555 ;
    RECT 313.16 28.845 313.37 28.915 ;
    RECT 312.7 28.125 312.91 28.195 ;
    RECT 312.7 28.485 312.91 28.555 ;
    RECT 312.7 28.845 312.91 28.915 ;
    RECT 309.84 28.125 310.05 28.195 ;
    RECT 309.84 28.485 310.05 28.555 ;
    RECT 309.84 28.845 310.05 28.915 ;
    RECT 309.38 28.125 309.59 28.195 ;
    RECT 309.38 28.485 309.59 28.555 ;
    RECT 309.38 28.845 309.59 28.915 ;
    RECT 306.52 28.125 306.73 28.195 ;
    RECT 306.52 28.485 306.73 28.555 ;
    RECT 306.52 28.845 306.73 28.915 ;
    RECT 306.06 28.125 306.27 28.195 ;
    RECT 306.06 28.485 306.27 28.555 ;
    RECT 306.06 28.845 306.27 28.915 ;
    RECT 303.2 27.405 303.41 27.475 ;
    RECT 303.2 27.765 303.41 27.835 ;
    RECT 303.2 28.125 303.41 28.195 ;
    RECT 302.74 27.405 302.95 27.475 ;
    RECT 302.74 27.765 302.95 27.835 ;
    RECT 302.74 28.125 302.95 28.195 ;
    RECT 372.92 27.405 373.13 27.475 ;
    RECT 372.92 27.765 373.13 27.835 ;
    RECT 372.92 28.125 373.13 28.195 ;
    RECT 372.46 27.405 372.67 27.475 ;
    RECT 372.46 27.765 372.67 27.835 ;
    RECT 372.46 28.125 372.67 28.195 ;
    RECT 369.6 27.405 369.81 27.475 ;
    RECT 369.6 27.765 369.81 27.835 ;
    RECT 369.6 28.125 369.81 28.195 ;
    RECT 369.14 27.405 369.35 27.475 ;
    RECT 369.14 27.765 369.35 27.835 ;
    RECT 369.14 28.125 369.35 28.195 ;
    RECT 200.605 27.765 200.675 27.835 ;
    RECT 299.88 27.405 300.09 27.475 ;
    RECT 299.88 27.765 300.09 27.835 ;
    RECT 299.88 28.125 300.09 28.195 ;
    RECT 299.42 27.405 299.63 27.475 ;
    RECT 299.42 27.765 299.63 27.835 ;
    RECT 299.42 28.125 299.63 28.195 ;
    RECT 296.56 27.405 296.77 27.475 ;
    RECT 296.56 27.765 296.77 27.835 ;
    RECT 296.56 28.125 296.77 28.195 ;
    RECT 296.1 27.405 296.31 27.475 ;
    RECT 296.1 27.765 296.31 27.835 ;
    RECT 296.1 28.125 296.31 28.195 ;
    RECT 293.24 27.405 293.45 27.475 ;
    RECT 293.24 27.765 293.45 27.835 ;
    RECT 293.24 28.125 293.45 28.195 ;
    RECT 292.78 27.405 292.99 27.475 ;
    RECT 292.78 27.765 292.99 27.835 ;
    RECT 292.78 28.125 292.99 28.195 ;
    RECT 289.92 27.405 290.13 27.475 ;
    RECT 289.92 27.765 290.13 27.835 ;
    RECT 289.92 28.125 290.13 28.195 ;
    RECT 289.46 27.405 289.67 27.475 ;
    RECT 289.46 27.765 289.67 27.835 ;
    RECT 289.46 28.125 289.67 28.195 ;
    RECT 286.6 27.405 286.81 27.475 ;
    RECT 286.6 27.765 286.81 27.835 ;
    RECT 286.6 28.125 286.81 28.195 ;
    RECT 286.14 27.405 286.35 27.475 ;
    RECT 286.14 27.765 286.35 27.835 ;
    RECT 286.14 28.125 286.35 28.195 ;
    RECT 283.28 27.405 283.49 27.475 ;
    RECT 283.28 27.765 283.49 27.835 ;
    RECT 283.28 28.125 283.49 28.195 ;
    RECT 282.82 27.405 283.03 27.475 ;
    RECT 282.82 27.765 283.03 27.835 ;
    RECT 282.82 28.125 283.03 28.195 ;
    RECT 279.96 27.405 280.17 27.475 ;
    RECT 279.96 27.765 280.17 27.835 ;
    RECT 279.96 28.125 280.17 28.195 ;
    RECT 279.5 27.405 279.71 27.475 ;
    RECT 279.5 27.765 279.71 27.835 ;
    RECT 279.5 28.125 279.71 28.195 ;
    RECT 276.64 27.405 276.85 27.475 ;
    RECT 276.64 27.765 276.85 27.835 ;
    RECT 276.64 28.125 276.85 28.195 ;
    RECT 276.18 27.405 276.39 27.475 ;
    RECT 276.18 27.765 276.39 27.835 ;
    RECT 276.18 28.125 276.39 28.195 ;
    RECT 273.32 27.405 273.53 27.475 ;
    RECT 273.32 27.765 273.53 27.835 ;
    RECT 273.32 28.125 273.53 28.195 ;
    RECT 272.86 27.405 273.07 27.475 ;
    RECT 272.86 27.765 273.07 27.835 ;
    RECT 272.86 28.125 273.07 28.195 ;
    RECT 270.0 27.405 270.21 27.475 ;
    RECT 270.0 27.765 270.21 27.835 ;
    RECT 270.0 28.125 270.21 28.195 ;
    RECT 269.54 27.405 269.75 27.475 ;
    RECT 269.54 27.765 269.75 27.835 ;
    RECT 269.54 28.125 269.75 28.195 ;
    RECT 233.48 27.405 233.69 27.475 ;
    RECT 233.48 27.765 233.69 27.835 ;
    RECT 233.48 28.125 233.69 28.195 ;
    RECT 233.02 27.405 233.23 27.475 ;
    RECT 233.02 27.765 233.23 27.835 ;
    RECT 233.02 28.125 233.23 28.195 ;
    RECT 230.16 27.405 230.37 27.475 ;
    RECT 230.16 27.765 230.37 27.835 ;
    RECT 230.16 28.125 230.37 28.195 ;
    RECT 229.7 27.405 229.91 27.475 ;
    RECT 229.7 27.765 229.91 27.835 ;
    RECT 229.7 28.125 229.91 28.195 ;
    RECT 366.28 27.405 366.49 27.475 ;
    RECT 366.28 27.765 366.49 27.835 ;
    RECT 366.28 28.125 366.49 28.195 ;
    RECT 365.82 27.405 366.03 27.475 ;
    RECT 365.82 27.765 366.03 27.835 ;
    RECT 365.82 28.125 366.03 28.195 ;
    RECT 226.84 27.405 227.05 27.475 ;
    RECT 226.84 27.765 227.05 27.835 ;
    RECT 226.84 28.125 227.05 28.195 ;
    RECT 226.38 27.405 226.59 27.475 ;
    RECT 226.38 27.765 226.59 27.835 ;
    RECT 226.38 28.125 226.59 28.195 ;
    RECT 362.96 27.405 363.17 27.475 ;
    RECT 362.96 27.765 363.17 27.835 ;
    RECT 362.96 28.125 363.17 28.195 ;
    RECT 362.5 27.405 362.71 27.475 ;
    RECT 362.5 27.765 362.71 27.835 ;
    RECT 362.5 28.125 362.71 28.195 ;
    RECT 223.52 27.405 223.73 27.475 ;
    RECT 223.52 27.765 223.73 27.835 ;
    RECT 223.52 28.125 223.73 28.195 ;
    RECT 223.06 27.405 223.27 27.475 ;
    RECT 223.06 27.765 223.27 27.835 ;
    RECT 223.06 28.125 223.27 28.195 ;
    RECT 359.64 27.405 359.85 27.475 ;
    RECT 359.64 27.765 359.85 27.835 ;
    RECT 359.64 28.125 359.85 28.195 ;
    RECT 359.18 27.405 359.39 27.475 ;
    RECT 359.18 27.765 359.39 27.835 ;
    RECT 359.18 28.125 359.39 28.195 ;
    RECT 220.2 27.405 220.41 27.475 ;
    RECT 220.2 27.765 220.41 27.835 ;
    RECT 220.2 28.125 220.41 28.195 ;
    RECT 219.74 27.405 219.95 27.475 ;
    RECT 219.74 27.765 219.95 27.835 ;
    RECT 219.74 28.125 219.95 28.195 ;
    RECT 356.32 27.405 356.53 27.475 ;
    RECT 356.32 27.765 356.53 27.835 ;
    RECT 356.32 28.125 356.53 28.195 ;
    RECT 355.86 27.405 356.07 27.475 ;
    RECT 355.86 27.765 356.07 27.835 ;
    RECT 355.86 28.125 356.07 28.195 ;
    RECT 353.0 27.405 353.21 27.475 ;
    RECT 353.0 27.765 353.21 27.835 ;
    RECT 353.0 28.125 353.21 28.195 ;
    RECT 352.54 27.405 352.75 27.475 ;
    RECT 352.54 27.765 352.75 27.835 ;
    RECT 352.54 28.125 352.75 28.195 ;
    RECT 216.88 27.405 217.09 27.475 ;
    RECT 216.88 27.765 217.09 27.835 ;
    RECT 216.88 28.125 217.09 28.195 ;
    RECT 216.42 27.405 216.63 27.475 ;
    RECT 216.42 27.765 216.63 27.835 ;
    RECT 216.42 28.125 216.63 28.195 ;
    RECT 349.68 27.405 349.89 27.475 ;
    RECT 349.68 27.765 349.89 27.835 ;
    RECT 349.68 28.125 349.89 28.195 ;
    RECT 349.22 27.405 349.43 27.475 ;
    RECT 349.22 27.765 349.43 27.835 ;
    RECT 349.22 28.125 349.43 28.195 ;
    RECT 213.56 27.405 213.77 27.475 ;
    RECT 213.56 27.765 213.77 27.835 ;
    RECT 213.56 28.125 213.77 28.195 ;
    RECT 213.1 27.405 213.31 27.475 ;
    RECT 213.1 27.765 213.31 27.835 ;
    RECT 213.1 28.125 213.31 28.195 ;
    RECT 346.36 27.405 346.57 27.475 ;
    RECT 346.36 27.765 346.57 27.835 ;
    RECT 346.36 28.125 346.57 28.195 ;
    RECT 345.9 27.405 346.11 27.475 ;
    RECT 345.9 27.765 346.11 27.835 ;
    RECT 345.9 28.125 346.11 28.195 ;
    RECT 210.24 27.405 210.45 27.475 ;
    RECT 210.24 27.765 210.45 27.835 ;
    RECT 210.24 28.125 210.45 28.195 ;
    RECT 209.78 27.405 209.99 27.475 ;
    RECT 209.78 27.765 209.99 27.835 ;
    RECT 209.78 28.125 209.99 28.195 ;
    RECT 343.04 27.405 343.25 27.475 ;
    RECT 343.04 27.765 343.25 27.835 ;
    RECT 343.04 28.125 343.25 28.195 ;
    RECT 342.58 27.405 342.79 27.475 ;
    RECT 342.58 27.765 342.79 27.835 ;
    RECT 342.58 28.125 342.79 28.195 ;
    RECT 206.92 27.405 207.13 27.475 ;
    RECT 206.92 27.765 207.13 27.835 ;
    RECT 206.92 28.125 207.13 28.195 ;
    RECT 206.46 27.405 206.67 27.475 ;
    RECT 206.46 27.765 206.67 27.835 ;
    RECT 206.46 28.125 206.67 28.195 ;
    RECT 339.72 27.405 339.93 27.475 ;
    RECT 339.72 27.765 339.93 27.835 ;
    RECT 339.72 28.125 339.93 28.195 ;
    RECT 339.26 27.405 339.47 27.475 ;
    RECT 339.26 27.765 339.47 27.835 ;
    RECT 339.26 28.125 339.47 28.195 ;
    RECT 203.6 27.405 203.81 27.475 ;
    RECT 203.6 27.765 203.81 27.835 ;
    RECT 203.6 28.125 203.81 28.195 ;
    RECT 203.14 27.405 203.35 27.475 ;
    RECT 203.14 27.765 203.35 27.835 ;
    RECT 203.14 28.125 203.35 28.195 ;
    RECT 336.4 27.405 336.61 27.475 ;
    RECT 336.4 27.765 336.61 27.835 ;
    RECT 336.4 28.125 336.61 28.195 ;
    RECT 335.94 27.405 336.15 27.475 ;
    RECT 335.94 27.765 336.15 27.835 ;
    RECT 335.94 28.125 336.15 28.195 ;
    RECT 266.68 27.405 266.89 27.475 ;
    RECT 266.68 27.765 266.89 27.835 ;
    RECT 266.68 28.125 266.89 28.195 ;
    RECT 266.22 27.405 266.43 27.475 ;
    RECT 266.22 27.765 266.43 27.835 ;
    RECT 266.22 28.125 266.43 28.195 ;
    RECT 263.36 27.405 263.57 27.475 ;
    RECT 263.36 27.765 263.57 27.835 ;
    RECT 263.36 28.125 263.57 28.195 ;
    RECT 262.9 27.405 263.11 27.475 ;
    RECT 262.9 27.765 263.11 27.835 ;
    RECT 262.9 28.125 263.11 28.195 ;
    RECT 260.04 27.405 260.25 27.475 ;
    RECT 260.04 27.765 260.25 27.835 ;
    RECT 260.04 28.125 260.25 28.195 ;
    RECT 259.58 27.405 259.79 27.475 ;
    RECT 259.58 27.765 259.79 27.835 ;
    RECT 259.58 28.125 259.79 28.195 ;
    RECT 256.72 27.405 256.93 27.475 ;
    RECT 256.72 27.765 256.93 27.835 ;
    RECT 256.72 28.125 256.93 28.195 ;
    RECT 256.26 27.405 256.47 27.475 ;
    RECT 256.26 27.765 256.47 27.835 ;
    RECT 256.26 28.125 256.47 28.195 ;
    RECT 253.4 27.405 253.61 27.475 ;
    RECT 253.4 27.765 253.61 27.835 ;
    RECT 253.4 28.125 253.61 28.195 ;
    RECT 252.94 27.405 253.15 27.475 ;
    RECT 252.94 27.765 253.15 27.835 ;
    RECT 252.94 28.125 253.15 28.195 ;
    RECT 250.08 27.405 250.29 27.475 ;
    RECT 250.08 27.765 250.29 27.835 ;
    RECT 250.08 28.125 250.29 28.195 ;
    RECT 249.62 27.405 249.83 27.475 ;
    RECT 249.62 27.765 249.83 27.835 ;
    RECT 249.62 28.125 249.83 28.195 ;
    RECT 246.76 27.405 246.97 27.475 ;
    RECT 246.76 27.765 246.97 27.835 ;
    RECT 246.76 28.125 246.97 28.195 ;
    RECT 246.3 27.405 246.51 27.475 ;
    RECT 246.3 27.765 246.51 27.835 ;
    RECT 246.3 28.125 246.51 28.195 ;
    RECT 243.44 27.405 243.65 27.475 ;
    RECT 243.44 27.765 243.65 27.835 ;
    RECT 243.44 28.125 243.65 28.195 ;
    RECT 242.98 27.405 243.19 27.475 ;
    RECT 242.98 27.765 243.19 27.835 ;
    RECT 242.98 28.125 243.19 28.195 ;
    RECT 240.12 27.405 240.33 27.475 ;
    RECT 240.12 27.765 240.33 27.835 ;
    RECT 240.12 28.125 240.33 28.195 ;
    RECT 239.66 27.405 239.87 27.475 ;
    RECT 239.66 27.765 239.87 27.835 ;
    RECT 239.66 28.125 239.87 28.195 ;
    RECT 236.8 27.405 237.01 27.475 ;
    RECT 236.8 27.765 237.01 27.835 ;
    RECT 236.8 28.125 237.01 28.195 ;
    RECT 236.34 27.405 236.55 27.475 ;
    RECT 236.34 27.765 236.55 27.835 ;
    RECT 236.34 28.125 236.55 28.195 ;
    RECT 374.15 27.765 374.22 27.835 ;
    RECT 333.08 27.405 333.29 27.475 ;
    RECT 333.08 27.765 333.29 27.835 ;
    RECT 333.08 28.125 333.29 28.195 ;
    RECT 332.62 27.405 332.83 27.475 ;
    RECT 332.62 27.765 332.83 27.835 ;
    RECT 332.62 28.125 332.83 28.195 ;
    RECT 329.76 27.405 329.97 27.475 ;
    RECT 329.76 27.765 329.97 27.835 ;
    RECT 329.76 28.125 329.97 28.195 ;
    RECT 329.3 27.405 329.51 27.475 ;
    RECT 329.3 27.765 329.51 27.835 ;
    RECT 329.3 28.125 329.51 28.195 ;
    RECT 326.44 27.405 326.65 27.475 ;
    RECT 326.44 27.765 326.65 27.835 ;
    RECT 326.44 28.125 326.65 28.195 ;
    RECT 325.98 27.405 326.19 27.475 ;
    RECT 325.98 27.765 326.19 27.835 ;
    RECT 325.98 28.125 326.19 28.195 ;
    RECT 323.12 27.405 323.33 27.475 ;
    RECT 323.12 27.765 323.33 27.835 ;
    RECT 323.12 28.125 323.33 28.195 ;
    RECT 322.66 27.405 322.87 27.475 ;
    RECT 322.66 27.765 322.87 27.835 ;
    RECT 322.66 28.125 322.87 28.195 ;
    RECT 319.8 27.405 320.01 27.475 ;
    RECT 319.8 27.765 320.01 27.835 ;
    RECT 319.8 28.125 320.01 28.195 ;
    RECT 319.34 27.405 319.55 27.475 ;
    RECT 319.34 27.765 319.55 27.835 ;
    RECT 319.34 28.125 319.55 28.195 ;
    RECT 316.48 27.405 316.69 27.475 ;
    RECT 316.48 27.765 316.69 27.835 ;
    RECT 316.48 28.125 316.69 28.195 ;
    RECT 316.02 27.405 316.23 27.475 ;
    RECT 316.02 27.765 316.23 27.835 ;
    RECT 316.02 28.125 316.23 28.195 ;
    RECT 313.16 27.405 313.37 27.475 ;
    RECT 313.16 27.765 313.37 27.835 ;
    RECT 313.16 28.125 313.37 28.195 ;
    RECT 312.7 27.405 312.91 27.475 ;
    RECT 312.7 27.765 312.91 27.835 ;
    RECT 312.7 28.125 312.91 28.195 ;
    RECT 309.84 27.405 310.05 27.475 ;
    RECT 309.84 27.765 310.05 27.835 ;
    RECT 309.84 28.125 310.05 28.195 ;
    RECT 309.38 27.405 309.59 27.475 ;
    RECT 309.38 27.765 309.59 27.835 ;
    RECT 309.38 28.125 309.59 28.195 ;
    RECT 306.52 27.405 306.73 27.475 ;
    RECT 306.52 27.765 306.73 27.835 ;
    RECT 306.52 28.125 306.73 28.195 ;
    RECT 306.06 27.405 306.27 27.475 ;
    RECT 306.06 27.765 306.27 27.835 ;
    RECT 306.06 28.125 306.27 28.195 ;
    RECT 303.2 26.685 303.41 26.755 ;
    RECT 303.2 27.045 303.41 27.115 ;
    RECT 303.2 27.405 303.41 27.475 ;
    RECT 302.74 26.685 302.95 26.755 ;
    RECT 302.74 27.045 302.95 27.115 ;
    RECT 302.74 27.405 302.95 27.475 ;
    RECT 372.92 26.685 373.13 26.755 ;
    RECT 372.92 27.045 373.13 27.115 ;
    RECT 372.92 27.405 373.13 27.475 ;
    RECT 372.46 26.685 372.67 26.755 ;
    RECT 372.46 27.045 372.67 27.115 ;
    RECT 372.46 27.405 372.67 27.475 ;
    RECT 369.6 26.685 369.81 26.755 ;
    RECT 369.6 27.045 369.81 27.115 ;
    RECT 369.6 27.405 369.81 27.475 ;
    RECT 369.14 26.685 369.35 26.755 ;
    RECT 369.14 27.045 369.35 27.115 ;
    RECT 369.14 27.405 369.35 27.475 ;
    RECT 200.605 27.045 200.675 27.115 ;
    RECT 299.88 26.685 300.09 26.755 ;
    RECT 299.88 27.045 300.09 27.115 ;
    RECT 299.88 27.405 300.09 27.475 ;
    RECT 299.42 26.685 299.63 26.755 ;
    RECT 299.42 27.045 299.63 27.115 ;
    RECT 299.42 27.405 299.63 27.475 ;
    RECT 296.56 26.685 296.77 26.755 ;
    RECT 296.56 27.045 296.77 27.115 ;
    RECT 296.56 27.405 296.77 27.475 ;
    RECT 296.1 26.685 296.31 26.755 ;
    RECT 296.1 27.045 296.31 27.115 ;
    RECT 296.1 27.405 296.31 27.475 ;
    RECT 293.24 26.685 293.45 26.755 ;
    RECT 293.24 27.045 293.45 27.115 ;
    RECT 293.24 27.405 293.45 27.475 ;
    RECT 292.78 26.685 292.99 26.755 ;
    RECT 292.78 27.045 292.99 27.115 ;
    RECT 292.78 27.405 292.99 27.475 ;
    RECT 289.92 26.685 290.13 26.755 ;
    RECT 289.92 27.045 290.13 27.115 ;
    RECT 289.92 27.405 290.13 27.475 ;
    RECT 289.46 26.685 289.67 26.755 ;
    RECT 289.46 27.045 289.67 27.115 ;
    RECT 289.46 27.405 289.67 27.475 ;
    RECT 286.6 26.685 286.81 26.755 ;
    RECT 286.6 27.045 286.81 27.115 ;
    RECT 286.6 27.405 286.81 27.475 ;
    RECT 286.14 26.685 286.35 26.755 ;
    RECT 286.14 27.045 286.35 27.115 ;
    RECT 286.14 27.405 286.35 27.475 ;
    RECT 283.28 26.685 283.49 26.755 ;
    RECT 283.28 27.045 283.49 27.115 ;
    RECT 283.28 27.405 283.49 27.475 ;
    RECT 282.82 26.685 283.03 26.755 ;
    RECT 282.82 27.045 283.03 27.115 ;
    RECT 282.82 27.405 283.03 27.475 ;
    RECT 279.96 26.685 280.17 26.755 ;
    RECT 279.96 27.045 280.17 27.115 ;
    RECT 279.96 27.405 280.17 27.475 ;
    RECT 279.5 26.685 279.71 26.755 ;
    RECT 279.5 27.045 279.71 27.115 ;
    RECT 279.5 27.405 279.71 27.475 ;
    RECT 276.64 26.685 276.85 26.755 ;
    RECT 276.64 27.045 276.85 27.115 ;
    RECT 276.64 27.405 276.85 27.475 ;
    RECT 276.18 26.685 276.39 26.755 ;
    RECT 276.18 27.045 276.39 27.115 ;
    RECT 276.18 27.405 276.39 27.475 ;
    RECT 273.32 26.685 273.53 26.755 ;
    RECT 273.32 27.045 273.53 27.115 ;
    RECT 273.32 27.405 273.53 27.475 ;
    RECT 272.86 26.685 273.07 26.755 ;
    RECT 272.86 27.045 273.07 27.115 ;
    RECT 272.86 27.405 273.07 27.475 ;
    RECT 270.0 26.685 270.21 26.755 ;
    RECT 270.0 27.045 270.21 27.115 ;
    RECT 270.0 27.405 270.21 27.475 ;
    RECT 269.54 26.685 269.75 26.755 ;
    RECT 269.54 27.045 269.75 27.115 ;
    RECT 269.54 27.405 269.75 27.475 ;
    RECT 233.48 26.685 233.69 26.755 ;
    RECT 233.48 27.045 233.69 27.115 ;
    RECT 233.48 27.405 233.69 27.475 ;
    RECT 233.02 26.685 233.23 26.755 ;
    RECT 233.02 27.045 233.23 27.115 ;
    RECT 233.02 27.405 233.23 27.475 ;
    RECT 230.16 26.685 230.37 26.755 ;
    RECT 230.16 27.045 230.37 27.115 ;
    RECT 230.16 27.405 230.37 27.475 ;
    RECT 229.7 26.685 229.91 26.755 ;
    RECT 229.7 27.045 229.91 27.115 ;
    RECT 229.7 27.405 229.91 27.475 ;
    RECT 366.28 26.685 366.49 26.755 ;
    RECT 366.28 27.045 366.49 27.115 ;
    RECT 366.28 27.405 366.49 27.475 ;
    RECT 365.82 26.685 366.03 26.755 ;
    RECT 365.82 27.045 366.03 27.115 ;
    RECT 365.82 27.405 366.03 27.475 ;
    RECT 226.84 26.685 227.05 26.755 ;
    RECT 226.84 27.045 227.05 27.115 ;
    RECT 226.84 27.405 227.05 27.475 ;
    RECT 226.38 26.685 226.59 26.755 ;
    RECT 226.38 27.045 226.59 27.115 ;
    RECT 226.38 27.405 226.59 27.475 ;
    RECT 362.96 26.685 363.17 26.755 ;
    RECT 362.96 27.045 363.17 27.115 ;
    RECT 362.96 27.405 363.17 27.475 ;
    RECT 362.5 26.685 362.71 26.755 ;
    RECT 362.5 27.045 362.71 27.115 ;
    RECT 362.5 27.405 362.71 27.475 ;
    RECT 223.52 26.685 223.73 26.755 ;
    RECT 223.52 27.045 223.73 27.115 ;
    RECT 223.52 27.405 223.73 27.475 ;
    RECT 223.06 26.685 223.27 26.755 ;
    RECT 223.06 27.045 223.27 27.115 ;
    RECT 223.06 27.405 223.27 27.475 ;
    RECT 359.64 26.685 359.85 26.755 ;
    RECT 359.64 27.045 359.85 27.115 ;
    RECT 359.64 27.405 359.85 27.475 ;
    RECT 359.18 26.685 359.39 26.755 ;
    RECT 359.18 27.045 359.39 27.115 ;
    RECT 359.18 27.405 359.39 27.475 ;
    RECT 220.2 26.685 220.41 26.755 ;
    RECT 220.2 27.045 220.41 27.115 ;
    RECT 220.2 27.405 220.41 27.475 ;
    RECT 219.74 26.685 219.95 26.755 ;
    RECT 219.74 27.045 219.95 27.115 ;
    RECT 219.74 27.405 219.95 27.475 ;
    RECT 356.32 26.685 356.53 26.755 ;
    RECT 356.32 27.045 356.53 27.115 ;
    RECT 356.32 27.405 356.53 27.475 ;
    RECT 355.86 26.685 356.07 26.755 ;
    RECT 355.86 27.045 356.07 27.115 ;
    RECT 355.86 27.405 356.07 27.475 ;
    RECT 353.0 26.685 353.21 26.755 ;
    RECT 353.0 27.045 353.21 27.115 ;
    RECT 353.0 27.405 353.21 27.475 ;
    RECT 352.54 26.685 352.75 26.755 ;
    RECT 352.54 27.045 352.75 27.115 ;
    RECT 352.54 27.405 352.75 27.475 ;
    RECT 216.88 26.685 217.09 26.755 ;
    RECT 216.88 27.045 217.09 27.115 ;
    RECT 216.88 27.405 217.09 27.475 ;
    RECT 216.42 26.685 216.63 26.755 ;
    RECT 216.42 27.045 216.63 27.115 ;
    RECT 216.42 27.405 216.63 27.475 ;
    RECT 349.68 26.685 349.89 26.755 ;
    RECT 349.68 27.045 349.89 27.115 ;
    RECT 349.68 27.405 349.89 27.475 ;
    RECT 349.22 26.685 349.43 26.755 ;
    RECT 349.22 27.045 349.43 27.115 ;
    RECT 349.22 27.405 349.43 27.475 ;
    RECT 213.56 26.685 213.77 26.755 ;
    RECT 213.56 27.045 213.77 27.115 ;
    RECT 213.56 27.405 213.77 27.475 ;
    RECT 213.1 26.685 213.31 26.755 ;
    RECT 213.1 27.045 213.31 27.115 ;
    RECT 213.1 27.405 213.31 27.475 ;
    RECT 346.36 26.685 346.57 26.755 ;
    RECT 346.36 27.045 346.57 27.115 ;
    RECT 346.36 27.405 346.57 27.475 ;
    RECT 345.9 26.685 346.11 26.755 ;
    RECT 345.9 27.045 346.11 27.115 ;
    RECT 345.9 27.405 346.11 27.475 ;
    RECT 210.24 26.685 210.45 26.755 ;
    RECT 210.24 27.045 210.45 27.115 ;
    RECT 210.24 27.405 210.45 27.475 ;
    RECT 209.78 26.685 209.99 26.755 ;
    RECT 209.78 27.045 209.99 27.115 ;
    RECT 209.78 27.405 209.99 27.475 ;
    RECT 343.04 26.685 343.25 26.755 ;
    RECT 343.04 27.045 343.25 27.115 ;
    RECT 343.04 27.405 343.25 27.475 ;
    RECT 342.58 26.685 342.79 26.755 ;
    RECT 342.58 27.045 342.79 27.115 ;
    RECT 342.58 27.405 342.79 27.475 ;
    RECT 206.92 26.685 207.13 26.755 ;
    RECT 206.92 27.045 207.13 27.115 ;
    RECT 206.92 27.405 207.13 27.475 ;
    RECT 206.46 26.685 206.67 26.755 ;
    RECT 206.46 27.045 206.67 27.115 ;
    RECT 206.46 27.405 206.67 27.475 ;
    RECT 339.72 26.685 339.93 26.755 ;
    RECT 339.72 27.045 339.93 27.115 ;
    RECT 339.72 27.405 339.93 27.475 ;
    RECT 339.26 26.685 339.47 26.755 ;
    RECT 339.26 27.045 339.47 27.115 ;
    RECT 339.26 27.405 339.47 27.475 ;
    RECT 203.6 26.685 203.81 26.755 ;
    RECT 203.6 27.045 203.81 27.115 ;
    RECT 203.6 27.405 203.81 27.475 ;
    RECT 203.14 26.685 203.35 26.755 ;
    RECT 203.14 27.045 203.35 27.115 ;
    RECT 203.14 27.405 203.35 27.475 ;
    RECT 336.4 26.685 336.61 26.755 ;
    RECT 336.4 27.045 336.61 27.115 ;
    RECT 336.4 27.405 336.61 27.475 ;
    RECT 335.94 26.685 336.15 26.755 ;
    RECT 335.94 27.045 336.15 27.115 ;
    RECT 335.94 27.405 336.15 27.475 ;
    RECT 266.68 26.685 266.89 26.755 ;
    RECT 266.68 27.045 266.89 27.115 ;
    RECT 266.68 27.405 266.89 27.475 ;
    RECT 266.22 26.685 266.43 26.755 ;
    RECT 266.22 27.045 266.43 27.115 ;
    RECT 266.22 27.405 266.43 27.475 ;
    RECT 263.36 26.685 263.57 26.755 ;
    RECT 263.36 27.045 263.57 27.115 ;
    RECT 263.36 27.405 263.57 27.475 ;
    RECT 262.9 26.685 263.11 26.755 ;
    RECT 262.9 27.045 263.11 27.115 ;
    RECT 262.9 27.405 263.11 27.475 ;
    RECT 260.04 26.685 260.25 26.755 ;
    RECT 260.04 27.045 260.25 27.115 ;
    RECT 260.04 27.405 260.25 27.475 ;
    RECT 259.58 26.685 259.79 26.755 ;
    RECT 259.58 27.045 259.79 27.115 ;
    RECT 259.58 27.405 259.79 27.475 ;
    RECT 256.72 26.685 256.93 26.755 ;
    RECT 256.72 27.045 256.93 27.115 ;
    RECT 256.72 27.405 256.93 27.475 ;
    RECT 256.26 26.685 256.47 26.755 ;
    RECT 256.26 27.045 256.47 27.115 ;
    RECT 256.26 27.405 256.47 27.475 ;
    RECT 253.4 26.685 253.61 26.755 ;
    RECT 253.4 27.045 253.61 27.115 ;
    RECT 253.4 27.405 253.61 27.475 ;
    RECT 252.94 26.685 253.15 26.755 ;
    RECT 252.94 27.045 253.15 27.115 ;
    RECT 252.94 27.405 253.15 27.475 ;
    RECT 250.08 26.685 250.29 26.755 ;
    RECT 250.08 27.045 250.29 27.115 ;
    RECT 250.08 27.405 250.29 27.475 ;
    RECT 249.62 26.685 249.83 26.755 ;
    RECT 249.62 27.045 249.83 27.115 ;
    RECT 249.62 27.405 249.83 27.475 ;
    RECT 246.76 26.685 246.97 26.755 ;
    RECT 246.76 27.045 246.97 27.115 ;
    RECT 246.76 27.405 246.97 27.475 ;
    RECT 246.3 26.685 246.51 26.755 ;
    RECT 246.3 27.045 246.51 27.115 ;
    RECT 246.3 27.405 246.51 27.475 ;
    RECT 243.44 26.685 243.65 26.755 ;
    RECT 243.44 27.045 243.65 27.115 ;
    RECT 243.44 27.405 243.65 27.475 ;
    RECT 242.98 26.685 243.19 26.755 ;
    RECT 242.98 27.045 243.19 27.115 ;
    RECT 242.98 27.405 243.19 27.475 ;
    RECT 240.12 26.685 240.33 26.755 ;
    RECT 240.12 27.045 240.33 27.115 ;
    RECT 240.12 27.405 240.33 27.475 ;
    RECT 239.66 26.685 239.87 26.755 ;
    RECT 239.66 27.045 239.87 27.115 ;
    RECT 239.66 27.405 239.87 27.475 ;
    RECT 236.8 26.685 237.01 26.755 ;
    RECT 236.8 27.045 237.01 27.115 ;
    RECT 236.8 27.405 237.01 27.475 ;
    RECT 236.34 26.685 236.55 26.755 ;
    RECT 236.34 27.045 236.55 27.115 ;
    RECT 236.34 27.405 236.55 27.475 ;
    RECT 374.15 27.045 374.22 27.115 ;
    RECT 333.08 26.685 333.29 26.755 ;
    RECT 333.08 27.045 333.29 27.115 ;
    RECT 333.08 27.405 333.29 27.475 ;
    RECT 332.62 26.685 332.83 26.755 ;
    RECT 332.62 27.045 332.83 27.115 ;
    RECT 332.62 27.405 332.83 27.475 ;
    RECT 329.76 26.685 329.97 26.755 ;
    RECT 329.76 27.045 329.97 27.115 ;
    RECT 329.76 27.405 329.97 27.475 ;
    RECT 329.3 26.685 329.51 26.755 ;
    RECT 329.3 27.045 329.51 27.115 ;
    RECT 329.3 27.405 329.51 27.475 ;
    RECT 326.44 26.685 326.65 26.755 ;
    RECT 326.44 27.045 326.65 27.115 ;
    RECT 326.44 27.405 326.65 27.475 ;
    RECT 325.98 26.685 326.19 26.755 ;
    RECT 325.98 27.045 326.19 27.115 ;
    RECT 325.98 27.405 326.19 27.475 ;
    RECT 323.12 26.685 323.33 26.755 ;
    RECT 323.12 27.045 323.33 27.115 ;
    RECT 323.12 27.405 323.33 27.475 ;
    RECT 322.66 26.685 322.87 26.755 ;
    RECT 322.66 27.045 322.87 27.115 ;
    RECT 322.66 27.405 322.87 27.475 ;
    RECT 319.8 26.685 320.01 26.755 ;
    RECT 319.8 27.045 320.01 27.115 ;
    RECT 319.8 27.405 320.01 27.475 ;
    RECT 319.34 26.685 319.55 26.755 ;
    RECT 319.34 27.045 319.55 27.115 ;
    RECT 319.34 27.405 319.55 27.475 ;
    RECT 316.48 26.685 316.69 26.755 ;
    RECT 316.48 27.045 316.69 27.115 ;
    RECT 316.48 27.405 316.69 27.475 ;
    RECT 316.02 26.685 316.23 26.755 ;
    RECT 316.02 27.045 316.23 27.115 ;
    RECT 316.02 27.405 316.23 27.475 ;
    RECT 313.16 26.685 313.37 26.755 ;
    RECT 313.16 27.045 313.37 27.115 ;
    RECT 313.16 27.405 313.37 27.475 ;
    RECT 312.7 26.685 312.91 26.755 ;
    RECT 312.7 27.045 312.91 27.115 ;
    RECT 312.7 27.405 312.91 27.475 ;
    RECT 309.84 26.685 310.05 26.755 ;
    RECT 309.84 27.045 310.05 27.115 ;
    RECT 309.84 27.405 310.05 27.475 ;
    RECT 309.38 26.685 309.59 26.755 ;
    RECT 309.38 27.045 309.59 27.115 ;
    RECT 309.38 27.405 309.59 27.475 ;
    RECT 306.52 26.685 306.73 26.755 ;
    RECT 306.52 27.045 306.73 27.115 ;
    RECT 306.52 27.405 306.73 27.475 ;
    RECT 306.06 26.685 306.27 26.755 ;
    RECT 306.06 27.045 306.27 27.115 ;
    RECT 306.06 27.405 306.27 27.475 ;
    RECT 303.2 25.965 303.41 26.035 ;
    RECT 303.2 26.325 303.41 26.395 ;
    RECT 303.2 26.685 303.41 26.755 ;
    RECT 302.74 25.965 302.95 26.035 ;
    RECT 302.74 26.325 302.95 26.395 ;
    RECT 302.74 26.685 302.95 26.755 ;
    RECT 372.92 25.965 373.13 26.035 ;
    RECT 372.92 26.325 373.13 26.395 ;
    RECT 372.92 26.685 373.13 26.755 ;
    RECT 372.46 25.965 372.67 26.035 ;
    RECT 372.46 26.325 372.67 26.395 ;
    RECT 372.46 26.685 372.67 26.755 ;
    RECT 369.6 25.965 369.81 26.035 ;
    RECT 369.6 26.325 369.81 26.395 ;
    RECT 369.6 26.685 369.81 26.755 ;
    RECT 369.14 25.965 369.35 26.035 ;
    RECT 369.14 26.325 369.35 26.395 ;
    RECT 369.14 26.685 369.35 26.755 ;
    RECT 200.605 26.325 200.675 26.395 ;
    RECT 299.88 25.965 300.09 26.035 ;
    RECT 299.88 26.325 300.09 26.395 ;
    RECT 299.88 26.685 300.09 26.755 ;
    RECT 299.42 25.965 299.63 26.035 ;
    RECT 299.42 26.325 299.63 26.395 ;
    RECT 299.42 26.685 299.63 26.755 ;
    RECT 296.56 25.965 296.77 26.035 ;
    RECT 296.56 26.325 296.77 26.395 ;
    RECT 296.56 26.685 296.77 26.755 ;
    RECT 296.1 25.965 296.31 26.035 ;
    RECT 296.1 26.325 296.31 26.395 ;
    RECT 296.1 26.685 296.31 26.755 ;
    RECT 293.24 25.965 293.45 26.035 ;
    RECT 293.24 26.325 293.45 26.395 ;
    RECT 293.24 26.685 293.45 26.755 ;
    RECT 292.78 25.965 292.99 26.035 ;
    RECT 292.78 26.325 292.99 26.395 ;
    RECT 292.78 26.685 292.99 26.755 ;
    RECT 289.92 25.965 290.13 26.035 ;
    RECT 289.92 26.325 290.13 26.395 ;
    RECT 289.92 26.685 290.13 26.755 ;
    RECT 289.46 25.965 289.67 26.035 ;
    RECT 289.46 26.325 289.67 26.395 ;
    RECT 289.46 26.685 289.67 26.755 ;
    RECT 286.6 25.965 286.81 26.035 ;
    RECT 286.6 26.325 286.81 26.395 ;
    RECT 286.6 26.685 286.81 26.755 ;
    RECT 286.14 25.965 286.35 26.035 ;
    RECT 286.14 26.325 286.35 26.395 ;
    RECT 286.14 26.685 286.35 26.755 ;
    RECT 283.28 25.965 283.49 26.035 ;
    RECT 283.28 26.325 283.49 26.395 ;
    RECT 283.28 26.685 283.49 26.755 ;
    RECT 282.82 25.965 283.03 26.035 ;
    RECT 282.82 26.325 283.03 26.395 ;
    RECT 282.82 26.685 283.03 26.755 ;
    RECT 279.96 25.965 280.17 26.035 ;
    RECT 279.96 26.325 280.17 26.395 ;
    RECT 279.96 26.685 280.17 26.755 ;
    RECT 279.5 25.965 279.71 26.035 ;
    RECT 279.5 26.325 279.71 26.395 ;
    RECT 279.5 26.685 279.71 26.755 ;
    RECT 276.64 25.965 276.85 26.035 ;
    RECT 276.64 26.325 276.85 26.395 ;
    RECT 276.64 26.685 276.85 26.755 ;
    RECT 276.18 25.965 276.39 26.035 ;
    RECT 276.18 26.325 276.39 26.395 ;
    RECT 276.18 26.685 276.39 26.755 ;
    RECT 273.32 25.965 273.53 26.035 ;
    RECT 273.32 26.325 273.53 26.395 ;
    RECT 273.32 26.685 273.53 26.755 ;
    RECT 272.86 25.965 273.07 26.035 ;
    RECT 272.86 26.325 273.07 26.395 ;
    RECT 272.86 26.685 273.07 26.755 ;
    RECT 270.0 25.965 270.21 26.035 ;
    RECT 270.0 26.325 270.21 26.395 ;
    RECT 270.0 26.685 270.21 26.755 ;
    RECT 269.54 25.965 269.75 26.035 ;
    RECT 269.54 26.325 269.75 26.395 ;
    RECT 269.54 26.685 269.75 26.755 ;
    RECT 233.48 25.965 233.69 26.035 ;
    RECT 233.48 26.325 233.69 26.395 ;
    RECT 233.48 26.685 233.69 26.755 ;
    RECT 233.02 25.965 233.23 26.035 ;
    RECT 233.02 26.325 233.23 26.395 ;
    RECT 233.02 26.685 233.23 26.755 ;
    RECT 230.16 25.965 230.37 26.035 ;
    RECT 230.16 26.325 230.37 26.395 ;
    RECT 230.16 26.685 230.37 26.755 ;
    RECT 229.7 25.965 229.91 26.035 ;
    RECT 229.7 26.325 229.91 26.395 ;
    RECT 229.7 26.685 229.91 26.755 ;
    RECT 366.28 25.965 366.49 26.035 ;
    RECT 366.28 26.325 366.49 26.395 ;
    RECT 366.28 26.685 366.49 26.755 ;
    RECT 365.82 25.965 366.03 26.035 ;
    RECT 365.82 26.325 366.03 26.395 ;
    RECT 365.82 26.685 366.03 26.755 ;
    RECT 226.84 25.965 227.05 26.035 ;
    RECT 226.84 26.325 227.05 26.395 ;
    RECT 226.84 26.685 227.05 26.755 ;
    RECT 226.38 25.965 226.59 26.035 ;
    RECT 226.38 26.325 226.59 26.395 ;
    RECT 226.38 26.685 226.59 26.755 ;
    RECT 362.96 25.965 363.17 26.035 ;
    RECT 362.96 26.325 363.17 26.395 ;
    RECT 362.96 26.685 363.17 26.755 ;
    RECT 362.5 25.965 362.71 26.035 ;
    RECT 362.5 26.325 362.71 26.395 ;
    RECT 362.5 26.685 362.71 26.755 ;
    RECT 223.52 25.965 223.73 26.035 ;
    RECT 223.52 26.325 223.73 26.395 ;
    RECT 223.52 26.685 223.73 26.755 ;
    RECT 223.06 25.965 223.27 26.035 ;
    RECT 223.06 26.325 223.27 26.395 ;
    RECT 223.06 26.685 223.27 26.755 ;
    RECT 359.64 25.965 359.85 26.035 ;
    RECT 359.64 26.325 359.85 26.395 ;
    RECT 359.64 26.685 359.85 26.755 ;
    RECT 359.18 25.965 359.39 26.035 ;
    RECT 359.18 26.325 359.39 26.395 ;
    RECT 359.18 26.685 359.39 26.755 ;
    RECT 220.2 25.965 220.41 26.035 ;
    RECT 220.2 26.325 220.41 26.395 ;
    RECT 220.2 26.685 220.41 26.755 ;
    RECT 219.74 25.965 219.95 26.035 ;
    RECT 219.74 26.325 219.95 26.395 ;
    RECT 219.74 26.685 219.95 26.755 ;
    RECT 356.32 25.965 356.53 26.035 ;
    RECT 356.32 26.325 356.53 26.395 ;
    RECT 356.32 26.685 356.53 26.755 ;
    RECT 355.86 25.965 356.07 26.035 ;
    RECT 355.86 26.325 356.07 26.395 ;
    RECT 355.86 26.685 356.07 26.755 ;
    RECT 353.0 25.965 353.21 26.035 ;
    RECT 353.0 26.325 353.21 26.395 ;
    RECT 353.0 26.685 353.21 26.755 ;
    RECT 352.54 25.965 352.75 26.035 ;
    RECT 352.54 26.325 352.75 26.395 ;
    RECT 352.54 26.685 352.75 26.755 ;
    RECT 216.88 25.965 217.09 26.035 ;
    RECT 216.88 26.325 217.09 26.395 ;
    RECT 216.88 26.685 217.09 26.755 ;
    RECT 216.42 25.965 216.63 26.035 ;
    RECT 216.42 26.325 216.63 26.395 ;
    RECT 216.42 26.685 216.63 26.755 ;
    RECT 349.68 25.965 349.89 26.035 ;
    RECT 349.68 26.325 349.89 26.395 ;
    RECT 349.68 26.685 349.89 26.755 ;
    RECT 349.22 25.965 349.43 26.035 ;
    RECT 349.22 26.325 349.43 26.395 ;
    RECT 349.22 26.685 349.43 26.755 ;
    RECT 213.56 25.965 213.77 26.035 ;
    RECT 213.56 26.325 213.77 26.395 ;
    RECT 213.56 26.685 213.77 26.755 ;
    RECT 213.1 25.965 213.31 26.035 ;
    RECT 213.1 26.325 213.31 26.395 ;
    RECT 213.1 26.685 213.31 26.755 ;
    RECT 346.36 25.965 346.57 26.035 ;
    RECT 346.36 26.325 346.57 26.395 ;
    RECT 346.36 26.685 346.57 26.755 ;
    RECT 345.9 25.965 346.11 26.035 ;
    RECT 345.9 26.325 346.11 26.395 ;
    RECT 345.9 26.685 346.11 26.755 ;
    RECT 210.24 25.965 210.45 26.035 ;
    RECT 210.24 26.325 210.45 26.395 ;
    RECT 210.24 26.685 210.45 26.755 ;
    RECT 209.78 25.965 209.99 26.035 ;
    RECT 209.78 26.325 209.99 26.395 ;
    RECT 209.78 26.685 209.99 26.755 ;
    RECT 343.04 25.965 343.25 26.035 ;
    RECT 343.04 26.325 343.25 26.395 ;
    RECT 343.04 26.685 343.25 26.755 ;
    RECT 342.58 25.965 342.79 26.035 ;
    RECT 342.58 26.325 342.79 26.395 ;
    RECT 342.58 26.685 342.79 26.755 ;
    RECT 206.92 25.965 207.13 26.035 ;
    RECT 206.92 26.325 207.13 26.395 ;
    RECT 206.92 26.685 207.13 26.755 ;
    RECT 206.46 25.965 206.67 26.035 ;
    RECT 206.46 26.325 206.67 26.395 ;
    RECT 206.46 26.685 206.67 26.755 ;
    RECT 339.72 25.965 339.93 26.035 ;
    RECT 339.72 26.325 339.93 26.395 ;
    RECT 339.72 26.685 339.93 26.755 ;
    RECT 339.26 25.965 339.47 26.035 ;
    RECT 339.26 26.325 339.47 26.395 ;
    RECT 339.26 26.685 339.47 26.755 ;
    RECT 203.6 25.965 203.81 26.035 ;
    RECT 203.6 26.325 203.81 26.395 ;
    RECT 203.6 26.685 203.81 26.755 ;
    RECT 203.14 25.965 203.35 26.035 ;
    RECT 203.14 26.325 203.35 26.395 ;
    RECT 203.14 26.685 203.35 26.755 ;
    RECT 336.4 25.965 336.61 26.035 ;
    RECT 336.4 26.325 336.61 26.395 ;
    RECT 336.4 26.685 336.61 26.755 ;
    RECT 335.94 25.965 336.15 26.035 ;
    RECT 335.94 26.325 336.15 26.395 ;
    RECT 335.94 26.685 336.15 26.755 ;
    RECT 266.68 25.965 266.89 26.035 ;
    RECT 266.68 26.325 266.89 26.395 ;
    RECT 266.68 26.685 266.89 26.755 ;
    RECT 266.22 25.965 266.43 26.035 ;
    RECT 266.22 26.325 266.43 26.395 ;
    RECT 266.22 26.685 266.43 26.755 ;
    RECT 263.36 25.965 263.57 26.035 ;
    RECT 263.36 26.325 263.57 26.395 ;
    RECT 263.36 26.685 263.57 26.755 ;
    RECT 262.9 25.965 263.11 26.035 ;
    RECT 262.9 26.325 263.11 26.395 ;
    RECT 262.9 26.685 263.11 26.755 ;
    RECT 260.04 25.965 260.25 26.035 ;
    RECT 260.04 26.325 260.25 26.395 ;
    RECT 260.04 26.685 260.25 26.755 ;
    RECT 259.58 25.965 259.79 26.035 ;
    RECT 259.58 26.325 259.79 26.395 ;
    RECT 259.58 26.685 259.79 26.755 ;
    RECT 256.72 25.965 256.93 26.035 ;
    RECT 256.72 26.325 256.93 26.395 ;
    RECT 256.72 26.685 256.93 26.755 ;
    RECT 256.26 25.965 256.47 26.035 ;
    RECT 256.26 26.325 256.47 26.395 ;
    RECT 256.26 26.685 256.47 26.755 ;
    RECT 253.4 25.965 253.61 26.035 ;
    RECT 253.4 26.325 253.61 26.395 ;
    RECT 253.4 26.685 253.61 26.755 ;
    RECT 252.94 25.965 253.15 26.035 ;
    RECT 252.94 26.325 253.15 26.395 ;
    RECT 252.94 26.685 253.15 26.755 ;
    RECT 250.08 25.965 250.29 26.035 ;
    RECT 250.08 26.325 250.29 26.395 ;
    RECT 250.08 26.685 250.29 26.755 ;
    RECT 249.62 25.965 249.83 26.035 ;
    RECT 249.62 26.325 249.83 26.395 ;
    RECT 249.62 26.685 249.83 26.755 ;
    RECT 246.76 25.965 246.97 26.035 ;
    RECT 246.76 26.325 246.97 26.395 ;
    RECT 246.76 26.685 246.97 26.755 ;
    RECT 246.3 25.965 246.51 26.035 ;
    RECT 246.3 26.325 246.51 26.395 ;
    RECT 246.3 26.685 246.51 26.755 ;
    RECT 243.44 25.965 243.65 26.035 ;
    RECT 243.44 26.325 243.65 26.395 ;
    RECT 243.44 26.685 243.65 26.755 ;
    RECT 242.98 25.965 243.19 26.035 ;
    RECT 242.98 26.325 243.19 26.395 ;
    RECT 242.98 26.685 243.19 26.755 ;
    RECT 240.12 25.965 240.33 26.035 ;
    RECT 240.12 26.325 240.33 26.395 ;
    RECT 240.12 26.685 240.33 26.755 ;
    RECT 239.66 25.965 239.87 26.035 ;
    RECT 239.66 26.325 239.87 26.395 ;
    RECT 239.66 26.685 239.87 26.755 ;
    RECT 236.8 25.965 237.01 26.035 ;
    RECT 236.8 26.325 237.01 26.395 ;
    RECT 236.8 26.685 237.01 26.755 ;
    RECT 236.34 25.965 236.55 26.035 ;
    RECT 236.34 26.325 236.55 26.395 ;
    RECT 236.34 26.685 236.55 26.755 ;
    RECT 374.15 26.325 374.22 26.395 ;
    RECT 333.08 25.965 333.29 26.035 ;
    RECT 333.08 26.325 333.29 26.395 ;
    RECT 333.08 26.685 333.29 26.755 ;
    RECT 332.62 25.965 332.83 26.035 ;
    RECT 332.62 26.325 332.83 26.395 ;
    RECT 332.62 26.685 332.83 26.755 ;
    RECT 329.76 25.965 329.97 26.035 ;
    RECT 329.76 26.325 329.97 26.395 ;
    RECT 329.76 26.685 329.97 26.755 ;
    RECT 329.3 25.965 329.51 26.035 ;
    RECT 329.3 26.325 329.51 26.395 ;
    RECT 329.3 26.685 329.51 26.755 ;
    RECT 326.44 25.965 326.65 26.035 ;
    RECT 326.44 26.325 326.65 26.395 ;
    RECT 326.44 26.685 326.65 26.755 ;
    RECT 325.98 25.965 326.19 26.035 ;
    RECT 325.98 26.325 326.19 26.395 ;
    RECT 325.98 26.685 326.19 26.755 ;
    RECT 323.12 25.965 323.33 26.035 ;
    RECT 323.12 26.325 323.33 26.395 ;
    RECT 323.12 26.685 323.33 26.755 ;
    RECT 322.66 25.965 322.87 26.035 ;
    RECT 322.66 26.325 322.87 26.395 ;
    RECT 322.66 26.685 322.87 26.755 ;
    RECT 319.8 25.965 320.01 26.035 ;
    RECT 319.8 26.325 320.01 26.395 ;
    RECT 319.8 26.685 320.01 26.755 ;
    RECT 319.34 25.965 319.55 26.035 ;
    RECT 319.34 26.325 319.55 26.395 ;
    RECT 319.34 26.685 319.55 26.755 ;
    RECT 316.48 25.965 316.69 26.035 ;
    RECT 316.48 26.325 316.69 26.395 ;
    RECT 316.48 26.685 316.69 26.755 ;
    RECT 316.02 25.965 316.23 26.035 ;
    RECT 316.02 26.325 316.23 26.395 ;
    RECT 316.02 26.685 316.23 26.755 ;
    RECT 313.16 25.965 313.37 26.035 ;
    RECT 313.16 26.325 313.37 26.395 ;
    RECT 313.16 26.685 313.37 26.755 ;
    RECT 312.7 25.965 312.91 26.035 ;
    RECT 312.7 26.325 312.91 26.395 ;
    RECT 312.7 26.685 312.91 26.755 ;
    RECT 309.84 25.965 310.05 26.035 ;
    RECT 309.84 26.325 310.05 26.395 ;
    RECT 309.84 26.685 310.05 26.755 ;
    RECT 309.38 25.965 309.59 26.035 ;
    RECT 309.38 26.325 309.59 26.395 ;
    RECT 309.38 26.685 309.59 26.755 ;
    RECT 306.52 25.965 306.73 26.035 ;
    RECT 306.52 26.325 306.73 26.395 ;
    RECT 306.52 26.685 306.73 26.755 ;
    RECT 306.06 25.965 306.27 26.035 ;
    RECT 306.06 26.325 306.27 26.395 ;
    RECT 306.06 26.685 306.27 26.755 ;
    RECT 303.2 35.325 303.41 35.395 ;
    RECT 303.2 35.685 303.41 35.755 ;
    RECT 303.2 36.045 303.41 36.115 ;
    RECT 302.74 35.325 302.95 35.395 ;
    RECT 302.74 35.685 302.95 35.755 ;
    RECT 302.74 36.045 302.95 36.115 ;
    RECT 372.92 35.325 373.13 35.395 ;
    RECT 372.92 35.685 373.13 35.755 ;
    RECT 372.92 36.045 373.13 36.115 ;
    RECT 372.46 35.325 372.67 35.395 ;
    RECT 372.46 35.685 372.67 35.755 ;
    RECT 372.46 36.045 372.67 36.115 ;
    RECT 369.6 35.325 369.81 35.395 ;
    RECT 369.6 35.685 369.81 35.755 ;
    RECT 369.6 36.045 369.81 36.115 ;
    RECT 369.14 35.325 369.35 35.395 ;
    RECT 369.14 35.685 369.35 35.755 ;
    RECT 369.14 36.045 369.35 36.115 ;
    RECT 299.88 35.325 300.09 35.395 ;
    RECT 299.88 35.685 300.09 35.755 ;
    RECT 299.88 36.045 300.09 36.115 ;
    RECT 299.42 35.325 299.63 35.395 ;
    RECT 299.42 35.685 299.63 35.755 ;
    RECT 299.42 36.045 299.63 36.115 ;
    RECT 296.56 35.325 296.77 35.395 ;
    RECT 296.56 35.685 296.77 35.755 ;
    RECT 296.56 36.045 296.77 36.115 ;
    RECT 296.1 35.325 296.31 35.395 ;
    RECT 296.1 35.685 296.31 35.755 ;
    RECT 296.1 36.045 296.31 36.115 ;
    RECT 293.24 35.325 293.45 35.395 ;
    RECT 293.24 35.685 293.45 35.755 ;
    RECT 293.24 36.045 293.45 36.115 ;
    RECT 292.78 35.325 292.99 35.395 ;
    RECT 292.78 35.685 292.99 35.755 ;
    RECT 292.78 36.045 292.99 36.115 ;
    RECT 289.92 35.325 290.13 35.395 ;
    RECT 289.92 35.685 290.13 35.755 ;
    RECT 289.92 36.045 290.13 36.115 ;
    RECT 289.46 35.325 289.67 35.395 ;
    RECT 289.46 35.685 289.67 35.755 ;
    RECT 289.46 36.045 289.67 36.115 ;
    RECT 286.6 35.325 286.81 35.395 ;
    RECT 286.6 35.685 286.81 35.755 ;
    RECT 286.6 36.045 286.81 36.115 ;
    RECT 286.14 35.325 286.35 35.395 ;
    RECT 286.14 35.685 286.35 35.755 ;
    RECT 286.14 36.045 286.35 36.115 ;
    RECT 283.28 35.325 283.49 35.395 ;
    RECT 283.28 35.685 283.49 35.755 ;
    RECT 283.28 36.045 283.49 36.115 ;
    RECT 282.82 35.325 283.03 35.395 ;
    RECT 282.82 35.685 283.03 35.755 ;
    RECT 282.82 36.045 283.03 36.115 ;
    RECT 279.96 35.325 280.17 35.395 ;
    RECT 279.96 35.685 280.17 35.755 ;
    RECT 279.96 36.045 280.17 36.115 ;
    RECT 279.5 35.325 279.71 35.395 ;
    RECT 279.5 35.685 279.71 35.755 ;
    RECT 279.5 36.045 279.71 36.115 ;
    RECT 276.64 35.325 276.85 35.395 ;
    RECT 276.64 35.685 276.85 35.755 ;
    RECT 276.64 36.045 276.85 36.115 ;
    RECT 276.18 35.325 276.39 35.395 ;
    RECT 276.18 35.685 276.39 35.755 ;
    RECT 276.18 36.045 276.39 36.115 ;
    RECT 273.32 35.325 273.53 35.395 ;
    RECT 273.32 35.685 273.53 35.755 ;
    RECT 273.32 36.045 273.53 36.115 ;
    RECT 272.86 35.325 273.07 35.395 ;
    RECT 272.86 35.685 273.07 35.755 ;
    RECT 272.86 36.045 273.07 36.115 ;
    RECT 270.0 35.325 270.21 35.395 ;
    RECT 270.0 35.685 270.21 35.755 ;
    RECT 270.0 36.045 270.21 36.115 ;
    RECT 269.54 35.325 269.75 35.395 ;
    RECT 269.54 35.685 269.75 35.755 ;
    RECT 269.54 36.045 269.75 36.115 ;
    RECT 233.48 35.325 233.69 35.395 ;
    RECT 233.48 35.685 233.69 35.755 ;
    RECT 233.48 36.045 233.69 36.115 ;
    RECT 233.02 35.325 233.23 35.395 ;
    RECT 233.02 35.685 233.23 35.755 ;
    RECT 233.02 36.045 233.23 36.115 ;
    RECT 230.16 35.325 230.37 35.395 ;
    RECT 230.16 35.685 230.37 35.755 ;
    RECT 230.16 36.045 230.37 36.115 ;
    RECT 229.7 35.325 229.91 35.395 ;
    RECT 229.7 35.685 229.91 35.755 ;
    RECT 229.7 36.045 229.91 36.115 ;
    RECT 366.28 35.325 366.49 35.395 ;
    RECT 366.28 35.685 366.49 35.755 ;
    RECT 366.28 36.045 366.49 36.115 ;
    RECT 365.82 35.325 366.03 35.395 ;
    RECT 365.82 35.685 366.03 35.755 ;
    RECT 365.82 36.045 366.03 36.115 ;
    RECT 374.15 35.685 374.22 35.755 ;
    RECT 226.84 35.325 227.05 35.395 ;
    RECT 226.84 35.685 227.05 35.755 ;
    RECT 226.84 36.045 227.05 36.115 ;
    RECT 226.38 35.325 226.59 35.395 ;
    RECT 226.38 35.685 226.59 35.755 ;
    RECT 226.38 36.045 226.59 36.115 ;
    RECT 362.96 35.325 363.17 35.395 ;
    RECT 362.96 35.685 363.17 35.755 ;
    RECT 362.96 36.045 363.17 36.115 ;
    RECT 362.5 35.325 362.71 35.395 ;
    RECT 362.5 35.685 362.71 35.755 ;
    RECT 362.5 36.045 362.71 36.115 ;
    RECT 223.52 35.325 223.73 35.395 ;
    RECT 223.52 35.685 223.73 35.755 ;
    RECT 223.52 36.045 223.73 36.115 ;
    RECT 223.06 35.325 223.27 35.395 ;
    RECT 223.06 35.685 223.27 35.755 ;
    RECT 223.06 36.045 223.27 36.115 ;
    RECT 359.64 35.325 359.85 35.395 ;
    RECT 359.64 35.685 359.85 35.755 ;
    RECT 359.64 36.045 359.85 36.115 ;
    RECT 359.18 35.325 359.39 35.395 ;
    RECT 359.18 35.685 359.39 35.755 ;
    RECT 359.18 36.045 359.39 36.115 ;
    RECT 220.2 35.325 220.41 35.395 ;
    RECT 220.2 35.685 220.41 35.755 ;
    RECT 220.2 36.045 220.41 36.115 ;
    RECT 219.74 35.325 219.95 35.395 ;
    RECT 219.74 35.685 219.95 35.755 ;
    RECT 219.74 36.045 219.95 36.115 ;
    RECT 356.32 35.325 356.53 35.395 ;
    RECT 356.32 35.685 356.53 35.755 ;
    RECT 356.32 36.045 356.53 36.115 ;
    RECT 355.86 35.325 356.07 35.395 ;
    RECT 355.86 35.685 356.07 35.755 ;
    RECT 355.86 36.045 356.07 36.115 ;
    RECT 353.0 35.325 353.21 35.395 ;
    RECT 353.0 35.685 353.21 35.755 ;
    RECT 353.0 36.045 353.21 36.115 ;
    RECT 352.54 35.325 352.75 35.395 ;
    RECT 352.54 35.685 352.75 35.755 ;
    RECT 352.54 36.045 352.75 36.115 ;
    RECT 216.88 35.325 217.09 35.395 ;
    RECT 216.88 35.685 217.09 35.755 ;
    RECT 216.88 36.045 217.09 36.115 ;
    RECT 216.42 35.325 216.63 35.395 ;
    RECT 216.42 35.685 216.63 35.755 ;
    RECT 216.42 36.045 216.63 36.115 ;
    RECT 349.68 35.325 349.89 35.395 ;
    RECT 349.68 35.685 349.89 35.755 ;
    RECT 349.68 36.045 349.89 36.115 ;
    RECT 349.22 35.325 349.43 35.395 ;
    RECT 349.22 35.685 349.43 35.755 ;
    RECT 349.22 36.045 349.43 36.115 ;
    RECT 213.56 35.325 213.77 35.395 ;
    RECT 213.56 35.685 213.77 35.755 ;
    RECT 213.56 36.045 213.77 36.115 ;
    RECT 213.1 35.325 213.31 35.395 ;
    RECT 213.1 35.685 213.31 35.755 ;
    RECT 213.1 36.045 213.31 36.115 ;
    RECT 346.36 35.325 346.57 35.395 ;
    RECT 346.36 35.685 346.57 35.755 ;
    RECT 346.36 36.045 346.57 36.115 ;
    RECT 345.9 35.325 346.11 35.395 ;
    RECT 345.9 35.685 346.11 35.755 ;
    RECT 345.9 36.045 346.11 36.115 ;
    RECT 210.24 35.325 210.45 35.395 ;
    RECT 210.24 35.685 210.45 35.755 ;
    RECT 210.24 36.045 210.45 36.115 ;
    RECT 209.78 35.325 209.99 35.395 ;
    RECT 209.78 35.685 209.99 35.755 ;
    RECT 209.78 36.045 209.99 36.115 ;
    RECT 343.04 35.325 343.25 35.395 ;
    RECT 343.04 35.685 343.25 35.755 ;
    RECT 343.04 36.045 343.25 36.115 ;
    RECT 342.58 35.325 342.79 35.395 ;
    RECT 342.58 35.685 342.79 35.755 ;
    RECT 342.58 36.045 342.79 36.115 ;
    RECT 206.92 35.325 207.13 35.395 ;
    RECT 206.92 35.685 207.13 35.755 ;
    RECT 206.92 36.045 207.13 36.115 ;
    RECT 206.46 35.325 206.67 35.395 ;
    RECT 206.46 35.685 206.67 35.755 ;
    RECT 206.46 36.045 206.67 36.115 ;
    RECT 339.72 35.325 339.93 35.395 ;
    RECT 339.72 35.685 339.93 35.755 ;
    RECT 339.72 36.045 339.93 36.115 ;
    RECT 339.26 35.325 339.47 35.395 ;
    RECT 339.26 35.685 339.47 35.755 ;
    RECT 339.26 36.045 339.47 36.115 ;
    RECT 203.6 35.325 203.81 35.395 ;
    RECT 203.6 35.685 203.81 35.755 ;
    RECT 203.6 36.045 203.81 36.115 ;
    RECT 203.14 35.325 203.35 35.395 ;
    RECT 203.14 35.685 203.35 35.755 ;
    RECT 203.14 36.045 203.35 36.115 ;
    RECT 336.4 35.325 336.61 35.395 ;
    RECT 336.4 35.685 336.61 35.755 ;
    RECT 336.4 36.045 336.61 36.115 ;
    RECT 335.94 35.325 336.15 35.395 ;
    RECT 335.94 35.685 336.15 35.755 ;
    RECT 335.94 36.045 336.15 36.115 ;
    RECT 266.68 35.325 266.89 35.395 ;
    RECT 266.68 35.685 266.89 35.755 ;
    RECT 266.68 36.045 266.89 36.115 ;
    RECT 266.22 35.325 266.43 35.395 ;
    RECT 266.22 35.685 266.43 35.755 ;
    RECT 266.22 36.045 266.43 36.115 ;
    RECT 263.36 35.325 263.57 35.395 ;
    RECT 263.36 35.685 263.57 35.755 ;
    RECT 263.36 36.045 263.57 36.115 ;
    RECT 262.9 35.325 263.11 35.395 ;
    RECT 262.9 35.685 263.11 35.755 ;
    RECT 262.9 36.045 263.11 36.115 ;
    RECT 260.04 35.325 260.25 35.395 ;
    RECT 260.04 35.685 260.25 35.755 ;
    RECT 260.04 36.045 260.25 36.115 ;
    RECT 259.58 35.325 259.79 35.395 ;
    RECT 259.58 35.685 259.79 35.755 ;
    RECT 259.58 36.045 259.79 36.115 ;
    RECT 256.72 35.325 256.93 35.395 ;
    RECT 256.72 35.685 256.93 35.755 ;
    RECT 256.72 36.045 256.93 36.115 ;
    RECT 256.26 35.325 256.47 35.395 ;
    RECT 256.26 35.685 256.47 35.755 ;
    RECT 256.26 36.045 256.47 36.115 ;
    RECT 253.4 35.325 253.61 35.395 ;
    RECT 253.4 35.685 253.61 35.755 ;
    RECT 253.4 36.045 253.61 36.115 ;
    RECT 252.94 35.325 253.15 35.395 ;
    RECT 252.94 35.685 253.15 35.755 ;
    RECT 252.94 36.045 253.15 36.115 ;
    RECT 250.08 35.325 250.29 35.395 ;
    RECT 250.08 35.685 250.29 35.755 ;
    RECT 250.08 36.045 250.29 36.115 ;
    RECT 249.62 35.325 249.83 35.395 ;
    RECT 249.62 35.685 249.83 35.755 ;
    RECT 249.62 36.045 249.83 36.115 ;
    RECT 246.76 35.325 246.97 35.395 ;
    RECT 246.76 35.685 246.97 35.755 ;
    RECT 246.76 36.045 246.97 36.115 ;
    RECT 246.3 35.325 246.51 35.395 ;
    RECT 246.3 35.685 246.51 35.755 ;
    RECT 246.3 36.045 246.51 36.115 ;
    RECT 243.44 35.325 243.65 35.395 ;
    RECT 243.44 35.685 243.65 35.755 ;
    RECT 243.44 36.045 243.65 36.115 ;
    RECT 242.98 35.325 243.19 35.395 ;
    RECT 242.98 35.685 243.19 35.755 ;
    RECT 242.98 36.045 243.19 36.115 ;
    RECT 240.12 35.325 240.33 35.395 ;
    RECT 240.12 35.685 240.33 35.755 ;
    RECT 240.12 36.045 240.33 36.115 ;
    RECT 239.66 35.325 239.87 35.395 ;
    RECT 239.66 35.685 239.87 35.755 ;
    RECT 239.66 36.045 239.87 36.115 ;
    RECT 236.8 35.325 237.01 35.395 ;
    RECT 236.8 35.685 237.01 35.755 ;
    RECT 236.8 36.045 237.01 36.115 ;
    RECT 236.34 35.325 236.55 35.395 ;
    RECT 236.34 35.685 236.55 35.755 ;
    RECT 236.34 36.045 236.55 36.115 ;
    RECT 200.605 35.685 200.675 35.755 ;
    RECT 333.08 35.325 333.29 35.395 ;
    RECT 333.08 35.685 333.29 35.755 ;
    RECT 333.08 36.045 333.29 36.115 ;
    RECT 332.62 35.325 332.83 35.395 ;
    RECT 332.62 35.685 332.83 35.755 ;
    RECT 332.62 36.045 332.83 36.115 ;
    RECT 329.76 35.325 329.97 35.395 ;
    RECT 329.76 35.685 329.97 35.755 ;
    RECT 329.76 36.045 329.97 36.115 ;
    RECT 329.3 35.325 329.51 35.395 ;
    RECT 329.3 35.685 329.51 35.755 ;
    RECT 329.3 36.045 329.51 36.115 ;
    RECT 326.44 35.325 326.65 35.395 ;
    RECT 326.44 35.685 326.65 35.755 ;
    RECT 326.44 36.045 326.65 36.115 ;
    RECT 325.98 35.325 326.19 35.395 ;
    RECT 325.98 35.685 326.19 35.755 ;
    RECT 325.98 36.045 326.19 36.115 ;
    RECT 323.12 35.325 323.33 35.395 ;
    RECT 323.12 35.685 323.33 35.755 ;
    RECT 323.12 36.045 323.33 36.115 ;
    RECT 322.66 35.325 322.87 35.395 ;
    RECT 322.66 35.685 322.87 35.755 ;
    RECT 322.66 36.045 322.87 36.115 ;
    RECT 319.8 35.325 320.01 35.395 ;
    RECT 319.8 35.685 320.01 35.755 ;
    RECT 319.8 36.045 320.01 36.115 ;
    RECT 319.34 35.325 319.55 35.395 ;
    RECT 319.34 35.685 319.55 35.755 ;
    RECT 319.34 36.045 319.55 36.115 ;
    RECT 316.48 35.325 316.69 35.395 ;
    RECT 316.48 35.685 316.69 35.755 ;
    RECT 316.48 36.045 316.69 36.115 ;
    RECT 316.02 35.325 316.23 35.395 ;
    RECT 316.02 35.685 316.23 35.755 ;
    RECT 316.02 36.045 316.23 36.115 ;
    RECT 313.16 35.325 313.37 35.395 ;
    RECT 313.16 35.685 313.37 35.755 ;
    RECT 313.16 36.045 313.37 36.115 ;
    RECT 312.7 35.325 312.91 35.395 ;
    RECT 312.7 35.685 312.91 35.755 ;
    RECT 312.7 36.045 312.91 36.115 ;
    RECT 309.84 35.325 310.05 35.395 ;
    RECT 309.84 35.685 310.05 35.755 ;
    RECT 309.84 36.045 310.05 36.115 ;
    RECT 309.38 35.325 309.59 35.395 ;
    RECT 309.38 35.685 309.59 35.755 ;
    RECT 309.38 36.045 309.59 36.115 ;
    RECT 306.52 35.325 306.73 35.395 ;
    RECT 306.52 35.685 306.73 35.755 ;
    RECT 306.52 36.045 306.73 36.115 ;
    RECT 306.06 35.325 306.27 35.395 ;
    RECT 306.06 35.685 306.27 35.755 ;
    RECT 306.06 36.045 306.27 36.115 ;
    RECT 328.81 59.605 329.02 59.675 ;
    RECT 292.78 59.345 292.99 59.415 ;
    RECT 279.01 59.605 279.22 59.675 ;
    RECT 293.24 59.345 293.45 59.415 ;
    RECT 345.9 59.345 346.11 59.415 ;
    RECT 346.36 59.345 346.57 59.415 ;
    RECT 358.69 59.865 358.9 59.935 ;
    RECT 298.93 59.865 299.14 59.935 ;
    RECT 368.65 59.865 368.86 59.935 ;
    RECT 225.89 59.605 226.1 59.675 ;
    RECT 308.89 59.865 309.1 59.935 ;
    RECT 219.74 59.345 219.95 59.415 ;
    RECT 325.49 59.605 325.7 59.675 ;
    RECT 265.73 59.605 265.94 59.675 ;
    RECT 289.46 59.345 289.67 59.415 ;
    RECT 289.92 59.345 290.13 59.415 ;
    RECT 249.13 59.865 249.34 59.935 ;
    RECT 220.2 59.345 220.41 59.415 ;
    RECT 342.58 59.345 342.79 59.415 ;
    RECT 343.04 59.345 343.25 59.415 ;
    RECT 355.37 59.865 355.58 59.935 ;
    RECT 295.61 59.865 295.82 59.935 ;
    RECT 305.57 59.865 305.78 59.935 ;
    RECT 262.41 59.605 262.62 59.675 ;
    RECT 286.14 59.345 286.35 59.415 ;
    RECT 245.81 59.865 246.02 59.935 ;
    RECT 332.62 59.345 332.83 59.415 ;
    RECT 333.08 59.345 333.29 59.415 ;
    RECT 222.57 59.605 222.78 59.675 ;
    RECT 216.42 59.345 216.63 59.415 ;
    RECT 216.88 59.345 217.09 59.415 ;
    RECT 322.17 59.605 322.38 59.675 ;
    RECT 339.26 59.345 339.47 59.415 ;
    RECT 352.05 59.865 352.26 59.935 ;
    RECT 339.72 59.345 339.93 59.415 ;
    RECT 292.29 59.865 292.5 59.935 ;
    RECT 286.6 59.345 286.81 59.415 ;
    RECT 302.25 59.865 302.46 59.935 ;
    RECT 259.09 59.605 259.3 59.675 ;
    RECT 242.49 59.865 242.7 59.935 ;
    RECT 329.3 59.345 329.51 59.415 ;
    RECT 329.76 59.345 329.97 59.415 ;
    RECT 219.25 59.605 219.46 59.675 ;
    RECT 213.1 59.345 213.31 59.415 ;
    RECT 213.56 59.345 213.77 59.415 ;
    RECT 318.85 59.605 319.06 59.675 ;
    RECT 335.94 59.345 336.15 59.415 ;
    RECT 288.97 59.865 289.18 59.935 ;
    RECT 282.82 59.345 283.03 59.415 ;
    RECT 283.28 59.345 283.49 59.415 ;
    RECT 239.17 59.865 239.38 59.935 ;
    RECT 348.73 59.865 348.94 59.935 ;
    RECT 325.98 59.345 326.19 59.415 ;
    RECT 336.4 59.345 336.61 59.415 ;
    RECT 326.44 59.345 326.65 59.415 ;
    RECT 215.93 59.605 216.14 59.675 ;
    RECT 365.33 59.605 365.54 59.675 ;
    RECT 209.78 59.345 209.99 59.415 ;
    RECT 315.53 59.605 315.74 59.675 ;
    RECT 210.24 59.345 210.45 59.415 ;
    RECT 255.77 59.605 255.98 59.675 ;
    RECT 285.65 59.865 285.86 59.935 ;
    RECT 279.5 59.345 279.71 59.415 ;
    RECT 279.96 59.345 280.17 59.415 ;
    RECT 235.85 59.865 236.06 59.935 ;
    RECT 345.41 59.865 345.62 59.935 ;
    RECT 322.66 59.345 322.87 59.415 ;
    RECT 323.12 59.345 323.33 59.415 ;
    RECT 212.61 59.605 212.82 59.675 ;
    RECT 362.01 59.605 362.22 59.675 ;
    RECT 371.97 59.605 372.18 59.675 ;
    RECT 312.21 59.605 312.42 59.675 ;
    RECT 206.46 59.345 206.67 59.415 ;
    RECT 252.45 59.605 252.66 59.675 ;
    RECT 206.92 59.345 207.13 59.415 ;
    RECT 233.935 60.125 234.155 60.195 ;
    RECT 276.18 59.345 276.39 59.415 ;
    RECT 230.615 60.125 230.835 60.195 ;
    RECT 276.64 59.345 276.85 59.415 ;
    RECT 227.295 60.125 227.515 60.195 ;
    RECT 223.975 60.125 224.195 60.195 ;
    RECT 220.655 60.125 220.875 60.195 ;
    RECT 217.335 60.125 217.555 60.195 ;
    RECT 214.015 60.125 214.235 60.195 ;
    RECT 210.695 60.125 210.915 60.195 ;
    RECT 207.375 60.125 207.595 60.195 ;
    RECT 204.055 60.125 204.275 60.195 ;
    RECT 342.09 59.865 342.3 59.935 ;
    RECT 282.33 59.865 282.54 59.935 ;
    RECT 319.34 59.345 319.55 59.415 ;
    RECT 209.29 59.605 209.5 59.675 ;
    RECT 266.22 59.345 266.43 59.415 ;
    RECT 266.68 59.345 266.89 59.415 ;
    RECT 358.69 59.605 358.9 59.675 ;
    RECT 368.65 59.605 368.86 59.675 ;
    RECT 308.89 59.605 309.1 59.675 ;
    RECT 249.13 59.605 249.34 59.675 ;
    RECT 203.14 59.345 203.35 59.415 ;
    RECT 272.86 59.345 273.07 59.415 ;
    RECT 273.32 59.345 273.53 59.415 ;
    RECT 319.8 59.345 320.01 59.415 ;
    RECT 232.53 59.865 232.74 59.935 ;
    RECT 373.375 60.125 373.595 60.195 ;
    RECT 370.055 60.125 370.275 60.195 ;
    RECT 203.6 59.345 203.81 59.415 ;
    RECT 372.46 59.345 372.67 59.415 ;
    RECT 338.77 59.865 338.98 59.935 ;
    RECT 372.92 59.345 373.13 59.415 ;
    RECT 279.01 59.865 279.22 59.935 ;
    RECT 205.97 59.605 206.18 59.675 ;
    RECT 262.9 59.345 263.11 59.415 ;
    RECT 263.36 59.345 263.57 59.415 ;
    RECT 305.57 59.605 305.78 59.675 ;
    RECT 245.81 59.605 246.02 59.675 ;
    RECT 366.735 60.125 366.955 60.195 ;
    RECT 363.415 60.125 363.635 60.195 ;
    RECT 360.095 60.125 360.315 60.195 ;
    RECT 269.54 59.345 269.75 59.415 ;
    RECT 356.775 60.125 356.995 60.195 ;
    RECT 353.455 60.125 353.675 60.195 ;
    RECT 350.135 60.125 350.355 60.195 ;
    RECT 346.815 60.125 347.035 60.195 ;
    RECT 343.495 60.125 343.715 60.195 ;
    RECT 340.175 60.125 340.395 60.195 ;
    RECT 316.02 59.345 316.23 59.415 ;
    RECT 229.21 59.865 229.42 59.935 ;
    RECT 336.855 60.125 337.075 60.195 ;
    RECT 316.48 59.345 316.69 59.415 ;
    RECT 355.37 59.605 355.58 59.675 ;
    RECT 335.45 59.865 335.66 59.935 ;
    RECT 369.14 59.345 369.35 59.415 ;
    RECT 275.69 59.865 275.9 59.935 ;
    RECT 202.65 59.605 202.86 59.675 ;
    RECT 259.58 59.345 259.79 59.415 ;
    RECT 270.0 59.345 270.21 59.415 ;
    RECT 260.04 59.345 260.25 59.415 ;
    RECT 302.25 59.605 302.46 59.675 ;
    RECT 242.49 59.605 242.7 59.675 ;
    RECT 333.535 60.125 333.755 60.195 ;
    RECT 330.215 60.125 330.435 60.195 ;
    RECT 326.895 60.125 327.115 60.195 ;
    RECT 323.575 60.125 323.795 60.195 ;
    RECT 320.255 60.125 320.475 60.195 ;
    RECT 316.935 60.125 317.155 60.195 ;
    RECT 313.615 60.125 313.835 60.195 ;
    RECT 310.295 60.125 310.515 60.195 ;
    RECT 306.975 60.125 307.195 60.195 ;
    RECT 303.655 60.125 303.875 60.195 ;
    RECT 369.6 59.345 369.81 59.415 ;
    RECT 225.89 59.865 226.1 59.935 ;
    RECT 312.7 59.345 312.91 59.415 ;
    RECT 313.16 59.345 313.37 59.415 ;
    RECT 352.05 59.605 352.26 59.675 ;
    RECT 272.37 59.865 272.58 59.935 ;
    RECT 256.26 59.345 256.47 59.415 ;
    RECT 256.72 59.345 256.93 59.415 ;
    RECT 300.335 60.125 300.555 60.195 ;
    RECT 297.015 60.125 297.235 60.195 ;
    RECT 293.695 60.125 293.915 60.195 ;
    RECT 239.17 59.605 239.38 59.675 ;
    RECT 290.375 60.125 290.595 60.195 ;
    RECT 287.055 60.125 287.275 60.195 ;
    RECT 283.735 60.125 283.955 60.195 ;
    RECT 280.415 60.125 280.635 60.195 ;
    RECT 277.095 60.125 277.315 60.195 ;
    RECT 273.775 60.125 273.995 60.195 ;
    RECT 270.455 60.125 270.675 60.195 ;
    RECT 222.57 59.865 222.78 59.935 ;
    RECT 309.38 59.345 309.59 59.415 ;
    RECT 309.84 59.345 310.05 59.415 ;
    RECT 348.73 59.605 348.94 59.675 ;
    RECT 269.05 59.865 269.26 59.935 ;
    RECT 267.135 60.125 267.355 60.195 ;
    RECT 263.815 60.125 264.035 60.195 ;
    RECT 260.495 60.125 260.715 60.195 ;
    RECT 257.175 60.125 257.395 60.195 ;
    RECT 252.94 59.345 253.15 59.415 ;
    RECT 253.855 60.125 254.075 60.195 ;
    RECT 250.535 60.125 250.755 60.195 ;
    RECT 247.215 60.125 247.435 60.195 ;
    RECT 235.85 59.605 236.06 59.675 ;
    RECT 243.895 60.125 244.115 60.195 ;
    RECT 240.575 60.125 240.795 60.195 ;
    RECT 237.255 60.125 237.475 60.195 ;
    RECT 219.25 59.865 219.46 59.935 ;
    RECT 306.06 59.345 306.27 59.415 ;
    RECT 345.41 59.605 345.62 59.675 ;
    RECT 306.52 59.345 306.73 59.415 ;
    RECT 253.4 59.345 253.61 59.415 ;
    RECT 332.13 59.865 332.34 59.935 ;
    RECT 298.93 59.605 299.14 59.675 ;
    RECT 365.82 59.345 366.03 59.415 ;
    RECT 342.09 59.605 342.3 59.675 ;
    RECT 302.74 59.345 302.95 59.415 ;
    RECT 366.28 59.345 366.49 59.415 ;
    RECT 249.62 59.345 249.83 59.415 ;
    RECT 250.08 59.345 250.29 59.415 ;
    RECT 328.81 59.865 329.02 59.935 ;
    RECT 215.93 59.865 216.14 59.935 ;
    RECT 295.61 59.605 295.82 59.675 ;
    RECT 303.2 59.345 303.41 59.415 ;
    RECT 338.77 59.605 338.98 59.675 ;
    RECT 362.5 59.345 362.71 59.415 ;
    RECT 362.96 59.345 363.17 59.415 ;
    RECT 246.3 59.345 246.51 59.415 ;
    RECT 246.76 59.345 246.97 59.415 ;
    RECT 325.49 59.865 325.7 59.935 ;
    RECT 265.73 59.865 265.94 59.935 ;
    RECT 212.61 59.865 212.82 59.935 ;
    RECT 292.29 59.605 292.5 59.675 ;
    RECT 335.45 59.605 335.66 59.675 ;
    RECT 275.69 59.605 275.9 59.675 ;
    RECT 359.18 59.345 359.39 59.415 ;
    RECT 359.64 59.345 359.85 59.415 ;
    RECT 242.98 59.345 243.19 59.415 ;
    RECT 243.44 59.345 243.65 59.415 ;
    RECT 322.17 59.865 322.38 59.935 ;
    RECT 262.41 59.865 262.62 59.935 ;
    RECT 209.29 59.865 209.5 59.935 ;
    RECT 233.02 59.345 233.23 59.415 ;
    RECT 233.48 59.345 233.69 59.415 ;
    RECT 272.37 59.605 272.58 59.675 ;
    RECT 355.86 59.345 356.07 59.415 ;
    RECT 356.32 59.345 356.53 59.415 ;
    RECT 239.66 59.345 239.87 59.415 ;
    RECT 240.12 59.345 240.33 59.415 ;
    RECT 288.97 59.605 289.18 59.675 ;
    RECT 318.85 59.865 319.06 59.935 ;
    RECT 259.09 59.865 259.3 59.935 ;
    RECT 205.97 59.865 206.18 59.935 ;
    RECT 229.7 59.345 229.91 59.415 ;
    RECT 230.16 59.345 230.37 59.415 ;
    RECT 269.05 59.605 269.26 59.675 ;
    RECT 352.54 59.345 352.75 59.415 ;
    RECT 299.42 59.345 299.63 59.415 ;
    RECT 236.34 59.345 236.55 59.415 ;
    RECT 299.88 59.345 300.09 59.415 ;
    RECT 285.65 59.605 285.86 59.675 ;
    RECT 255.77 59.865 255.98 59.935 ;
    RECT 202.65 59.865 202.86 59.935 ;
    RECT 353.0 59.345 353.21 59.415 ;
    RECT 236.8 59.345 237.01 59.415 ;
    RECT 365.33 59.865 365.54 59.935 ;
    RECT 374.36 59.605 374.43 59.675 ;
    RECT 374.15 59.345 374.22 59.415 ;
    RECT 232.53 59.605 232.74 59.675 ;
    RECT 315.53 59.865 315.74 59.935 ;
    RECT 226.38 59.345 226.59 59.415 ;
    RECT 226.84 59.345 227.05 59.415 ;
    RECT 200.395 59.605 200.465 59.675 ;
    RECT 200.605 59.345 200.675 59.415 ;
    RECT 332.13 59.605 332.34 59.675 ;
    RECT 296.1 59.345 296.31 59.415 ;
    RECT 296.56 59.345 296.77 59.415 ;
    RECT 282.33 59.605 282.54 59.675 ;
    RECT 252.45 59.865 252.66 59.935 ;
    RECT 349.22 59.345 349.43 59.415 ;
    RECT 349.68 59.345 349.89 59.415 ;
    RECT 362.01 59.865 362.22 59.935 ;
    RECT 371.97 59.865 372.18 59.935 ;
    RECT 229.21 59.605 229.42 59.675 ;
    RECT 312.21 59.865 312.42 59.935 ;
    RECT 223.06 59.345 223.27 59.415 ;
    RECT 223.52 59.345 223.73 59.415 ;
    RECT 303.2 25.245 303.41 25.315 ;
    RECT 303.2 25.605 303.41 25.675 ;
    RECT 303.2 25.965 303.41 26.035 ;
    RECT 302.74 25.245 302.95 25.315 ;
    RECT 302.74 25.605 302.95 25.675 ;
    RECT 302.74 25.965 302.95 26.035 ;
    RECT 372.92 25.245 373.13 25.315 ;
    RECT 372.92 25.605 373.13 25.675 ;
    RECT 372.92 25.965 373.13 26.035 ;
    RECT 372.46 25.245 372.67 25.315 ;
    RECT 372.46 25.605 372.67 25.675 ;
    RECT 372.46 25.965 372.67 26.035 ;
    RECT 369.6 25.245 369.81 25.315 ;
    RECT 369.6 25.605 369.81 25.675 ;
    RECT 369.6 25.965 369.81 26.035 ;
    RECT 369.14 25.245 369.35 25.315 ;
    RECT 369.14 25.605 369.35 25.675 ;
    RECT 369.14 25.965 369.35 26.035 ;
    RECT 200.605 25.605 200.675 25.675 ;
    RECT 299.88 25.245 300.09 25.315 ;
    RECT 299.88 25.605 300.09 25.675 ;
    RECT 299.88 25.965 300.09 26.035 ;
    RECT 299.42 25.245 299.63 25.315 ;
    RECT 299.42 25.605 299.63 25.675 ;
    RECT 299.42 25.965 299.63 26.035 ;
    RECT 296.56 25.245 296.77 25.315 ;
    RECT 296.56 25.605 296.77 25.675 ;
    RECT 296.56 25.965 296.77 26.035 ;
    RECT 296.1 25.245 296.31 25.315 ;
    RECT 296.1 25.605 296.31 25.675 ;
    RECT 296.1 25.965 296.31 26.035 ;
    RECT 293.24 25.245 293.45 25.315 ;
    RECT 293.24 25.605 293.45 25.675 ;
    RECT 293.24 25.965 293.45 26.035 ;
    RECT 292.78 25.245 292.99 25.315 ;
    RECT 292.78 25.605 292.99 25.675 ;
    RECT 292.78 25.965 292.99 26.035 ;
    RECT 289.92 25.245 290.13 25.315 ;
    RECT 289.92 25.605 290.13 25.675 ;
    RECT 289.92 25.965 290.13 26.035 ;
    RECT 289.46 25.245 289.67 25.315 ;
    RECT 289.46 25.605 289.67 25.675 ;
    RECT 289.46 25.965 289.67 26.035 ;
    RECT 286.6 25.245 286.81 25.315 ;
    RECT 286.6 25.605 286.81 25.675 ;
    RECT 286.6 25.965 286.81 26.035 ;
    RECT 286.14 25.245 286.35 25.315 ;
    RECT 286.14 25.605 286.35 25.675 ;
    RECT 286.14 25.965 286.35 26.035 ;
    RECT 283.28 25.245 283.49 25.315 ;
    RECT 283.28 25.605 283.49 25.675 ;
    RECT 283.28 25.965 283.49 26.035 ;
    RECT 282.82 25.245 283.03 25.315 ;
    RECT 282.82 25.605 283.03 25.675 ;
    RECT 282.82 25.965 283.03 26.035 ;
    RECT 279.96 25.245 280.17 25.315 ;
    RECT 279.96 25.605 280.17 25.675 ;
    RECT 279.96 25.965 280.17 26.035 ;
    RECT 279.5 25.245 279.71 25.315 ;
    RECT 279.5 25.605 279.71 25.675 ;
    RECT 279.5 25.965 279.71 26.035 ;
    RECT 276.64 25.245 276.85 25.315 ;
    RECT 276.64 25.605 276.85 25.675 ;
    RECT 276.64 25.965 276.85 26.035 ;
    RECT 276.18 25.245 276.39 25.315 ;
    RECT 276.18 25.605 276.39 25.675 ;
    RECT 276.18 25.965 276.39 26.035 ;
    RECT 273.32 25.245 273.53 25.315 ;
    RECT 273.32 25.605 273.53 25.675 ;
    RECT 273.32 25.965 273.53 26.035 ;
    RECT 272.86 25.245 273.07 25.315 ;
    RECT 272.86 25.605 273.07 25.675 ;
    RECT 272.86 25.965 273.07 26.035 ;
    RECT 270.0 25.245 270.21 25.315 ;
    RECT 270.0 25.605 270.21 25.675 ;
    RECT 270.0 25.965 270.21 26.035 ;
    RECT 269.54 25.245 269.75 25.315 ;
    RECT 269.54 25.605 269.75 25.675 ;
    RECT 269.54 25.965 269.75 26.035 ;
    RECT 233.48 25.245 233.69 25.315 ;
    RECT 233.48 25.605 233.69 25.675 ;
    RECT 233.48 25.965 233.69 26.035 ;
    RECT 233.02 25.245 233.23 25.315 ;
    RECT 233.02 25.605 233.23 25.675 ;
    RECT 233.02 25.965 233.23 26.035 ;
    RECT 230.16 25.245 230.37 25.315 ;
    RECT 230.16 25.605 230.37 25.675 ;
    RECT 230.16 25.965 230.37 26.035 ;
    RECT 229.7 25.245 229.91 25.315 ;
    RECT 229.7 25.605 229.91 25.675 ;
    RECT 229.7 25.965 229.91 26.035 ;
    RECT 366.28 25.245 366.49 25.315 ;
    RECT 366.28 25.605 366.49 25.675 ;
    RECT 366.28 25.965 366.49 26.035 ;
    RECT 365.82 25.245 366.03 25.315 ;
    RECT 365.82 25.605 366.03 25.675 ;
    RECT 365.82 25.965 366.03 26.035 ;
    RECT 226.84 25.245 227.05 25.315 ;
    RECT 226.84 25.605 227.05 25.675 ;
    RECT 226.84 25.965 227.05 26.035 ;
    RECT 226.38 25.245 226.59 25.315 ;
    RECT 226.38 25.605 226.59 25.675 ;
    RECT 226.38 25.965 226.59 26.035 ;
    RECT 362.96 25.245 363.17 25.315 ;
    RECT 362.96 25.605 363.17 25.675 ;
    RECT 362.96 25.965 363.17 26.035 ;
    RECT 362.5 25.245 362.71 25.315 ;
    RECT 362.5 25.605 362.71 25.675 ;
    RECT 362.5 25.965 362.71 26.035 ;
    RECT 223.52 25.245 223.73 25.315 ;
    RECT 223.52 25.605 223.73 25.675 ;
    RECT 223.52 25.965 223.73 26.035 ;
    RECT 223.06 25.245 223.27 25.315 ;
    RECT 223.06 25.605 223.27 25.675 ;
    RECT 223.06 25.965 223.27 26.035 ;
    RECT 359.64 25.245 359.85 25.315 ;
    RECT 359.64 25.605 359.85 25.675 ;
    RECT 359.64 25.965 359.85 26.035 ;
    RECT 359.18 25.245 359.39 25.315 ;
    RECT 359.18 25.605 359.39 25.675 ;
    RECT 359.18 25.965 359.39 26.035 ;
    RECT 220.2 25.245 220.41 25.315 ;
    RECT 220.2 25.605 220.41 25.675 ;
    RECT 220.2 25.965 220.41 26.035 ;
    RECT 219.74 25.245 219.95 25.315 ;
    RECT 219.74 25.605 219.95 25.675 ;
    RECT 219.74 25.965 219.95 26.035 ;
    RECT 356.32 25.245 356.53 25.315 ;
    RECT 356.32 25.605 356.53 25.675 ;
    RECT 356.32 25.965 356.53 26.035 ;
    RECT 355.86 25.245 356.07 25.315 ;
    RECT 355.86 25.605 356.07 25.675 ;
    RECT 355.86 25.965 356.07 26.035 ;
    RECT 353.0 25.245 353.21 25.315 ;
    RECT 353.0 25.605 353.21 25.675 ;
    RECT 353.0 25.965 353.21 26.035 ;
    RECT 352.54 25.245 352.75 25.315 ;
    RECT 352.54 25.605 352.75 25.675 ;
    RECT 352.54 25.965 352.75 26.035 ;
    RECT 216.88 25.245 217.09 25.315 ;
    RECT 216.88 25.605 217.09 25.675 ;
    RECT 216.88 25.965 217.09 26.035 ;
    RECT 216.42 25.245 216.63 25.315 ;
    RECT 216.42 25.605 216.63 25.675 ;
    RECT 216.42 25.965 216.63 26.035 ;
    RECT 349.68 25.245 349.89 25.315 ;
    RECT 349.68 25.605 349.89 25.675 ;
    RECT 349.68 25.965 349.89 26.035 ;
    RECT 349.22 25.245 349.43 25.315 ;
    RECT 349.22 25.605 349.43 25.675 ;
    RECT 349.22 25.965 349.43 26.035 ;
    RECT 213.56 25.245 213.77 25.315 ;
    RECT 213.56 25.605 213.77 25.675 ;
    RECT 213.56 25.965 213.77 26.035 ;
    RECT 213.1 25.245 213.31 25.315 ;
    RECT 213.1 25.605 213.31 25.675 ;
    RECT 213.1 25.965 213.31 26.035 ;
    RECT 346.36 25.245 346.57 25.315 ;
    RECT 346.36 25.605 346.57 25.675 ;
    RECT 346.36 25.965 346.57 26.035 ;
    RECT 345.9 25.245 346.11 25.315 ;
    RECT 345.9 25.605 346.11 25.675 ;
    RECT 345.9 25.965 346.11 26.035 ;
    RECT 210.24 25.245 210.45 25.315 ;
    RECT 210.24 25.605 210.45 25.675 ;
    RECT 210.24 25.965 210.45 26.035 ;
    RECT 209.78 25.245 209.99 25.315 ;
    RECT 209.78 25.605 209.99 25.675 ;
    RECT 209.78 25.965 209.99 26.035 ;
    RECT 343.04 25.245 343.25 25.315 ;
    RECT 343.04 25.605 343.25 25.675 ;
    RECT 343.04 25.965 343.25 26.035 ;
    RECT 342.58 25.245 342.79 25.315 ;
    RECT 342.58 25.605 342.79 25.675 ;
    RECT 342.58 25.965 342.79 26.035 ;
    RECT 206.92 25.245 207.13 25.315 ;
    RECT 206.92 25.605 207.13 25.675 ;
    RECT 206.92 25.965 207.13 26.035 ;
    RECT 206.46 25.245 206.67 25.315 ;
    RECT 206.46 25.605 206.67 25.675 ;
    RECT 206.46 25.965 206.67 26.035 ;
    RECT 339.72 25.245 339.93 25.315 ;
    RECT 339.72 25.605 339.93 25.675 ;
    RECT 339.72 25.965 339.93 26.035 ;
    RECT 339.26 25.245 339.47 25.315 ;
    RECT 339.26 25.605 339.47 25.675 ;
    RECT 339.26 25.965 339.47 26.035 ;
    RECT 203.6 25.245 203.81 25.315 ;
    RECT 203.6 25.605 203.81 25.675 ;
    RECT 203.6 25.965 203.81 26.035 ;
    RECT 203.14 25.245 203.35 25.315 ;
    RECT 203.14 25.605 203.35 25.675 ;
    RECT 203.14 25.965 203.35 26.035 ;
    RECT 336.4 25.245 336.61 25.315 ;
    RECT 336.4 25.605 336.61 25.675 ;
    RECT 336.4 25.965 336.61 26.035 ;
    RECT 335.94 25.245 336.15 25.315 ;
    RECT 335.94 25.605 336.15 25.675 ;
    RECT 335.94 25.965 336.15 26.035 ;
    RECT 266.68 25.245 266.89 25.315 ;
    RECT 266.68 25.605 266.89 25.675 ;
    RECT 266.68 25.965 266.89 26.035 ;
    RECT 266.22 25.245 266.43 25.315 ;
    RECT 266.22 25.605 266.43 25.675 ;
    RECT 266.22 25.965 266.43 26.035 ;
    RECT 263.36 25.245 263.57 25.315 ;
    RECT 263.36 25.605 263.57 25.675 ;
    RECT 263.36 25.965 263.57 26.035 ;
    RECT 262.9 25.245 263.11 25.315 ;
    RECT 262.9 25.605 263.11 25.675 ;
    RECT 262.9 25.965 263.11 26.035 ;
    RECT 260.04 25.245 260.25 25.315 ;
    RECT 260.04 25.605 260.25 25.675 ;
    RECT 260.04 25.965 260.25 26.035 ;
    RECT 259.58 25.245 259.79 25.315 ;
    RECT 259.58 25.605 259.79 25.675 ;
    RECT 259.58 25.965 259.79 26.035 ;
    RECT 256.72 25.245 256.93 25.315 ;
    RECT 256.72 25.605 256.93 25.675 ;
    RECT 256.72 25.965 256.93 26.035 ;
    RECT 256.26 25.245 256.47 25.315 ;
    RECT 256.26 25.605 256.47 25.675 ;
    RECT 256.26 25.965 256.47 26.035 ;
    RECT 253.4 25.245 253.61 25.315 ;
    RECT 253.4 25.605 253.61 25.675 ;
    RECT 253.4 25.965 253.61 26.035 ;
    RECT 252.94 25.245 253.15 25.315 ;
    RECT 252.94 25.605 253.15 25.675 ;
    RECT 252.94 25.965 253.15 26.035 ;
    RECT 250.08 25.245 250.29 25.315 ;
    RECT 250.08 25.605 250.29 25.675 ;
    RECT 250.08 25.965 250.29 26.035 ;
    RECT 249.62 25.245 249.83 25.315 ;
    RECT 249.62 25.605 249.83 25.675 ;
    RECT 249.62 25.965 249.83 26.035 ;
    RECT 246.76 25.245 246.97 25.315 ;
    RECT 246.76 25.605 246.97 25.675 ;
    RECT 246.76 25.965 246.97 26.035 ;
    RECT 246.3 25.245 246.51 25.315 ;
    RECT 246.3 25.605 246.51 25.675 ;
    RECT 246.3 25.965 246.51 26.035 ;
    RECT 243.44 25.245 243.65 25.315 ;
    RECT 243.44 25.605 243.65 25.675 ;
    RECT 243.44 25.965 243.65 26.035 ;
    RECT 242.98 25.245 243.19 25.315 ;
    RECT 242.98 25.605 243.19 25.675 ;
    RECT 242.98 25.965 243.19 26.035 ;
    RECT 240.12 25.245 240.33 25.315 ;
    RECT 240.12 25.605 240.33 25.675 ;
    RECT 240.12 25.965 240.33 26.035 ;
    RECT 239.66 25.245 239.87 25.315 ;
    RECT 239.66 25.605 239.87 25.675 ;
    RECT 239.66 25.965 239.87 26.035 ;
    RECT 236.8 25.245 237.01 25.315 ;
    RECT 236.8 25.605 237.01 25.675 ;
    RECT 236.8 25.965 237.01 26.035 ;
    RECT 236.34 25.245 236.55 25.315 ;
    RECT 236.34 25.605 236.55 25.675 ;
    RECT 236.34 25.965 236.55 26.035 ;
    RECT 374.15 25.605 374.22 25.675 ;
    RECT 333.08 25.245 333.29 25.315 ;
    RECT 333.08 25.605 333.29 25.675 ;
    RECT 333.08 25.965 333.29 26.035 ;
    RECT 332.62 25.245 332.83 25.315 ;
    RECT 332.62 25.605 332.83 25.675 ;
    RECT 332.62 25.965 332.83 26.035 ;
    RECT 329.76 25.245 329.97 25.315 ;
    RECT 329.76 25.605 329.97 25.675 ;
    RECT 329.76 25.965 329.97 26.035 ;
    RECT 329.3 25.245 329.51 25.315 ;
    RECT 329.3 25.605 329.51 25.675 ;
    RECT 329.3 25.965 329.51 26.035 ;
    RECT 326.44 25.245 326.65 25.315 ;
    RECT 326.44 25.605 326.65 25.675 ;
    RECT 326.44 25.965 326.65 26.035 ;
    RECT 325.98 25.245 326.19 25.315 ;
    RECT 325.98 25.605 326.19 25.675 ;
    RECT 325.98 25.965 326.19 26.035 ;
    RECT 323.12 25.245 323.33 25.315 ;
    RECT 323.12 25.605 323.33 25.675 ;
    RECT 323.12 25.965 323.33 26.035 ;
    RECT 322.66 25.245 322.87 25.315 ;
    RECT 322.66 25.605 322.87 25.675 ;
    RECT 322.66 25.965 322.87 26.035 ;
    RECT 319.8 25.245 320.01 25.315 ;
    RECT 319.8 25.605 320.01 25.675 ;
    RECT 319.8 25.965 320.01 26.035 ;
    RECT 319.34 25.245 319.55 25.315 ;
    RECT 319.34 25.605 319.55 25.675 ;
    RECT 319.34 25.965 319.55 26.035 ;
    RECT 316.48 25.245 316.69 25.315 ;
    RECT 316.48 25.605 316.69 25.675 ;
    RECT 316.48 25.965 316.69 26.035 ;
    RECT 316.02 25.245 316.23 25.315 ;
    RECT 316.02 25.605 316.23 25.675 ;
    RECT 316.02 25.965 316.23 26.035 ;
    RECT 313.16 25.245 313.37 25.315 ;
    RECT 313.16 25.605 313.37 25.675 ;
    RECT 313.16 25.965 313.37 26.035 ;
    RECT 312.7 25.245 312.91 25.315 ;
    RECT 312.7 25.605 312.91 25.675 ;
    RECT 312.7 25.965 312.91 26.035 ;
    RECT 309.84 25.245 310.05 25.315 ;
    RECT 309.84 25.605 310.05 25.675 ;
    RECT 309.84 25.965 310.05 26.035 ;
    RECT 309.38 25.245 309.59 25.315 ;
    RECT 309.38 25.605 309.59 25.675 ;
    RECT 309.38 25.965 309.59 26.035 ;
    RECT 306.52 25.245 306.73 25.315 ;
    RECT 306.52 25.605 306.73 25.675 ;
    RECT 306.52 25.965 306.73 26.035 ;
    RECT 306.06 25.245 306.27 25.315 ;
    RECT 306.06 25.605 306.27 25.675 ;
    RECT 306.06 25.965 306.27 26.035 ;
    RECT 303.2 24.525 303.41 24.595 ;
    RECT 303.2 24.885 303.41 24.955 ;
    RECT 303.2 25.245 303.41 25.315 ;
    RECT 302.74 24.525 302.95 24.595 ;
    RECT 302.74 24.885 302.95 24.955 ;
    RECT 302.74 25.245 302.95 25.315 ;
    RECT 372.92 24.525 373.13 24.595 ;
    RECT 372.92 24.885 373.13 24.955 ;
    RECT 372.92 25.245 373.13 25.315 ;
    RECT 372.46 24.525 372.67 24.595 ;
    RECT 372.46 24.885 372.67 24.955 ;
    RECT 372.46 25.245 372.67 25.315 ;
    RECT 369.6 24.525 369.81 24.595 ;
    RECT 369.6 24.885 369.81 24.955 ;
    RECT 369.6 25.245 369.81 25.315 ;
    RECT 369.14 24.525 369.35 24.595 ;
    RECT 369.14 24.885 369.35 24.955 ;
    RECT 369.14 25.245 369.35 25.315 ;
    RECT 200.605 24.885 200.675 24.955 ;
    RECT 299.88 24.525 300.09 24.595 ;
    RECT 299.88 24.885 300.09 24.955 ;
    RECT 299.88 25.245 300.09 25.315 ;
    RECT 299.42 24.525 299.63 24.595 ;
    RECT 299.42 24.885 299.63 24.955 ;
    RECT 299.42 25.245 299.63 25.315 ;
    RECT 296.56 24.525 296.77 24.595 ;
    RECT 296.56 24.885 296.77 24.955 ;
    RECT 296.56 25.245 296.77 25.315 ;
    RECT 296.1 24.525 296.31 24.595 ;
    RECT 296.1 24.885 296.31 24.955 ;
    RECT 296.1 25.245 296.31 25.315 ;
    RECT 293.24 24.525 293.45 24.595 ;
    RECT 293.24 24.885 293.45 24.955 ;
    RECT 293.24 25.245 293.45 25.315 ;
    RECT 292.78 24.525 292.99 24.595 ;
    RECT 292.78 24.885 292.99 24.955 ;
    RECT 292.78 25.245 292.99 25.315 ;
    RECT 289.92 24.525 290.13 24.595 ;
    RECT 289.92 24.885 290.13 24.955 ;
    RECT 289.92 25.245 290.13 25.315 ;
    RECT 289.46 24.525 289.67 24.595 ;
    RECT 289.46 24.885 289.67 24.955 ;
    RECT 289.46 25.245 289.67 25.315 ;
    RECT 286.6 24.525 286.81 24.595 ;
    RECT 286.6 24.885 286.81 24.955 ;
    RECT 286.6 25.245 286.81 25.315 ;
    RECT 286.14 24.525 286.35 24.595 ;
    RECT 286.14 24.885 286.35 24.955 ;
    RECT 286.14 25.245 286.35 25.315 ;
    RECT 283.28 24.525 283.49 24.595 ;
    RECT 283.28 24.885 283.49 24.955 ;
    RECT 283.28 25.245 283.49 25.315 ;
    RECT 282.82 24.525 283.03 24.595 ;
    RECT 282.82 24.885 283.03 24.955 ;
    RECT 282.82 25.245 283.03 25.315 ;
    RECT 279.96 24.525 280.17 24.595 ;
    RECT 279.96 24.885 280.17 24.955 ;
    RECT 279.96 25.245 280.17 25.315 ;
    RECT 279.5 24.525 279.71 24.595 ;
    RECT 279.5 24.885 279.71 24.955 ;
    RECT 279.5 25.245 279.71 25.315 ;
    RECT 276.64 24.525 276.85 24.595 ;
    RECT 276.64 24.885 276.85 24.955 ;
    RECT 276.64 25.245 276.85 25.315 ;
    RECT 276.18 24.525 276.39 24.595 ;
    RECT 276.18 24.885 276.39 24.955 ;
    RECT 276.18 25.245 276.39 25.315 ;
    RECT 273.32 24.525 273.53 24.595 ;
    RECT 273.32 24.885 273.53 24.955 ;
    RECT 273.32 25.245 273.53 25.315 ;
    RECT 272.86 24.525 273.07 24.595 ;
    RECT 272.86 24.885 273.07 24.955 ;
    RECT 272.86 25.245 273.07 25.315 ;
    RECT 270.0 24.525 270.21 24.595 ;
    RECT 270.0 24.885 270.21 24.955 ;
    RECT 270.0 25.245 270.21 25.315 ;
    RECT 269.54 24.525 269.75 24.595 ;
    RECT 269.54 24.885 269.75 24.955 ;
    RECT 269.54 25.245 269.75 25.315 ;
    RECT 233.48 24.525 233.69 24.595 ;
    RECT 233.48 24.885 233.69 24.955 ;
    RECT 233.48 25.245 233.69 25.315 ;
    RECT 233.02 24.525 233.23 24.595 ;
    RECT 233.02 24.885 233.23 24.955 ;
    RECT 233.02 25.245 233.23 25.315 ;
    RECT 230.16 24.525 230.37 24.595 ;
    RECT 230.16 24.885 230.37 24.955 ;
    RECT 230.16 25.245 230.37 25.315 ;
    RECT 229.7 24.525 229.91 24.595 ;
    RECT 229.7 24.885 229.91 24.955 ;
    RECT 229.7 25.245 229.91 25.315 ;
    RECT 366.28 24.525 366.49 24.595 ;
    RECT 366.28 24.885 366.49 24.955 ;
    RECT 366.28 25.245 366.49 25.315 ;
    RECT 365.82 24.525 366.03 24.595 ;
    RECT 365.82 24.885 366.03 24.955 ;
    RECT 365.82 25.245 366.03 25.315 ;
    RECT 226.84 24.525 227.05 24.595 ;
    RECT 226.84 24.885 227.05 24.955 ;
    RECT 226.84 25.245 227.05 25.315 ;
    RECT 226.38 24.525 226.59 24.595 ;
    RECT 226.38 24.885 226.59 24.955 ;
    RECT 226.38 25.245 226.59 25.315 ;
    RECT 362.96 24.525 363.17 24.595 ;
    RECT 362.96 24.885 363.17 24.955 ;
    RECT 362.96 25.245 363.17 25.315 ;
    RECT 362.5 24.525 362.71 24.595 ;
    RECT 362.5 24.885 362.71 24.955 ;
    RECT 362.5 25.245 362.71 25.315 ;
    RECT 223.52 24.525 223.73 24.595 ;
    RECT 223.52 24.885 223.73 24.955 ;
    RECT 223.52 25.245 223.73 25.315 ;
    RECT 223.06 24.525 223.27 24.595 ;
    RECT 223.06 24.885 223.27 24.955 ;
    RECT 223.06 25.245 223.27 25.315 ;
    RECT 359.64 24.525 359.85 24.595 ;
    RECT 359.64 24.885 359.85 24.955 ;
    RECT 359.64 25.245 359.85 25.315 ;
    RECT 359.18 24.525 359.39 24.595 ;
    RECT 359.18 24.885 359.39 24.955 ;
    RECT 359.18 25.245 359.39 25.315 ;
    RECT 220.2 24.525 220.41 24.595 ;
    RECT 220.2 24.885 220.41 24.955 ;
    RECT 220.2 25.245 220.41 25.315 ;
    RECT 219.74 24.525 219.95 24.595 ;
    RECT 219.74 24.885 219.95 24.955 ;
    RECT 219.74 25.245 219.95 25.315 ;
    RECT 356.32 24.525 356.53 24.595 ;
    RECT 356.32 24.885 356.53 24.955 ;
    RECT 356.32 25.245 356.53 25.315 ;
    RECT 355.86 24.525 356.07 24.595 ;
    RECT 355.86 24.885 356.07 24.955 ;
    RECT 355.86 25.245 356.07 25.315 ;
    RECT 353.0 24.525 353.21 24.595 ;
    RECT 353.0 24.885 353.21 24.955 ;
    RECT 353.0 25.245 353.21 25.315 ;
    RECT 352.54 24.525 352.75 24.595 ;
    RECT 352.54 24.885 352.75 24.955 ;
    RECT 352.54 25.245 352.75 25.315 ;
    RECT 216.88 24.525 217.09 24.595 ;
    RECT 216.88 24.885 217.09 24.955 ;
    RECT 216.88 25.245 217.09 25.315 ;
    RECT 216.42 24.525 216.63 24.595 ;
    RECT 216.42 24.885 216.63 24.955 ;
    RECT 216.42 25.245 216.63 25.315 ;
    RECT 349.68 24.525 349.89 24.595 ;
    RECT 349.68 24.885 349.89 24.955 ;
    RECT 349.68 25.245 349.89 25.315 ;
    RECT 349.22 24.525 349.43 24.595 ;
    RECT 349.22 24.885 349.43 24.955 ;
    RECT 349.22 25.245 349.43 25.315 ;
    RECT 213.56 24.525 213.77 24.595 ;
    RECT 213.56 24.885 213.77 24.955 ;
    RECT 213.56 25.245 213.77 25.315 ;
    RECT 213.1 24.525 213.31 24.595 ;
    RECT 213.1 24.885 213.31 24.955 ;
    RECT 213.1 25.245 213.31 25.315 ;
    RECT 346.36 24.525 346.57 24.595 ;
    RECT 346.36 24.885 346.57 24.955 ;
    RECT 346.36 25.245 346.57 25.315 ;
    RECT 345.9 24.525 346.11 24.595 ;
    RECT 345.9 24.885 346.11 24.955 ;
    RECT 345.9 25.245 346.11 25.315 ;
    RECT 210.24 24.525 210.45 24.595 ;
    RECT 210.24 24.885 210.45 24.955 ;
    RECT 210.24 25.245 210.45 25.315 ;
    RECT 209.78 24.525 209.99 24.595 ;
    RECT 209.78 24.885 209.99 24.955 ;
    RECT 209.78 25.245 209.99 25.315 ;
    RECT 343.04 24.525 343.25 24.595 ;
    RECT 343.04 24.885 343.25 24.955 ;
    RECT 343.04 25.245 343.25 25.315 ;
    RECT 342.58 24.525 342.79 24.595 ;
    RECT 342.58 24.885 342.79 24.955 ;
    RECT 342.58 25.245 342.79 25.315 ;
    RECT 206.92 24.525 207.13 24.595 ;
    RECT 206.92 24.885 207.13 24.955 ;
    RECT 206.92 25.245 207.13 25.315 ;
    RECT 206.46 24.525 206.67 24.595 ;
    RECT 206.46 24.885 206.67 24.955 ;
    RECT 206.46 25.245 206.67 25.315 ;
    RECT 339.72 24.525 339.93 24.595 ;
    RECT 339.72 24.885 339.93 24.955 ;
    RECT 339.72 25.245 339.93 25.315 ;
    RECT 339.26 24.525 339.47 24.595 ;
    RECT 339.26 24.885 339.47 24.955 ;
    RECT 339.26 25.245 339.47 25.315 ;
    RECT 203.6 24.525 203.81 24.595 ;
    RECT 203.6 24.885 203.81 24.955 ;
    RECT 203.6 25.245 203.81 25.315 ;
    RECT 203.14 24.525 203.35 24.595 ;
    RECT 203.14 24.885 203.35 24.955 ;
    RECT 203.14 25.245 203.35 25.315 ;
    RECT 336.4 24.525 336.61 24.595 ;
    RECT 336.4 24.885 336.61 24.955 ;
    RECT 336.4 25.245 336.61 25.315 ;
    RECT 335.94 24.525 336.15 24.595 ;
    RECT 335.94 24.885 336.15 24.955 ;
    RECT 335.94 25.245 336.15 25.315 ;
    RECT 266.68 24.525 266.89 24.595 ;
    RECT 266.68 24.885 266.89 24.955 ;
    RECT 266.68 25.245 266.89 25.315 ;
    RECT 266.22 24.525 266.43 24.595 ;
    RECT 266.22 24.885 266.43 24.955 ;
    RECT 266.22 25.245 266.43 25.315 ;
    RECT 263.36 24.525 263.57 24.595 ;
    RECT 263.36 24.885 263.57 24.955 ;
    RECT 263.36 25.245 263.57 25.315 ;
    RECT 262.9 24.525 263.11 24.595 ;
    RECT 262.9 24.885 263.11 24.955 ;
    RECT 262.9 25.245 263.11 25.315 ;
    RECT 260.04 24.525 260.25 24.595 ;
    RECT 260.04 24.885 260.25 24.955 ;
    RECT 260.04 25.245 260.25 25.315 ;
    RECT 259.58 24.525 259.79 24.595 ;
    RECT 259.58 24.885 259.79 24.955 ;
    RECT 259.58 25.245 259.79 25.315 ;
    RECT 256.72 24.525 256.93 24.595 ;
    RECT 256.72 24.885 256.93 24.955 ;
    RECT 256.72 25.245 256.93 25.315 ;
    RECT 256.26 24.525 256.47 24.595 ;
    RECT 256.26 24.885 256.47 24.955 ;
    RECT 256.26 25.245 256.47 25.315 ;
    RECT 253.4 24.525 253.61 24.595 ;
    RECT 253.4 24.885 253.61 24.955 ;
    RECT 253.4 25.245 253.61 25.315 ;
    RECT 252.94 24.525 253.15 24.595 ;
    RECT 252.94 24.885 253.15 24.955 ;
    RECT 252.94 25.245 253.15 25.315 ;
    RECT 250.08 24.525 250.29 24.595 ;
    RECT 250.08 24.885 250.29 24.955 ;
    RECT 250.08 25.245 250.29 25.315 ;
    RECT 249.62 24.525 249.83 24.595 ;
    RECT 249.62 24.885 249.83 24.955 ;
    RECT 249.62 25.245 249.83 25.315 ;
    RECT 246.76 24.525 246.97 24.595 ;
    RECT 246.76 24.885 246.97 24.955 ;
    RECT 246.76 25.245 246.97 25.315 ;
    RECT 246.3 24.525 246.51 24.595 ;
    RECT 246.3 24.885 246.51 24.955 ;
    RECT 246.3 25.245 246.51 25.315 ;
    RECT 243.44 24.525 243.65 24.595 ;
    RECT 243.44 24.885 243.65 24.955 ;
    RECT 243.44 25.245 243.65 25.315 ;
    RECT 242.98 24.525 243.19 24.595 ;
    RECT 242.98 24.885 243.19 24.955 ;
    RECT 242.98 25.245 243.19 25.315 ;
    RECT 240.12 24.525 240.33 24.595 ;
    RECT 240.12 24.885 240.33 24.955 ;
    RECT 240.12 25.245 240.33 25.315 ;
    RECT 239.66 24.525 239.87 24.595 ;
    RECT 239.66 24.885 239.87 24.955 ;
    RECT 239.66 25.245 239.87 25.315 ;
    RECT 236.8 24.525 237.01 24.595 ;
    RECT 236.8 24.885 237.01 24.955 ;
    RECT 236.8 25.245 237.01 25.315 ;
    RECT 236.34 24.525 236.55 24.595 ;
    RECT 236.34 24.885 236.55 24.955 ;
    RECT 236.34 25.245 236.55 25.315 ;
    RECT 374.15 24.885 374.22 24.955 ;
    RECT 333.08 24.525 333.29 24.595 ;
    RECT 333.08 24.885 333.29 24.955 ;
    RECT 333.08 25.245 333.29 25.315 ;
    RECT 332.62 24.525 332.83 24.595 ;
    RECT 332.62 24.885 332.83 24.955 ;
    RECT 332.62 25.245 332.83 25.315 ;
    RECT 329.76 24.525 329.97 24.595 ;
    RECT 329.76 24.885 329.97 24.955 ;
    RECT 329.76 25.245 329.97 25.315 ;
    RECT 329.3 24.525 329.51 24.595 ;
    RECT 329.3 24.885 329.51 24.955 ;
    RECT 329.3 25.245 329.51 25.315 ;
    RECT 326.44 24.525 326.65 24.595 ;
    RECT 326.44 24.885 326.65 24.955 ;
    RECT 326.44 25.245 326.65 25.315 ;
    RECT 325.98 24.525 326.19 24.595 ;
    RECT 325.98 24.885 326.19 24.955 ;
    RECT 325.98 25.245 326.19 25.315 ;
    RECT 323.12 24.525 323.33 24.595 ;
    RECT 323.12 24.885 323.33 24.955 ;
    RECT 323.12 25.245 323.33 25.315 ;
    RECT 322.66 24.525 322.87 24.595 ;
    RECT 322.66 24.885 322.87 24.955 ;
    RECT 322.66 25.245 322.87 25.315 ;
    RECT 319.8 24.525 320.01 24.595 ;
    RECT 319.8 24.885 320.01 24.955 ;
    RECT 319.8 25.245 320.01 25.315 ;
    RECT 319.34 24.525 319.55 24.595 ;
    RECT 319.34 24.885 319.55 24.955 ;
    RECT 319.34 25.245 319.55 25.315 ;
    RECT 316.48 24.525 316.69 24.595 ;
    RECT 316.48 24.885 316.69 24.955 ;
    RECT 316.48 25.245 316.69 25.315 ;
    RECT 316.02 24.525 316.23 24.595 ;
    RECT 316.02 24.885 316.23 24.955 ;
    RECT 316.02 25.245 316.23 25.315 ;
    RECT 313.16 24.525 313.37 24.595 ;
    RECT 313.16 24.885 313.37 24.955 ;
    RECT 313.16 25.245 313.37 25.315 ;
    RECT 312.7 24.525 312.91 24.595 ;
    RECT 312.7 24.885 312.91 24.955 ;
    RECT 312.7 25.245 312.91 25.315 ;
    RECT 309.84 24.525 310.05 24.595 ;
    RECT 309.84 24.885 310.05 24.955 ;
    RECT 309.84 25.245 310.05 25.315 ;
    RECT 309.38 24.525 309.59 24.595 ;
    RECT 309.38 24.885 309.59 24.955 ;
    RECT 309.38 25.245 309.59 25.315 ;
    RECT 306.52 24.525 306.73 24.595 ;
    RECT 306.52 24.885 306.73 24.955 ;
    RECT 306.52 25.245 306.73 25.315 ;
    RECT 306.06 24.525 306.27 24.595 ;
    RECT 306.06 24.885 306.27 24.955 ;
    RECT 306.06 25.245 306.27 25.315 ;
    RECT 303.2 23.805 303.41 23.875 ;
    RECT 303.2 24.165 303.41 24.235 ;
    RECT 303.2 24.525 303.41 24.595 ;
    RECT 302.74 23.805 302.95 23.875 ;
    RECT 302.74 24.165 302.95 24.235 ;
    RECT 302.74 24.525 302.95 24.595 ;
    RECT 372.92 23.805 373.13 23.875 ;
    RECT 372.92 24.165 373.13 24.235 ;
    RECT 372.92 24.525 373.13 24.595 ;
    RECT 372.46 23.805 372.67 23.875 ;
    RECT 372.46 24.165 372.67 24.235 ;
    RECT 372.46 24.525 372.67 24.595 ;
    RECT 369.6 23.805 369.81 23.875 ;
    RECT 369.6 24.165 369.81 24.235 ;
    RECT 369.6 24.525 369.81 24.595 ;
    RECT 369.14 23.805 369.35 23.875 ;
    RECT 369.14 24.165 369.35 24.235 ;
    RECT 369.14 24.525 369.35 24.595 ;
    RECT 200.605 24.165 200.675 24.235 ;
    RECT 299.88 23.805 300.09 23.875 ;
    RECT 299.88 24.165 300.09 24.235 ;
    RECT 299.88 24.525 300.09 24.595 ;
    RECT 299.42 23.805 299.63 23.875 ;
    RECT 299.42 24.165 299.63 24.235 ;
    RECT 299.42 24.525 299.63 24.595 ;
    RECT 296.56 23.805 296.77 23.875 ;
    RECT 296.56 24.165 296.77 24.235 ;
    RECT 296.56 24.525 296.77 24.595 ;
    RECT 296.1 23.805 296.31 23.875 ;
    RECT 296.1 24.165 296.31 24.235 ;
    RECT 296.1 24.525 296.31 24.595 ;
    RECT 293.24 23.805 293.45 23.875 ;
    RECT 293.24 24.165 293.45 24.235 ;
    RECT 293.24 24.525 293.45 24.595 ;
    RECT 292.78 23.805 292.99 23.875 ;
    RECT 292.78 24.165 292.99 24.235 ;
    RECT 292.78 24.525 292.99 24.595 ;
    RECT 289.92 23.805 290.13 23.875 ;
    RECT 289.92 24.165 290.13 24.235 ;
    RECT 289.92 24.525 290.13 24.595 ;
    RECT 289.46 23.805 289.67 23.875 ;
    RECT 289.46 24.165 289.67 24.235 ;
    RECT 289.46 24.525 289.67 24.595 ;
    RECT 286.6 23.805 286.81 23.875 ;
    RECT 286.6 24.165 286.81 24.235 ;
    RECT 286.6 24.525 286.81 24.595 ;
    RECT 286.14 23.805 286.35 23.875 ;
    RECT 286.14 24.165 286.35 24.235 ;
    RECT 286.14 24.525 286.35 24.595 ;
    RECT 283.28 23.805 283.49 23.875 ;
    RECT 283.28 24.165 283.49 24.235 ;
    RECT 283.28 24.525 283.49 24.595 ;
    RECT 282.82 23.805 283.03 23.875 ;
    RECT 282.82 24.165 283.03 24.235 ;
    RECT 282.82 24.525 283.03 24.595 ;
    RECT 279.96 23.805 280.17 23.875 ;
    RECT 279.96 24.165 280.17 24.235 ;
    RECT 279.96 24.525 280.17 24.595 ;
    RECT 279.5 23.805 279.71 23.875 ;
    RECT 279.5 24.165 279.71 24.235 ;
    RECT 279.5 24.525 279.71 24.595 ;
    RECT 276.64 23.805 276.85 23.875 ;
    RECT 276.64 24.165 276.85 24.235 ;
    RECT 276.64 24.525 276.85 24.595 ;
    RECT 276.18 23.805 276.39 23.875 ;
    RECT 276.18 24.165 276.39 24.235 ;
    RECT 276.18 24.525 276.39 24.595 ;
    RECT 273.32 23.805 273.53 23.875 ;
    RECT 273.32 24.165 273.53 24.235 ;
    RECT 273.32 24.525 273.53 24.595 ;
    RECT 272.86 23.805 273.07 23.875 ;
    RECT 272.86 24.165 273.07 24.235 ;
    RECT 272.86 24.525 273.07 24.595 ;
    RECT 270.0 23.805 270.21 23.875 ;
    RECT 270.0 24.165 270.21 24.235 ;
    RECT 270.0 24.525 270.21 24.595 ;
    RECT 269.54 23.805 269.75 23.875 ;
    RECT 269.54 24.165 269.75 24.235 ;
    RECT 269.54 24.525 269.75 24.595 ;
    RECT 233.48 23.805 233.69 23.875 ;
    RECT 233.48 24.165 233.69 24.235 ;
    RECT 233.48 24.525 233.69 24.595 ;
    RECT 233.02 23.805 233.23 23.875 ;
    RECT 233.02 24.165 233.23 24.235 ;
    RECT 233.02 24.525 233.23 24.595 ;
    RECT 230.16 23.805 230.37 23.875 ;
    RECT 230.16 24.165 230.37 24.235 ;
    RECT 230.16 24.525 230.37 24.595 ;
    RECT 229.7 23.805 229.91 23.875 ;
    RECT 229.7 24.165 229.91 24.235 ;
    RECT 229.7 24.525 229.91 24.595 ;
    RECT 366.28 23.805 366.49 23.875 ;
    RECT 366.28 24.165 366.49 24.235 ;
    RECT 366.28 24.525 366.49 24.595 ;
    RECT 365.82 23.805 366.03 23.875 ;
    RECT 365.82 24.165 366.03 24.235 ;
    RECT 365.82 24.525 366.03 24.595 ;
    RECT 226.84 23.805 227.05 23.875 ;
    RECT 226.84 24.165 227.05 24.235 ;
    RECT 226.84 24.525 227.05 24.595 ;
    RECT 226.38 23.805 226.59 23.875 ;
    RECT 226.38 24.165 226.59 24.235 ;
    RECT 226.38 24.525 226.59 24.595 ;
    RECT 362.96 23.805 363.17 23.875 ;
    RECT 362.96 24.165 363.17 24.235 ;
    RECT 362.96 24.525 363.17 24.595 ;
    RECT 362.5 23.805 362.71 23.875 ;
    RECT 362.5 24.165 362.71 24.235 ;
    RECT 362.5 24.525 362.71 24.595 ;
    RECT 223.52 23.805 223.73 23.875 ;
    RECT 223.52 24.165 223.73 24.235 ;
    RECT 223.52 24.525 223.73 24.595 ;
    RECT 223.06 23.805 223.27 23.875 ;
    RECT 223.06 24.165 223.27 24.235 ;
    RECT 223.06 24.525 223.27 24.595 ;
    RECT 359.64 23.805 359.85 23.875 ;
    RECT 359.64 24.165 359.85 24.235 ;
    RECT 359.64 24.525 359.85 24.595 ;
    RECT 359.18 23.805 359.39 23.875 ;
    RECT 359.18 24.165 359.39 24.235 ;
    RECT 359.18 24.525 359.39 24.595 ;
    RECT 220.2 23.805 220.41 23.875 ;
    RECT 220.2 24.165 220.41 24.235 ;
    RECT 220.2 24.525 220.41 24.595 ;
    RECT 219.74 23.805 219.95 23.875 ;
    RECT 219.74 24.165 219.95 24.235 ;
    RECT 219.74 24.525 219.95 24.595 ;
    RECT 356.32 23.805 356.53 23.875 ;
    RECT 356.32 24.165 356.53 24.235 ;
    RECT 356.32 24.525 356.53 24.595 ;
    RECT 355.86 23.805 356.07 23.875 ;
    RECT 355.86 24.165 356.07 24.235 ;
    RECT 355.86 24.525 356.07 24.595 ;
    RECT 353.0 23.805 353.21 23.875 ;
    RECT 353.0 24.165 353.21 24.235 ;
    RECT 353.0 24.525 353.21 24.595 ;
    RECT 352.54 23.805 352.75 23.875 ;
    RECT 352.54 24.165 352.75 24.235 ;
    RECT 352.54 24.525 352.75 24.595 ;
    RECT 216.88 23.805 217.09 23.875 ;
    RECT 216.88 24.165 217.09 24.235 ;
    RECT 216.88 24.525 217.09 24.595 ;
    RECT 216.42 23.805 216.63 23.875 ;
    RECT 216.42 24.165 216.63 24.235 ;
    RECT 216.42 24.525 216.63 24.595 ;
    RECT 349.68 23.805 349.89 23.875 ;
    RECT 349.68 24.165 349.89 24.235 ;
    RECT 349.68 24.525 349.89 24.595 ;
    RECT 349.22 23.805 349.43 23.875 ;
    RECT 349.22 24.165 349.43 24.235 ;
    RECT 349.22 24.525 349.43 24.595 ;
    RECT 213.56 23.805 213.77 23.875 ;
    RECT 213.56 24.165 213.77 24.235 ;
    RECT 213.56 24.525 213.77 24.595 ;
    RECT 213.1 23.805 213.31 23.875 ;
    RECT 213.1 24.165 213.31 24.235 ;
    RECT 213.1 24.525 213.31 24.595 ;
    RECT 346.36 23.805 346.57 23.875 ;
    RECT 346.36 24.165 346.57 24.235 ;
    RECT 346.36 24.525 346.57 24.595 ;
    RECT 345.9 23.805 346.11 23.875 ;
    RECT 345.9 24.165 346.11 24.235 ;
    RECT 345.9 24.525 346.11 24.595 ;
    RECT 210.24 23.805 210.45 23.875 ;
    RECT 210.24 24.165 210.45 24.235 ;
    RECT 210.24 24.525 210.45 24.595 ;
    RECT 209.78 23.805 209.99 23.875 ;
    RECT 209.78 24.165 209.99 24.235 ;
    RECT 209.78 24.525 209.99 24.595 ;
    RECT 343.04 23.805 343.25 23.875 ;
    RECT 343.04 24.165 343.25 24.235 ;
    RECT 343.04 24.525 343.25 24.595 ;
    RECT 342.58 23.805 342.79 23.875 ;
    RECT 342.58 24.165 342.79 24.235 ;
    RECT 342.58 24.525 342.79 24.595 ;
    RECT 206.92 23.805 207.13 23.875 ;
    RECT 206.92 24.165 207.13 24.235 ;
    RECT 206.92 24.525 207.13 24.595 ;
    RECT 206.46 23.805 206.67 23.875 ;
    RECT 206.46 24.165 206.67 24.235 ;
    RECT 206.46 24.525 206.67 24.595 ;
    RECT 339.72 23.805 339.93 23.875 ;
    RECT 339.72 24.165 339.93 24.235 ;
    RECT 339.72 24.525 339.93 24.595 ;
    RECT 339.26 23.805 339.47 23.875 ;
    RECT 339.26 24.165 339.47 24.235 ;
    RECT 339.26 24.525 339.47 24.595 ;
    RECT 203.6 23.805 203.81 23.875 ;
    RECT 203.6 24.165 203.81 24.235 ;
    RECT 203.6 24.525 203.81 24.595 ;
    RECT 203.14 23.805 203.35 23.875 ;
    RECT 203.14 24.165 203.35 24.235 ;
    RECT 203.14 24.525 203.35 24.595 ;
    RECT 336.4 23.805 336.61 23.875 ;
    RECT 336.4 24.165 336.61 24.235 ;
    RECT 336.4 24.525 336.61 24.595 ;
    RECT 335.94 23.805 336.15 23.875 ;
    RECT 335.94 24.165 336.15 24.235 ;
    RECT 335.94 24.525 336.15 24.595 ;
    RECT 266.68 23.805 266.89 23.875 ;
    RECT 266.68 24.165 266.89 24.235 ;
    RECT 266.68 24.525 266.89 24.595 ;
    RECT 266.22 23.805 266.43 23.875 ;
    RECT 266.22 24.165 266.43 24.235 ;
    RECT 266.22 24.525 266.43 24.595 ;
    RECT 263.36 23.805 263.57 23.875 ;
    RECT 263.36 24.165 263.57 24.235 ;
    RECT 263.36 24.525 263.57 24.595 ;
    RECT 262.9 23.805 263.11 23.875 ;
    RECT 262.9 24.165 263.11 24.235 ;
    RECT 262.9 24.525 263.11 24.595 ;
    RECT 260.04 23.805 260.25 23.875 ;
    RECT 260.04 24.165 260.25 24.235 ;
    RECT 260.04 24.525 260.25 24.595 ;
    RECT 259.58 23.805 259.79 23.875 ;
    RECT 259.58 24.165 259.79 24.235 ;
    RECT 259.58 24.525 259.79 24.595 ;
    RECT 256.72 23.805 256.93 23.875 ;
    RECT 256.72 24.165 256.93 24.235 ;
    RECT 256.72 24.525 256.93 24.595 ;
    RECT 256.26 23.805 256.47 23.875 ;
    RECT 256.26 24.165 256.47 24.235 ;
    RECT 256.26 24.525 256.47 24.595 ;
    RECT 253.4 23.805 253.61 23.875 ;
    RECT 253.4 24.165 253.61 24.235 ;
    RECT 253.4 24.525 253.61 24.595 ;
    RECT 252.94 23.805 253.15 23.875 ;
    RECT 252.94 24.165 253.15 24.235 ;
    RECT 252.94 24.525 253.15 24.595 ;
    RECT 250.08 23.805 250.29 23.875 ;
    RECT 250.08 24.165 250.29 24.235 ;
    RECT 250.08 24.525 250.29 24.595 ;
    RECT 249.62 23.805 249.83 23.875 ;
    RECT 249.62 24.165 249.83 24.235 ;
    RECT 249.62 24.525 249.83 24.595 ;
    RECT 246.76 23.805 246.97 23.875 ;
    RECT 246.76 24.165 246.97 24.235 ;
    RECT 246.76 24.525 246.97 24.595 ;
    RECT 246.3 23.805 246.51 23.875 ;
    RECT 246.3 24.165 246.51 24.235 ;
    RECT 246.3 24.525 246.51 24.595 ;
    RECT 243.44 23.805 243.65 23.875 ;
    RECT 243.44 24.165 243.65 24.235 ;
    RECT 243.44 24.525 243.65 24.595 ;
    RECT 242.98 23.805 243.19 23.875 ;
    RECT 242.98 24.165 243.19 24.235 ;
    RECT 242.98 24.525 243.19 24.595 ;
    RECT 240.12 23.805 240.33 23.875 ;
    RECT 240.12 24.165 240.33 24.235 ;
    RECT 240.12 24.525 240.33 24.595 ;
    RECT 239.66 23.805 239.87 23.875 ;
    RECT 239.66 24.165 239.87 24.235 ;
    RECT 239.66 24.525 239.87 24.595 ;
    RECT 236.8 23.805 237.01 23.875 ;
    RECT 236.8 24.165 237.01 24.235 ;
    RECT 236.8 24.525 237.01 24.595 ;
    RECT 236.34 23.805 236.55 23.875 ;
    RECT 236.34 24.165 236.55 24.235 ;
    RECT 236.34 24.525 236.55 24.595 ;
    RECT 374.15 24.165 374.22 24.235 ;
    RECT 333.08 23.805 333.29 23.875 ;
    RECT 333.08 24.165 333.29 24.235 ;
    RECT 333.08 24.525 333.29 24.595 ;
    RECT 332.62 23.805 332.83 23.875 ;
    RECT 332.62 24.165 332.83 24.235 ;
    RECT 332.62 24.525 332.83 24.595 ;
    RECT 329.76 23.805 329.97 23.875 ;
    RECT 329.76 24.165 329.97 24.235 ;
    RECT 329.76 24.525 329.97 24.595 ;
    RECT 329.3 23.805 329.51 23.875 ;
    RECT 329.3 24.165 329.51 24.235 ;
    RECT 329.3 24.525 329.51 24.595 ;
    RECT 326.44 23.805 326.65 23.875 ;
    RECT 326.44 24.165 326.65 24.235 ;
    RECT 326.44 24.525 326.65 24.595 ;
    RECT 325.98 23.805 326.19 23.875 ;
    RECT 325.98 24.165 326.19 24.235 ;
    RECT 325.98 24.525 326.19 24.595 ;
    RECT 323.12 23.805 323.33 23.875 ;
    RECT 323.12 24.165 323.33 24.235 ;
    RECT 323.12 24.525 323.33 24.595 ;
    RECT 322.66 23.805 322.87 23.875 ;
    RECT 322.66 24.165 322.87 24.235 ;
    RECT 322.66 24.525 322.87 24.595 ;
    RECT 319.8 23.805 320.01 23.875 ;
    RECT 319.8 24.165 320.01 24.235 ;
    RECT 319.8 24.525 320.01 24.595 ;
    RECT 319.34 23.805 319.55 23.875 ;
    RECT 319.34 24.165 319.55 24.235 ;
    RECT 319.34 24.525 319.55 24.595 ;
    RECT 316.48 23.805 316.69 23.875 ;
    RECT 316.48 24.165 316.69 24.235 ;
    RECT 316.48 24.525 316.69 24.595 ;
    RECT 316.02 23.805 316.23 23.875 ;
    RECT 316.02 24.165 316.23 24.235 ;
    RECT 316.02 24.525 316.23 24.595 ;
    RECT 313.16 23.805 313.37 23.875 ;
    RECT 313.16 24.165 313.37 24.235 ;
    RECT 313.16 24.525 313.37 24.595 ;
    RECT 312.7 23.805 312.91 23.875 ;
    RECT 312.7 24.165 312.91 24.235 ;
    RECT 312.7 24.525 312.91 24.595 ;
    RECT 309.84 23.805 310.05 23.875 ;
    RECT 309.84 24.165 310.05 24.235 ;
    RECT 309.84 24.525 310.05 24.595 ;
    RECT 309.38 23.805 309.59 23.875 ;
    RECT 309.38 24.165 309.59 24.235 ;
    RECT 309.38 24.525 309.59 24.595 ;
    RECT 306.52 23.805 306.73 23.875 ;
    RECT 306.52 24.165 306.73 24.235 ;
    RECT 306.52 24.525 306.73 24.595 ;
    RECT 306.06 23.805 306.27 23.875 ;
    RECT 306.06 24.165 306.27 24.235 ;
    RECT 306.06 24.525 306.27 24.595 ;
    RECT 303.2 23.085 303.41 23.155 ;
    RECT 303.2 23.445 303.41 23.515 ;
    RECT 303.2 23.805 303.41 23.875 ;
    RECT 302.74 23.085 302.95 23.155 ;
    RECT 302.74 23.445 302.95 23.515 ;
    RECT 302.74 23.805 302.95 23.875 ;
    RECT 372.92 23.085 373.13 23.155 ;
    RECT 372.92 23.445 373.13 23.515 ;
    RECT 372.92 23.805 373.13 23.875 ;
    RECT 372.46 23.085 372.67 23.155 ;
    RECT 372.46 23.445 372.67 23.515 ;
    RECT 372.46 23.805 372.67 23.875 ;
    RECT 369.6 23.085 369.81 23.155 ;
    RECT 369.6 23.445 369.81 23.515 ;
    RECT 369.6 23.805 369.81 23.875 ;
    RECT 369.14 23.085 369.35 23.155 ;
    RECT 369.14 23.445 369.35 23.515 ;
    RECT 369.14 23.805 369.35 23.875 ;
    RECT 200.605 23.445 200.675 23.515 ;
    RECT 299.88 23.085 300.09 23.155 ;
    RECT 299.88 23.445 300.09 23.515 ;
    RECT 299.88 23.805 300.09 23.875 ;
    RECT 299.42 23.085 299.63 23.155 ;
    RECT 299.42 23.445 299.63 23.515 ;
    RECT 299.42 23.805 299.63 23.875 ;
    RECT 296.56 23.085 296.77 23.155 ;
    RECT 296.56 23.445 296.77 23.515 ;
    RECT 296.56 23.805 296.77 23.875 ;
    RECT 296.1 23.085 296.31 23.155 ;
    RECT 296.1 23.445 296.31 23.515 ;
    RECT 296.1 23.805 296.31 23.875 ;
    RECT 293.24 23.085 293.45 23.155 ;
    RECT 293.24 23.445 293.45 23.515 ;
    RECT 293.24 23.805 293.45 23.875 ;
    RECT 292.78 23.085 292.99 23.155 ;
    RECT 292.78 23.445 292.99 23.515 ;
    RECT 292.78 23.805 292.99 23.875 ;
    RECT 289.92 23.085 290.13 23.155 ;
    RECT 289.92 23.445 290.13 23.515 ;
    RECT 289.92 23.805 290.13 23.875 ;
    RECT 289.46 23.085 289.67 23.155 ;
    RECT 289.46 23.445 289.67 23.515 ;
    RECT 289.46 23.805 289.67 23.875 ;
    RECT 286.6 23.085 286.81 23.155 ;
    RECT 286.6 23.445 286.81 23.515 ;
    RECT 286.6 23.805 286.81 23.875 ;
    RECT 286.14 23.085 286.35 23.155 ;
    RECT 286.14 23.445 286.35 23.515 ;
    RECT 286.14 23.805 286.35 23.875 ;
    RECT 283.28 23.085 283.49 23.155 ;
    RECT 283.28 23.445 283.49 23.515 ;
    RECT 283.28 23.805 283.49 23.875 ;
    RECT 282.82 23.085 283.03 23.155 ;
    RECT 282.82 23.445 283.03 23.515 ;
    RECT 282.82 23.805 283.03 23.875 ;
    RECT 279.96 23.085 280.17 23.155 ;
    RECT 279.96 23.445 280.17 23.515 ;
    RECT 279.96 23.805 280.17 23.875 ;
    RECT 279.5 23.085 279.71 23.155 ;
    RECT 279.5 23.445 279.71 23.515 ;
    RECT 279.5 23.805 279.71 23.875 ;
    RECT 276.64 23.085 276.85 23.155 ;
    RECT 276.64 23.445 276.85 23.515 ;
    RECT 276.64 23.805 276.85 23.875 ;
    RECT 276.18 23.085 276.39 23.155 ;
    RECT 276.18 23.445 276.39 23.515 ;
    RECT 276.18 23.805 276.39 23.875 ;
    RECT 273.32 23.085 273.53 23.155 ;
    RECT 273.32 23.445 273.53 23.515 ;
    RECT 273.32 23.805 273.53 23.875 ;
    RECT 272.86 23.085 273.07 23.155 ;
    RECT 272.86 23.445 273.07 23.515 ;
    RECT 272.86 23.805 273.07 23.875 ;
    RECT 270.0 23.085 270.21 23.155 ;
    RECT 270.0 23.445 270.21 23.515 ;
    RECT 270.0 23.805 270.21 23.875 ;
    RECT 269.54 23.085 269.75 23.155 ;
    RECT 269.54 23.445 269.75 23.515 ;
    RECT 269.54 23.805 269.75 23.875 ;
    RECT 233.48 23.085 233.69 23.155 ;
    RECT 233.48 23.445 233.69 23.515 ;
    RECT 233.48 23.805 233.69 23.875 ;
    RECT 233.02 23.085 233.23 23.155 ;
    RECT 233.02 23.445 233.23 23.515 ;
    RECT 233.02 23.805 233.23 23.875 ;
    RECT 230.16 23.085 230.37 23.155 ;
    RECT 230.16 23.445 230.37 23.515 ;
    RECT 230.16 23.805 230.37 23.875 ;
    RECT 229.7 23.085 229.91 23.155 ;
    RECT 229.7 23.445 229.91 23.515 ;
    RECT 229.7 23.805 229.91 23.875 ;
    RECT 366.28 23.085 366.49 23.155 ;
    RECT 366.28 23.445 366.49 23.515 ;
    RECT 366.28 23.805 366.49 23.875 ;
    RECT 365.82 23.085 366.03 23.155 ;
    RECT 365.82 23.445 366.03 23.515 ;
    RECT 365.82 23.805 366.03 23.875 ;
    RECT 226.84 23.085 227.05 23.155 ;
    RECT 226.84 23.445 227.05 23.515 ;
    RECT 226.84 23.805 227.05 23.875 ;
    RECT 226.38 23.085 226.59 23.155 ;
    RECT 226.38 23.445 226.59 23.515 ;
    RECT 226.38 23.805 226.59 23.875 ;
    RECT 362.96 23.085 363.17 23.155 ;
    RECT 362.96 23.445 363.17 23.515 ;
    RECT 362.96 23.805 363.17 23.875 ;
    RECT 362.5 23.085 362.71 23.155 ;
    RECT 362.5 23.445 362.71 23.515 ;
    RECT 362.5 23.805 362.71 23.875 ;
    RECT 223.52 23.085 223.73 23.155 ;
    RECT 223.52 23.445 223.73 23.515 ;
    RECT 223.52 23.805 223.73 23.875 ;
    RECT 223.06 23.085 223.27 23.155 ;
    RECT 223.06 23.445 223.27 23.515 ;
    RECT 223.06 23.805 223.27 23.875 ;
    RECT 359.64 23.085 359.85 23.155 ;
    RECT 359.64 23.445 359.85 23.515 ;
    RECT 359.64 23.805 359.85 23.875 ;
    RECT 359.18 23.085 359.39 23.155 ;
    RECT 359.18 23.445 359.39 23.515 ;
    RECT 359.18 23.805 359.39 23.875 ;
    RECT 220.2 23.085 220.41 23.155 ;
    RECT 220.2 23.445 220.41 23.515 ;
    RECT 220.2 23.805 220.41 23.875 ;
    RECT 219.74 23.085 219.95 23.155 ;
    RECT 219.74 23.445 219.95 23.515 ;
    RECT 219.74 23.805 219.95 23.875 ;
    RECT 356.32 23.085 356.53 23.155 ;
    RECT 356.32 23.445 356.53 23.515 ;
    RECT 356.32 23.805 356.53 23.875 ;
    RECT 355.86 23.085 356.07 23.155 ;
    RECT 355.86 23.445 356.07 23.515 ;
    RECT 355.86 23.805 356.07 23.875 ;
    RECT 353.0 23.085 353.21 23.155 ;
    RECT 353.0 23.445 353.21 23.515 ;
    RECT 353.0 23.805 353.21 23.875 ;
    RECT 352.54 23.085 352.75 23.155 ;
    RECT 352.54 23.445 352.75 23.515 ;
    RECT 352.54 23.805 352.75 23.875 ;
    RECT 216.88 23.085 217.09 23.155 ;
    RECT 216.88 23.445 217.09 23.515 ;
    RECT 216.88 23.805 217.09 23.875 ;
    RECT 216.42 23.085 216.63 23.155 ;
    RECT 216.42 23.445 216.63 23.515 ;
    RECT 216.42 23.805 216.63 23.875 ;
    RECT 349.68 23.085 349.89 23.155 ;
    RECT 349.68 23.445 349.89 23.515 ;
    RECT 349.68 23.805 349.89 23.875 ;
    RECT 349.22 23.085 349.43 23.155 ;
    RECT 349.22 23.445 349.43 23.515 ;
    RECT 349.22 23.805 349.43 23.875 ;
    RECT 213.56 23.085 213.77 23.155 ;
    RECT 213.56 23.445 213.77 23.515 ;
    RECT 213.56 23.805 213.77 23.875 ;
    RECT 213.1 23.085 213.31 23.155 ;
    RECT 213.1 23.445 213.31 23.515 ;
    RECT 213.1 23.805 213.31 23.875 ;
    RECT 346.36 23.085 346.57 23.155 ;
    RECT 346.36 23.445 346.57 23.515 ;
    RECT 346.36 23.805 346.57 23.875 ;
    RECT 345.9 23.085 346.11 23.155 ;
    RECT 345.9 23.445 346.11 23.515 ;
    RECT 345.9 23.805 346.11 23.875 ;
    RECT 210.24 23.085 210.45 23.155 ;
    RECT 210.24 23.445 210.45 23.515 ;
    RECT 210.24 23.805 210.45 23.875 ;
    RECT 209.78 23.085 209.99 23.155 ;
    RECT 209.78 23.445 209.99 23.515 ;
    RECT 209.78 23.805 209.99 23.875 ;
    RECT 343.04 23.085 343.25 23.155 ;
    RECT 343.04 23.445 343.25 23.515 ;
    RECT 343.04 23.805 343.25 23.875 ;
    RECT 342.58 23.085 342.79 23.155 ;
    RECT 342.58 23.445 342.79 23.515 ;
    RECT 342.58 23.805 342.79 23.875 ;
    RECT 206.92 23.085 207.13 23.155 ;
    RECT 206.92 23.445 207.13 23.515 ;
    RECT 206.92 23.805 207.13 23.875 ;
    RECT 206.46 23.085 206.67 23.155 ;
    RECT 206.46 23.445 206.67 23.515 ;
    RECT 206.46 23.805 206.67 23.875 ;
    RECT 339.72 23.085 339.93 23.155 ;
    RECT 339.72 23.445 339.93 23.515 ;
    RECT 339.72 23.805 339.93 23.875 ;
    RECT 339.26 23.085 339.47 23.155 ;
    RECT 339.26 23.445 339.47 23.515 ;
    RECT 339.26 23.805 339.47 23.875 ;
    RECT 203.6 23.085 203.81 23.155 ;
    RECT 203.6 23.445 203.81 23.515 ;
    RECT 203.6 23.805 203.81 23.875 ;
    RECT 203.14 23.085 203.35 23.155 ;
    RECT 203.14 23.445 203.35 23.515 ;
    RECT 203.14 23.805 203.35 23.875 ;
    RECT 336.4 23.085 336.61 23.155 ;
    RECT 336.4 23.445 336.61 23.515 ;
    RECT 336.4 23.805 336.61 23.875 ;
    RECT 335.94 23.085 336.15 23.155 ;
    RECT 335.94 23.445 336.15 23.515 ;
    RECT 335.94 23.805 336.15 23.875 ;
    RECT 266.68 23.085 266.89 23.155 ;
    RECT 266.68 23.445 266.89 23.515 ;
    RECT 266.68 23.805 266.89 23.875 ;
    RECT 266.22 23.085 266.43 23.155 ;
    RECT 266.22 23.445 266.43 23.515 ;
    RECT 266.22 23.805 266.43 23.875 ;
    RECT 263.36 23.085 263.57 23.155 ;
    RECT 263.36 23.445 263.57 23.515 ;
    RECT 263.36 23.805 263.57 23.875 ;
    RECT 262.9 23.085 263.11 23.155 ;
    RECT 262.9 23.445 263.11 23.515 ;
    RECT 262.9 23.805 263.11 23.875 ;
    RECT 260.04 23.085 260.25 23.155 ;
    RECT 260.04 23.445 260.25 23.515 ;
    RECT 260.04 23.805 260.25 23.875 ;
    RECT 259.58 23.085 259.79 23.155 ;
    RECT 259.58 23.445 259.79 23.515 ;
    RECT 259.58 23.805 259.79 23.875 ;
    RECT 256.72 23.085 256.93 23.155 ;
    RECT 256.72 23.445 256.93 23.515 ;
    RECT 256.72 23.805 256.93 23.875 ;
    RECT 256.26 23.085 256.47 23.155 ;
    RECT 256.26 23.445 256.47 23.515 ;
    RECT 256.26 23.805 256.47 23.875 ;
    RECT 253.4 23.085 253.61 23.155 ;
    RECT 253.4 23.445 253.61 23.515 ;
    RECT 253.4 23.805 253.61 23.875 ;
    RECT 252.94 23.085 253.15 23.155 ;
    RECT 252.94 23.445 253.15 23.515 ;
    RECT 252.94 23.805 253.15 23.875 ;
    RECT 250.08 23.085 250.29 23.155 ;
    RECT 250.08 23.445 250.29 23.515 ;
    RECT 250.08 23.805 250.29 23.875 ;
    RECT 249.62 23.085 249.83 23.155 ;
    RECT 249.62 23.445 249.83 23.515 ;
    RECT 249.62 23.805 249.83 23.875 ;
    RECT 246.76 23.085 246.97 23.155 ;
    RECT 246.76 23.445 246.97 23.515 ;
    RECT 246.76 23.805 246.97 23.875 ;
    RECT 246.3 23.085 246.51 23.155 ;
    RECT 246.3 23.445 246.51 23.515 ;
    RECT 246.3 23.805 246.51 23.875 ;
    RECT 243.44 23.085 243.65 23.155 ;
    RECT 243.44 23.445 243.65 23.515 ;
    RECT 243.44 23.805 243.65 23.875 ;
    RECT 242.98 23.085 243.19 23.155 ;
    RECT 242.98 23.445 243.19 23.515 ;
    RECT 242.98 23.805 243.19 23.875 ;
    RECT 240.12 23.085 240.33 23.155 ;
    RECT 240.12 23.445 240.33 23.515 ;
    RECT 240.12 23.805 240.33 23.875 ;
    RECT 239.66 23.085 239.87 23.155 ;
    RECT 239.66 23.445 239.87 23.515 ;
    RECT 239.66 23.805 239.87 23.875 ;
    RECT 236.8 23.085 237.01 23.155 ;
    RECT 236.8 23.445 237.01 23.515 ;
    RECT 236.8 23.805 237.01 23.875 ;
    RECT 236.34 23.085 236.55 23.155 ;
    RECT 236.34 23.445 236.55 23.515 ;
    RECT 236.34 23.805 236.55 23.875 ;
    RECT 374.15 23.445 374.22 23.515 ;
    RECT 333.08 23.085 333.29 23.155 ;
    RECT 333.08 23.445 333.29 23.515 ;
    RECT 333.08 23.805 333.29 23.875 ;
    RECT 332.62 23.085 332.83 23.155 ;
    RECT 332.62 23.445 332.83 23.515 ;
    RECT 332.62 23.805 332.83 23.875 ;
    RECT 329.76 23.085 329.97 23.155 ;
    RECT 329.76 23.445 329.97 23.515 ;
    RECT 329.76 23.805 329.97 23.875 ;
    RECT 329.3 23.085 329.51 23.155 ;
    RECT 329.3 23.445 329.51 23.515 ;
    RECT 329.3 23.805 329.51 23.875 ;
    RECT 326.44 23.085 326.65 23.155 ;
    RECT 326.44 23.445 326.65 23.515 ;
    RECT 326.44 23.805 326.65 23.875 ;
    RECT 325.98 23.085 326.19 23.155 ;
    RECT 325.98 23.445 326.19 23.515 ;
    RECT 325.98 23.805 326.19 23.875 ;
    RECT 323.12 23.085 323.33 23.155 ;
    RECT 323.12 23.445 323.33 23.515 ;
    RECT 323.12 23.805 323.33 23.875 ;
    RECT 322.66 23.085 322.87 23.155 ;
    RECT 322.66 23.445 322.87 23.515 ;
    RECT 322.66 23.805 322.87 23.875 ;
    RECT 319.8 23.085 320.01 23.155 ;
    RECT 319.8 23.445 320.01 23.515 ;
    RECT 319.8 23.805 320.01 23.875 ;
    RECT 319.34 23.085 319.55 23.155 ;
    RECT 319.34 23.445 319.55 23.515 ;
    RECT 319.34 23.805 319.55 23.875 ;
    RECT 316.48 23.085 316.69 23.155 ;
    RECT 316.48 23.445 316.69 23.515 ;
    RECT 316.48 23.805 316.69 23.875 ;
    RECT 316.02 23.085 316.23 23.155 ;
    RECT 316.02 23.445 316.23 23.515 ;
    RECT 316.02 23.805 316.23 23.875 ;
    RECT 313.16 23.085 313.37 23.155 ;
    RECT 313.16 23.445 313.37 23.515 ;
    RECT 313.16 23.805 313.37 23.875 ;
    RECT 312.7 23.085 312.91 23.155 ;
    RECT 312.7 23.445 312.91 23.515 ;
    RECT 312.7 23.805 312.91 23.875 ;
    RECT 309.84 23.085 310.05 23.155 ;
    RECT 309.84 23.445 310.05 23.515 ;
    RECT 309.84 23.805 310.05 23.875 ;
    RECT 309.38 23.085 309.59 23.155 ;
    RECT 309.38 23.445 309.59 23.515 ;
    RECT 309.38 23.805 309.59 23.875 ;
    RECT 306.52 23.085 306.73 23.155 ;
    RECT 306.52 23.445 306.73 23.515 ;
    RECT 306.52 23.805 306.73 23.875 ;
    RECT 306.06 23.085 306.27 23.155 ;
    RECT 306.06 23.445 306.27 23.515 ;
    RECT 306.06 23.805 306.27 23.875 ;
    RECT 303.2 22.365 303.41 22.435 ;
    RECT 303.2 22.725 303.41 22.795 ;
    RECT 303.2 23.085 303.41 23.155 ;
    RECT 302.74 22.365 302.95 22.435 ;
    RECT 302.74 22.725 302.95 22.795 ;
    RECT 302.74 23.085 302.95 23.155 ;
    RECT 372.92 22.365 373.13 22.435 ;
    RECT 372.92 22.725 373.13 22.795 ;
    RECT 372.92 23.085 373.13 23.155 ;
    RECT 372.46 22.365 372.67 22.435 ;
    RECT 372.46 22.725 372.67 22.795 ;
    RECT 372.46 23.085 372.67 23.155 ;
    RECT 369.6 22.365 369.81 22.435 ;
    RECT 369.6 22.725 369.81 22.795 ;
    RECT 369.6 23.085 369.81 23.155 ;
    RECT 369.14 22.365 369.35 22.435 ;
    RECT 369.14 22.725 369.35 22.795 ;
    RECT 369.14 23.085 369.35 23.155 ;
    RECT 200.605 22.725 200.675 22.795 ;
    RECT 299.88 22.365 300.09 22.435 ;
    RECT 299.88 22.725 300.09 22.795 ;
    RECT 299.88 23.085 300.09 23.155 ;
    RECT 299.42 22.365 299.63 22.435 ;
    RECT 299.42 22.725 299.63 22.795 ;
    RECT 299.42 23.085 299.63 23.155 ;
    RECT 296.56 22.365 296.77 22.435 ;
    RECT 296.56 22.725 296.77 22.795 ;
    RECT 296.56 23.085 296.77 23.155 ;
    RECT 296.1 22.365 296.31 22.435 ;
    RECT 296.1 22.725 296.31 22.795 ;
    RECT 296.1 23.085 296.31 23.155 ;
    RECT 293.24 22.365 293.45 22.435 ;
    RECT 293.24 22.725 293.45 22.795 ;
    RECT 293.24 23.085 293.45 23.155 ;
    RECT 292.78 22.365 292.99 22.435 ;
    RECT 292.78 22.725 292.99 22.795 ;
    RECT 292.78 23.085 292.99 23.155 ;
    RECT 289.92 22.365 290.13 22.435 ;
    RECT 289.92 22.725 290.13 22.795 ;
    RECT 289.92 23.085 290.13 23.155 ;
    RECT 289.46 22.365 289.67 22.435 ;
    RECT 289.46 22.725 289.67 22.795 ;
    RECT 289.46 23.085 289.67 23.155 ;
    RECT 286.6 22.365 286.81 22.435 ;
    RECT 286.6 22.725 286.81 22.795 ;
    RECT 286.6 23.085 286.81 23.155 ;
    RECT 286.14 22.365 286.35 22.435 ;
    RECT 286.14 22.725 286.35 22.795 ;
    RECT 286.14 23.085 286.35 23.155 ;
    RECT 283.28 22.365 283.49 22.435 ;
    RECT 283.28 22.725 283.49 22.795 ;
    RECT 283.28 23.085 283.49 23.155 ;
    RECT 282.82 22.365 283.03 22.435 ;
    RECT 282.82 22.725 283.03 22.795 ;
    RECT 282.82 23.085 283.03 23.155 ;
    RECT 279.96 22.365 280.17 22.435 ;
    RECT 279.96 22.725 280.17 22.795 ;
    RECT 279.96 23.085 280.17 23.155 ;
    RECT 279.5 22.365 279.71 22.435 ;
    RECT 279.5 22.725 279.71 22.795 ;
    RECT 279.5 23.085 279.71 23.155 ;
    RECT 276.64 22.365 276.85 22.435 ;
    RECT 276.64 22.725 276.85 22.795 ;
    RECT 276.64 23.085 276.85 23.155 ;
    RECT 276.18 22.365 276.39 22.435 ;
    RECT 276.18 22.725 276.39 22.795 ;
    RECT 276.18 23.085 276.39 23.155 ;
    RECT 273.32 22.365 273.53 22.435 ;
    RECT 273.32 22.725 273.53 22.795 ;
    RECT 273.32 23.085 273.53 23.155 ;
    RECT 272.86 22.365 273.07 22.435 ;
    RECT 272.86 22.725 273.07 22.795 ;
    RECT 272.86 23.085 273.07 23.155 ;
    RECT 270.0 22.365 270.21 22.435 ;
    RECT 270.0 22.725 270.21 22.795 ;
    RECT 270.0 23.085 270.21 23.155 ;
    RECT 269.54 22.365 269.75 22.435 ;
    RECT 269.54 22.725 269.75 22.795 ;
    RECT 269.54 23.085 269.75 23.155 ;
    RECT 233.48 22.365 233.69 22.435 ;
    RECT 233.48 22.725 233.69 22.795 ;
    RECT 233.48 23.085 233.69 23.155 ;
    RECT 233.02 22.365 233.23 22.435 ;
    RECT 233.02 22.725 233.23 22.795 ;
    RECT 233.02 23.085 233.23 23.155 ;
    RECT 230.16 22.365 230.37 22.435 ;
    RECT 230.16 22.725 230.37 22.795 ;
    RECT 230.16 23.085 230.37 23.155 ;
    RECT 229.7 22.365 229.91 22.435 ;
    RECT 229.7 22.725 229.91 22.795 ;
    RECT 229.7 23.085 229.91 23.155 ;
    RECT 366.28 22.365 366.49 22.435 ;
    RECT 366.28 22.725 366.49 22.795 ;
    RECT 366.28 23.085 366.49 23.155 ;
    RECT 365.82 22.365 366.03 22.435 ;
    RECT 365.82 22.725 366.03 22.795 ;
    RECT 365.82 23.085 366.03 23.155 ;
    RECT 226.84 22.365 227.05 22.435 ;
    RECT 226.84 22.725 227.05 22.795 ;
    RECT 226.84 23.085 227.05 23.155 ;
    RECT 226.38 22.365 226.59 22.435 ;
    RECT 226.38 22.725 226.59 22.795 ;
    RECT 226.38 23.085 226.59 23.155 ;
    RECT 362.96 22.365 363.17 22.435 ;
    RECT 362.96 22.725 363.17 22.795 ;
    RECT 362.96 23.085 363.17 23.155 ;
    RECT 362.5 22.365 362.71 22.435 ;
    RECT 362.5 22.725 362.71 22.795 ;
    RECT 362.5 23.085 362.71 23.155 ;
    RECT 223.52 22.365 223.73 22.435 ;
    RECT 223.52 22.725 223.73 22.795 ;
    RECT 223.52 23.085 223.73 23.155 ;
    RECT 223.06 22.365 223.27 22.435 ;
    RECT 223.06 22.725 223.27 22.795 ;
    RECT 223.06 23.085 223.27 23.155 ;
    RECT 359.64 22.365 359.85 22.435 ;
    RECT 359.64 22.725 359.85 22.795 ;
    RECT 359.64 23.085 359.85 23.155 ;
    RECT 359.18 22.365 359.39 22.435 ;
    RECT 359.18 22.725 359.39 22.795 ;
    RECT 359.18 23.085 359.39 23.155 ;
    RECT 220.2 22.365 220.41 22.435 ;
    RECT 220.2 22.725 220.41 22.795 ;
    RECT 220.2 23.085 220.41 23.155 ;
    RECT 219.74 22.365 219.95 22.435 ;
    RECT 219.74 22.725 219.95 22.795 ;
    RECT 219.74 23.085 219.95 23.155 ;
    RECT 356.32 22.365 356.53 22.435 ;
    RECT 356.32 22.725 356.53 22.795 ;
    RECT 356.32 23.085 356.53 23.155 ;
    RECT 355.86 22.365 356.07 22.435 ;
    RECT 355.86 22.725 356.07 22.795 ;
    RECT 355.86 23.085 356.07 23.155 ;
    RECT 353.0 22.365 353.21 22.435 ;
    RECT 353.0 22.725 353.21 22.795 ;
    RECT 353.0 23.085 353.21 23.155 ;
    RECT 352.54 22.365 352.75 22.435 ;
    RECT 352.54 22.725 352.75 22.795 ;
    RECT 352.54 23.085 352.75 23.155 ;
    RECT 216.88 22.365 217.09 22.435 ;
    RECT 216.88 22.725 217.09 22.795 ;
    RECT 216.88 23.085 217.09 23.155 ;
    RECT 216.42 22.365 216.63 22.435 ;
    RECT 216.42 22.725 216.63 22.795 ;
    RECT 216.42 23.085 216.63 23.155 ;
    RECT 349.68 22.365 349.89 22.435 ;
    RECT 349.68 22.725 349.89 22.795 ;
    RECT 349.68 23.085 349.89 23.155 ;
    RECT 349.22 22.365 349.43 22.435 ;
    RECT 349.22 22.725 349.43 22.795 ;
    RECT 349.22 23.085 349.43 23.155 ;
    RECT 213.56 22.365 213.77 22.435 ;
    RECT 213.56 22.725 213.77 22.795 ;
    RECT 213.56 23.085 213.77 23.155 ;
    RECT 213.1 22.365 213.31 22.435 ;
    RECT 213.1 22.725 213.31 22.795 ;
    RECT 213.1 23.085 213.31 23.155 ;
    RECT 346.36 22.365 346.57 22.435 ;
    RECT 346.36 22.725 346.57 22.795 ;
    RECT 346.36 23.085 346.57 23.155 ;
    RECT 345.9 22.365 346.11 22.435 ;
    RECT 345.9 22.725 346.11 22.795 ;
    RECT 345.9 23.085 346.11 23.155 ;
    RECT 210.24 22.365 210.45 22.435 ;
    RECT 210.24 22.725 210.45 22.795 ;
    RECT 210.24 23.085 210.45 23.155 ;
    RECT 209.78 22.365 209.99 22.435 ;
    RECT 209.78 22.725 209.99 22.795 ;
    RECT 209.78 23.085 209.99 23.155 ;
    RECT 343.04 22.365 343.25 22.435 ;
    RECT 343.04 22.725 343.25 22.795 ;
    RECT 343.04 23.085 343.25 23.155 ;
    RECT 342.58 22.365 342.79 22.435 ;
    RECT 342.58 22.725 342.79 22.795 ;
    RECT 342.58 23.085 342.79 23.155 ;
    RECT 206.92 22.365 207.13 22.435 ;
    RECT 206.92 22.725 207.13 22.795 ;
    RECT 206.92 23.085 207.13 23.155 ;
    RECT 206.46 22.365 206.67 22.435 ;
    RECT 206.46 22.725 206.67 22.795 ;
    RECT 206.46 23.085 206.67 23.155 ;
    RECT 339.72 22.365 339.93 22.435 ;
    RECT 339.72 22.725 339.93 22.795 ;
    RECT 339.72 23.085 339.93 23.155 ;
    RECT 339.26 22.365 339.47 22.435 ;
    RECT 339.26 22.725 339.47 22.795 ;
    RECT 339.26 23.085 339.47 23.155 ;
    RECT 203.6 22.365 203.81 22.435 ;
    RECT 203.6 22.725 203.81 22.795 ;
    RECT 203.6 23.085 203.81 23.155 ;
    RECT 203.14 22.365 203.35 22.435 ;
    RECT 203.14 22.725 203.35 22.795 ;
    RECT 203.14 23.085 203.35 23.155 ;
    RECT 336.4 22.365 336.61 22.435 ;
    RECT 336.4 22.725 336.61 22.795 ;
    RECT 336.4 23.085 336.61 23.155 ;
    RECT 335.94 22.365 336.15 22.435 ;
    RECT 335.94 22.725 336.15 22.795 ;
    RECT 335.94 23.085 336.15 23.155 ;
    RECT 266.68 22.365 266.89 22.435 ;
    RECT 266.68 22.725 266.89 22.795 ;
    RECT 266.68 23.085 266.89 23.155 ;
    RECT 266.22 22.365 266.43 22.435 ;
    RECT 266.22 22.725 266.43 22.795 ;
    RECT 266.22 23.085 266.43 23.155 ;
    RECT 263.36 22.365 263.57 22.435 ;
    RECT 263.36 22.725 263.57 22.795 ;
    RECT 263.36 23.085 263.57 23.155 ;
    RECT 262.9 22.365 263.11 22.435 ;
    RECT 262.9 22.725 263.11 22.795 ;
    RECT 262.9 23.085 263.11 23.155 ;
    RECT 260.04 22.365 260.25 22.435 ;
    RECT 260.04 22.725 260.25 22.795 ;
    RECT 260.04 23.085 260.25 23.155 ;
    RECT 259.58 22.365 259.79 22.435 ;
    RECT 259.58 22.725 259.79 22.795 ;
    RECT 259.58 23.085 259.79 23.155 ;
    RECT 256.72 22.365 256.93 22.435 ;
    RECT 256.72 22.725 256.93 22.795 ;
    RECT 256.72 23.085 256.93 23.155 ;
    RECT 256.26 22.365 256.47 22.435 ;
    RECT 256.26 22.725 256.47 22.795 ;
    RECT 256.26 23.085 256.47 23.155 ;
    RECT 253.4 22.365 253.61 22.435 ;
    RECT 253.4 22.725 253.61 22.795 ;
    RECT 253.4 23.085 253.61 23.155 ;
    RECT 252.94 22.365 253.15 22.435 ;
    RECT 252.94 22.725 253.15 22.795 ;
    RECT 252.94 23.085 253.15 23.155 ;
    RECT 250.08 22.365 250.29 22.435 ;
    RECT 250.08 22.725 250.29 22.795 ;
    RECT 250.08 23.085 250.29 23.155 ;
    RECT 249.62 22.365 249.83 22.435 ;
    RECT 249.62 22.725 249.83 22.795 ;
    RECT 249.62 23.085 249.83 23.155 ;
    RECT 246.76 22.365 246.97 22.435 ;
    RECT 246.76 22.725 246.97 22.795 ;
    RECT 246.76 23.085 246.97 23.155 ;
    RECT 246.3 22.365 246.51 22.435 ;
    RECT 246.3 22.725 246.51 22.795 ;
    RECT 246.3 23.085 246.51 23.155 ;
    RECT 243.44 22.365 243.65 22.435 ;
    RECT 243.44 22.725 243.65 22.795 ;
    RECT 243.44 23.085 243.65 23.155 ;
    RECT 242.98 22.365 243.19 22.435 ;
    RECT 242.98 22.725 243.19 22.795 ;
    RECT 242.98 23.085 243.19 23.155 ;
    RECT 240.12 22.365 240.33 22.435 ;
    RECT 240.12 22.725 240.33 22.795 ;
    RECT 240.12 23.085 240.33 23.155 ;
    RECT 239.66 22.365 239.87 22.435 ;
    RECT 239.66 22.725 239.87 22.795 ;
    RECT 239.66 23.085 239.87 23.155 ;
    RECT 236.8 22.365 237.01 22.435 ;
    RECT 236.8 22.725 237.01 22.795 ;
    RECT 236.8 23.085 237.01 23.155 ;
    RECT 236.34 22.365 236.55 22.435 ;
    RECT 236.34 22.725 236.55 22.795 ;
    RECT 236.34 23.085 236.55 23.155 ;
    RECT 374.15 22.725 374.22 22.795 ;
    RECT 333.08 22.365 333.29 22.435 ;
    RECT 333.08 22.725 333.29 22.795 ;
    RECT 333.08 23.085 333.29 23.155 ;
    RECT 332.62 22.365 332.83 22.435 ;
    RECT 332.62 22.725 332.83 22.795 ;
    RECT 332.62 23.085 332.83 23.155 ;
    RECT 329.76 22.365 329.97 22.435 ;
    RECT 329.76 22.725 329.97 22.795 ;
    RECT 329.76 23.085 329.97 23.155 ;
    RECT 329.3 22.365 329.51 22.435 ;
    RECT 329.3 22.725 329.51 22.795 ;
    RECT 329.3 23.085 329.51 23.155 ;
    RECT 326.44 22.365 326.65 22.435 ;
    RECT 326.44 22.725 326.65 22.795 ;
    RECT 326.44 23.085 326.65 23.155 ;
    RECT 325.98 22.365 326.19 22.435 ;
    RECT 325.98 22.725 326.19 22.795 ;
    RECT 325.98 23.085 326.19 23.155 ;
    RECT 323.12 22.365 323.33 22.435 ;
    RECT 323.12 22.725 323.33 22.795 ;
    RECT 323.12 23.085 323.33 23.155 ;
    RECT 322.66 22.365 322.87 22.435 ;
    RECT 322.66 22.725 322.87 22.795 ;
    RECT 322.66 23.085 322.87 23.155 ;
    RECT 319.8 22.365 320.01 22.435 ;
    RECT 319.8 22.725 320.01 22.795 ;
    RECT 319.8 23.085 320.01 23.155 ;
    RECT 319.34 22.365 319.55 22.435 ;
    RECT 319.34 22.725 319.55 22.795 ;
    RECT 319.34 23.085 319.55 23.155 ;
    RECT 316.48 22.365 316.69 22.435 ;
    RECT 316.48 22.725 316.69 22.795 ;
    RECT 316.48 23.085 316.69 23.155 ;
    RECT 316.02 22.365 316.23 22.435 ;
    RECT 316.02 22.725 316.23 22.795 ;
    RECT 316.02 23.085 316.23 23.155 ;
    RECT 313.16 22.365 313.37 22.435 ;
    RECT 313.16 22.725 313.37 22.795 ;
    RECT 313.16 23.085 313.37 23.155 ;
    RECT 312.7 22.365 312.91 22.435 ;
    RECT 312.7 22.725 312.91 22.795 ;
    RECT 312.7 23.085 312.91 23.155 ;
    RECT 309.84 22.365 310.05 22.435 ;
    RECT 309.84 22.725 310.05 22.795 ;
    RECT 309.84 23.085 310.05 23.155 ;
    RECT 309.38 22.365 309.59 22.435 ;
    RECT 309.38 22.725 309.59 22.795 ;
    RECT 309.38 23.085 309.59 23.155 ;
    RECT 306.52 22.365 306.73 22.435 ;
    RECT 306.52 22.725 306.73 22.795 ;
    RECT 306.52 23.085 306.73 23.155 ;
    RECT 306.06 22.365 306.27 22.435 ;
    RECT 306.06 22.725 306.27 22.795 ;
    RECT 306.06 23.085 306.27 23.155 ;
    RECT 303.2 21.645 303.41 21.715 ;
    RECT 303.2 22.005 303.41 22.075 ;
    RECT 303.2 22.365 303.41 22.435 ;
    RECT 302.74 21.645 302.95 21.715 ;
    RECT 302.74 22.005 302.95 22.075 ;
    RECT 302.74 22.365 302.95 22.435 ;
    RECT 372.92 21.645 373.13 21.715 ;
    RECT 372.92 22.005 373.13 22.075 ;
    RECT 372.92 22.365 373.13 22.435 ;
    RECT 372.46 21.645 372.67 21.715 ;
    RECT 372.46 22.005 372.67 22.075 ;
    RECT 372.46 22.365 372.67 22.435 ;
    RECT 369.6 21.645 369.81 21.715 ;
    RECT 369.6 22.005 369.81 22.075 ;
    RECT 369.6 22.365 369.81 22.435 ;
    RECT 369.14 21.645 369.35 21.715 ;
    RECT 369.14 22.005 369.35 22.075 ;
    RECT 369.14 22.365 369.35 22.435 ;
    RECT 200.605 22.005 200.675 22.075 ;
    RECT 299.88 21.645 300.09 21.715 ;
    RECT 299.88 22.005 300.09 22.075 ;
    RECT 299.88 22.365 300.09 22.435 ;
    RECT 299.42 21.645 299.63 21.715 ;
    RECT 299.42 22.005 299.63 22.075 ;
    RECT 299.42 22.365 299.63 22.435 ;
    RECT 296.56 21.645 296.77 21.715 ;
    RECT 296.56 22.005 296.77 22.075 ;
    RECT 296.56 22.365 296.77 22.435 ;
    RECT 296.1 21.645 296.31 21.715 ;
    RECT 296.1 22.005 296.31 22.075 ;
    RECT 296.1 22.365 296.31 22.435 ;
    RECT 293.24 21.645 293.45 21.715 ;
    RECT 293.24 22.005 293.45 22.075 ;
    RECT 293.24 22.365 293.45 22.435 ;
    RECT 292.78 21.645 292.99 21.715 ;
    RECT 292.78 22.005 292.99 22.075 ;
    RECT 292.78 22.365 292.99 22.435 ;
    RECT 289.92 21.645 290.13 21.715 ;
    RECT 289.92 22.005 290.13 22.075 ;
    RECT 289.92 22.365 290.13 22.435 ;
    RECT 289.46 21.645 289.67 21.715 ;
    RECT 289.46 22.005 289.67 22.075 ;
    RECT 289.46 22.365 289.67 22.435 ;
    RECT 286.6 21.645 286.81 21.715 ;
    RECT 286.6 22.005 286.81 22.075 ;
    RECT 286.6 22.365 286.81 22.435 ;
    RECT 286.14 21.645 286.35 21.715 ;
    RECT 286.14 22.005 286.35 22.075 ;
    RECT 286.14 22.365 286.35 22.435 ;
    RECT 283.28 21.645 283.49 21.715 ;
    RECT 283.28 22.005 283.49 22.075 ;
    RECT 283.28 22.365 283.49 22.435 ;
    RECT 282.82 21.645 283.03 21.715 ;
    RECT 282.82 22.005 283.03 22.075 ;
    RECT 282.82 22.365 283.03 22.435 ;
    RECT 279.96 21.645 280.17 21.715 ;
    RECT 279.96 22.005 280.17 22.075 ;
    RECT 279.96 22.365 280.17 22.435 ;
    RECT 279.5 21.645 279.71 21.715 ;
    RECT 279.5 22.005 279.71 22.075 ;
    RECT 279.5 22.365 279.71 22.435 ;
    RECT 276.64 21.645 276.85 21.715 ;
    RECT 276.64 22.005 276.85 22.075 ;
    RECT 276.64 22.365 276.85 22.435 ;
    RECT 276.18 21.645 276.39 21.715 ;
    RECT 276.18 22.005 276.39 22.075 ;
    RECT 276.18 22.365 276.39 22.435 ;
    RECT 273.32 21.645 273.53 21.715 ;
    RECT 273.32 22.005 273.53 22.075 ;
    RECT 273.32 22.365 273.53 22.435 ;
    RECT 272.86 21.645 273.07 21.715 ;
    RECT 272.86 22.005 273.07 22.075 ;
    RECT 272.86 22.365 273.07 22.435 ;
    RECT 270.0 21.645 270.21 21.715 ;
    RECT 270.0 22.005 270.21 22.075 ;
    RECT 270.0 22.365 270.21 22.435 ;
    RECT 269.54 21.645 269.75 21.715 ;
    RECT 269.54 22.005 269.75 22.075 ;
    RECT 269.54 22.365 269.75 22.435 ;
    RECT 233.48 21.645 233.69 21.715 ;
    RECT 233.48 22.005 233.69 22.075 ;
    RECT 233.48 22.365 233.69 22.435 ;
    RECT 233.02 21.645 233.23 21.715 ;
    RECT 233.02 22.005 233.23 22.075 ;
    RECT 233.02 22.365 233.23 22.435 ;
    RECT 230.16 21.645 230.37 21.715 ;
    RECT 230.16 22.005 230.37 22.075 ;
    RECT 230.16 22.365 230.37 22.435 ;
    RECT 229.7 21.645 229.91 21.715 ;
    RECT 229.7 22.005 229.91 22.075 ;
    RECT 229.7 22.365 229.91 22.435 ;
    RECT 366.28 21.645 366.49 21.715 ;
    RECT 366.28 22.005 366.49 22.075 ;
    RECT 366.28 22.365 366.49 22.435 ;
    RECT 365.82 21.645 366.03 21.715 ;
    RECT 365.82 22.005 366.03 22.075 ;
    RECT 365.82 22.365 366.03 22.435 ;
    RECT 226.84 21.645 227.05 21.715 ;
    RECT 226.84 22.005 227.05 22.075 ;
    RECT 226.84 22.365 227.05 22.435 ;
    RECT 226.38 21.645 226.59 21.715 ;
    RECT 226.38 22.005 226.59 22.075 ;
    RECT 226.38 22.365 226.59 22.435 ;
    RECT 362.96 21.645 363.17 21.715 ;
    RECT 362.96 22.005 363.17 22.075 ;
    RECT 362.96 22.365 363.17 22.435 ;
    RECT 362.5 21.645 362.71 21.715 ;
    RECT 362.5 22.005 362.71 22.075 ;
    RECT 362.5 22.365 362.71 22.435 ;
    RECT 223.52 21.645 223.73 21.715 ;
    RECT 223.52 22.005 223.73 22.075 ;
    RECT 223.52 22.365 223.73 22.435 ;
    RECT 223.06 21.645 223.27 21.715 ;
    RECT 223.06 22.005 223.27 22.075 ;
    RECT 223.06 22.365 223.27 22.435 ;
    RECT 359.64 21.645 359.85 21.715 ;
    RECT 359.64 22.005 359.85 22.075 ;
    RECT 359.64 22.365 359.85 22.435 ;
    RECT 359.18 21.645 359.39 21.715 ;
    RECT 359.18 22.005 359.39 22.075 ;
    RECT 359.18 22.365 359.39 22.435 ;
    RECT 220.2 21.645 220.41 21.715 ;
    RECT 220.2 22.005 220.41 22.075 ;
    RECT 220.2 22.365 220.41 22.435 ;
    RECT 219.74 21.645 219.95 21.715 ;
    RECT 219.74 22.005 219.95 22.075 ;
    RECT 219.74 22.365 219.95 22.435 ;
    RECT 356.32 21.645 356.53 21.715 ;
    RECT 356.32 22.005 356.53 22.075 ;
    RECT 356.32 22.365 356.53 22.435 ;
    RECT 355.86 21.645 356.07 21.715 ;
    RECT 355.86 22.005 356.07 22.075 ;
    RECT 355.86 22.365 356.07 22.435 ;
    RECT 353.0 21.645 353.21 21.715 ;
    RECT 353.0 22.005 353.21 22.075 ;
    RECT 353.0 22.365 353.21 22.435 ;
    RECT 352.54 21.645 352.75 21.715 ;
    RECT 352.54 22.005 352.75 22.075 ;
    RECT 352.54 22.365 352.75 22.435 ;
    RECT 216.88 21.645 217.09 21.715 ;
    RECT 216.88 22.005 217.09 22.075 ;
    RECT 216.88 22.365 217.09 22.435 ;
    RECT 216.42 21.645 216.63 21.715 ;
    RECT 216.42 22.005 216.63 22.075 ;
    RECT 216.42 22.365 216.63 22.435 ;
    RECT 349.68 21.645 349.89 21.715 ;
    RECT 349.68 22.005 349.89 22.075 ;
    RECT 349.68 22.365 349.89 22.435 ;
    RECT 349.22 21.645 349.43 21.715 ;
    RECT 349.22 22.005 349.43 22.075 ;
    RECT 349.22 22.365 349.43 22.435 ;
    RECT 213.56 21.645 213.77 21.715 ;
    RECT 213.56 22.005 213.77 22.075 ;
    RECT 213.56 22.365 213.77 22.435 ;
    RECT 213.1 21.645 213.31 21.715 ;
    RECT 213.1 22.005 213.31 22.075 ;
    RECT 213.1 22.365 213.31 22.435 ;
    RECT 346.36 21.645 346.57 21.715 ;
    RECT 346.36 22.005 346.57 22.075 ;
    RECT 346.36 22.365 346.57 22.435 ;
    RECT 345.9 21.645 346.11 21.715 ;
    RECT 345.9 22.005 346.11 22.075 ;
    RECT 345.9 22.365 346.11 22.435 ;
    RECT 210.24 21.645 210.45 21.715 ;
    RECT 210.24 22.005 210.45 22.075 ;
    RECT 210.24 22.365 210.45 22.435 ;
    RECT 209.78 21.645 209.99 21.715 ;
    RECT 209.78 22.005 209.99 22.075 ;
    RECT 209.78 22.365 209.99 22.435 ;
    RECT 343.04 21.645 343.25 21.715 ;
    RECT 343.04 22.005 343.25 22.075 ;
    RECT 343.04 22.365 343.25 22.435 ;
    RECT 342.58 21.645 342.79 21.715 ;
    RECT 342.58 22.005 342.79 22.075 ;
    RECT 342.58 22.365 342.79 22.435 ;
    RECT 206.92 21.645 207.13 21.715 ;
    RECT 206.92 22.005 207.13 22.075 ;
    RECT 206.92 22.365 207.13 22.435 ;
    RECT 206.46 21.645 206.67 21.715 ;
    RECT 206.46 22.005 206.67 22.075 ;
    RECT 206.46 22.365 206.67 22.435 ;
    RECT 339.72 21.645 339.93 21.715 ;
    RECT 339.72 22.005 339.93 22.075 ;
    RECT 339.72 22.365 339.93 22.435 ;
    RECT 339.26 21.645 339.47 21.715 ;
    RECT 339.26 22.005 339.47 22.075 ;
    RECT 339.26 22.365 339.47 22.435 ;
    RECT 203.6 21.645 203.81 21.715 ;
    RECT 203.6 22.005 203.81 22.075 ;
    RECT 203.6 22.365 203.81 22.435 ;
    RECT 203.14 21.645 203.35 21.715 ;
    RECT 203.14 22.005 203.35 22.075 ;
    RECT 203.14 22.365 203.35 22.435 ;
    RECT 336.4 21.645 336.61 21.715 ;
    RECT 336.4 22.005 336.61 22.075 ;
    RECT 336.4 22.365 336.61 22.435 ;
    RECT 335.94 21.645 336.15 21.715 ;
    RECT 335.94 22.005 336.15 22.075 ;
    RECT 335.94 22.365 336.15 22.435 ;
    RECT 266.68 21.645 266.89 21.715 ;
    RECT 266.68 22.005 266.89 22.075 ;
    RECT 266.68 22.365 266.89 22.435 ;
    RECT 266.22 21.645 266.43 21.715 ;
    RECT 266.22 22.005 266.43 22.075 ;
    RECT 266.22 22.365 266.43 22.435 ;
    RECT 263.36 21.645 263.57 21.715 ;
    RECT 263.36 22.005 263.57 22.075 ;
    RECT 263.36 22.365 263.57 22.435 ;
    RECT 262.9 21.645 263.11 21.715 ;
    RECT 262.9 22.005 263.11 22.075 ;
    RECT 262.9 22.365 263.11 22.435 ;
    RECT 260.04 21.645 260.25 21.715 ;
    RECT 260.04 22.005 260.25 22.075 ;
    RECT 260.04 22.365 260.25 22.435 ;
    RECT 259.58 21.645 259.79 21.715 ;
    RECT 259.58 22.005 259.79 22.075 ;
    RECT 259.58 22.365 259.79 22.435 ;
    RECT 256.72 21.645 256.93 21.715 ;
    RECT 256.72 22.005 256.93 22.075 ;
    RECT 256.72 22.365 256.93 22.435 ;
    RECT 256.26 21.645 256.47 21.715 ;
    RECT 256.26 22.005 256.47 22.075 ;
    RECT 256.26 22.365 256.47 22.435 ;
    RECT 253.4 21.645 253.61 21.715 ;
    RECT 253.4 22.005 253.61 22.075 ;
    RECT 253.4 22.365 253.61 22.435 ;
    RECT 252.94 21.645 253.15 21.715 ;
    RECT 252.94 22.005 253.15 22.075 ;
    RECT 252.94 22.365 253.15 22.435 ;
    RECT 250.08 21.645 250.29 21.715 ;
    RECT 250.08 22.005 250.29 22.075 ;
    RECT 250.08 22.365 250.29 22.435 ;
    RECT 249.62 21.645 249.83 21.715 ;
    RECT 249.62 22.005 249.83 22.075 ;
    RECT 249.62 22.365 249.83 22.435 ;
    RECT 246.76 21.645 246.97 21.715 ;
    RECT 246.76 22.005 246.97 22.075 ;
    RECT 246.76 22.365 246.97 22.435 ;
    RECT 246.3 21.645 246.51 21.715 ;
    RECT 246.3 22.005 246.51 22.075 ;
    RECT 246.3 22.365 246.51 22.435 ;
    RECT 243.44 21.645 243.65 21.715 ;
    RECT 243.44 22.005 243.65 22.075 ;
    RECT 243.44 22.365 243.65 22.435 ;
    RECT 242.98 21.645 243.19 21.715 ;
    RECT 242.98 22.005 243.19 22.075 ;
    RECT 242.98 22.365 243.19 22.435 ;
    RECT 240.12 21.645 240.33 21.715 ;
    RECT 240.12 22.005 240.33 22.075 ;
    RECT 240.12 22.365 240.33 22.435 ;
    RECT 239.66 21.645 239.87 21.715 ;
    RECT 239.66 22.005 239.87 22.075 ;
    RECT 239.66 22.365 239.87 22.435 ;
    RECT 236.8 21.645 237.01 21.715 ;
    RECT 236.8 22.005 237.01 22.075 ;
    RECT 236.8 22.365 237.01 22.435 ;
    RECT 236.34 21.645 236.55 21.715 ;
    RECT 236.34 22.005 236.55 22.075 ;
    RECT 236.34 22.365 236.55 22.435 ;
    RECT 374.15 22.005 374.22 22.075 ;
    RECT 333.08 21.645 333.29 21.715 ;
    RECT 333.08 22.005 333.29 22.075 ;
    RECT 333.08 22.365 333.29 22.435 ;
    RECT 332.62 21.645 332.83 21.715 ;
    RECT 332.62 22.005 332.83 22.075 ;
    RECT 332.62 22.365 332.83 22.435 ;
    RECT 329.76 21.645 329.97 21.715 ;
    RECT 329.76 22.005 329.97 22.075 ;
    RECT 329.76 22.365 329.97 22.435 ;
    RECT 329.3 21.645 329.51 21.715 ;
    RECT 329.3 22.005 329.51 22.075 ;
    RECT 329.3 22.365 329.51 22.435 ;
    RECT 326.44 21.645 326.65 21.715 ;
    RECT 326.44 22.005 326.65 22.075 ;
    RECT 326.44 22.365 326.65 22.435 ;
    RECT 325.98 21.645 326.19 21.715 ;
    RECT 325.98 22.005 326.19 22.075 ;
    RECT 325.98 22.365 326.19 22.435 ;
    RECT 323.12 21.645 323.33 21.715 ;
    RECT 323.12 22.005 323.33 22.075 ;
    RECT 323.12 22.365 323.33 22.435 ;
    RECT 322.66 21.645 322.87 21.715 ;
    RECT 322.66 22.005 322.87 22.075 ;
    RECT 322.66 22.365 322.87 22.435 ;
    RECT 319.8 21.645 320.01 21.715 ;
    RECT 319.8 22.005 320.01 22.075 ;
    RECT 319.8 22.365 320.01 22.435 ;
    RECT 319.34 21.645 319.55 21.715 ;
    RECT 319.34 22.005 319.55 22.075 ;
    RECT 319.34 22.365 319.55 22.435 ;
    RECT 316.48 21.645 316.69 21.715 ;
    RECT 316.48 22.005 316.69 22.075 ;
    RECT 316.48 22.365 316.69 22.435 ;
    RECT 316.02 21.645 316.23 21.715 ;
    RECT 316.02 22.005 316.23 22.075 ;
    RECT 316.02 22.365 316.23 22.435 ;
    RECT 313.16 21.645 313.37 21.715 ;
    RECT 313.16 22.005 313.37 22.075 ;
    RECT 313.16 22.365 313.37 22.435 ;
    RECT 312.7 21.645 312.91 21.715 ;
    RECT 312.7 22.005 312.91 22.075 ;
    RECT 312.7 22.365 312.91 22.435 ;
    RECT 309.84 21.645 310.05 21.715 ;
    RECT 309.84 22.005 310.05 22.075 ;
    RECT 309.84 22.365 310.05 22.435 ;
    RECT 309.38 21.645 309.59 21.715 ;
    RECT 309.38 22.005 309.59 22.075 ;
    RECT 309.38 22.365 309.59 22.435 ;
    RECT 306.52 21.645 306.73 21.715 ;
    RECT 306.52 22.005 306.73 22.075 ;
    RECT 306.52 22.365 306.73 22.435 ;
    RECT 306.06 21.645 306.27 21.715 ;
    RECT 306.06 22.005 306.27 22.075 ;
    RECT 306.06 22.365 306.27 22.435 ;
    RECT 303.2 20.925 303.41 20.995 ;
    RECT 303.2 21.285 303.41 21.355 ;
    RECT 303.2 21.645 303.41 21.715 ;
    RECT 302.74 20.925 302.95 20.995 ;
    RECT 302.74 21.285 302.95 21.355 ;
    RECT 302.74 21.645 302.95 21.715 ;
    RECT 372.92 20.925 373.13 20.995 ;
    RECT 372.92 21.285 373.13 21.355 ;
    RECT 372.92 21.645 373.13 21.715 ;
    RECT 372.46 20.925 372.67 20.995 ;
    RECT 372.46 21.285 372.67 21.355 ;
    RECT 372.46 21.645 372.67 21.715 ;
    RECT 369.6 20.925 369.81 20.995 ;
    RECT 369.6 21.285 369.81 21.355 ;
    RECT 369.6 21.645 369.81 21.715 ;
    RECT 369.14 20.925 369.35 20.995 ;
    RECT 369.14 21.285 369.35 21.355 ;
    RECT 369.14 21.645 369.35 21.715 ;
    RECT 200.605 21.285 200.675 21.355 ;
    RECT 299.88 20.925 300.09 20.995 ;
    RECT 299.88 21.285 300.09 21.355 ;
    RECT 299.88 21.645 300.09 21.715 ;
    RECT 299.42 20.925 299.63 20.995 ;
    RECT 299.42 21.285 299.63 21.355 ;
    RECT 299.42 21.645 299.63 21.715 ;
    RECT 296.56 20.925 296.77 20.995 ;
    RECT 296.56 21.285 296.77 21.355 ;
    RECT 296.56 21.645 296.77 21.715 ;
    RECT 296.1 20.925 296.31 20.995 ;
    RECT 296.1 21.285 296.31 21.355 ;
    RECT 296.1 21.645 296.31 21.715 ;
    RECT 293.24 20.925 293.45 20.995 ;
    RECT 293.24 21.285 293.45 21.355 ;
    RECT 293.24 21.645 293.45 21.715 ;
    RECT 292.78 20.925 292.99 20.995 ;
    RECT 292.78 21.285 292.99 21.355 ;
    RECT 292.78 21.645 292.99 21.715 ;
    RECT 289.92 20.925 290.13 20.995 ;
    RECT 289.92 21.285 290.13 21.355 ;
    RECT 289.92 21.645 290.13 21.715 ;
    RECT 289.46 20.925 289.67 20.995 ;
    RECT 289.46 21.285 289.67 21.355 ;
    RECT 289.46 21.645 289.67 21.715 ;
    RECT 286.6 20.925 286.81 20.995 ;
    RECT 286.6 21.285 286.81 21.355 ;
    RECT 286.6 21.645 286.81 21.715 ;
    RECT 286.14 20.925 286.35 20.995 ;
    RECT 286.14 21.285 286.35 21.355 ;
    RECT 286.14 21.645 286.35 21.715 ;
    RECT 283.28 20.925 283.49 20.995 ;
    RECT 283.28 21.285 283.49 21.355 ;
    RECT 283.28 21.645 283.49 21.715 ;
    RECT 282.82 20.925 283.03 20.995 ;
    RECT 282.82 21.285 283.03 21.355 ;
    RECT 282.82 21.645 283.03 21.715 ;
    RECT 279.96 20.925 280.17 20.995 ;
    RECT 279.96 21.285 280.17 21.355 ;
    RECT 279.96 21.645 280.17 21.715 ;
    RECT 279.5 20.925 279.71 20.995 ;
    RECT 279.5 21.285 279.71 21.355 ;
    RECT 279.5 21.645 279.71 21.715 ;
    RECT 276.64 20.925 276.85 20.995 ;
    RECT 276.64 21.285 276.85 21.355 ;
    RECT 276.64 21.645 276.85 21.715 ;
    RECT 276.18 20.925 276.39 20.995 ;
    RECT 276.18 21.285 276.39 21.355 ;
    RECT 276.18 21.645 276.39 21.715 ;
    RECT 273.32 20.925 273.53 20.995 ;
    RECT 273.32 21.285 273.53 21.355 ;
    RECT 273.32 21.645 273.53 21.715 ;
    RECT 272.86 20.925 273.07 20.995 ;
    RECT 272.86 21.285 273.07 21.355 ;
    RECT 272.86 21.645 273.07 21.715 ;
    RECT 270.0 20.925 270.21 20.995 ;
    RECT 270.0 21.285 270.21 21.355 ;
    RECT 270.0 21.645 270.21 21.715 ;
    RECT 269.54 20.925 269.75 20.995 ;
    RECT 269.54 21.285 269.75 21.355 ;
    RECT 269.54 21.645 269.75 21.715 ;
    RECT 233.48 20.925 233.69 20.995 ;
    RECT 233.48 21.285 233.69 21.355 ;
    RECT 233.48 21.645 233.69 21.715 ;
    RECT 233.02 20.925 233.23 20.995 ;
    RECT 233.02 21.285 233.23 21.355 ;
    RECT 233.02 21.645 233.23 21.715 ;
    RECT 230.16 20.925 230.37 20.995 ;
    RECT 230.16 21.285 230.37 21.355 ;
    RECT 230.16 21.645 230.37 21.715 ;
    RECT 229.7 20.925 229.91 20.995 ;
    RECT 229.7 21.285 229.91 21.355 ;
    RECT 229.7 21.645 229.91 21.715 ;
    RECT 366.28 20.925 366.49 20.995 ;
    RECT 366.28 21.285 366.49 21.355 ;
    RECT 366.28 21.645 366.49 21.715 ;
    RECT 365.82 20.925 366.03 20.995 ;
    RECT 365.82 21.285 366.03 21.355 ;
    RECT 365.82 21.645 366.03 21.715 ;
    RECT 226.84 20.925 227.05 20.995 ;
    RECT 226.84 21.285 227.05 21.355 ;
    RECT 226.84 21.645 227.05 21.715 ;
    RECT 226.38 20.925 226.59 20.995 ;
    RECT 226.38 21.285 226.59 21.355 ;
    RECT 226.38 21.645 226.59 21.715 ;
    RECT 362.96 20.925 363.17 20.995 ;
    RECT 362.96 21.285 363.17 21.355 ;
    RECT 362.96 21.645 363.17 21.715 ;
    RECT 362.5 20.925 362.71 20.995 ;
    RECT 362.5 21.285 362.71 21.355 ;
    RECT 362.5 21.645 362.71 21.715 ;
    RECT 223.52 20.925 223.73 20.995 ;
    RECT 223.52 21.285 223.73 21.355 ;
    RECT 223.52 21.645 223.73 21.715 ;
    RECT 223.06 20.925 223.27 20.995 ;
    RECT 223.06 21.285 223.27 21.355 ;
    RECT 223.06 21.645 223.27 21.715 ;
    RECT 359.64 20.925 359.85 20.995 ;
    RECT 359.64 21.285 359.85 21.355 ;
    RECT 359.64 21.645 359.85 21.715 ;
    RECT 359.18 20.925 359.39 20.995 ;
    RECT 359.18 21.285 359.39 21.355 ;
    RECT 359.18 21.645 359.39 21.715 ;
    RECT 220.2 20.925 220.41 20.995 ;
    RECT 220.2 21.285 220.41 21.355 ;
    RECT 220.2 21.645 220.41 21.715 ;
    RECT 219.74 20.925 219.95 20.995 ;
    RECT 219.74 21.285 219.95 21.355 ;
    RECT 219.74 21.645 219.95 21.715 ;
    RECT 356.32 20.925 356.53 20.995 ;
    RECT 356.32 21.285 356.53 21.355 ;
    RECT 356.32 21.645 356.53 21.715 ;
    RECT 355.86 20.925 356.07 20.995 ;
    RECT 355.86 21.285 356.07 21.355 ;
    RECT 355.86 21.645 356.07 21.715 ;
    RECT 353.0 20.925 353.21 20.995 ;
    RECT 353.0 21.285 353.21 21.355 ;
    RECT 353.0 21.645 353.21 21.715 ;
    RECT 352.54 20.925 352.75 20.995 ;
    RECT 352.54 21.285 352.75 21.355 ;
    RECT 352.54 21.645 352.75 21.715 ;
    RECT 216.88 20.925 217.09 20.995 ;
    RECT 216.88 21.285 217.09 21.355 ;
    RECT 216.88 21.645 217.09 21.715 ;
    RECT 216.42 20.925 216.63 20.995 ;
    RECT 216.42 21.285 216.63 21.355 ;
    RECT 216.42 21.645 216.63 21.715 ;
    RECT 349.68 20.925 349.89 20.995 ;
    RECT 349.68 21.285 349.89 21.355 ;
    RECT 349.68 21.645 349.89 21.715 ;
    RECT 349.22 20.925 349.43 20.995 ;
    RECT 349.22 21.285 349.43 21.355 ;
    RECT 349.22 21.645 349.43 21.715 ;
    RECT 213.56 20.925 213.77 20.995 ;
    RECT 213.56 21.285 213.77 21.355 ;
    RECT 213.56 21.645 213.77 21.715 ;
    RECT 213.1 20.925 213.31 20.995 ;
    RECT 213.1 21.285 213.31 21.355 ;
    RECT 213.1 21.645 213.31 21.715 ;
    RECT 346.36 20.925 346.57 20.995 ;
    RECT 346.36 21.285 346.57 21.355 ;
    RECT 346.36 21.645 346.57 21.715 ;
    RECT 345.9 20.925 346.11 20.995 ;
    RECT 345.9 21.285 346.11 21.355 ;
    RECT 345.9 21.645 346.11 21.715 ;
    RECT 210.24 20.925 210.45 20.995 ;
    RECT 210.24 21.285 210.45 21.355 ;
    RECT 210.24 21.645 210.45 21.715 ;
    RECT 209.78 20.925 209.99 20.995 ;
    RECT 209.78 21.285 209.99 21.355 ;
    RECT 209.78 21.645 209.99 21.715 ;
    RECT 343.04 20.925 343.25 20.995 ;
    RECT 343.04 21.285 343.25 21.355 ;
    RECT 343.04 21.645 343.25 21.715 ;
    RECT 342.58 20.925 342.79 20.995 ;
    RECT 342.58 21.285 342.79 21.355 ;
    RECT 342.58 21.645 342.79 21.715 ;
    RECT 206.92 20.925 207.13 20.995 ;
    RECT 206.92 21.285 207.13 21.355 ;
    RECT 206.92 21.645 207.13 21.715 ;
    RECT 206.46 20.925 206.67 20.995 ;
    RECT 206.46 21.285 206.67 21.355 ;
    RECT 206.46 21.645 206.67 21.715 ;
    RECT 339.72 20.925 339.93 20.995 ;
    RECT 339.72 21.285 339.93 21.355 ;
    RECT 339.72 21.645 339.93 21.715 ;
    RECT 339.26 20.925 339.47 20.995 ;
    RECT 339.26 21.285 339.47 21.355 ;
    RECT 339.26 21.645 339.47 21.715 ;
    RECT 203.6 20.925 203.81 20.995 ;
    RECT 203.6 21.285 203.81 21.355 ;
    RECT 203.6 21.645 203.81 21.715 ;
    RECT 203.14 20.925 203.35 20.995 ;
    RECT 203.14 21.285 203.35 21.355 ;
    RECT 203.14 21.645 203.35 21.715 ;
    RECT 336.4 20.925 336.61 20.995 ;
    RECT 336.4 21.285 336.61 21.355 ;
    RECT 336.4 21.645 336.61 21.715 ;
    RECT 335.94 20.925 336.15 20.995 ;
    RECT 335.94 21.285 336.15 21.355 ;
    RECT 335.94 21.645 336.15 21.715 ;
    RECT 266.68 20.925 266.89 20.995 ;
    RECT 266.68 21.285 266.89 21.355 ;
    RECT 266.68 21.645 266.89 21.715 ;
    RECT 266.22 20.925 266.43 20.995 ;
    RECT 266.22 21.285 266.43 21.355 ;
    RECT 266.22 21.645 266.43 21.715 ;
    RECT 263.36 20.925 263.57 20.995 ;
    RECT 263.36 21.285 263.57 21.355 ;
    RECT 263.36 21.645 263.57 21.715 ;
    RECT 262.9 20.925 263.11 20.995 ;
    RECT 262.9 21.285 263.11 21.355 ;
    RECT 262.9 21.645 263.11 21.715 ;
    RECT 260.04 20.925 260.25 20.995 ;
    RECT 260.04 21.285 260.25 21.355 ;
    RECT 260.04 21.645 260.25 21.715 ;
    RECT 259.58 20.925 259.79 20.995 ;
    RECT 259.58 21.285 259.79 21.355 ;
    RECT 259.58 21.645 259.79 21.715 ;
    RECT 256.72 20.925 256.93 20.995 ;
    RECT 256.72 21.285 256.93 21.355 ;
    RECT 256.72 21.645 256.93 21.715 ;
    RECT 256.26 20.925 256.47 20.995 ;
    RECT 256.26 21.285 256.47 21.355 ;
    RECT 256.26 21.645 256.47 21.715 ;
    RECT 253.4 20.925 253.61 20.995 ;
    RECT 253.4 21.285 253.61 21.355 ;
    RECT 253.4 21.645 253.61 21.715 ;
    RECT 252.94 20.925 253.15 20.995 ;
    RECT 252.94 21.285 253.15 21.355 ;
    RECT 252.94 21.645 253.15 21.715 ;
    RECT 250.08 20.925 250.29 20.995 ;
    RECT 250.08 21.285 250.29 21.355 ;
    RECT 250.08 21.645 250.29 21.715 ;
    RECT 249.62 20.925 249.83 20.995 ;
    RECT 249.62 21.285 249.83 21.355 ;
    RECT 249.62 21.645 249.83 21.715 ;
    RECT 246.76 20.925 246.97 20.995 ;
    RECT 246.76 21.285 246.97 21.355 ;
    RECT 246.76 21.645 246.97 21.715 ;
    RECT 246.3 20.925 246.51 20.995 ;
    RECT 246.3 21.285 246.51 21.355 ;
    RECT 246.3 21.645 246.51 21.715 ;
    RECT 243.44 20.925 243.65 20.995 ;
    RECT 243.44 21.285 243.65 21.355 ;
    RECT 243.44 21.645 243.65 21.715 ;
    RECT 242.98 20.925 243.19 20.995 ;
    RECT 242.98 21.285 243.19 21.355 ;
    RECT 242.98 21.645 243.19 21.715 ;
    RECT 240.12 20.925 240.33 20.995 ;
    RECT 240.12 21.285 240.33 21.355 ;
    RECT 240.12 21.645 240.33 21.715 ;
    RECT 239.66 20.925 239.87 20.995 ;
    RECT 239.66 21.285 239.87 21.355 ;
    RECT 239.66 21.645 239.87 21.715 ;
    RECT 236.8 20.925 237.01 20.995 ;
    RECT 236.8 21.285 237.01 21.355 ;
    RECT 236.8 21.645 237.01 21.715 ;
    RECT 236.34 20.925 236.55 20.995 ;
    RECT 236.34 21.285 236.55 21.355 ;
    RECT 236.34 21.645 236.55 21.715 ;
    RECT 374.15 21.285 374.22 21.355 ;
    RECT 333.08 20.925 333.29 20.995 ;
    RECT 333.08 21.285 333.29 21.355 ;
    RECT 333.08 21.645 333.29 21.715 ;
    RECT 332.62 20.925 332.83 20.995 ;
    RECT 332.62 21.285 332.83 21.355 ;
    RECT 332.62 21.645 332.83 21.715 ;
    RECT 329.76 20.925 329.97 20.995 ;
    RECT 329.76 21.285 329.97 21.355 ;
    RECT 329.76 21.645 329.97 21.715 ;
    RECT 329.3 20.925 329.51 20.995 ;
    RECT 329.3 21.285 329.51 21.355 ;
    RECT 329.3 21.645 329.51 21.715 ;
    RECT 326.44 20.925 326.65 20.995 ;
    RECT 326.44 21.285 326.65 21.355 ;
    RECT 326.44 21.645 326.65 21.715 ;
    RECT 325.98 20.925 326.19 20.995 ;
    RECT 325.98 21.285 326.19 21.355 ;
    RECT 325.98 21.645 326.19 21.715 ;
    RECT 323.12 20.925 323.33 20.995 ;
    RECT 323.12 21.285 323.33 21.355 ;
    RECT 323.12 21.645 323.33 21.715 ;
    RECT 322.66 20.925 322.87 20.995 ;
    RECT 322.66 21.285 322.87 21.355 ;
    RECT 322.66 21.645 322.87 21.715 ;
    RECT 319.8 20.925 320.01 20.995 ;
    RECT 319.8 21.285 320.01 21.355 ;
    RECT 319.8 21.645 320.01 21.715 ;
    RECT 319.34 20.925 319.55 20.995 ;
    RECT 319.34 21.285 319.55 21.355 ;
    RECT 319.34 21.645 319.55 21.715 ;
    RECT 316.48 20.925 316.69 20.995 ;
    RECT 316.48 21.285 316.69 21.355 ;
    RECT 316.48 21.645 316.69 21.715 ;
    RECT 316.02 20.925 316.23 20.995 ;
    RECT 316.02 21.285 316.23 21.355 ;
    RECT 316.02 21.645 316.23 21.715 ;
    RECT 313.16 20.925 313.37 20.995 ;
    RECT 313.16 21.285 313.37 21.355 ;
    RECT 313.16 21.645 313.37 21.715 ;
    RECT 312.7 20.925 312.91 20.995 ;
    RECT 312.7 21.285 312.91 21.355 ;
    RECT 312.7 21.645 312.91 21.715 ;
    RECT 309.84 20.925 310.05 20.995 ;
    RECT 309.84 21.285 310.05 21.355 ;
    RECT 309.84 21.645 310.05 21.715 ;
    RECT 309.38 20.925 309.59 20.995 ;
    RECT 309.38 21.285 309.59 21.355 ;
    RECT 309.38 21.645 309.59 21.715 ;
    RECT 306.52 20.925 306.73 20.995 ;
    RECT 306.52 21.285 306.73 21.355 ;
    RECT 306.52 21.645 306.73 21.715 ;
    RECT 306.06 20.925 306.27 20.995 ;
    RECT 306.06 21.285 306.27 21.355 ;
    RECT 306.06 21.645 306.27 21.715 ;
    RECT 303.2 34.605 303.41 34.675 ;
    RECT 303.2 34.965 303.41 35.035 ;
    RECT 303.2 35.325 303.41 35.395 ;
    RECT 302.74 34.605 302.95 34.675 ;
    RECT 302.74 34.965 302.95 35.035 ;
    RECT 302.74 35.325 302.95 35.395 ;
    RECT 200.605 34.965 200.675 35.035 ;
    RECT 372.92 34.605 373.13 34.675 ;
    RECT 372.92 34.965 373.13 35.035 ;
    RECT 372.92 35.325 373.13 35.395 ;
    RECT 372.46 34.605 372.67 34.675 ;
    RECT 372.46 34.965 372.67 35.035 ;
    RECT 372.46 35.325 372.67 35.395 ;
    RECT 369.6 34.605 369.81 34.675 ;
    RECT 369.6 34.965 369.81 35.035 ;
    RECT 369.6 35.325 369.81 35.395 ;
    RECT 369.14 34.605 369.35 34.675 ;
    RECT 369.14 34.965 369.35 35.035 ;
    RECT 369.14 35.325 369.35 35.395 ;
    RECT 299.88 34.605 300.09 34.675 ;
    RECT 299.88 34.965 300.09 35.035 ;
    RECT 299.88 35.325 300.09 35.395 ;
    RECT 299.42 34.605 299.63 34.675 ;
    RECT 299.42 34.965 299.63 35.035 ;
    RECT 299.42 35.325 299.63 35.395 ;
    RECT 296.56 34.605 296.77 34.675 ;
    RECT 296.56 34.965 296.77 35.035 ;
    RECT 296.56 35.325 296.77 35.395 ;
    RECT 296.1 34.605 296.31 34.675 ;
    RECT 296.1 34.965 296.31 35.035 ;
    RECT 296.1 35.325 296.31 35.395 ;
    RECT 293.24 34.605 293.45 34.675 ;
    RECT 293.24 34.965 293.45 35.035 ;
    RECT 293.24 35.325 293.45 35.395 ;
    RECT 292.78 34.605 292.99 34.675 ;
    RECT 292.78 34.965 292.99 35.035 ;
    RECT 292.78 35.325 292.99 35.395 ;
    RECT 289.92 34.605 290.13 34.675 ;
    RECT 289.92 34.965 290.13 35.035 ;
    RECT 289.92 35.325 290.13 35.395 ;
    RECT 289.46 34.605 289.67 34.675 ;
    RECT 289.46 34.965 289.67 35.035 ;
    RECT 289.46 35.325 289.67 35.395 ;
    RECT 286.6 34.605 286.81 34.675 ;
    RECT 286.6 34.965 286.81 35.035 ;
    RECT 286.6 35.325 286.81 35.395 ;
    RECT 286.14 34.605 286.35 34.675 ;
    RECT 286.14 34.965 286.35 35.035 ;
    RECT 286.14 35.325 286.35 35.395 ;
    RECT 283.28 34.605 283.49 34.675 ;
    RECT 283.28 34.965 283.49 35.035 ;
    RECT 283.28 35.325 283.49 35.395 ;
    RECT 282.82 34.605 283.03 34.675 ;
    RECT 282.82 34.965 283.03 35.035 ;
    RECT 282.82 35.325 283.03 35.395 ;
    RECT 279.96 34.605 280.17 34.675 ;
    RECT 279.96 34.965 280.17 35.035 ;
    RECT 279.96 35.325 280.17 35.395 ;
    RECT 279.5 34.605 279.71 34.675 ;
    RECT 279.5 34.965 279.71 35.035 ;
    RECT 279.5 35.325 279.71 35.395 ;
    RECT 276.64 34.605 276.85 34.675 ;
    RECT 276.64 34.965 276.85 35.035 ;
    RECT 276.64 35.325 276.85 35.395 ;
    RECT 276.18 34.605 276.39 34.675 ;
    RECT 276.18 34.965 276.39 35.035 ;
    RECT 276.18 35.325 276.39 35.395 ;
    RECT 273.32 34.605 273.53 34.675 ;
    RECT 273.32 34.965 273.53 35.035 ;
    RECT 273.32 35.325 273.53 35.395 ;
    RECT 272.86 34.605 273.07 34.675 ;
    RECT 272.86 34.965 273.07 35.035 ;
    RECT 272.86 35.325 273.07 35.395 ;
    RECT 270.0 34.605 270.21 34.675 ;
    RECT 270.0 34.965 270.21 35.035 ;
    RECT 270.0 35.325 270.21 35.395 ;
    RECT 269.54 34.605 269.75 34.675 ;
    RECT 269.54 34.965 269.75 35.035 ;
    RECT 269.54 35.325 269.75 35.395 ;
    RECT 233.48 34.605 233.69 34.675 ;
    RECT 233.48 34.965 233.69 35.035 ;
    RECT 233.48 35.325 233.69 35.395 ;
    RECT 233.02 34.605 233.23 34.675 ;
    RECT 233.02 34.965 233.23 35.035 ;
    RECT 233.02 35.325 233.23 35.395 ;
    RECT 230.16 34.605 230.37 34.675 ;
    RECT 230.16 34.965 230.37 35.035 ;
    RECT 230.16 35.325 230.37 35.395 ;
    RECT 229.7 34.605 229.91 34.675 ;
    RECT 229.7 34.965 229.91 35.035 ;
    RECT 229.7 35.325 229.91 35.395 ;
    RECT 366.28 34.605 366.49 34.675 ;
    RECT 366.28 34.965 366.49 35.035 ;
    RECT 366.28 35.325 366.49 35.395 ;
    RECT 365.82 34.605 366.03 34.675 ;
    RECT 365.82 34.965 366.03 35.035 ;
    RECT 365.82 35.325 366.03 35.395 ;
    RECT 226.84 34.605 227.05 34.675 ;
    RECT 226.84 34.965 227.05 35.035 ;
    RECT 226.84 35.325 227.05 35.395 ;
    RECT 226.38 34.605 226.59 34.675 ;
    RECT 226.38 34.965 226.59 35.035 ;
    RECT 226.38 35.325 226.59 35.395 ;
    RECT 362.96 34.605 363.17 34.675 ;
    RECT 362.96 34.965 363.17 35.035 ;
    RECT 362.96 35.325 363.17 35.395 ;
    RECT 362.5 34.605 362.71 34.675 ;
    RECT 362.5 34.965 362.71 35.035 ;
    RECT 362.5 35.325 362.71 35.395 ;
    RECT 223.52 34.605 223.73 34.675 ;
    RECT 223.52 34.965 223.73 35.035 ;
    RECT 223.52 35.325 223.73 35.395 ;
    RECT 223.06 34.605 223.27 34.675 ;
    RECT 223.06 34.965 223.27 35.035 ;
    RECT 223.06 35.325 223.27 35.395 ;
    RECT 359.64 34.605 359.85 34.675 ;
    RECT 359.64 34.965 359.85 35.035 ;
    RECT 359.64 35.325 359.85 35.395 ;
    RECT 359.18 34.605 359.39 34.675 ;
    RECT 359.18 34.965 359.39 35.035 ;
    RECT 359.18 35.325 359.39 35.395 ;
    RECT 220.2 34.605 220.41 34.675 ;
    RECT 220.2 34.965 220.41 35.035 ;
    RECT 220.2 35.325 220.41 35.395 ;
    RECT 219.74 34.605 219.95 34.675 ;
    RECT 219.74 34.965 219.95 35.035 ;
    RECT 219.74 35.325 219.95 35.395 ;
    RECT 356.32 34.605 356.53 34.675 ;
    RECT 356.32 34.965 356.53 35.035 ;
    RECT 356.32 35.325 356.53 35.395 ;
    RECT 355.86 34.605 356.07 34.675 ;
    RECT 355.86 34.965 356.07 35.035 ;
    RECT 355.86 35.325 356.07 35.395 ;
    RECT 374.15 34.965 374.22 35.035 ;
    RECT 353.0 34.605 353.21 34.675 ;
    RECT 353.0 34.965 353.21 35.035 ;
    RECT 353.0 35.325 353.21 35.395 ;
    RECT 352.54 34.605 352.75 34.675 ;
    RECT 352.54 34.965 352.75 35.035 ;
    RECT 352.54 35.325 352.75 35.395 ;
    RECT 216.88 34.605 217.09 34.675 ;
    RECT 216.88 34.965 217.09 35.035 ;
    RECT 216.88 35.325 217.09 35.395 ;
    RECT 216.42 34.605 216.63 34.675 ;
    RECT 216.42 34.965 216.63 35.035 ;
    RECT 216.42 35.325 216.63 35.395 ;
    RECT 349.68 34.605 349.89 34.675 ;
    RECT 349.68 34.965 349.89 35.035 ;
    RECT 349.68 35.325 349.89 35.395 ;
    RECT 349.22 34.605 349.43 34.675 ;
    RECT 349.22 34.965 349.43 35.035 ;
    RECT 349.22 35.325 349.43 35.395 ;
    RECT 213.56 34.605 213.77 34.675 ;
    RECT 213.56 34.965 213.77 35.035 ;
    RECT 213.56 35.325 213.77 35.395 ;
    RECT 213.1 34.605 213.31 34.675 ;
    RECT 213.1 34.965 213.31 35.035 ;
    RECT 213.1 35.325 213.31 35.395 ;
    RECT 346.36 34.605 346.57 34.675 ;
    RECT 346.36 34.965 346.57 35.035 ;
    RECT 346.36 35.325 346.57 35.395 ;
    RECT 345.9 34.605 346.11 34.675 ;
    RECT 345.9 34.965 346.11 35.035 ;
    RECT 345.9 35.325 346.11 35.395 ;
    RECT 210.24 34.605 210.45 34.675 ;
    RECT 210.24 34.965 210.45 35.035 ;
    RECT 210.24 35.325 210.45 35.395 ;
    RECT 209.78 34.605 209.99 34.675 ;
    RECT 209.78 34.965 209.99 35.035 ;
    RECT 209.78 35.325 209.99 35.395 ;
    RECT 343.04 34.605 343.25 34.675 ;
    RECT 343.04 34.965 343.25 35.035 ;
    RECT 343.04 35.325 343.25 35.395 ;
    RECT 342.58 34.605 342.79 34.675 ;
    RECT 342.58 34.965 342.79 35.035 ;
    RECT 342.58 35.325 342.79 35.395 ;
    RECT 206.92 34.605 207.13 34.675 ;
    RECT 206.92 34.965 207.13 35.035 ;
    RECT 206.92 35.325 207.13 35.395 ;
    RECT 206.46 34.605 206.67 34.675 ;
    RECT 206.46 34.965 206.67 35.035 ;
    RECT 206.46 35.325 206.67 35.395 ;
    RECT 339.72 34.605 339.93 34.675 ;
    RECT 339.72 34.965 339.93 35.035 ;
    RECT 339.72 35.325 339.93 35.395 ;
    RECT 339.26 34.605 339.47 34.675 ;
    RECT 339.26 34.965 339.47 35.035 ;
    RECT 339.26 35.325 339.47 35.395 ;
    RECT 203.6 34.605 203.81 34.675 ;
    RECT 203.6 34.965 203.81 35.035 ;
    RECT 203.6 35.325 203.81 35.395 ;
    RECT 203.14 34.605 203.35 34.675 ;
    RECT 203.14 34.965 203.35 35.035 ;
    RECT 203.14 35.325 203.35 35.395 ;
    RECT 336.4 34.605 336.61 34.675 ;
    RECT 336.4 34.965 336.61 35.035 ;
    RECT 336.4 35.325 336.61 35.395 ;
    RECT 335.94 34.605 336.15 34.675 ;
    RECT 335.94 34.965 336.15 35.035 ;
    RECT 335.94 35.325 336.15 35.395 ;
    RECT 266.68 34.605 266.89 34.675 ;
    RECT 266.68 34.965 266.89 35.035 ;
    RECT 266.68 35.325 266.89 35.395 ;
    RECT 266.22 34.605 266.43 34.675 ;
    RECT 266.22 34.965 266.43 35.035 ;
    RECT 266.22 35.325 266.43 35.395 ;
    RECT 263.36 34.605 263.57 34.675 ;
    RECT 263.36 34.965 263.57 35.035 ;
    RECT 263.36 35.325 263.57 35.395 ;
    RECT 262.9 34.605 263.11 34.675 ;
    RECT 262.9 34.965 263.11 35.035 ;
    RECT 262.9 35.325 263.11 35.395 ;
    RECT 260.04 34.605 260.25 34.675 ;
    RECT 260.04 34.965 260.25 35.035 ;
    RECT 260.04 35.325 260.25 35.395 ;
    RECT 259.58 34.605 259.79 34.675 ;
    RECT 259.58 34.965 259.79 35.035 ;
    RECT 259.58 35.325 259.79 35.395 ;
    RECT 256.72 34.605 256.93 34.675 ;
    RECT 256.72 34.965 256.93 35.035 ;
    RECT 256.72 35.325 256.93 35.395 ;
    RECT 256.26 34.605 256.47 34.675 ;
    RECT 256.26 34.965 256.47 35.035 ;
    RECT 256.26 35.325 256.47 35.395 ;
    RECT 253.4 34.605 253.61 34.675 ;
    RECT 253.4 34.965 253.61 35.035 ;
    RECT 253.4 35.325 253.61 35.395 ;
    RECT 252.94 34.605 253.15 34.675 ;
    RECT 252.94 34.965 253.15 35.035 ;
    RECT 252.94 35.325 253.15 35.395 ;
    RECT 250.08 34.605 250.29 34.675 ;
    RECT 250.08 34.965 250.29 35.035 ;
    RECT 250.08 35.325 250.29 35.395 ;
    RECT 249.62 34.605 249.83 34.675 ;
    RECT 249.62 34.965 249.83 35.035 ;
    RECT 249.62 35.325 249.83 35.395 ;
    RECT 246.76 34.605 246.97 34.675 ;
    RECT 246.76 34.965 246.97 35.035 ;
    RECT 246.76 35.325 246.97 35.395 ;
    RECT 246.3 34.605 246.51 34.675 ;
    RECT 246.3 34.965 246.51 35.035 ;
    RECT 246.3 35.325 246.51 35.395 ;
    RECT 243.44 34.605 243.65 34.675 ;
    RECT 243.44 34.965 243.65 35.035 ;
    RECT 243.44 35.325 243.65 35.395 ;
    RECT 242.98 34.605 243.19 34.675 ;
    RECT 242.98 34.965 243.19 35.035 ;
    RECT 242.98 35.325 243.19 35.395 ;
    RECT 240.12 34.605 240.33 34.675 ;
    RECT 240.12 34.965 240.33 35.035 ;
    RECT 240.12 35.325 240.33 35.395 ;
    RECT 239.66 34.605 239.87 34.675 ;
    RECT 239.66 34.965 239.87 35.035 ;
    RECT 239.66 35.325 239.87 35.395 ;
    RECT 236.8 34.605 237.01 34.675 ;
    RECT 236.8 34.965 237.01 35.035 ;
    RECT 236.8 35.325 237.01 35.395 ;
    RECT 236.34 34.605 236.55 34.675 ;
    RECT 236.34 34.965 236.55 35.035 ;
    RECT 236.34 35.325 236.55 35.395 ;
    RECT 333.08 34.605 333.29 34.675 ;
    RECT 333.08 34.965 333.29 35.035 ;
    RECT 333.08 35.325 333.29 35.395 ;
    RECT 332.62 34.605 332.83 34.675 ;
    RECT 332.62 34.965 332.83 35.035 ;
    RECT 332.62 35.325 332.83 35.395 ;
    RECT 329.76 34.605 329.97 34.675 ;
    RECT 329.76 34.965 329.97 35.035 ;
    RECT 329.76 35.325 329.97 35.395 ;
    RECT 329.3 34.605 329.51 34.675 ;
    RECT 329.3 34.965 329.51 35.035 ;
    RECT 329.3 35.325 329.51 35.395 ;
    RECT 326.44 34.605 326.65 34.675 ;
    RECT 326.44 34.965 326.65 35.035 ;
    RECT 326.44 35.325 326.65 35.395 ;
    RECT 325.98 34.605 326.19 34.675 ;
    RECT 325.98 34.965 326.19 35.035 ;
    RECT 325.98 35.325 326.19 35.395 ;
    RECT 323.12 34.605 323.33 34.675 ;
    RECT 323.12 34.965 323.33 35.035 ;
    RECT 323.12 35.325 323.33 35.395 ;
    RECT 322.66 34.605 322.87 34.675 ;
    RECT 322.66 34.965 322.87 35.035 ;
    RECT 322.66 35.325 322.87 35.395 ;
    RECT 319.8 34.605 320.01 34.675 ;
    RECT 319.8 34.965 320.01 35.035 ;
    RECT 319.8 35.325 320.01 35.395 ;
    RECT 319.34 34.605 319.55 34.675 ;
    RECT 319.34 34.965 319.55 35.035 ;
    RECT 319.34 35.325 319.55 35.395 ;
    RECT 316.48 34.605 316.69 34.675 ;
    RECT 316.48 34.965 316.69 35.035 ;
    RECT 316.48 35.325 316.69 35.395 ;
    RECT 316.02 34.605 316.23 34.675 ;
    RECT 316.02 34.965 316.23 35.035 ;
    RECT 316.02 35.325 316.23 35.395 ;
    RECT 313.16 34.605 313.37 34.675 ;
    RECT 313.16 34.965 313.37 35.035 ;
    RECT 313.16 35.325 313.37 35.395 ;
    RECT 312.7 34.605 312.91 34.675 ;
    RECT 312.7 34.965 312.91 35.035 ;
    RECT 312.7 35.325 312.91 35.395 ;
    RECT 309.84 34.605 310.05 34.675 ;
    RECT 309.84 34.965 310.05 35.035 ;
    RECT 309.84 35.325 310.05 35.395 ;
    RECT 309.38 34.605 309.59 34.675 ;
    RECT 309.38 34.965 309.59 35.035 ;
    RECT 309.38 35.325 309.59 35.395 ;
    RECT 306.52 34.605 306.73 34.675 ;
    RECT 306.52 34.965 306.73 35.035 ;
    RECT 306.52 35.325 306.73 35.395 ;
    RECT 306.06 34.605 306.27 34.675 ;
    RECT 306.06 34.965 306.27 35.035 ;
    RECT 306.06 35.325 306.27 35.395 ;
    RECT 303.2 20.205 303.41 20.275 ;
    RECT 303.2 20.565 303.41 20.635 ;
    RECT 303.2 20.925 303.41 20.995 ;
    RECT 302.74 20.205 302.95 20.275 ;
    RECT 302.74 20.565 302.95 20.635 ;
    RECT 302.74 20.925 302.95 20.995 ;
    RECT 372.92 20.205 373.13 20.275 ;
    RECT 372.92 20.565 373.13 20.635 ;
    RECT 372.92 20.925 373.13 20.995 ;
    RECT 372.46 20.205 372.67 20.275 ;
    RECT 372.46 20.565 372.67 20.635 ;
    RECT 372.46 20.925 372.67 20.995 ;
    RECT 369.6 20.205 369.81 20.275 ;
    RECT 369.6 20.565 369.81 20.635 ;
    RECT 369.6 20.925 369.81 20.995 ;
    RECT 369.14 20.205 369.35 20.275 ;
    RECT 369.14 20.565 369.35 20.635 ;
    RECT 369.14 20.925 369.35 20.995 ;
    RECT 200.605 20.565 200.675 20.635 ;
    RECT 299.88 20.205 300.09 20.275 ;
    RECT 299.88 20.565 300.09 20.635 ;
    RECT 299.88 20.925 300.09 20.995 ;
    RECT 299.42 20.205 299.63 20.275 ;
    RECT 299.42 20.565 299.63 20.635 ;
    RECT 299.42 20.925 299.63 20.995 ;
    RECT 296.56 20.205 296.77 20.275 ;
    RECT 296.56 20.565 296.77 20.635 ;
    RECT 296.56 20.925 296.77 20.995 ;
    RECT 296.1 20.205 296.31 20.275 ;
    RECT 296.1 20.565 296.31 20.635 ;
    RECT 296.1 20.925 296.31 20.995 ;
    RECT 293.24 20.205 293.45 20.275 ;
    RECT 293.24 20.565 293.45 20.635 ;
    RECT 293.24 20.925 293.45 20.995 ;
    RECT 292.78 20.205 292.99 20.275 ;
    RECT 292.78 20.565 292.99 20.635 ;
    RECT 292.78 20.925 292.99 20.995 ;
    RECT 289.92 20.205 290.13 20.275 ;
    RECT 289.92 20.565 290.13 20.635 ;
    RECT 289.92 20.925 290.13 20.995 ;
    RECT 289.46 20.205 289.67 20.275 ;
    RECT 289.46 20.565 289.67 20.635 ;
    RECT 289.46 20.925 289.67 20.995 ;
    RECT 286.6 20.205 286.81 20.275 ;
    RECT 286.6 20.565 286.81 20.635 ;
    RECT 286.6 20.925 286.81 20.995 ;
    RECT 286.14 20.205 286.35 20.275 ;
    RECT 286.14 20.565 286.35 20.635 ;
    RECT 286.14 20.925 286.35 20.995 ;
    RECT 283.28 20.205 283.49 20.275 ;
    RECT 283.28 20.565 283.49 20.635 ;
    RECT 283.28 20.925 283.49 20.995 ;
    RECT 282.82 20.205 283.03 20.275 ;
    RECT 282.82 20.565 283.03 20.635 ;
    RECT 282.82 20.925 283.03 20.995 ;
    RECT 279.96 20.205 280.17 20.275 ;
    RECT 279.96 20.565 280.17 20.635 ;
    RECT 279.96 20.925 280.17 20.995 ;
    RECT 279.5 20.205 279.71 20.275 ;
    RECT 279.5 20.565 279.71 20.635 ;
    RECT 279.5 20.925 279.71 20.995 ;
    RECT 276.64 20.205 276.85 20.275 ;
    RECT 276.64 20.565 276.85 20.635 ;
    RECT 276.64 20.925 276.85 20.995 ;
    RECT 276.18 20.205 276.39 20.275 ;
    RECT 276.18 20.565 276.39 20.635 ;
    RECT 276.18 20.925 276.39 20.995 ;
    RECT 273.32 20.205 273.53 20.275 ;
    RECT 273.32 20.565 273.53 20.635 ;
    RECT 273.32 20.925 273.53 20.995 ;
    RECT 272.86 20.205 273.07 20.275 ;
    RECT 272.86 20.565 273.07 20.635 ;
    RECT 272.86 20.925 273.07 20.995 ;
    RECT 270.0 20.205 270.21 20.275 ;
    RECT 270.0 20.565 270.21 20.635 ;
    RECT 270.0 20.925 270.21 20.995 ;
    RECT 269.54 20.205 269.75 20.275 ;
    RECT 269.54 20.565 269.75 20.635 ;
    RECT 269.54 20.925 269.75 20.995 ;
    RECT 233.48 20.205 233.69 20.275 ;
    RECT 233.48 20.565 233.69 20.635 ;
    RECT 233.48 20.925 233.69 20.995 ;
    RECT 233.02 20.205 233.23 20.275 ;
    RECT 233.02 20.565 233.23 20.635 ;
    RECT 233.02 20.925 233.23 20.995 ;
    RECT 230.16 20.205 230.37 20.275 ;
    RECT 230.16 20.565 230.37 20.635 ;
    RECT 230.16 20.925 230.37 20.995 ;
    RECT 229.7 20.205 229.91 20.275 ;
    RECT 229.7 20.565 229.91 20.635 ;
    RECT 229.7 20.925 229.91 20.995 ;
    RECT 366.28 20.205 366.49 20.275 ;
    RECT 366.28 20.565 366.49 20.635 ;
    RECT 366.28 20.925 366.49 20.995 ;
    RECT 365.82 20.205 366.03 20.275 ;
    RECT 365.82 20.565 366.03 20.635 ;
    RECT 365.82 20.925 366.03 20.995 ;
    RECT 226.84 20.205 227.05 20.275 ;
    RECT 226.84 20.565 227.05 20.635 ;
    RECT 226.84 20.925 227.05 20.995 ;
    RECT 226.38 20.205 226.59 20.275 ;
    RECT 226.38 20.565 226.59 20.635 ;
    RECT 226.38 20.925 226.59 20.995 ;
    RECT 362.96 20.205 363.17 20.275 ;
    RECT 362.96 20.565 363.17 20.635 ;
    RECT 362.96 20.925 363.17 20.995 ;
    RECT 362.5 20.205 362.71 20.275 ;
    RECT 362.5 20.565 362.71 20.635 ;
    RECT 362.5 20.925 362.71 20.995 ;
    RECT 223.52 20.205 223.73 20.275 ;
    RECT 223.52 20.565 223.73 20.635 ;
    RECT 223.52 20.925 223.73 20.995 ;
    RECT 223.06 20.205 223.27 20.275 ;
    RECT 223.06 20.565 223.27 20.635 ;
    RECT 223.06 20.925 223.27 20.995 ;
    RECT 359.64 20.205 359.85 20.275 ;
    RECT 359.64 20.565 359.85 20.635 ;
    RECT 359.64 20.925 359.85 20.995 ;
    RECT 359.18 20.205 359.39 20.275 ;
    RECT 359.18 20.565 359.39 20.635 ;
    RECT 359.18 20.925 359.39 20.995 ;
    RECT 220.2 20.205 220.41 20.275 ;
    RECT 220.2 20.565 220.41 20.635 ;
    RECT 220.2 20.925 220.41 20.995 ;
    RECT 219.74 20.205 219.95 20.275 ;
    RECT 219.74 20.565 219.95 20.635 ;
    RECT 219.74 20.925 219.95 20.995 ;
    RECT 356.32 20.205 356.53 20.275 ;
    RECT 356.32 20.565 356.53 20.635 ;
    RECT 356.32 20.925 356.53 20.995 ;
    RECT 355.86 20.205 356.07 20.275 ;
    RECT 355.86 20.565 356.07 20.635 ;
    RECT 355.86 20.925 356.07 20.995 ;
    RECT 353.0 20.205 353.21 20.275 ;
    RECT 353.0 20.565 353.21 20.635 ;
    RECT 353.0 20.925 353.21 20.995 ;
    RECT 352.54 20.205 352.75 20.275 ;
    RECT 352.54 20.565 352.75 20.635 ;
    RECT 352.54 20.925 352.75 20.995 ;
    RECT 216.88 20.205 217.09 20.275 ;
    RECT 216.88 20.565 217.09 20.635 ;
    RECT 216.88 20.925 217.09 20.995 ;
    RECT 216.42 20.205 216.63 20.275 ;
    RECT 216.42 20.565 216.63 20.635 ;
    RECT 216.42 20.925 216.63 20.995 ;
    RECT 349.68 20.205 349.89 20.275 ;
    RECT 349.68 20.565 349.89 20.635 ;
    RECT 349.68 20.925 349.89 20.995 ;
    RECT 349.22 20.205 349.43 20.275 ;
    RECT 349.22 20.565 349.43 20.635 ;
    RECT 349.22 20.925 349.43 20.995 ;
    RECT 213.56 20.205 213.77 20.275 ;
    RECT 213.56 20.565 213.77 20.635 ;
    RECT 213.56 20.925 213.77 20.995 ;
    RECT 213.1 20.205 213.31 20.275 ;
    RECT 213.1 20.565 213.31 20.635 ;
    RECT 213.1 20.925 213.31 20.995 ;
    RECT 346.36 20.205 346.57 20.275 ;
    RECT 346.36 20.565 346.57 20.635 ;
    RECT 346.36 20.925 346.57 20.995 ;
    RECT 345.9 20.205 346.11 20.275 ;
    RECT 345.9 20.565 346.11 20.635 ;
    RECT 345.9 20.925 346.11 20.995 ;
    RECT 210.24 20.205 210.45 20.275 ;
    RECT 210.24 20.565 210.45 20.635 ;
    RECT 210.24 20.925 210.45 20.995 ;
    RECT 209.78 20.205 209.99 20.275 ;
    RECT 209.78 20.565 209.99 20.635 ;
    RECT 209.78 20.925 209.99 20.995 ;
    RECT 343.04 20.205 343.25 20.275 ;
    RECT 343.04 20.565 343.25 20.635 ;
    RECT 343.04 20.925 343.25 20.995 ;
    RECT 342.58 20.205 342.79 20.275 ;
    RECT 342.58 20.565 342.79 20.635 ;
    RECT 342.58 20.925 342.79 20.995 ;
    RECT 206.92 20.205 207.13 20.275 ;
    RECT 206.92 20.565 207.13 20.635 ;
    RECT 206.92 20.925 207.13 20.995 ;
    RECT 206.46 20.205 206.67 20.275 ;
    RECT 206.46 20.565 206.67 20.635 ;
    RECT 206.46 20.925 206.67 20.995 ;
    RECT 339.72 20.205 339.93 20.275 ;
    RECT 339.72 20.565 339.93 20.635 ;
    RECT 339.72 20.925 339.93 20.995 ;
    RECT 339.26 20.205 339.47 20.275 ;
    RECT 339.26 20.565 339.47 20.635 ;
    RECT 339.26 20.925 339.47 20.995 ;
    RECT 203.6 20.205 203.81 20.275 ;
    RECT 203.6 20.565 203.81 20.635 ;
    RECT 203.6 20.925 203.81 20.995 ;
    RECT 203.14 20.205 203.35 20.275 ;
    RECT 203.14 20.565 203.35 20.635 ;
    RECT 203.14 20.925 203.35 20.995 ;
    RECT 336.4 20.205 336.61 20.275 ;
    RECT 336.4 20.565 336.61 20.635 ;
    RECT 336.4 20.925 336.61 20.995 ;
    RECT 335.94 20.205 336.15 20.275 ;
    RECT 335.94 20.565 336.15 20.635 ;
    RECT 335.94 20.925 336.15 20.995 ;
    RECT 266.68 20.205 266.89 20.275 ;
    RECT 266.68 20.565 266.89 20.635 ;
    RECT 266.68 20.925 266.89 20.995 ;
    RECT 266.22 20.205 266.43 20.275 ;
    RECT 266.22 20.565 266.43 20.635 ;
    RECT 266.22 20.925 266.43 20.995 ;
    RECT 263.36 20.205 263.57 20.275 ;
    RECT 263.36 20.565 263.57 20.635 ;
    RECT 263.36 20.925 263.57 20.995 ;
    RECT 262.9 20.205 263.11 20.275 ;
    RECT 262.9 20.565 263.11 20.635 ;
    RECT 262.9 20.925 263.11 20.995 ;
    RECT 260.04 20.205 260.25 20.275 ;
    RECT 260.04 20.565 260.25 20.635 ;
    RECT 260.04 20.925 260.25 20.995 ;
    RECT 259.58 20.205 259.79 20.275 ;
    RECT 259.58 20.565 259.79 20.635 ;
    RECT 259.58 20.925 259.79 20.995 ;
    RECT 256.72 20.205 256.93 20.275 ;
    RECT 256.72 20.565 256.93 20.635 ;
    RECT 256.72 20.925 256.93 20.995 ;
    RECT 256.26 20.205 256.47 20.275 ;
    RECT 256.26 20.565 256.47 20.635 ;
    RECT 256.26 20.925 256.47 20.995 ;
    RECT 253.4 20.205 253.61 20.275 ;
    RECT 253.4 20.565 253.61 20.635 ;
    RECT 253.4 20.925 253.61 20.995 ;
    RECT 252.94 20.205 253.15 20.275 ;
    RECT 252.94 20.565 253.15 20.635 ;
    RECT 252.94 20.925 253.15 20.995 ;
    RECT 250.08 20.205 250.29 20.275 ;
    RECT 250.08 20.565 250.29 20.635 ;
    RECT 250.08 20.925 250.29 20.995 ;
    RECT 249.62 20.205 249.83 20.275 ;
    RECT 249.62 20.565 249.83 20.635 ;
    RECT 249.62 20.925 249.83 20.995 ;
    RECT 246.76 20.205 246.97 20.275 ;
    RECT 246.76 20.565 246.97 20.635 ;
    RECT 246.76 20.925 246.97 20.995 ;
    RECT 246.3 20.205 246.51 20.275 ;
    RECT 246.3 20.565 246.51 20.635 ;
    RECT 246.3 20.925 246.51 20.995 ;
    RECT 243.44 20.205 243.65 20.275 ;
    RECT 243.44 20.565 243.65 20.635 ;
    RECT 243.44 20.925 243.65 20.995 ;
    RECT 242.98 20.205 243.19 20.275 ;
    RECT 242.98 20.565 243.19 20.635 ;
    RECT 242.98 20.925 243.19 20.995 ;
    RECT 240.12 20.205 240.33 20.275 ;
    RECT 240.12 20.565 240.33 20.635 ;
    RECT 240.12 20.925 240.33 20.995 ;
    RECT 239.66 20.205 239.87 20.275 ;
    RECT 239.66 20.565 239.87 20.635 ;
    RECT 239.66 20.925 239.87 20.995 ;
    RECT 236.8 20.205 237.01 20.275 ;
    RECT 236.8 20.565 237.01 20.635 ;
    RECT 236.8 20.925 237.01 20.995 ;
    RECT 236.34 20.205 236.55 20.275 ;
    RECT 236.34 20.565 236.55 20.635 ;
    RECT 236.34 20.925 236.55 20.995 ;
    RECT 374.15 20.565 374.22 20.635 ;
    RECT 333.08 20.205 333.29 20.275 ;
    RECT 333.08 20.565 333.29 20.635 ;
    RECT 333.08 20.925 333.29 20.995 ;
    RECT 332.62 20.205 332.83 20.275 ;
    RECT 332.62 20.565 332.83 20.635 ;
    RECT 332.62 20.925 332.83 20.995 ;
    RECT 329.76 20.205 329.97 20.275 ;
    RECT 329.76 20.565 329.97 20.635 ;
    RECT 329.76 20.925 329.97 20.995 ;
    RECT 329.3 20.205 329.51 20.275 ;
    RECT 329.3 20.565 329.51 20.635 ;
    RECT 329.3 20.925 329.51 20.995 ;
    RECT 326.44 20.205 326.65 20.275 ;
    RECT 326.44 20.565 326.65 20.635 ;
    RECT 326.44 20.925 326.65 20.995 ;
    RECT 325.98 20.205 326.19 20.275 ;
    RECT 325.98 20.565 326.19 20.635 ;
    RECT 325.98 20.925 326.19 20.995 ;
    RECT 323.12 20.205 323.33 20.275 ;
    RECT 323.12 20.565 323.33 20.635 ;
    RECT 323.12 20.925 323.33 20.995 ;
    RECT 322.66 20.205 322.87 20.275 ;
    RECT 322.66 20.565 322.87 20.635 ;
    RECT 322.66 20.925 322.87 20.995 ;
    RECT 319.8 20.205 320.01 20.275 ;
    RECT 319.8 20.565 320.01 20.635 ;
    RECT 319.8 20.925 320.01 20.995 ;
    RECT 319.34 20.205 319.55 20.275 ;
    RECT 319.34 20.565 319.55 20.635 ;
    RECT 319.34 20.925 319.55 20.995 ;
    RECT 316.48 20.205 316.69 20.275 ;
    RECT 316.48 20.565 316.69 20.635 ;
    RECT 316.48 20.925 316.69 20.995 ;
    RECT 316.02 20.205 316.23 20.275 ;
    RECT 316.02 20.565 316.23 20.635 ;
    RECT 316.02 20.925 316.23 20.995 ;
    RECT 313.16 20.205 313.37 20.275 ;
    RECT 313.16 20.565 313.37 20.635 ;
    RECT 313.16 20.925 313.37 20.995 ;
    RECT 312.7 20.205 312.91 20.275 ;
    RECT 312.7 20.565 312.91 20.635 ;
    RECT 312.7 20.925 312.91 20.995 ;
    RECT 309.84 20.205 310.05 20.275 ;
    RECT 309.84 20.565 310.05 20.635 ;
    RECT 309.84 20.925 310.05 20.995 ;
    RECT 309.38 20.205 309.59 20.275 ;
    RECT 309.38 20.565 309.59 20.635 ;
    RECT 309.38 20.925 309.59 20.995 ;
    RECT 306.52 20.205 306.73 20.275 ;
    RECT 306.52 20.565 306.73 20.635 ;
    RECT 306.52 20.925 306.73 20.995 ;
    RECT 306.06 20.205 306.27 20.275 ;
    RECT 306.06 20.565 306.27 20.635 ;
    RECT 306.06 20.925 306.27 20.995 ;
    RECT 303.2 33.885 303.41 33.955 ;
    RECT 303.2 34.245 303.41 34.315 ;
    RECT 303.2 34.605 303.41 34.675 ;
    RECT 302.74 33.885 302.95 33.955 ;
    RECT 302.74 34.245 302.95 34.315 ;
    RECT 302.74 34.605 302.95 34.675 ;
    RECT 200.605 34.245 200.675 34.315 ;
    RECT 372.92 33.885 373.13 33.955 ;
    RECT 372.92 34.245 373.13 34.315 ;
    RECT 372.92 34.605 373.13 34.675 ;
    RECT 372.46 33.885 372.67 33.955 ;
    RECT 372.46 34.245 372.67 34.315 ;
    RECT 372.46 34.605 372.67 34.675 ;
    RECT 369.6 33.885 369.81 33.955 ;
    RECT 369.6 34.245 369.81 34.315 ;
    RECT 369.6 34.605 369.81 34.675 ;
    RECT 369.14 33.885 369.35 33.955 ;
    RECT 369.14 34.245 369.35 34.315 ;
    RECT 369.14 34.605 369.35 34.675 ;
    RECT 299.88 33.885 300.09 33.955 ;
    RECT 299.88 34.245 300.09 34.315 ;
    RECT 299.88 34.605 300.09 34.675 ;
    RECT 299.42 33.885 299.63 33.955 ;
    RECT 299.42 34.245 299.63 34.315 ;
    RECT 299.42 34.605 299.63 34.675 ;
    RECT 296.56 33.885 296.77 33.955 ;
    RECT 296.56 34.245 296.77 34.315 ;
    RECT 296.56 34.605 296.77 34.675 ;
    RECT 296.1 33.885 296.31 33.955 ;
    RECT 296.1 34.245 296.31 34.315 ;
    RECT 296.1 34.605 296.31 34.675 ;
    RECT 293.24 33.885 293.45 33.955 ;
    RECT 293.24 34.245 293.45 34.315 ;
    RECT 293.24 34.605 293.45 34.675 ;
    RECT 292.78 33.885 292.99 33.955 ;
    RECT 292.78 34.245 292.99 34.315 ;
    RECT 292.78 34.605 292.99 34.675 ;
    RECT 289.92 33.885 290.13 33.955 ;
    RECT 289.92 34.245 290.13 34.315 ;
    RECT 289.92 34.605 290.13 34.675 ;
    RECT 289.46 33.885 289.67 33.955 ;
    RECT 289.46 34.245 289.67 34.315 ;
    RECT 289.46 34.605 289.67 34.675 ;
    RECT 286.6 33.885 286.81 33.955 ;
    RECT 286.6 34.245 286.81 34.315 ;
    RECT 286.6 34.605 286.81 34.675 ;
    RECT 286.14 33.885 286.35 33.955 ;
    RECT 286.14 34.245 286.35 34.315 ;
    RECT 286.14 34.605 286.35 34.675 ;
    RECT 283.28 33.885 283.49 33.955 ;
    RECT 283.28 34.245 283.49 34.315 ;
    RECT 283.28 34.605 283.49 34.675 ;
    RECT 282.82 33.885 283.03 33.955 ;
    RECT 282.82 34.245 283.03 34.315 ;
    RECT 282.82 34.605 283.03 34.675 ;
    RECT 279.96 33.885 280.17 33.955 ;
    RECT 279.96 34.245 280.17 34.315 ;
    RECT 279.96 34.605 280.17 34.675 ;
    RECT 279.5 33.885 279.71 33.955 ;
    RECT 279.5 34.245 279.71 34.315 ;
    RECT 279.5 34.605 279.71 34.675 ;
    RECT 276.64 33.885 276.85 33.955 ;
    RECT 276.64 34.245 276.85 34.315 ;
    RECT 276.64 34.605 276.85 34.675 ;
    RECT 276.18 33.885 276.39 33.955 ;
    RECT 276.18 34.245 276.39 34.315 ;
    RECT 276.18 34.605 276.39 34.675 ;
    RECT 273.32 33.885 273.53 33.955 ;
    RECT 273.32 34.245 273.53 34.315 ;
    RECT 273.32 34.605 273.53 34.675 ;
    RECT 272.86 33.885 273.07 33.955 ;
    RECT 272.86 34.245 273.07 34.315 ;
    RECT 272.86 34.605 273.07 34.675 ;
    RECT 270.0 33.885 270.21 33.955 ;
    RECT 270.0 34.245 270.21 34.315 ;
    RECT 270.0 34.605 270.21 34.675 ;
    RECT 269.54 33.885 269.75 33.955 ;
    RECT 269.54 34.245 269.75 34.315 ;
    RECT 269.54 34.605 269.75 34.675 ;
    RECT 233.48 33.885 233.69 33.955 ;
    RECT 233.48 34.245 233.69 34.315 ;
    RECT 233.48 34.605 233.69 34.675 ;
    RECT 233.02 33.885 233.23 33.955 ;
    RECT 233.02 34.245 233.23 34.315 ;
    RECT 233.02 34.605 233.23 34.675 ;
    RECT 230.16 33.885 230.37 33.955 ;
    RECT 230.16 34.245 230.37 34.315 ;
    RECT 230.16 34.605 230.37 34.675 ;
    RECT 229.7 33.885 229.91 33.955 ;
    RECT 229.7 34.245 229.91 34.315 ;
    RECT 229.7 34.605 229.91 34.675 ;
    RECT 366.28 33.885 366.49 33.955 ;
    RECT 366.28 34.245 366.49 34.315 ;
    RECT 366.28 34.605 366.49 34.675 ;
    RECT 365.82 33.885 366.03 33.955 ;
    RECT 365.82 34.245 366.03 34.315 ;
    RECT 365.82 34.605 366.03 34.675 ;
    RECT 226.84 33.885 227.05 33.955 ;
    RECT 226.84 34.245 227.05 34.315 ;
    RECT 226.84 34.605 227.05 34.675 ;
    RECT 226.38 33.885 226.59 33.955 ;
    RECT 226.38 34.245 226.59 34.315 ;
    RECT 226.38 34.605 226.59 34.675 ;
    RECT 362.96 33.885 363.17 33.955 ;
    RECT 362.96 34.245 363.17 34.315 ;
    RECT 362.96 34.605 363.17 34.675 ;
    RECT 362.5 33.885 362.71 33.955 ;
    RECT 362.5 34.245 362.71 34.315 ;
    RECT 362.5 34.605 362.71 34.675 ;
    RECT 223.52 33.885 223.73 33.955 ;
    RECT 223.52 34.245 223.73 34.315 ;
    RECT 223.52 34.605 223.73 34.675 ;
    RECT 223.06 33.885 223.27 33.955 ;
    RECT 223.06 34.245 223.27 34.315 ;
    RECT 223.06 34.605 223.27 34.675 ;
    RECT 359.64 33.885 359.85 33.955 ;
    RECT 359.64 34.245 359.85 34.315 ;
    RECT 359.64 34.605 359.85 34.675 ;
    RECT 359.18 33.885 359.39 33.955 ;
    RECT 359.18 34.245 359.39 34.315 ;
    RECT 359.18 34.605 359.39 34.675 ;
    RECT 220.2 33.885 220.41 33.955 ;
    RECT 220.2 34.245 220.41 34.315 ;
    RECT 220.2 34.605 220.41 34.675 ;
    RECT 219.74 33.885 219.95 33.955 ;
    RECT 219.74 34.245 219.95 34.315 ;
    RECT 219.74 34.605 219.95 34.675 ;
    RECT 356.32 33.885 356.53 33.955 ;
    RECT 356.32 34.245 356.53 34.315 ;
    RECT 356.32 34.605 356.53 34.675 ;
    RECT 355.86 33.885 356.07 33.955 ;
    RECT 355.86 34.245 356.07 34.315 ;
    RECT 355.86 34.605 356.07 34.675 ;
    RECT 353.0 33.885 353.21 33.955 ;
    RECT 353.0 34.245 353.21 34.315 ;
    RECT 353.0 34.605 353.21 34.675 ;
    RECT 352.54 33.885 352.75 33.955 ;
    RECT 352.54 34.245 352.75 34.315 ;
    RECT 352.54 34.605 352.75 34.675 ;
    RECT 216.88 33.885 217.09 33.955 ;
    RECT 216.88 34.245 217.09 34.315 ;
    RECT 216.88 34.605 217.09 34.675 ;
    RECT 216.42 33.885 216.63 33.955 ;
    RECT 216.42 34.245 216.63 34.315 ;
    RECT 216.42 34.605 216.63 34.675 ;
    RECT 349.68 33.885 349.89 33.955 ;
    RECT 349.68 34.245 349.89 34.315 ;
    RECT 349.68 34.605 349.89 34.675 ;
    RECT 349.22 33.885 349.43 33.955 ;
    RECT 349.22 34.245 349.43 34.315 ;
    RECT 349.22 34.605 349.43 34.675 ;
    RECT 213.56 33.885 213.77 33.955 ;
    RECT 213.56 34.245 213.77 34.315 ;
    RECT 213.56 34.605 213.77 34.675 ;
    RECT 213.1 33.885 213.31 33.955 ;
    RECT 213.1 34.245 213.31 34.315 ;
    RECT 213.1 34.605 213.31 34.675 ;
    RECT 346.36 33.885 346.57 33.955 ;
    RECT 346.36 34.245 346.57 34.315 ;
    RECT 346.36 34.605 346.57 34.675 ;
    RECT 345.9 33.885 346.11 33.955 ;
    RECT 345.9 34.245 346.11 34.315 ;
    RECT 345.9 34.605 346.11 34.675 ;
    RECT 210.24 33.885 210.45 33.955 ;
    RECT 210.24 34.245 210.45 34.315 ;
    RECT 210.24 34.605 210.45 34.675 ;
    RECT 209.78 33.885 209.99 33.955 ;
    RECT 209.78 34.245 209.99 34.315 ;
    RECT 209.78 34.605 209.99 34.675 ;
    RECT 343.04 33.885 343.25 33.955 ;
    RECT 343.04 34.245 343.25 34.315 ;
    RECT 343.04 34.605 343.25 34.675 ;
    RECT 342.58 33.885 342.79 33.955 ;
    RECT 342.58 34.245 342.79 34.315 ;
    RECT 342.58 34.605 342.79 34.675 ;
    RECT 206.92 33.885 207.13 33.955 ;
    RECT 206.92 34.245 207.13 34.315 ;
    RECT 206.92 34.605 207.13 34.675 ;
    RECT 206.46 33.885 206.67 33.955 ;
    RECT 206.46 34.245 206.67 34.315 ;
    RECT 206.46 34.605 206.67 34.675 ;
    RECT 339.72 33.885 339.93 33.955 ;
    RECT 339.72 34.245 339.93 34.315 ;
    RECT 339.72 34.605 339.93 34.675 ;
    RECT 339.26 33.885 339.47 33.955 ;
    RECT 339.26 34.245 339.47 34.315 ;
    RECT 339.26 34.605 339.47 34.675 ;
    RECT 203.6 33.885 203.81 33.955 ;
    RECT 203.6 34.245 203.81 34.315 ;
    RECT 203.6 34.605 203.81 34.675 ;
    RECT 203.14 33.885 203.35 33.955 ;
    RECT 203.14 34.245 203.35 34.315 ;
    RECT 203.14 34.605 203.35 34.675 ;
    RECT 336.4 33.885 336.61 33.955 ;
    RECT 336.4 34.245 336.61 34.315 ;
    RECT 336.4 34.605 336.61 34.675 ;
    RECT 335.94 33.885 336.15 33.955 ;
    RECT 335.94 34.245 336.15 34.315 ;
    RECT 335.94 34.605 336.15 34.675 ;
    RECT 266.68 33.885 266.89 33.955 ;
    RECT 266.68 34.245 266.89 34.315 ;
    RECT 266.68 34.605 266.89 34.675 ;
    RECT 266.22 33.885 266.43 33.955 ;
    RECT 266.22 34.245 266.43 34.315 ;
    RECT 266.22 34.605 266.43 34.675 ;
    RECT 263.36 33.885 263.57 33.955 ;
    RECT 263.36 34.245 263.57 34.315 ;
    RECT 263.36 34.605 263.57 34.675 ;
    RECT 262.9 33.885 263.11 33.955 ;
    RECT 262.9 34.245 263.11 34.315 ;
    RECT 262.9 34.605 263.11 34.675 ;
    RECT 260.04 33.885 260.25 33.955 ;
    RECT 260.04 34.245 260.25 34.315 ;
    RECT 260.04 34.605 260.25 34.675 ;
    RECT 259.58 33.885 259.79 33.955 ;
    RECT 259.58 34.245 259.79 34.315 ;
    RECT 259.58 34.605 259.79 34.675 ;
    RECT 256.72 33.885 256.93 33.955 ;
    RECT 256.72 34.245 256.93 34.315 ;
    RECT 256.72 34.605 256.93 34.675 ;
    RECT 256.26 33.885 256.47 33.955 ;
    RECT 256.26 34.245 256.47 34.315 ;
    RECT 256.26 34.605 256.47 34.675 ;
    RECT 253.4 33.885 253.61 33.955 ;
    RECT 253.4 34.245 253.61 34.315 ;
    RECT 253.4 34.605 253.61 34.675 ;
    RECT 252.94 33.885 253.15 33.955 ;
    RECT 252.94 34.245 253.15 34.315 ;
    RECT 252.94 34.605 253.15 34.675 ;
    RECT 250.08 33.885 250.29 33.955 ;
    RECT 250.08 34.245 250.29 34.315 ;
    RECT 250.08 34.605 250.29 34.675 ;
    RECT 249.62 33.885 249.83 33.955 ;
    RECT 249.62 34.245 249.83 34.315 ;
    RECT 249.62 34.605 249.83 34.675 ;
    RECT 246.76 33.885 246.97 33.955 ;
    RECT 246.76 34.245 246.97 34.315 ;
    RECT 246.76 34.605 246.97 34.675 ;
    RECT 246.3 33.885 246.51 33.955 ;
    RECT 246.3 34.245 246.51 34.315 ;
    RECT 246.3 34.605 246.51 34.675 ;
    RECT 243.44 33.885 243.65 33.955 ;
    RECT 243.44 34.245 243.65 34.315 ;
    RECT 243.44 34.605 243.65 34.675 ;
    RECT 242.98 33.885 243.19 33.955 ;
    RECT 242.98 34.245 243.19 34.315 ;
    RECT 242.98 34.605 243.19 34.675 ;
    RECT 240.12 33.885 240.33 33.955 ;
    RECT 240.12 34.245 240.33 34.315 ;
    RECT 240.12 34.605 240.33 34.675 ;
    RECT 239.66 33.885 239.87 33.955 ;
    RECT 239.66 34.245 239.87 34.315 ;
    RECT 239.66 34.605 239.87 34.675 ;
    RECT 236.8 33.885 237.01 33.955 ;
    RECT 236.8 34.245 237.01 34.315 ;
    RECT 236.8 34.605 237.01 34.675 ;
    RECT 236.34 33.885 236.55 33.955 ;
    RECT 236.34 34.245 236.55 34.315 ;
    RECT 236.34 34.605 236.55 34.675 ;
    RECT 374.15 34.245 374.22 34.315 ;
    RECT 333.08 33.885 333.29 33.955 ;
    RECT 333.08 34.245 333.29 34.315 ;
    RECT 333.08 34.605 333.29 34.675 ;
    RECT 332.62 33.885 332.83 33.955 ;
    RECT 332.62 34.245 332.83 34.315 ;
    RECT 332.62 34.605 332.83 34.675 ;
    RECT 329.76 33.885 329.97 33.955 ;
    RECT 329.76 34.245 329.97 34.315 ;
    RECT 329.76 34.605 329.97 34.675 ;
    RECT 329.3 33.885 329.51 33.955 ;
    RECT 329.3 34.245 329.51 34.315 ;
    RECT 329.3 34.605 329.51 34.675 ;
    RECT 326.44 33.885 326.65 33.955 ;
    RECT 326.44 34.245 326.65 34.315 ;
    RECT 326.44 34.605 326.65 34.675 ;
    RECT 325.98 33.885 326.19 33.955 ;
    RECT 325.98 34.245 326.19 34.315 ;
    RECT 325.98 34.605 326.19 34.675 ;
    RECT 323.12 33.885 323.33 33.955 ;
    RECT 323.12 34.245 323.33 34.315 ;
    RECT 323.12 34.605 323.33 34.675 ;
    RECT 322.66 33.885 322.87 33.955 ;
    RECT 322.66 34.245 322.87 34.315 ;
    RECT 322.66 34.605 322.87 34.675 ;
    RECT 319.8 33.885 320.01 33.955 ;
    RECT 319.8 34.245 320.01 34.315 ;
    RECT 319.8 34.605 320.01 34.675 ;
    RECT 319.34 33.885 319.55 33.955 ;
    RECT 319.34 34.245 319.55 34.315 ;
    RECT 319.34 34.605 319.55 34.675 ;
    RECT 316.48 33.885 316.69 33.955 ;
    RECT 316.48 34.245 316.69 34.315 ;
    RECT 316.48 34.605 316.69 34.675 ;
    RECT 316.02 33.885 316.23 33.955 ;
    RECT 316.02 34.245 316.23 34.315 ;
    RECT 316.02 34.605 316.23 34.675 ;
    RECT 313.16 33.885 313.37 33.955 ;
    RECT 313.16 34.245 313.37 34.315 ;
    RECT 313.16 34.605 313.37 34.675 ;
    RECT 312.7 33.885 312.91 33.955 ;
    RECT 312.7 34.245 312.91 34.315 ;
    RECT 312.7 34.605 312.91 34.675 ;
    RECT 309.84 33.885 310.05 33.955 ;
    RECT 309.84 34.245 310.05 34.315 ;
    RECT 309.84 34.605 310.05 34.675 ;
    RECT 309.38 33.885 309.59 33.955 ;
    RECT 309.38 34.245 309.59 34.315 ;
    RECT 309.38 34.605 309.59 34.675 ;
    RECT 306.52 33.885 306.73 33.955 ;
    RECT 306.52 34.245 306.73 34.315 ;
    RECT 306.52 34.605 306.73 34.675 ;
    RECT 306.06 33.885 306.27 33.955 ;
    RECT 306.06 34.245 306.27 34.315 ;
    RECT 306.06 34.605 306.27 34.675 ;
    RECT 303.2 19.485 303.41 19.555 ;
    RECT 303.2 19.845 303.41 19.915 ;
    RECT 303.2 20.205 303.41 20.275 ;
    RECT 302.74 19.485 302.95 19.555 ;
    RECT 302.74 19.845 302.95 19.915 ;
    RECT 302.74 20.205 302.95 20.275 ;
    RECT 372.92 19.485 373.13 19.555 ;
    RECT 372.92 19.845 373.13 19.915 ;
    RECT 372.92 20.205 373.13 20.275 ;
    RECT 372.46 19.485 372.67 19.555 ;
    RECT 372.46 19.845 372.67 19.915 ;
    RECT 372.46 20.205 372.67 20.275 ;
    RECT 369.6 19.485 369.81 19.555 ;
    RECT 369.6 19.845 369.81 19.915 ;
    RECT 369.6 20.205 369.81 20.275 ;
    RECT 369.14 19.485 369.35 19.555 ;
    RECT 369.14 19.845 369.35 19.915 ;
    RECT 369.14 20.205 369.35 20.275 ;
    RECT 200.605 19.845 200.675 19.915 ;
    RECT 299.88 19.485 300.09 19.555 ;
    RECT 299.88 19.845 300.09 19.915 ;
    RECT 299.88 20.205 300.09 20.275 ;
    RECT 299.42 19.485 299.63 19.555 ;
    RECT 299.42 19.845 299.63 19.915 ;
    RECT 299.42 20.205 299.63 20.275 ;
    RECT 296.56 19.485 296.77 19.555 ;
    RECT 296.56 19.845 296.77 19.915 ;
    RECT 296.56 20.205 296.77 20.275 ;
    RECT 296.1 19.485 296.31 19.555 ;
    RECT 296.1 19.845 296.31 19.915 ;
    RECT 296.1 20.205 296.31 20.275 ;
    RECT 293.24 19.485 293.45 19.555 ;
    RECT 293.24 19.845 293.45 19.915 ;
    RECT 293.24 20.205 293.45 20.275 ;
    RECT 292.78 19.485 292.99 19.555 ;
    RECT 292.78 19.845 292.99 19.915 ;
    RECT 292.78 20.205 292.99 20.275 ;
    RECT 289.92 19.485 290.13 19.555 ;
    RECT 289.92 19.845 290.13 19.915 ;
    RECT 289.92 20.205 290.13 20.275 ;
    RECT 289.46 19.485 289.67 19.555 ;
    RECT 289.46 19.845 289.67 19.915 ;
    RECT 289.46 20.205 289.67 20.275 ;
    RECT 286.6 19.485 286.81 19.555 ;
    RECT 286.6 19.845 286.81 19.915 ;
    RECT 286.6 20.205 286.81 20.275 ;
    RECT 286.14 19.485 286.35 19.555 ;
    RECT 286.14 19.845 286.35 19.915 ;
    RECT 286.14 20.205 286.35 20.275 ;
    RECT 283.28 19.485 283.49 19.555 ;
    RECT 283.28 19.845 283.49 19.915 ;
    RECT 283.28 20.205 283.49 20.275 ;
    RECT 282.82 19.485 283.03 19.555 ;
    RECT 282.82 19.845 283.03 19.915 ;
    RECT 282.82 20.205 283.03 20.275 ;
    RECT 279.96 19.485 280.17 19.555 ;
    RECT 279.96 19.845 280.17 19.915 ;
    RECT 279.96 20.205 280.17 20.275 ;
    RECT 279.5 19.485 279.71 19.555 ;
    RECT 279.5 19.845 279.71 19.915 ;
    RECT 279.5 20.205 279.71 20.275 ;
    RECT 276.64 19.485 276.85 19.555 ;
    RECT 276.64 19.845 276.85 19.915 ;
    RECT 276.64 20.205 276.85 20.275 ;
    RECT 276.18 19.485 276.39 19.555 ;
    RECT 276.18 19.845 276.39 19.915 ;
    RECT 276.18 20.205 276.39 20.275 ;
    RECT 273.32 19.485 273.53 19.555 ;
    RECT 273.32 19.845 273.53 19.915 ;
    RECT 273.32 20.205 273.53 20.275 ;
    RECT 272.86 19.485 273.07 19.555 ;
    RECT 272.86 19.845 273.07 19.915 ;
    RECT 272.86 20.205 273.07 20.275 ;
    RECT 270.0 19.485 270.21 19.555 ;
    RECT 270.0 19.845 270.21 19.915 ;
    RECT 270.0 20.205 270.21 20.275 ;
    RECT 269.54 19.485 269.75 19.555 ;
    RECT 269.54 19.845 269.75 19.915 ;
    RECT 269.54 20.205 269.75 20.275 ;
    RECT 233.48 19.485 233.69 19.555 ;
    RECT 233.48 19.845 233.69 19.915 ;
    RECT 233.48 20.205 233.69 20.275 ;
    RECT 233.02 19.485 233.23 19.555 ;
    RECT 233.02 19.845 233.23 19.915 ;
    RECT 233.02 20.205 233.23 20.275 ;
    RECT 230.16 19.485 230.37 19.555 ;
    RECT 230.16 19.845 230.37 19.915 ;
    RECT 230.16 20.205 230.37 20.275 ;
    RECT 229.7 19.485 229.91 19.555 ;
    RECT 229.7 19.845 229.91 19.915 ;
    RECT 229.7 20.205 229.91 20.275 ;
    RECT 366.28 19.485 366.49 19.555 ;
    RECT 366.28 19.845 366.49 19.915 ;
    RECT 366.28 20.205 366.49 20.275 ;
    RECT 365.82 19.485 366.03 19.555 ;
    RECT 365.82 19.845 366.03 19.915 ;
    RECT 365.82 20.205 366.03 20.275 ;
    RECT 226.84 19.485 227.05 19.555 ;
    RECT 226.84 19.845 227.05 19.915 ;
    RECT 226.84 20.205 227.05 20.275 ;
    RECT 226.38 19.485 226.59 19.555 ;
    RECT 226.38 19.845 226.59 19.915 ;
    RECT 226.38 20.205 226.59 20.275 ;
    RECT 362.96 19.485 363.17 19.555 ;
    RECT 362.96 19.845 363.17 19.915 ;
    RECT 362.96 20.205 363.17 20.275 ;
    RECT 362.5 19.485 362.71 19.555 ;
    RECT 362.5 19.845 362.71 19.915 ;
    RECT 362.5 20.205 362.71 20.275 ;
    RECT 223.52 19.485 223.73 19.555 ;
    RECT 223.52 19.845 223.73 19.915 ;
    RECT 223.52 20.205 223.73 20.275 ;
    RECT 223.06 19.485 223.27 19.555 ;
    RECT 223.06 19.845 223.27 19.915 ;
    RECT 223.06 20.205 223.27 20.275 ;
    RECT 359.64 19.485 359.85 19.555 ;
    RECT 359.64 19.845 359.85 19.915 ;
    RECT 359.64 20.205 359.85 20.275 ;
    RECT 359.18 19.485 359.39 19.555 ;
    RECT 359.18 19.845 359.39 19.915 ;
    RECT 359.18 20.205 359.39 20.275 ;
    RECT 220.2 19.485 220.41 19.555 ;
    RECT 220.2 19.845 220.41 19.915 ;
    RECT 220.2 20.205 220.41 20.275 ;
    RECT 219.74 19.485 219.95 19.555 ;
    RECT 219.74 19.845 219.95 19.915 ;
    RECT 219.74 20.205 219.95 20.275 ;
    RECT 356.32 19.485 356.53 19.555 ;
    RECT 356.32 19.845 356.53 19.915 ;
    RECT 356.32 20.205 356.53 20.275 ;
    RECT 355.86 19.485 356.07 19.555 ;
    RECT 355.86 19.845 356.07 19.915 ;
    RECT 355.86 20.205 356.07 20.275 ;
    RECT 353.0 19.485 353.21 19.555 ;
    RECT 353.0 19.845 353.21 19.915 ;
    RECT 353.0 20.205 353.21 20.275 ;
    RECT 352.54 19.485 352.75 19.555 ;
    RECT 352.54 19.845 352.75 19.915 ;
    RECT 352.54 20.205 352.75 20.275 ;
    RECT 216.88 19.485 217.09 19.555 ;
    RECT 216.88 19.845 217.09 19.915 ;
    RECT 216.88 20.205 217.09 20.275 ;
    RECT 216.42 19.485 216.63 19.555 ;
    RECT 216.42 19.845 216.63 19.915 ;
    RECT 216.42 20.205 216.63 20.275 ;
    RECT 349.68 19.485 349.89 19.555 ;
    RECT 349.68 19.845 349.89 19.915 ;
    RECT 349.68 20.205 349.89 20.275 ;
    RECT 349.22 19.485 349.43 19.555 ;
    RECT 349.22 19.845 349.43 19.915 ;
    RECT 349.22 20.205 349.43 20.275 ;
    RECT 213.56 19.485 213.77 19.555 ;
    RECT 213.56 19.845 213.77 19.915 ;
    RECT 213.56 20.205 213.77 20.275 ;
    RECT 213.1 19.485 213.31 19.555 ;
    RECT 213.1 19.845 213.31 19.915 ;
    RECT 213.1 20.205 213.31 20.275 ;
    RECT 346.36 19.485 346.57 19.555 ;
    RECT 346.36 19.845 346.57 19.915 ;
    RECT 346.36 20.205 346.57 20.275 ;
    RECT 345.9 19.485 346.11 19.555 ;
    RECT 345.9 19.845 346.11 19.915 ;
    RECT 345.9 20.205 346.11 20.275 ;
    RECT 210.24 19.485 210.45 19.555 ;
    RECT 210.24 19.845 210.45 19.915 ;
    RECT 210.24 20.205 210.45 20.275 ;
    RECT 209.78 19.485 209.99 19.555 ;
    RECT 209.78 19.845 209.99 19.915 ;
    RECT 209.78 20.205 209.99 20.275 ;
    RECT 343.04 19.485 343.25 19.555 ;
    RECT 343.04 19.845 343.25 19.915 ;
    RECT 343.04 20.205 343.25 20.275 ;
    RECT 342.58 19.485 342.79 19.555 ;
    RECT 342.58 19.845 342.79 19.915 ;
    RECT 342.58 20.205 342.79 20.275 ;
    RECT 206.92 19.485 207.13 19.555 ;
    RECT 206.92 19.845 207.13 19.915 ;
    RECT 206.92 20.205 207.13 20.275 ;
    RECT 206.46 19.485 206.67 19.555 ;
    RECT 206.46 19.845 206.67 19.915 ;
    RECT 206.46 20.205 206.67 20.275 ;
    RECT 339.72 19.485 339.93 19.555 ;
    RECT 339.72 19.845 339.93 19.915 ;
    RECT 339.72 20.205 339.93 20.275 ;
    RECT 339.26 19.485 339.47 19.555 ;
    RECT 339.26 19.845 339.47 19.915 ;
    RECT 339.26 20.205 339.47 20.275 ;
    RECT 203.6 19.485 203.81 19.555 ;
    RECT 203.6 19.845 203.81 19.915 ;
    RECT 203.6 20.205 203.81 20.275 ;
    RECT 203.14 19.485 203.35 19.555 ;
    RECT 203.14 19.845 203.35 19.915 ;
    RECT 203.14 20.205 203.35 20.275 ;
    RECT 336.4 19.485 336.61 19.555 ;
    RECT 336.4 19.845 336.61 19.915 ;
    RECT 336.4 20.205 336.61 20.275 ;
    RECT 335.94 19.485 336.15 19.555 ;
    RECT 335.94 19.845 336.15 19.915 ;
    RECT 335.94 20.205 336.15 20.275 ;
    RECT 266.68 19.485 266.89 19.555 ;
    RECT 266.68 19.845 266.89 19.915 ;
    RECT 266.68 20.205 266.89 20.275 ;
    RECT 266.22 19.485 266.43 19.555 ;
    RECT 266.22 19.845 266.43 19.915 ;
    RECT 266.22 20.205 266.43 20.275 ;
    RECT 263.36 19.485 263.57 19.555 ;
    RECT 263.36 19.845 263.57 19.915 ;
    RECT 263.36 20.205 263.57 20.275 ;
    RECT 262.9 19.485 263.11 19.555 ;
    RECT 262.9 19.845 263.11 19.915 ;
    RECT 262.9 20.205 263.11 20.275 ;
    RECT 260.04 19.485 260.25 19.555 ;
    RECT 260.04 19.845 260.25 19.915 ;
    RECT 260.04 20.205 260.25 20.275 ;
    RECT 259.58 19.485 259.79 19.555 ;
    RECT 259.58 19.845 259.79 19.915 ;
    RECT 259.58 20.205 259.79 20.275 ;
    RECT 256.72 19.485 256.93 19.555 ;
    RECT 256.72 19.845 256.93 19.915 ;
    RECT 256.72 20.205 256.93 20.275 ;
    RECT 256.26 19.485 256.47 19.555 ;
    RECT 256.26 19.845 256.47 19.915 ;
    RECT 256.26 20.205 256.47 20.275 ;
    RECT 253.4 19.485 253.61 19.555 ;
    RECT 253.4 19.845 253.61 19.915 ;
    RECT 253.4 20.205 253.61 20.275 ;
    RECT 252.94 19.485 253.15 19.555 ;
    RECT 252.94 19.845 253.15 19.915 ;
    RECT 252.94 20.205 253.15 20.275 ;
    RECT 250.08 19.485 250.29 19.555 ;
    RECT 250.08 19.845 250.29 19.915 ;
    RECT 250.08 20.205 250.29 20.275 ;
    RECT 249.62 19.485 249.83 19.555 ;
    RECT 249.62 19.845 249.83 19.915 ;
    RECT 249.62 20.205 249.83 20.275 ;
    RECT 246.76 19.485 246.97 19.555 ;
    RECT 246.76 19.845 246.97 19.915 ;
    RECT 246.76 20.205 246.97 20.275 ;
    RECT 246.3 19.485 246.51 19.555 ;
    RECT 246.3 19.845 246.51 19.915 ;
    RECT 246.3 20.205 246.51 20.275 ;
    RECT 243.44 19.485 243.65 19.555 ;
    RECT 243.44 19.845 243.65 19.915 ;
    RECT 243.44 20.205 243.65 20.275 ;
    RECT 242.98 19.485 243.19 19.555 ;
    RECT 242.98 19.845 243.19 19.915 ;
    RECT 242.98 20.205 243.19 20.275 ;
    RECT 240.12 19.485 240.33 19.555 ;
    RECT 240.12 19.845 240.33 19.915 ;
    RECT 240.12 20.205 240.33 20.275 ;
    RECT 239.66 19.485 239.87 19.555 ;
    RECT 239.66 19.845 239.87 19.915 ;
    RECT 239.66 20.205 239.87 20.275 ;
    RECT 236.8 19.485 237.01 19.555 ;
    RECT 236.8 19.845 237.01 19.915 ;
    RECT 236.8 20.205 237.01 20.275 ;
    RECT 236.34 19.485 236.55 19.555 ;
    RECT 236.34 19.845 236.55 19.915 ;
    RECT 236.34 20.205 236.55 20.275 ;
    RECT 374.15 19.845 374.22 19.915 ;
    RECT 333.08 19.485 333.29 19.555 ;
    RECT 333.08 19.845 333.29 19.915 ;
    RECT 333.08 20.205 333.29 20.275 ;
    RECT 332.62 19.485 332.83 19.555 ;
    RECT 332.62 19.845 332.83 19.915 ;
    RECT 332.62 20.205 332.83 20.275 ;
    RECT 329.76 19.485 329.97 19.555 ;
    RECT 329.76 19.845 329.97 19.915 ;
    RECT 329.76 20.205 329.97 20.275 ;
    RECT 329.3 19.485 329.51 19.555 ;
    RECT 329.3 19.845 329.51 19.915 ;
    RECT 329.3 20.205 329.51 20.275 ;
    RECT 326.44 19.485 326.65 19.555 ;
    RECT 326.44 19.845 326.65 19.915 ;
    RECT 326.44 20.205 326.65 20.275 ;
    RECT 325.98 19.485 326.19 19.555 ;
    RECT 325.98 19.845 326.19 19.915 ;
    RECT 325.98 20.205 326.19 20.275 ;
    RECT 323.12 19.485 323.33 19.555 ;
    RECT 323.12 19.845 323.33 19.915 ;
    RECT 323.12 20.205 323.33 20.275 ;
    RECT 322.66 19.485 322.87 19.555 ;
    RECT 322.66 19.845 322.87 19.915 ;
    RECT 322.66 20.205 322.87 20.275 ;
    RECT 319.8 19.485 320.01 19.555 ;
    RECT 319.8 19.845 320.01 19.915 ;
    RECT 319.8 20.205 320.01 20.275 ;
    RECT 319.34 19.485 319.55 19.555 ;
    RECT 319.34 19.845 319.55 19.915 ;
    RECT 319.34 20.205 319.55 20.275 ;
    RECT 316.48 19.485 316.69 19.555 ;
    RECT 316.48 19.845 316.69 19.915 ;
    RECT 316.48 20.205 316.69 20.275 ;
    RECT 316.02 19.485 316.23 19.555 ;
    RECT 316.02 19.845 316.23 19.915 ;
    RECT 316.02 20.205 316.23 20.275 ;
    RECT 313.16 19.485 313.37 19.555 ;
    RECT 313.16 19.845 313.37 19.915 ;
    RECT 313.16 20.205 313.37 20.275 ;
    RECT 312.7 19.485 312.91 19.555 ;
    RECT 312.7 19.845 312.91 19.915 ;
    RECT 312.7 20.205 312.91 20.275 ;
    RECT 309.84 19.485 310.05 19.555 ;
    RECT 309.84 19.845 310.05 19.915 ;
    RECT 309.84 20.205 310.05 20.275 ;
    RECT 309.38 19.485 309.59 19.555 ;
    RECT 309.38 19.845 309.59 19.915 ;
    RECT 309.38 20.205 309.59 20.275 ;
    RECT 306.52 19.485 306.73 19.555 ;
    RECT 306.52 19.845 306.73 19.915 ;
    RECT 306.52 20.205 306.73 20.275 ;
    RECT 306.06 19.485 306.27 19.555 ;
    RECT 306.06 19.845 306.27 19.915 ;
    RECT 306.06 20.205 306.27 20.275 ;
    RECT 303.2 18.765 303.41 18.835 ;
    RECT 303.2 19.125 303.41 19.195 ;
    RECT 303.2 19.485 303.41 19.555 ;
    RECT 302.74 18.765 302.95 18.835 ;
    RECT 302.74 19.125 302.95 19.195 ;
    RECT 302.74 19.485 302.95 19.555 ;
    RECT 372.92 18.765 373.13 18.835 ;
    RECT 372.92 19.125 373.13 19.195 ;
    RECT 372.92 19.485 373.13 19.555 ;
    RECT 372.46 18.765 372.67 18.835 ;
    RECT 372.46 19.125 372.67 19.195 ;
    RECT 372.46 19.485 372.67 19.555 ;
    RECT 369.6 18.765 369.81 18.835 ;
    RECT 369.6 19.125 369.81 19.195 ;
    RECT 369.6 19.485 369.81 19.555 ;
    RECT 369.14 18.765 369.35 18.835 ;
    RECT 369.14 19.125 369.35 19.195 ;
    RECT 369.14 19.485 369.35 19.555 ;
    RECT 200.605 19.125 200.675 19.195 ;
    RECT 299.88 18.765 300.09 18.835 ;
    RECT 299.88 19.125 300.09 19.195 ;
    RECT 299.88 19.485 300.09 19.555 ;
    RECT 299.42 18.765 299.63 18.835 ;
    RECT 299.42 19.125 299.63 19.195 ;
    RECT 299.42 19.485 299.63 19.555 ;
    RECT 296.56 18.765 296.77 18.835 ;
    RECT 296.56 19.125 296.77 19.195 ;
    RECT 296.56 19.485 296.77 19.555 ;
    RECT 296.1 18.765 296.31 18.835 ;
    RECT 296.1 19.125 296.31 19.195 ;
    RECT 296.1 19.485 296.31 19.555 ;
    RECT 293.24 18.765 293.45 18.835 ;
    RECT 293.24 19.125 293.45 19.195 ;
    RECT 293.24 19.485 293.45 19.555 ;
    RECT 292.78 18.765 292.99 18.835 ;
    RECT 292.78 19.125 292.99 19.195 ;
    RECT 292.78 19.485 292.99 19.555 ;
    RECT 289.92 18.765 290.13 18.835 ;
    RECT 289.92 19.125 290.13 19.195 ;
    RECT 289.92 19.485 290.13 19.555 ;
    RECT 289.46 18.765 289.67 18.835 ;
    RECT 289.46 19.125 289.67 19.195 ;
    RECT 289.46 19.485 289.67 19.555 ;
    RECT 286.6 18.765 286.81 18.835 ;
    RECT 286.6 19.125 286.81 19.195 ;
    RECT 286.6 19.485 286.81 19.555 ;
    RECT 286.14 18.765 286.35 18.835 ;
    RECT 286.14 19.125 286.35 19.195 ;
    RECT 286.14 19.485 286.35 19.555 ;
    RECT 283.28 18.765 283.49 18.835 ;
    RECT 283.28 19.125 283.49 19.195 ;
    RECT 283.28 19.485 283.49 19.555 ;
    RECT 282.82 18.765 283.03 18.835 ;
    RECT 282.82 19.125 283.03 19.195 ;
    RECT 282.82 19.485 283.03 19.555 ;
    RECT 279.96 18.765 280.17 18.835 ;
    RECT 279.96 19.125 280.17 19.195 ;
    RECT 279.96 19.485 280.17 19.555 ;
    RECT 279.5 18.765 279.71 18.835 ;
    RECT 279.5 19.125 279.71 19.195 ;
    RECT 279.5 19.485 279.71 19.555 ;
    RECT 276.64 18.765 276.85 18.835 ;
    RECT 276.64 19.125 276.85 19.195 ;
    RECT 276.64 19.485 276.85 19.555 ;
    RECT 276.18 18.765 276.39 18.835 ;
    RECT 276.18 19.125 276.39 19.195 ;
    RECT 276.18 19.485 276.39 19.555 ;
    RECT 273.32 18.765 273.53 18.835 ;
    RECT 273.32 19.125 273.53 19.195 ;
    RECT 273.32 19.485 273.53 19.555 ;
    RECT 272.86 18.765 273.07 18.835 ;
    RECT 272.86 19.125 273.07 19.195 ;
    RECT 272.86 19.485 273.07 19.555 ;
    RECT 270.0 18.765 270.21 18.835 ;
    RECT 270.0 19.125 270.21 19.195 ;
    RECT 270.0 19.485 270.21 19.555 ;
    RECT 269.54 18.765 269.75 18.835 ;
    RECT 269.54 19.125 269.75 19.195 ;
    RECT 269.54 19.485 269.75 19.555 ;
    RECT 233.48 18.765 233.69 18.835 ;
    RECT 233.48 19.125 233.69 19.195 ;
    RECT 233.48 19.485 233.69 19.555 ;
    RECT 233.02 18.765 233.23 18.835 ;
    RECT 233.02 19.125 233.23 19.195 ;
    RECT 233.02 19.485 233.23 19.555 ;
    RECT 230.16 18.765 230.37 18.835 ;
    RECT 230.16 19.125 230.37 19.195 ;
    RECT 230.16 19.485 230.37 19.555 ;
    RECT 229.7 18.765 229.91 18.835 ;
    RECT 229.7 19.125 229.91 19.195 ;
    RECT 229.7 19.485 229.91 19.555 ;
    RECT 366.28 18.765 366.49 18.835 ;
    RECT 366.28 19.125 366.49 19.195 ;
    RECT 366.28 19.485 366.49 19.555 ;
    RECT 365.82 18.765 366.03 18.835 ;
    RECT 365.82 19.125 366.03 19.195 ;
    RECT 365.82 19.485 366.03 19.555 ;
    RECT 226.84 18.765 227.05 18.835 ;
    RECT 226.84 19.125 227.05 19.195 ;
    RECT 226.84 19.485 227.05 19.555 ;
    RECT 226.38 18.765 226.59 18.835 ;
    RECT 226.38 19.125 226.59 19.195 ;
    RECT 226.38 19.485 226.59 19.555 ;
    RECT 362.96 18.765 363.17 18.835 ;
    RECT 362.96 19.125 363.17 19.195 ;
    RECT 362.96 19.485 363.17 19.555 ;
    RECT 362.5 18.765 362.71 18.835 ;
    RECT 362.5 19.125 362.71 19.195 ;
    RECT 362.5 19.485 362.71 19.555 ;
    RECT 223.52 18.765 223.73 18.835 ;
    RECT 223.52 19.125 223.73 19.195 ;
    RECT 223.52 19.485 223.73 19.555 ;
    RECT 223.06 18.765 223.27 18.835 ;
    RECT 223.06 19.125 223.27 19.195 ;
    RECT 223.06 19.485 223.27 19.555 ;
    RECT 359.64 18.765 359.85 18.835 ;
    RECT 359.64 19.125 359.85 19.195 ;
    RECT 359.64 19.485 359.85 19.555 ;
    RECT 359.18 18.765 359.39 18.835 ;
    RECT 359.18 19.125 359.39 19.195 ;
    RECT 359.18 19.485 359.39 19.555 ;
    RECT 220.2 18.765 220.41 18.835 ;
    RECT 220.2 19.125 220.41 19.195 ;
    RECT 220.2 19.485 220.41 19.555 ;
    RECT 219.74 18.765 219.95 18.835 ;
    RECT 219.74 19.125 219.95 19.195 ;
    RECT 219.74 19.485 219.95 19.555 ;
    RECT 356.32 18.765 356.53 18.835 ;
    RECT 356.32 19.125 356.53 19.195 ;
    RECT 356.32 19.485 356.53 19.555 ;
    RECT 355.86 18.765 356.07 18.835 ;
    RECT 355.86 19.125 356.07 19.195 ;
    RECT 355.86 19.485 356.07 19.555 ;
    RECT 353.0 18.765 353.21 18.835 ;
    RECT 353.0 19.125 353.21 19.195 ;
    RECT 353.0 19.485 353.21 19.555 ;
    RECT 352.54 18.765 352.75 18.835 ;
    RECT 352.54 19.125 352.75 19.195 ;
    RECT 352.54 19.485 352.75 19.555 ;
    RECT 216.88 18.765 217.09 18.835 ;
    RECT 216.88 19.125 217.09 19.195 ;
    RECT 216.88 19.485 217.09 19.555 ;
    RECT 216.42 18.765 216.63 18.835 ;
    RECT 216.42 19.125 216.63 19.195 ;
    RECT 216.42 19.485 216.63 19.555 ;
    RECT 349.68 18.765 349.89 18.835 ;
    RECT 349.68 19.125 349.89 19.195 ;
    RECT 349.68 19.485 349.89 19.555 ;
    RECT 349.22 18.765 349.43 18.835 ;
    RECT 349.22 19.125 349.43 19.195 ;
    RECT 349.22 19.485 349.43 19.555 ;
    RECT 213.56 18.765 213.77 18.835 ;
    RECT 213.56 19.125 213.77 19.195 ;
    RECT 213.56 19.485 213.77 19.555 ;
    RECT 213.1 18.765 213.31 18.835 ;
    RECT 213.1 19.125 213.31 19.195 ;
    RECT 213.1 19.485 213.31 19.555 ;
    RECT 346.36 18.765 346.57 18.835 ;
    RECT 346.36 19.125 346.57 19.195 ;
    RECT 346.36 19.485 346.57 19.555 ;
    RECT 345.9 18.765 346.11 18.835 ;
    RECT 345.9 19.125 346.11 19.195 ;
    RECT 345.9 19.485 346.11 19.555 ;
    RECT 210.24 18.765 210.45 18.835 ;
    RECT 210.24 19.125 210.45 19.195 ;
    RECT 210.24 19.485 210.45 19.555 ;
    RECT 209.78 18.765 209.99 18.835 ;
    RECT 209.78 19.125 209.99 19.195 ;
    RECT 209.78 19.485 209.99 19.555 ;
    RECT 343.04 18.765 343.25 18.835 ;
    RECT 343.04 19.125 343.25 19.195 ;
    RECT 343.04 19.485 343.25 19.555 ;
    RECT 342.58 18.765 342.79 18.835 ;
    RECT 342.58 19.125 342.79 19.195 ;
    RECT 342.58 19.485 342.79 19.555 ;
    RECT 206.92 18.765 207.13 18.835 ;
    RECT 206.92 19.125 207.13 19.195 ;
    RECT 206.92 19.485 207.13 19.555 ;
    RECT 206.46 18.765 206.67 18.835 ;
    RECT 206.46 19.125 206.67 19.195 ;
    RECT 206.46 19.485 206.67 19.555 ;
    RECT 339.72 18.765 339.93 18.835 ;
    RECT 339.72 19.125 339.93 19.195 ;
    RECT 339.72 19.485 339.93 19.555 ;
    RECT 339.26 18.765 339.47 18.835 ;
    RECT 339.26 19.125 339.47 19.195 ;
    RECT 339.26 19.485 339.47 19.555 ;
    RECT 203.6 18.765 203.81 18.835 ;
    RECT 203.6 19.125 203.81 19.195 ;
    RECT 203.6 19.485 203.81 19.555 ;
    RECT 203.14 18.765 203.35 18.835 ;
    RECT 203.14 19.125 203.35 19.195 ;
    RECT 203.14 19.485 203.35 19.555 ;
    RECT 336.4 18.765 336.61 18.835 ;
    RECT 336.4 19.125 336.61 19.195 ;
    RECT 336.4 19.485 336.61 19.555 ;
    RECT 335.94 18.765 336.15 18.835 ;
    RECT 335.94 19.125 336.15 19.195 ;
    RECT 335.94 19.485 336.15 19.555 ;
    RECT 266.68 18.765 266.89 18.835 ;
    RECT 266.68 19.125 266.89 19.195 ;
    RECT 266.68 19.485 266.89 19.555 ;
    RECT 266.22 18.765 266.43 18.835 ;
    RECT 266.22 19.125 266.43 19.195 ;
    RECT 266.22 19.485 266.43 19.555 ;
    RECT 263.36 18.765 263.57 18.835 ;
    RECT 263.36 19.125 263.57 19.195 ;
    RECT 263.36 19.485 263.57 19.555 ;
    RECT 262.9 18.765 263.11 18.835 ;
    RECT 262.9 19.125 263.11 19.195 ;
    RECT 262.9 19.485 263.11 19.555 ;
    RECT 260.04 18.765 260.25 18.835 ;
    RECT 260.04 19.125 260.25 19.195 ;
    RECT 260.04 19.485 260.25 19.555 ;
    RECT 259.58 18.765 259.79 18.835 ;
    RECT 259.58 19.125 259.79 19.195 ;
    RECT 259.58 19.485 259.79 19.555 ;
    RECT 256.72 18.765 256.93 18.835 ;
    RECT 256.72 19.125 256.93 19.195 ;
    RECT 256.72 19.485 256.93 19.555 ;
    RECT 256.26 18.765 256.47 18.835 ;
    RECT 256.26 19.125 256.47 19.195 ;
    RECT 256.26 19.485 256.47 19.555 ;
    RECT 253.4 18.765 253.61 18.835 ;
    RECT 253.4 19.125 253.61 19.195 ;
    RECT 253.4 19.485 253.61 19.555 ;
    RECT 252.94 18.765 253.15 18.835 ;
    RECT 252.94 19.125 253.15 19.195 ;
    RECT 252.94 19.485 253.15 19.555 ;
    RECT 250.08 18.765 250.29 18.835 ;
    RECT 250.08 19.125 250.29 19.195 ;
    RECT 250.08 19.485 250.29 19.555 ;
    RECT 249.62 18.765 249.83 18.835 ;
    RECT 249.62 19.125 249.83 19.195 ;
    RECT 249.62 19.485 249.83 19.555 ;
    RECT 246.76 18.765 246.97 18.835 ;
    RECT 246.76 19.125 246.97 19.195 ;
    RECT 246.76 19.485 246.97 19.555 ;
    RECT 246.3 18.765 246.51 18.835 ;
    RECT 246.3 19.125 246.51 19.195 ;
    RECT 246.3 19.485 246.51 19.555 ;
    RECT 243.44 18.765 243.65 18.835 ;
    RECT 243.44 19.125 243.65 19.195 ;
    RECT 243.44 19.485 243.65 19.555 ;
    RECT 242.98 18.765 243.19 18.835 ;
    RECT 242.98 19.125 243.19 19.195 ;
    RECT 242.98 19.485 243.19 19.555 ;
    RECT 240.12 18.765 240.33 18.835 ;
    RECT 240.12 19.125 240.33 19.195 ;
    RECT 240.12 19.485 240.33 19.555 ;
    RECT 239.66 18.765 239.87 18.835 ;
    RECT 239.66 19.125 239.87 19.195 ;
    RECT 239.66 19.485 239.87 19.555 ;
    RECT 236.8 18.765 237.01 18.835 ;
    RECT 236.8 19.125 237.01 19.195 ;
    RECT 236.8 19.485 237.01 19.555 ;
    RECT 236.34 18.765 236.55 18.835 ;
    RECT 236.34 19.125 236.55 19.195 ;
    RECT 236.34 19.485 236.55 19.555 ;
    RECT 374.15 19.125 374.22 19.195 ;
    RECT 333.08 18.765 333.29 18.835 ;
    RECT 333.08 19.125 333.29 19.195 ;
    RECT 333.08 19.485 333.29 19.555 ;
    RECT 332.62 18.765 332.83 18.835 ;
    RECT 332.62 19.125 332.83 19.195 ;
    RECT 332.62 19.485 332.83 19.555 ;
    RECT 329.76 18.765 329.97 18.835 ;
    RECT 329.76 19.125 329.97 19.195 ;
    RECT 329.76 19.485 329.97 19.555 ;
    RECT 329.3 18.765 329.51 18.835 ;
    RECT 329.3 19.125 329.51 19.195 ;
    RECT 329.3 19.485 329.51 19.555 ;
    RECT 326.44 18.765 326.65 18.835 ;
    RECT 326.44 19.125 326.65 19.195 ;
    RECT 326.44 19.485 326.65 19.555 ;
    RECT 325.98 18.765 326.19 18.835 ;
    RECT 325.98 19.125 326.19 19.195 ;
    RECT 325.98 19.485 326.19 19.555 ;
    RECT 323.12 18.765 323.33 18.835 ;
    RECT 323.12 19.125 323.33 19.195 ;
    RECT 323.12 19.485 323.33 19.555 ;
    RECT 322.66 18.765 322.87 18.835 ;
    RECT 322.66 19.125 322.87 19.195 ;
    RECT 322.66 19.485 322.87 19.555 ;
    RECT 319.8 18.765 320.01 18.835 ;
    RECT 319.8 19.125 320.01 19.195 ;
    RECT 319.8 19.485 320.01 19.555 ;
    RECT 319.34 18.765 319.55 18.835 ;
    RECT 319.34 19.125 319.55 19.195 ;
    RECT 319.34 19.485 319.55 19.555 ;
    RECT 316.48 18.765 316.69 18.835 ;
    RECT 316.48 19.125 316.69 19.195 ;
    RECT 316.48 19.485 316.69 19.555 ;
    RECT 316.02 18.765 316.23 18.835 ;
    RECT 316.02 19.125 316.23 19.195 ;
    RECT 316.02 19.485 316.23 19.555 ;
    RECT 313.16 18.765 313.37 18.835 ;
    RECT 313.16 19.125 313.37 19.195 ;
    RECT 313.16 19.485 313.37 19.555 ;
    RECT 312.7 18.765 312.91 18.835 ;
    RECT 312.7 19.125 312.91 19.195 ;
    RECT 312.7 19.485 312.91 19.555 ;
    RECT 309.84 18.765 310.05 18.835 ;
    RECT 309.84 19.125 310.05 19.195 ;
    RECT 309.84 19.485 310.05 19.555 ;
    RECT 309.38 18.765 309.59 18.835 ;
    RECT 309.38 19.125 309.59 19.195 ;
    RECT 309.38 19.485 309.59 19.555 ;
    RECT 306.52 18.765 306.73 18.835 ;
    RECT 306.52 19.125 306.73 19.195 ;
    RECT 306.52 19.485 306.73 19.555 ;
    RECT 306.06 18.765 306.27 18.835 ;
    RECT 306.06 19.125 306.27 19.195 ;
    RECT 306.06 19.485 306.27 19.555 ;
    RECT 252.45 57.885 252.66 57.955 ;
    RECT 272.37 57.885 272.58 57.955 ;
    RECT 222.57 57.885 222.78 57.955 ;
    RECT 272.86 58.145 273.07 58.215 ;
    RECT 355.86 58.145 356.07 58.215 ;
    RECT 273.32 58.145 273.53 58.215 ;
    RECT 356.32 58.145 356.53 58.215 ;
    RECT 296.1 58.145 296.31 58.215 ;
    RECT 296.56 58.145 296.77 58.215 ;
    RECT 318.85 57.885 319.06 57.955 ;
    RECT 338.77 57.885 338.98 57.955 ;
    RECT 309.38 58.145 309.59 58.215 ;
    RECT 309.84 58.145 310.05 58.215 ;
    RECT 249.62 58.145 249.83 58.215 ;
    RECT 332.62 58.145 332.83 58.215 ;
    RECT 250.08 58.145 250.29 58.215 ;
    RECT 333.08 58.145 333.29 58.215 ;
    RECT 213.1 58.145 213.31 58.215 ;
    RECT 213.56 58.145 213.77 58.215 ;
    RECT 362.01 57.885 362.22 57.955 ;
    RECT 215.93 57.885 216.14 57.955 ;
    RECT 298.93 57.885 299.14 57.955 ;
    RECT 369.14 58.145 369.35 58.215 ;
    RECT 369.6 58.145 369.81 58.215 ;
    RECT 289.46 58.145 289.67 58.215 ;
    RECT 289.92 58.145 290.13 58.215 ;
    RECT 245.81 57.885 246.02 57.955 ;
    RECT 242.98 58.145 243.19 58.215 ;
    RECT 325.98 58.145 326.19 58.215 ;
    RECT 243.44 58.145 243.65 58.215 ;
    RECT 326.44 58.145 326.65 58.215 ;
    RECT 266.22 58.145 266.43 58.215 ;
    RECT 355.37 57.885 355.58 57.955 ;
    RECT 266.68 58.145 266.89 58.215 ;
    RECT 206.46 58.145 206.67 58.215 ;
    RECT 206.92 58.145 207.13 58.215 ;
    RECT 349.22 58.145 349.43 58.215 ;
    RECT 229.7 58.145 229.91 58.215 ;
    RECT 349.68 58.145 349.89 58.215 ;
    RECT 230.16 58.145 230.37 58.215 ;
    RECT 292.29 57.885 292.5 57.955 ;
    RECT 312.21 57.885 312.42 57.955 ;
    RECT 302.74 58.145 302.95 58.215 ;
    RECT 303.2 58.145 303.41 58.215 ;
    RECT 374.36 57.885 374.43 57.955 ;
    RECT 374.15 58.145 374.22 58.215 ;
    RECT 239.17 57.885 239.38 57.955 ;
    RECT 209.29 57.885 209.5 57.955 ;
    RECT 200.395 57.885 200.465 57.955 ;
    RECT 200.605 58.145 200.675 58.215 ;
    RECT 348.73 57.885 348.94 57.955 ;
    RECT 262.41 57.885 262.62 57.955 ;
    RECT 232.53 57.885 232.74 57.955 ;
    RECT 259.58 58.145 259.79 58.215 ;
    RECT 260.04 58.145 260.25 58.215 ;
    RECT 342.58 58.145 342.79 58.215 ;
    RECT 223.06 58.145 223.27 58.215 ;
    RECT 343.04 58.145 343.25 58.215 ;
    RECT 223.52 58.145 223.73 58.215 ;
    RECT 282.82 58.145 283.03 58.215 ;
    RECT 365.82 58.145 366.03 58.215 ;
    RECT 283.28 58.145 283.49 58.215 ;
    RECT 366.28 58.145 366.49 58.215 ;
    RECT 285.65 57.885 285.86 57.955 ;
    RECT 305.57 57.885 305.78 57.955 ;
    RECT 319.34 58.145 319.55 58.215 ;
    RECT 328.81 57.885 329.02 57.955 ;
    RECT 319.8 58.145 320.01 58.215 ;
    RECT 202.65 57.885 202.86 57.955 ;
    RECT 236.34 58.145 236.55 58.215 ;
    RECT 371.97 57.885 372.18 57.955 ;
    RECT 236.8 58.145 237.01 58.215 ;
    RECT 255.77 57.885 255.98 57.955 ;
    RECT 275.69 57.885 275.9 57.955 ;
    RECT 225.89 57.885 226.1 57.955 ;
    RECT 276.18 58.145 276.39 58.215 ;
    RECT 359.18 58.145 359.39 58.215 ;
    RECT 276.64 58.145 276.85 58.215 ;
    RECT 359.64 58.145 359.85 58.215 ;
    RECT 299.42 58.145 299.63 58.215 ;
    RECT 299.88 58.145 300.09 58.215 ;
    RECT 372.46 58.145 372.67 58.215 ;
    RECT 322.17 57.885 322.38 57.955 ;
    RECT 342.09 57.885 342.3 57.955 ;
    RECT 372.92 58.145 373.13 58.215 ;
    RECT 312.7 58.145 312.91 58.215 ;
    RECT 313.16 58.145 313.37 58.215 ;
    RECT 252.94 58.145 253.15 58.215 ;
    RECT 253.4 58.145 253.61 58.215 ;
    RECT 335.94 58.145 336.15 58.215 ;
    RECT 336.4 58.145 336.61 58.215 ;
    RECT 216.42 58.145 216.63 58.215 ;
    RECT 216.88 58.145 217.09 58.215 ;
    RECT 365.33 57.885 365.54 57.955 ;
    RECT 279.01 57.885 279.22 57.955 ;
    RECT 249.13 57.885 249.34 57.955 ;
    RECT 269.05 57.885 269.26 57.955 ;
    RECT 219.25 57.885 219.46 57.955 ;
    RECT 292.78 58.145 292.99 58.215 ;
    RECT 293.24 58.145 293.45 58.215 ;
    RECT 315.53 57.885 315.74 57.955 ;
    RECT 335.45 57.885 335.66 57.955 ;
    RECT 306.06 58.145 306.27 58.215 ;
    RECT 306.52 58.145 306.73 58.215 ;
    RECT 246.3 58.145 246.51 58.215 ;
    RECT 329.3 58.145 329.51 58.215 ;
    RECT 246.76 58.145 246.97 58.215 ;
    RECT 329.76 58.145 329.97 58.215 ;
    RECT 358.69 57.885 358.9 57.955 ;
    RECT 209.78 58.145 209.99 58.215 ;
    RECT 269.54 58.145 269.75 58.215 ;
    RECT 352.54 58.145 352.75 58.215 ;
    RECT 210.24 58.145 210.45 58.215 ;
    RECT 270.0 58.145 270.21 58.215 ;
    RECT 353.0 58.145 353.21 58.215 ;
    RECT 233.02 58.145 233.23 58.215 ;
    RECT 233.48 58.145 233.69 58.215 ;
    RECT 295.61 57.885 295.82 57.955 ;
    RECT 242.49 57.885 242.7 57.955 ;
    RECT 212.61 57.885 212.82 57.955 ;
    RECT 239.66 58.145 239.87 58.215 ;
    RECT 322.66 58.145 322.87 58.215 ;
    RECT 240.12 58.145 240.33 58.215 ;
    RECT 323.12 58.145 323.33 58.215 ;
    RECT 262.9 58.145 263.11 58.215 ;
    RECT 265.73 57.885 265.94 57.955 ;
    RECT 352.05 57.885 352.26 57.955 ;
    RECT 263.36 58.145 263.57 58.215 ;
    RECT 345.9 58.145 346.11 58.215 ;
    RECT 346.36 58.145 346.57 58.215 ;
    RECT 226.38 58.145 226.59 58.215 ;
    RECT 286.14 58.145 286.35 58.215 ;
    RECT 226.84 58.145 227.05 58.215 ;
    RECT 286.6 58.145 286.81 58.215 ;
    RECT 288.97 57.885 289.18 57.955 ;
    RECT 308.89 57.885 309.1 57.955 ;
    RECT 332.13 57.885 332.34 57.955 ;
    RECT 203.14 58.145 203.35 58.215 ;
    RECT 203.6 58.145 203.81 58.215 ;
    RECT 235.85 57.885 236.06 57.955 ;
    RECT 205.97 57.885 206.18 57.955 ;
    RECT 259.09 57.885 259.3 57.955 ;
    RECT 229.21 57.885 229.42 57.955 ;
    RECT 256.26 58.145 256.47 58.215 ;
    RECT 256.72 58.145 256.93 58.215 ;
    RECT 339.26 58.145 339.47 58.215 ;
    RECT 339.72 58.145 339.93 58.215 ;
    RECT 279.5 58.145 279.71 58.215 ;
    RECT 362.5 58.145 362.71 58.215 ;
    RECT 279.96 58.145 280.17 58.215 ;
    RECT 362.96 58.145 363.17 58.215 ;
    RECT 282.33 57.885 282.54 57.955 ;
    RECT 302.25 57.885 302.46 57.955 ;
    RECT 316.02 58.145 316.23 58.215 ;
    RECT 325.49 57.885 325.7 57.955 ;
    RECT 345.41 57.885 345.62 57.955 ;
    RECT 316.48 58.145 316.69 58.215 ;
    RECT 219.74 58.145 219.95 58.215 ;
    RECT 220.2 58.145 220.41 58.215 ;
    RECT 368.65 57.885 368.86 57.955 ;
    RECT 303.2 56.925 303.41 56.995 ;
    RECT 303.2 57.285 303.41 57.355 ;
    RECT 303.2 57.645 303.41 57.715 ;
    RECT 302.74 56.925 302.95 56.995 ;
    RECT 302.74 57.285 302.95 57.355 ;
    RECT 302.74 57.645 302.95 57.715 ;
    RECT 372.92 56.925 373.13 56.995 ;
    RECT 372.92 57.285 373.13 57.355 ;
    RECT 372.92 57.645 373.13 57.715 ;
    RECT 372.46 56.925 372.67 56.995 ;
    RECT 372.46 57.285 372.67 57.355 ;
    RECT 372.46 57.645 372.67 57.715 ;
    RECT 369.6 56.925 369.81 56.995 ;
    RECT 369.6 57.285 369.81 57.355 ;
    RECT 369.6 57.645 369.81 57.715 ;
    RECT 369.14 56.925 369.35 56.995 ;
    RECT 369.14 57.285 369.35 57.355 ;
    RECT 369.14 57.645 369.35 57.715 ;
    RECT 200.605 57.285 200.675 57.355 ;
    RECT 299.88 56.925 300.09 56.995 ;
    RECT 299.88 57.285 300.09 57.355 ;
    RECT 299.88 57.645 300.09 57.715 ;
    RECT 299.42 56.925 299.63 56.995 ;
    RECT 299.42 57.285 299.63 57.355 ;
    RECT 299.42 57.645 299.63 57.715 ;
    RECT 296.56 56.925 296.77 56.995 ;
    RECT 296.56 57.285 296.77 57.355 ;
    RECT 296.56 57.645 296.77 57.715 ;
    RECT 296.1 56.925 296.31 56.995 ;
    RECT 296.1 57.285 296.31 57.355 ;
    RECT 296.1 57.645 296.31 57.715 ;
    RECT 293.24 56.925 293.45 56.995 ;
    RECT 293.24 57.285 293.45 57.355 ;
    RECT 293.24 57.645 293.45 57.715 ;
    RECT 292.78 56.925 292.99 56.995 ;
    RECT 292.78 57.285 292.99 57.355 ;
    RECT 292.78 57.645 292.99 57.715 ;
    RECT 289.92 56.925 290.13 56.995 ;
    RECT 289.92 57.285 290.13 57.355 ;
    RECT 289.92 57.645 290.13 57.715 ;
    RECT 289.46 56.925 289.67 56.995 ;
    RECT 289.46 57.285 289.67 57.355 ;
    RECT 289.46 57.645 289.67 57.715 ;
    RECT 286.6 56.925 286.81 56.995 ;
    RECT 286.6 57.285 286.81 57.355 ;
    RECT 286.6 57.645 286.81 57.715 ;
    RECT 286.14 56.925 286.35 56.995 ;
    RECT 286.14 57.285 286.35 57.355 ;
    RECT 286.14 57.645 286.35 57.715 ;
    RECT 283.28 56.925 283.49 56.995 ;
    RECT 283.28 57.285 283.49 57.355 ;
    RECT 283.28 57.645 283.49 57.715 ;
    RECT 282.82 56.925 283.03 56.995 ;
    RECT 282.82 57.285 283.03 57.355 ;
    RECT 282.82 57.645 283.03 57.715 ;
    RECT 279.96 56.925 280.17 56.995 ;
    RECT 279.96 57.285 280.17 57.355 ;
    RECT 279.96 57.645 280.17 57.715 ;
    RECT 279.5 56.925 279.71 56.995 ;
    RECT 279.5 57.285 279.71 57.355 ;
    RECT 279.5 57.645 279.71 57.715 ;
    RECT 276.64 56.925 276.85 56.995 ;
    RECT 276.64 57.285 276.85 57.355 ;
    RECT 276.64 57.645 276.85 57.715 ;
    RECT 276.18 56.925 276.39 56.995 ;
    RECT 276.18 57.285 276.39 57.355 ;
    RECT 276.18 57.645 276.39 57.715 ;
    RECT 273.32 56.925 273.53 56.995 ;
    RECT 273.32 57.285 273.53 57.355 ;
    RECT 273.32 57.645 273.53 57.715 ;
    RECT 272.86 56.925 273.07 56.995 ;
    RECT 272.86 57.285 273.07 57.355 ;
    RECT 272.86 57.645 273.07 57.715 ;
    RECT 270.0 56.925 270.21 56.995 ;
    RECT 270.0 57.285 270.21 57.355 ;
    RECT 270.0 57.645 270.21 57.715 ;
    RECT 269.54 56.925 269.75 56.995 ;
    RECT 269.54 57.285 269.75 57.355 ;
    RECT 269.54 57.645 269.75 57.715 ;
    RECT 233.48 56.925 233.69 56.995 ;
    RECT 233.48 57.285 233.69 57.355 ;
    RECT 233.48 57.645 233.69 57.715 ;
    RECT 233.02 56.925 233.23 56.995 ;
    RECT 233.02 57.285 233.23 57.355 ;
    RECT 233.02 57.645 233.23 57.715 ;
    RECT 230.16 56.925 230.37 56.995 ;
    RECT 230.16 57.285 230.37 57.355 ;
    RECT 230.16 57.645 230.37 57.715 ;
    RECT 229.7 56.925 229.91 56.995 ;
    RECT 229.7 57.285 229.91 57.355 ;
    RECT 229.7 57.645 229.91 57.715 ;
    RECT 366.28 56.925 366.49 56.995 ;
    RECT 366.28 57.285 366.49 57.355 ;
    RECT 366.28 57.645 366.49 57.715 ;
    RECT 365.82 56.925 366.03 56.995 ;
    RECT 365.82 57.285 366.03 57.355 ;
    RECT 365.82 57.645 366.03 57.715 ;
    RECT 226.84 56.925 227.05 56.995 ;
    RECT 226.84 57.285 227.05 57.355 ;
    RECT 226.84 57.645 227.05 57.715 ;
    RECT 226.38 56.925 226.59 56.995 ;
    RECT 226.38 57.285 226.59 57.355 ;
    RECT 226.38 57.645 226.59 57.715 ;
    RECT 362.96 56.925 363.17 56.995 ;
    RECT 362.96 57.285 363.17 57.355 ;
    RECT 362.96 57.645 363.17 57.715 ;
    RECT 362.5 56.925 362.71 56.995 ;
    RECT 362.5 57.285 362.71 57.355 ;
    RECT 362.5 57.645 362.71 57.715 ;
    RECT 223.52 56.925 223.73 56.995 ;
    RECT 223.52 57.285 223.73 57.355 ;
    RECT 223.52 57.645 223.73 57.715 ;
    RECT 223.06 56.925 223.27 56.995 ;
    RECT 223.06 57.285 223.27 57.355 ;
    RECT 223.06 57.645 223.27 57.715 ;
    RECT 359.64 56.925 359.85 56.995 ;
    RECT 359.64 57.285 359.85 57.355 ;
    RECT 359.64 57.645 359.85 57.715 ;
    RECT 359.18 56.925 359.39 56.995 ;
    RECT 359.18 57.285 359.39 57.355 ;
    RECT 359.18 57.645 359.39 57.715 ;
    RECT 220.2 56.925 220.41 56.995 ;
    RECT 220.2 57.285 220.41 57.355 ;
    RECT 220.2 57.645 220.41 57.715 ;
    RECT 219.74 56.925 219.95 56.995 ;
    RECT 219.74 57.285 219.95 57.355 ;
    RECT 219.74 57.645 219.95 57.715 ;
    RECT 356.32 56.925 356.53 56.995 ;
    RECT 356.32 57.285 356.53 57.355 ;
    RECT 356.32 57.645 356.53 57.715 ;
    RECT 355.86 56.925 356.07 56.995 ;
    RECT 355.86 57.285 356.07 57.355 ;
    RECT 355.86 57.645 356.07 57.715 ;
    RECT 353.0 56.925 353.21 56.995 ;
    RECT 353.0 57.285 353.21 57.355 ;
    RECT 353.0 57.645 353.21 57.715 ;
    RECT 352.54 56.925 352.75 56.995 ;
    RECT 352.54 57.285 352.75 57.355 ;
    RECT 352.54 57.645 352.75 57.715 ;
    RECT 216.88 56.925 217.09 56.995 ;
    RECT 216.88 57.285 217.09 57.355 ;
    RECT 216.88 57.645 217.09 57.715 ;
    RECT 216.42 56.925 216.63 56.995 ;
    RECT 216.42 57.285 216.63 57.355 ;
    RECT 216.42 57.645 216.63 57.715 ;
    RECT 349.68 56.925 349.89 56.995 ;
    RECT 349.68 57.285 349.89 57.355 ;
    RECT 349.68 57.645 349.89 57.715 ;
    RECT 349.22 56.925 349.43 56.995 ;
    RECT 349.22 57.285 349.43 57.355 ;
    RECT 349.22 57.645 349.43 57.715 ;
    RECT 213.56 56.925 213.77 56.995 ;
    RECT 213.56 57.285 213.77 57.355 ;
    RECT 213.56 57.645 213.77 57.715 ;
    RECT 213.1 56.925 213.31 56.995 ;
    RECT 213.1 57.285 213.31 57.355 ;
    RECT 213.1 57.645 213.31 57.715 ;
    RECT 346.36 56.925 346.57 56.995 ;
    RECT 346.36 57.285 346.57 57.355 ;
    RECT 346.36 57.645 346.57 57.715 ;
    RECT 345.9 56.925 346.11 56.995 ;
    RECT 345.9 57.285 346.11 57.355 ;
    RECT 345.9 57.645 346.11 57.715 ;
    RECT 210.24 56.925 210.45 56.995 ;
    RECT 210.24 57.285 210.45 57.355 ;
    RECT 210.24 57.645 210.45 57.715 ;
    RECT 209.78 56.925 209.99 56.995 ;
    RECT 209.78 57.285 209.99 57.355 ;
    RECT 209.78 57.645 209.99 57.715 ;
    RECT 343.04 56.925 343.25 56.995 ;
    RECT 343.04 57.285 343.25 57.355 ;
    RECT 343.04 57.645 343.25 57.715 ;
    RECT 342.58 56.925 342.79 56.995 ;
    RECT 342.58 57.285 342.79 57.355 ;
    RECT 342.58 57.645 342.79 57.715 ;
    RECT 206.92 56.925 207.13 56.995 ;
    RECT 206.92 57.285 207.13 57.355 ;
    RECT 206.92 57.645 207.13 57.715 ;
    RECT 206.46 56.925 206.67 56.995 ;
    RECT 206.46 57.285 206.67 57.355 ;
    RECT 206.46 57.645 206.67 57.715 ;
    RECT 339.72 56.925 339.93 56.995 ;
    RECT 339.72 57.285 339.93 57.355 ;
    RECT 339.72 57.645 339.93 57.715 ;
    RECT 339.26 56.925 339.47 56.995 ;
    RECT 339.26 57.285 339.47 57.355 ;
    RECT 339.26 57.645 339.47 57.715 ;
    RECT 203.6 56.925 203.81 56.995 ;
    RECT 203.6 57.285 203.81 57.355 ;
    RECT 203.6 57.645 203.81 57.715 ;
    RECT 203.14 56.925 203.35 56.995 ;
    RECT 203.14 57.285 203.35 57.355 ;
    RECT 203.14 57.645 203.35 57.715 ;
    RECT 336.4 56.925 336.61 56.995 ;
    RECT 336.4 57.285 336.61 57.355 ;
    RECT 336.4 57.645 336.61 57.715 ;
    RECT 335.94 56.925 336.15 56.995 ;
    RECT 335.94 57.285 336.15 57.355 ;
    RECT 335.94 57.645 336.15 57.715 ;
    RECT 266.68 56.925 266.89 56.995 ;
    RECT 266.68 57.285 266.89 57.355 ;
    RECT 266.68 57.645 266.89 57.715 ;
    RECT 266.22 56.925 266.43 56.995 ;
    RECT 266.22 57.285 266.43 57.355 ;
    RECT 266.22 57.645 266.43 57.715 ;
    RECT 263.36 56.925 263.57 56.995 ;
    RECT 263.36 57.285 263.57 57.355 ;
    RECT 263.36 57.645 263.57 57.715 ;
    RECT 262.9 56.925 263.11 56.995 ;
    RECT 262.9 57.285 263.11 57.355 ;
    RECT 262.9 57.645 263.11 57.715 ;
    RECT 260.04 56.925 260.25 56.995 ;
    RECT 260.04 57.285 260.25 57.355 ;
    RECT 260.04 57.645 260.25 57.715 ;
    RECT 259.58 56.925 259.79 56.995 ;
    RECT 259.58 57.285 259.79 57.355 ;
    RECT 259.58 57.645 259.79 57.715 ;
    RECT 256.72 56.925 256.93 56.995 ;
    RECT 256.72 57.285 256.93 57.355 ;
    RECT 256.72 57.645 256.93 57.715 ;
    RECT 256.26 56.925 256.47 56.995 ;
    RECT 256.26 57.285 256.47 57.355 ;
    RECT 256.26 57.645 256.47 57.715 ;
    RECT 253.4 56.925 253.61 56.995 ;
    RECT 253.4 57.285 253.61 57.355 ;
    RECT 253.4 57.645 253.61 57.715 ;
    RECT 252.94 56.925 253.15 56.995 ;
    RECT 252.94 57.285 253.15 57.355 ;
    RECT 252.94 57.645 253.15 57.715 ;
    RECT 250.08 56.925 250.29 56.995 ;
    RECT 250.08 57.285 250.29 57.355 ;
    RECT 250.08 57.645 250.29 57.715 ;
    RECT 249.62 56.925 249.83 56.995 ;
    RECT 249.62 57.285 249.83 57.355 ;
    RECT 249.62 57.645 249.83 57.715 ;
    RECT 246.76 56.925 246.97 56.995 ;
    RECT 246.76 57.285 246.97 57.355 ;
    RECT 246.76 57.645 246.97 57.715 ;
    RECT 246.3 56.925 246.51 56.995 ;
    RECT 246.3 57.285 246.51 57.355 ;
    RECT 246.3 57.645 246.51 57.715 ;
    RECT 243.44 56.925 243.65 56.995 ;
    RECT 243.44 57.285 243.65 57.355 ;
    RECT 243.44 57.645 243.65 57.715 ;
    RECT 242.98 56.925 243.19 56.995 ;
    RECT 242.98 57.285 243.19 57.355 ;
    RECT 242.98 57.645 243.19 57.715 ;
    RECT 240.12 56.925 240.33 56.995 ;
    RECT 240.12 57.285 240.33 57.355 ;
    RECT 240.12 57.645 240.33 57.715 ;
    RECT 239.66 56.925 239.87 56.995 ;
    RECT 239.66 57.285 239.87 57.355 ;
    RECT 239.66 57.645 239.87 57.715 ;
    RECT 236.8 56.925 237.01 56.995 ;
    RECT 236.8 57.285 237.01 57.355 ;
    RECT 236.8 57.645 237.01 57.715 ;
    RECT 236.34 56.925 236.55 56.995 ;
    RECT 236.34 57.285 236.55 57.355 ;
    RECT 236.34 57.645 236.55 57.715 ;
    RECT 374.15 57.285 374.22 57.355 ;
    RECT 333.08 56.925 333.29 56.995 ;
    RECT 333.08 57.285 333.29 57.355 ;
    RECT 333.08 57.645 333.29 57.715 ;
    RECT 332.62 56.925 332.83 56.995 ;
    RECT 332.62 57.285 332.83 57.355 ;
    RECT 332.62 57.645 332.83 57.715 ;
    RECT 329.76 56.925 329.97 56.995 ;
    RECT 329.76 57.285 329.97 57.355 ;
    RECT 329.76 57.645 329.97 57.715 ;
    RECT 329.3 56.925 329.51 56.995 ;
    RECT 329.3 57.285 329.51 57.355 ;
    RECT 329.3 57.645 329.51 57.715 ;
    RECT 326.44 56.925 326.65 56.995 ;
    RECT 326.44 57.285 326.65 57.355 ;
    RECT 326.44 57.645 326.65 57.715 ;
    RECT 325.98 56.925 326.19 56.995 ;
    RECT 325.98 57.285 326.19 57.355 ;
    RECT 325.98 57.645 326.19 57.715 ;
    RECT 323.12 56.925 323.33 56.995 ;
    RECT 323.12 57.285 323.33 57.355 ;
    RECT 323.12 57.645 323.33 57.715 ;
    RECT 322.66 56.925 322.87 56.995 ;
    RECT 322.66 57.285 322.87 57.355 ;
    RECT 322.66 57.645 322.87 57.715 ;
    RECT 319.8 56.925 320.01 56.995 ;
    RECT 319.8 57.285 320.01 57.355 ;
    RECT 319.8 57.645 320.01 57.715 ;
    RECT 319.34 56.925 319.55 56.995 ;
    RECT 319.34 57.285 319.55 57.355 ;
    RECT 319.34 57.645 319.55 57.715 ;
    RECT 316.48 56.925 316.69 56.995 ;
    RECT 316.48 57.285 316.69 57.355 ;
    RECT 316.48 57.645 316.69 57.715 ;
    RECT 316.02 56.925 316.23 56.995 ;
    RECT 316.02 57.285 316.23 57.355 ;
    RECT 316.02 57.645 316.23 57.715 ;
    RECT 313.16 56.925 313.37 56.995 ;
    RECT 313.16 57.285 313.37 57.355 ;
    RECT 313.16 57.645 313.37 57.715 ;
    RECT 312.7 56.925 312.91 56.995 ;
    RECT 312.7 57.285 312.91 57.355 ;
    RECT 312.7 57.645 312.91 57.715 ;
    RECT 309.84 56.925 310.05 56.995 ;
    RECT 309.84 57.285 310.05 57.355 ;
    RECT 309.84 57.645 310.05 57.715 ;
    RECT 309.38 56.925 309.59 56.995 ;
    RECT 309.38 57.285 309.59 57.355 ;
    RECT 309.38 57.645 309.59 57.715 ;
    RECT 306.52 56.925 306.73 56.995 ;
    RECT 306.52 57.285 306.73 57.355 ;
    RECT 306.52 57.645 306.73 57.715 ;
    RECT 306.06 56.925 306.27 56.995 ;
    RECT 306.06 57.285 306.27 57.355 ;
    RECT 306.06 57.645 306.27 57.715 ;
    RECT 303.2 56.205 303.41 56.275 ;
    RECT 303.2 56.565 303.41 56.635 ;
    RECT 303.2 56.925 303.41 56.995 ;
    RECT 302.74 56.205 302.95 56.275 ;
    RECT 302.74 56.565 302.95 56.635 ;
    RECT 302.74 56.925 302.95 56.995 ;
    RECT 372.92 56.205 373.13 56.275 ;
    RECT 372.92 56.565 373.13 56.635 ;
    RECT 372.92 56.925 373.13 56.995 ;
    RECT 372.46 56.205 372.67 56.275 ;
    RECT 372.46 56.565 372.67 56.635 ;
    RECT 372.46 56.925 372.67 56.995 ;
    RECT 369.6 56.205 369.81 56.275 ;
    RECT 369.6 56.565 369.81 56.635 ;
    RECT 369.6 56.925 369.81 56.995 ;
    RECT 369.14 56.205 369.35 56.275 ;
    RECT 369.14 56.565 369.35 56.635 ;
    RECT 369.14 56.925 369.35 56.995 ;
    RECT 200.605 56.565 200.675 56.635 ;
    RECT 299.88 56.205 300.09 56.275 ;
    RECT 299.88 56.565 300.09 56.635 ;
    RECT 299.88 56.925 300.09 56.995 ;
    RECT 299.42 56.205 299.63 56.275 ;
    RECT 299.42 56.565 299.63 56.635 ;
    RECT 299.42 56.925 299.63 56.995 ;
    RECT 296.56 56.205 296.77 56.275 ;
    RECT 296.56 56.565 296.77 56.635 ;
    RECT 296.56 56.925 296.77 56.995 ;
    RECT 296.1 56.205 296.31 56.275 ;
    RECT 296.1 56.565 296.31 56.635 ;
    RECT 296.1 56.925 296.31 56.995 ;
    RECT 293.24 56.205 293.45 56.275 ;
    RECT 293.24 56.565 293.45 56.635 ;
    RECT 293.24 56.925 293.45 56.995 ;
    RECT 292.78 56.205 292.99 56.275 ;
    RECT 292.78 56.565 292.99 56.635 ;
    RECT 292.78 56.925 292.99 56.995 ;
    RECT 289.92 56.205 290.13 56.275 ;
    RECT 289.92 56.565 290.13 56.635 ;
    RECT 289.92 56.925 290.13 56.995 ;
    RECT 289.46 56.205 289.67 56.275 ;
    RECT 289.46 56.565 289.67 56.635 ;
    RECT 289.46 56.925 289.67 56.995 ;
    RECT 286.6 56.205 286.81 56.275 ;
    RECT 286.6 56.565 286.81 56.635 ;
    RECT 286.6 56.925 286.81 56.995 ;
    RECT 286.14 56.205 286.35 56.275 ;
    RECT 286.14 56.565 286.35 56.635 ;
    RECT 286.14 56.925 286.35 56.995 ;
    RECT 283.28 56.205 283.49 56.275 ;
    RECT 283.28 56.565 283.49 56.635 ;
    RECT 283.28 56.925 283.49 56.995 ;
    RECT 282.82 56.205 283.03 56.275 ;
    RECT 282.82 56.565 283.03 56.635 ;
    RECT 282.82 56.925 283.03 56.995 ;
    RECT 279.96 56.205 280.17 56.275 ;
    RECT 279.96 56.565 280.17 56.635 ;
    RECT 279.96 56.925 280.17 56.995 ;
    RECT 279.5 56.205 279.71 56.275 ;
    RECT 279.5 56.565 279.71 56.635 ;
    RECT 279.5 56.925 279.71 56.995 ;
    RECT 276.64 56.205 276.85 56.275 ;
    RECT 276.64 56.565 276.85 56.635 ;
    RECT 276.64 56.925 276.85 56.995 ;
    RECT 276.18 56.205 276.39 56.275 ;
    RECT 276.18 56.565 276.39 56.635 ;
    RECT 276.18 56.925 276.39 56.995 ;
    RECT 273.32 56.205 273.53 56.275 ;
    RECT 273.32 56.565 273.53 56.635 ;
    RECT 273.32 56.925 273.53 56.995 ;
    RECT 272.86 56.205 273.07 56.275 ;
    RECT 272.86 56.565 273.07 56.635 ;
    RECT 272.86 56.925 273.07 56.995 ;
    RECT 270.0 56.205 270.21 56.275 ;
    RECT 270.0 56.565 270.21 56.635 ;
    RECT 270.0 56.925 270.21 56.995 ;
    RECT 269.54 56.205 269.75 56.275 ;
    RECT 269.54 56.565 269.75 56.635 ;
    RECT 269.54 56.925 269.75 56.995 ;
    RECT 233.48 56.205 233.69 56.275 ;
    RECT 233.48 56.565 233.69 56.635 ;
    RECT 233.48 56.925 233.69 56.995 ;
    RECT 233.02 56.205 233.23 56.275 ;
    RECT 233.02 56.565 233.23 56.635 ;
    RECT 233.02 56.925 233.23 56.995 ;
    RECT 230.16 56.205 230.37 56.275 ;
    RECT 230.16 56.565 230.37 56.635 ;
    RECT 230.16 56.925 230.37 56.995 ;
    RECT 229.7 56.205 229.91 56.275 ;
    RECT 229.7 56.565 229.91 56.635 ;
    RECT 229.7 56.925 229.91 56.995 ;
    RECT 366.28 56.205 366.49 56.275 ;
    RECT 366.28 56.565 366.49 56.635 ;
    RECT 366.28 56.925 366.49 56.995 ;
    RECT 365.82 56.205 366.03 56.275 ;
    RECT 365.82 56.565 366.03 56.635 ;
    RECT 365.82 56.925 366.03 56.995 ;
    RECT 226.84 56.205 227.05 56.275 ;
    RECT 226.84 56.565 227.05 56.635 ;
    RECT 226.84 56.925 227.05 56.995 ;
    RECT 226.38 56.205 226.59 56.275 ;
    RECT 226.38 56.565 226.59 56.635 ;
    RECT 226.38 56.925 226.59 56.995 ;
    RECT 362.96 56.205 363.17 56.275 ;
    RECT 362.96 56.565 363.17 56.635 ;
    RECT 362.96 56.925 363.17 56.995 ;
    RECT 362.5 56.205 362.71 56.275 ;
    RECT 362.5 56.565 362.71 56.635 ;
    RECT 362.5 56.925 362.71 56.995 ;
    RECT 223.52 56.205 223.73 56.275 ;
    RECT 223.52 56.565 223.73 56.635 ;
    RECT 223.52 56.925 223.73 56.995 ;
    RECT 223.06 56.205 223.27 56.275 ;
    RECT 223.06 56.565 223.27 56.635 ;
    RECT 223.06 56.925 223.27 56.995 ;
    RECT 359.64 56.205 359.85 56.275 ;
    RECT 359.64 56.565 359.85 56.635 ;
    RECT 359.64 56.925 359.85 56.995 ;
    RECT 359.18 56.205 359.39 56.275 ;
    RECT 359.18 56.565 359.39 56.635 ;
    RECT 359.18 56.925 359.39 56.995 ;
    RECT 220.2 56.205 220.41 56.275 ;
    RECT 220.2 56.565 220.41 56.635 ;
    RECT 220.2 56.925 220.41 56.995 ;
    RECT 219.74 56.205 219.95 56.275 ;
    RECT 219.74 56.565 219.95 56.635 ;
    RECT 219.74 56.925 219.95 56.995 ;
    RECT 356.32 56.205 356.53 56.275 ;
    RECT 356.32 56.565 356.53 56.635 ;
    RECT 356.32 56.925 356.53 56.995 ;
    RECT 355.86 56.205 356.07 56.275 ;
    RECT 355.86 56.565 356.07 56.635 ;
    RECT 355.86 56.925 356.07 56.995 ;
    RECT 353.0 56.205 353.21 56.275 ;
    RECT 353.0 56.565 353.21 56.635 ;
    RECT 353.0 56.925 353.21 56.995 ;
    RECT 352.54 56.205 352.75 56.275 ;
    RECT 352.54 56.565 352.75 56.635 ;
    RECT 352.54 56.925 352.75 56.995 ;
    RECT 216.88 56.205 217.09 56.275 ;
    RECT 216.88 56.565 217.09 56.635 ;
    RECT 216.88 56.925 217.09 56.995 ;
    RECT 216.42 56.205 216.63 56.275 ;
    RECT 216.42 56.565 216.63 56.635 ;
    RECT 216.42 56.925 216.63 56.995 ;
    RECT 349.68 56.205 349.89 56.275 ;
    RECT 349.68 56.565 349.89 56.635 ;
    RECT 349.68 56.925 349.89 56.995 ;
    RECT 349.22 56.205 349.43 56.275 ;
    RECT 349.22 56.565 349.43 56.635 ;
    RECT 349.22 56.925 349.43 56.995 ;
    RECT 213.56 56.205 213.77 56.275 ;
    RECT 213.56 56.565 213.77 56.635 ;
    RECT 213.56 56.925 213.77 56.995 ;
    RECT 213.1 56.205 213.31 56.275 ;
    RECT 213.1 56.565 213.31 56.635 ;
    RECT 213.1 56.925 213.31 56.995 ;
    RECT 346.36 56.205 346.57 56.275 ;
    RECT 346.36 56.565 346.57 56.635 ;
    RECT 346.36 56.925 346.57 56.995 ;
    RECT 345.9 56.205 346.11 56.275 ;
    RECT 345.9 56.565 346.11 56.635 ;
    RECT 345.9 56.925 346.11 56.995 ;
    RECT 210.24 56.205 210.45 56.275 ;
    RECT 210.24 56.565 210.45 56.635 ;
    RECT 210.24 56.925 210.45 56.995 ;
    RECT 209.78 56.205 209.99 56.275 ;
    RECT 209.78 56.565 209.99 56.635 ;
    RECT 209.78 56.925 209.99 56.995 ;
    RECT 343.04 56.205 343.25 56.275 ;
    RECT 343.04 56.565 343.25 56.635 ;
    RECT 343.04 56.925 343.25 56.995 ;
    RECT 342.58 56.205 342.79 56.275 ;
    RECT 342.58 56.565 342.79 56.635 ;
    RECT 342.58 56.925 342.79 56.995 ;
    RECT 206.92 56.205 207.13 56.275 ;
    RECT 206.92 56.565 207.13 56.635 ;
    RECT 206.92 56.925 207.13 56.995 ;
    RECT 206.46 56.205 206.67 56.275 ;
    RECT 206.46 56.565 206.67 56.635 ;
    RECT 206.46 56.925 206.67 56.995 ;
    RECT 339.72 56.205 339.93 56.275 ;
    RECT 339.72 56.565 339.93 56.635 ;
    RECT 339.72 56.925 339.93 56.995 ;
    RECT 339.26 56.205 339.47 56.275 ;
    RECT 339.26 56.565 339.47 56.635 ;
    RECT 339.26 56.925 339.47 56.995 ;
    RECT 203.6 56.205 203.81 56.275 ;
    RECT 203.6 56.565 203.81 56.635 ;
    RECT 203.6 56.925 203.81 56.995 ;
    RECT 203.14 56.205 203.35 56.275 ;
    RECT 203.14 56.565 203.35 56.635 ;
    RECT 203.14 56.925 203.35 56.995 ;
    RECT 336.4 56.205 336.61 56.275 ;
    RECT 336.4 56.565 336.61 56.635 ;
    RECT 336.4 56.925 336.61 56.995 ;
    RECT 335.94 56.205 336.15 56.275 ;
    RECT 335.94 56.565 336.15 56.635 ;
    RECT 335.94 56.925 336.15 56.995 ;
    RECT 266.68 56.205 266.89 56.275 ;
    RECT 266.68 56.565 266.89 56.635 ;
    RECT 266.68 56.925 266.89 56.995 ;
    RECT 266.22 56.205 266.43 56.275 ;
    RECT 266.22 56.565 266.43 56.635 ;
    RECT 266.22 56.925 266.43 56.995 ;
    RECT 263.36 56.205 263.57 56.275 ;
    RECT 263.36 56.565 263.57 56.635 ;
    RECT 263.36 56.925 263.57 56.995 ;
    RECT 262.9 56.205 263.11 56.275 ;
    RECT 262.9 56.565 263.11 56.635 ;
    RECT 262.9 56.925 263.11 56.995 ;
    RECT 260.04 56.205 260.25 56.275 ;
    RECT 260.04 56.565 260.25 56.635 ;
    RECT 260.04 56.925 260.25 56.995 ;
    RECT 259.58 56.205 259.79 56.275 ;
    RECT 259.58 56.565 259.79 56.635 ;
    RECT 259.58 56.925 259.79 56.995 ;
    RECT 256.72 56.205 256.93 56.275 ;
    RECT 256.72 56.565 256.93 56.635 ;
    RECT 256.72 56.925 256.93 56.995 ;
    RECT 256.26 56.205 256.47 56.275 ;
    RECT 256.26 56.565 256.47 56.635 ;
    RECT 256.26 56.925 256.47 56.995 ;
    RECT 253.4 56.205 253.61 56.275 ;
    RECT 253.4 56.565 253.61 56.635 ;
    RECT 253.4 56.925 253.61 56.995 ;
    RECT 252.94 56.205 253.15 56.275 ;
    RECT 252.94 56.565 253.15 56.635 ;
    RECT 252.94 56.925 253.15 56.995 ;
    RECT 250.08 56.205 250.29 56.275 ;
    RECT 250.08 56.565 250.29 56.635 ;
    RECT 250.08 56.925 250.29 56.995 ;
    RECT 249.62 56.205 249.83 56.275 ;
    RECT 249.62 56.565 249.83 56.635 ;
    RECT 249.62 56.925 249.83 56.995 ;
    RECT 246.76 56.205 246.97 56.275 ;
    RECT 246.76 56.565 246.97 56.635 ;
    RECT 246.76 56.925 246.97 56.995 ;
    RECT 246.3 56.205 246.51 56.275 ;
    RECT 246.3 56.565 246.51 56.635 ;
    RECT 246.3 56.925 246.51 56.995 ;
    RECT 243.44 56.205 243.65 56.275 ;
    RECT 243.44 56.565 243.65 56.635 ;
    RECT 243.44 56.925 243.65 56.995 ;
    RECT 242.98 56.205 243.19 56.275 ;
    RECT 242.98 56.565 243.19 56.635 ;
    RECT 242.98 56.925 243.19 56.995 ;
    RECT 240.12 56.205 240.33 56.275 ;
    RECT 240.12 56.565 240.33 56.635 ;
    RECT 240.12 56.925 240.33 56.995 ;
    RECT 239.66 56.205 239.87 56.275 ;
    RECT 239.66 56.565 239.87 56.635 ;
    RECT 239.66 56.925 239.87 56.995 ;
    RECT 236.8 56.205 237.01 56.275 ;
    RECT 236.8 56.565 237.01 56.635 ;
    RECT 236.8 56.925 237.01 56.995 ;
    RECT 236.34 56.205 236.55 56.275 ;
    RECT 236.34 56.565 236.55 56.635 ;
    RECT 236.34 56.925 236.55 56.995 ;
    RECT 374.15 56.565 374.22 56.635 ;
    RECT 333.08 56.205 333.29 56.275 ;
    RECT 333.08 56.565 333.29 56.635 ;
    RECT 333.08 56.925 333.29 56.995 ;
    RECT 332.62 56.205 332.83 56.275 ;
    RECT 332.62 56.565 332.83 56.635 ;
    RECT 332.62 56.925 332.83 56.995 ;
    RECT 329.76 56.205 329.97 56.275 ;
    RECT 329.76 56.565 329.97 56.635 ;
    RECT 329.76 56.925 329.97 56.995 ;
    RECT 329.3 56.205 329.51 56.275 ;
    RECT 329.3 56.565 329.51 56.635 ;
    RECT 329.3 56.925 329.51 56.995 ;
    RECT 326.44 56.205 326.65 56.275 ;
    RECT 326.44 56.565 326.65 56.635 ;
    RECT 326.44 56.925 326.65 56.995 ;
    RECT 325.98 56.205 326.19 56.275 ;
    RECT 325.98 56.565 326.19 56.635 ;
    RECT 325.98 56.925 326.19 56.995 ;
    RECT 323.12 56.205 323.33 56.275 ;
    RECT 323.12 56.565 323.33 56.635 ;
    RECT 323.12 56.925 323.33 56.995 ;
    RECT 322.66 56.205 322.87 56.275 ;
    RECT 322.66 56.565 322.87 56.635 ;
    RECT 322.66 56.925 322.87 56.995 ;
    RECT 319.8 56.205 320.01 56.275 ;
    RECT 319.8 56.565 320.01 56.635 ;
    RECT 319.8 56.925 320.01 56.995 ;
    RECT 319.34 56.205 319.55 56.275 ;
    RECT 319.34 56.565 319.55 56.635 ;
    RECT 319.34 56.925 319.55 56.995 ;
    RECT 316.48 56.205 316.69 56.275 ;
    RECT 316.48 56.565 316.69 56.635 ;
    RECT 316.48 56.925 316.69 56.995 ;
    RECT 316.02 56.205 316.23 56.275 ;
    RECT 316.02 56.565 316.23 56.635 ;
    RECT 316.02 56.925 316.23 56.995 ;
    RECT 313.16 56.205 313.37 56.275 ;
    RECT 313.16 56.565 313.37 56.635 ;
    RECT 313.16 56.925 313.37 56.995 ;
    RECT 312.7 56.205 312.91 56.275 ;
    RECT 312.7 56.565 312.91 56.635 ;
    RECT 312.7 56.925 312.91 56.995 ;
    RECT 309.84 56.205 310.05 56.275 ;
    RECT 309.84 56.565 310.05 56.635 ;
    RECT 309.84 56.925 310.05 56.995 ;
    RECT 309.38 56.205 309.59 56.275 ;
    RECT 309.38 56.565 309.59 56.635 ;
    RECT 309.38 56.925 309.59 56.995 ;
    RECT 306.52 56.205 306.73 56.275 ;
    RECT 306.52 56.565 306.73 56.635 ;
    RECT 306.52 56.925 306.73 56.995 ;
    RECT 306.06 56.205 306.27 56.275 ;
    RECT 306.06 56.565 306.27 56.635 ;
    RECT 306.06 56.925 306.27 56.995 ;
    RECT 303.2 55.485 303.41 55.555 ;
    RECT 303.2 55.845 303.41 55.915 ;
    RECT 303.2 56.205 303.41 56.275 ;
    RECT 302.74 55.485 302.95 55.555 ;
    RECT 302.74 55.845 302.95 55.915 ;
    RECT 302.74 56.205 302.95 56.275 ;
    RECT 372.92 55.485 373.13 55.555 ;
    RECT 372.92 55.845 373.13 55.915 ;
    RECT 372.92 56.205 373.13 56.275 ;
    RECT 372.46 55.485 372.67 55.555 ;
    RECT 372.46 55.845 372.67 55.915 ;
    RECT 372.46 56.205 372.67 56.275 ;
    RECT 369.6 55.485 369.81 55.555 ;
    RECT 369.6 55.845 369.81 55.915 ;
    RECT 369.6 56.205 369.81 56.275 ;
    RECT 369.14 55.485 369.35 55.555 ;
    RECT 369.14 55.845 369.35 55.915 ;
    RECT 369.14 56.205 369.35 56.275 ;
    RECT 200.605 55.845 200.675 55.915 ;
    RECT 299.88 55.485 300.09 55.555 ;
    RECT 299.88 55.845 300.09 55.915 ;
    RECT 299.88 56.205 300.09 56.275 ;
    RECT 299.42 55.485 299.63 55.555 ;
    RECT 299.42 55.845 299.63 55.915 ;
    RECT 299.42 56.205 299.63 56.275 ;
    RECT 296.56 55.485 296.77 55.555 ;
    RECT 296.56 55.845 296.77 55.915 ;
    RECT 296.56 56.205 296.77 56.275 ;
    RECT 296.1 55.485 296.31 55.555 ;
    RECT 296.1 55.845 296.31 55.915 ;
    RECT 296.1 56.205 296.31 56.275 ;
    RECT 293.24 55.485 293.45 55.555 ;
    RECT 293.24 55.845 293.45 55.915 ;
    RECT 293.24 56.205 293.45 56.275 ;
    RECT 292.78 55.485 292.99 55.555 ;
    RECT 292.78 55.845 292.99 55.915 ;
    RECT 292.78 56.205 292.99 56.275 ;
    RECT 289.92 55.485 290.13 55.555 ;
    RECT 289.92 55.845 290.13 55.915 ;
    RECT 289.92 56.205 290.13 56.275 ;
    RECT 289.46 55.485 289.67 55.555 ;
    RECT 289.46 55.845 289.67 55.915 ;
    RECT 289.46 56.205 289.67 56.275 ;
    RECT 286.6 55.485 286.81 55.555 ;
    RECT 286.6 55.845 286.81 55.915 ;
    RECT 286.6 56.205 286.81 56.275 ;
    RECT 286.14 55.485 286.35 55.555 ;
    RECT 286.14 55.845 286.35 55.915 ;
    RECT 286.14 56.205 286.35 56.275 ;
    RECT 283.28 55.485 283.49 55.555 ;
    RECT 283.28 55.845 283.49 55.915 ;
    RECT 283.28 56.205 283.49 56.275 ;
    RECT 282.82 55.485 283.03 55.555 ;
    RECT 282.82 55.845 283.03 55.915 ;
    RECT 282.82 56.205 283.03 56.275 ;
    RECT 279.96 55.485 280.17 55.555 ;
    RECT 279.96 55.845 280.17 55.915 ;
    RECT 279.96 56.205 280.17 56.275 ;
    RECT 279.5 55.485 279.71 55.555 ;
    RECT 279.5 55.845 279.71 55.915 ;
    RECT 279.5 56.205 279.71 56.275 ;
    RECT 276.64 55.485 276.85 55.555 ;
    RECT 276.64 55.845 276.85 55.915 ;
    RECT 276.64 56.205 276.85 56.275 ;
    RECT 276.18 55.485 276.39 55.555 ;
    RECT 276.18 55.845 276.39 55.915 ;
    RECT 276.18 56.205 276.39 56.275 ;
    RECT 273.32 55.485 273.53 55.555 ;
    RECT 273.32 55.845 273.53 55.915 ;
    RECT 273.32 56.205 273.53 56.275 ;
    RECT 272.86 55.485 273.07 55.555 ;
    RECT 272.86 55.845 273.07 55.915 ;
    RECT 272.86 56.205 273.07 56.275 ;
    RECT 270.0 55.485 270.21 55.555 ;
    RECT 270.0 55.845 270.21 55.915 ;
    RECT 270.0 56.205 270.21 56.275 ;
    RECT 269.54 55.485 269.75 55.555 ;
    RECT 269.54 55.845 269.75 55.915 ;
    RECT 269.54 56.205 269.75 56.275 ;
    RECT 233.48 55.485 233.69 55.555 ;
    RECT 233.48 55.845 233.69 55.915 ;
    RECT 233.48 56.205 233.69 56.275 ;
    RECT 233.02 55.485 233.23 55.555 ;
    RECT 233.02 55.845 233.23 55.915 ;
    RECT 233.02 56.205 233.23 56.275 ;
    RECT 230.16 55.485 230.37 55.555 ;
    RECT 230.16 55.845 230.37 55.915 ;
    RECT 230.16 56.205 230.37 56.275 ;
    RECT 229.7 55.485 229.91 55.555 ;
    RECT 229.7 55.845 229.91 55.915 ;
    RECT 229.7 56.205 229.91 56.275 ;
    RECT 366.28 55.485 366.49 55.555 ;
    RECT 366.28 55.845 366.49 55.915 ;
    RECT 366.28 56.205 366.49 56.275 ;
    RECT 365.82 55.485 366.03 55.555 ;
    RECT 365.82 55.845 366.03 55.915 ;
    RECT 365.82 56.205 366.03 56.275 ;
    RECT 226.84 55.485 227.05 55.555 ;
    RECT 226.84 55.845 227.05 55.915 ;
    RECT 226.84 56.205 227.05 56.275 ;
    RECT 226.38 55.485 226.59 55.555 ;
    RECT 226.38 55.845 226.59 55.915 ;
    RECT 226.38 56.205 226.59 56.275 ;
    RECT 362.96 55.485 363.17 55.555 ;
    RECT 362.96 55.845 363.17 55.915 ;
    RECT 362.96 56.205 363.17 56.275 ;
    RECT 362.5 55.485 362.71 55.555 ;
    RECT 362.5 55.845 362.71 55.915 ;
    RECT 362.5 56.205 362.71 56.275 ;
    RECT 223.52 55.485 223.73 55.555 ;
    RECT 223.52 55.845 223.73 55.915 ;
    RECT 223.52 56.205 223.73 56.275 ;
    RECT 223.06 55.485 223.27 55.555 ;
    RECT 223.06 55.845 223.27 55.915 ;
    RECT 223.06 56.205 223.27 56.275 ;
    RECT 359.64 55.485 359.85 55.555 ;
    RECT 359.64 55.845 359.85 55.915 ;
    RECT 359.64 56.205 359.85 56.275 ;
    RECT 359.18 55.485 359.39 55.555 ;
    RECT 359.18 55.845 359.39 55.915 ;
    RECT 359.18 56.205 359.39 56.275 ;
    RECT 220.2 55.485 220.41 55.555 ;
    RECT 220.2 55.845 220.41 55.915 ;
    RECT 220.2 56.205 220.41 56.275 ;
    RECT 219.74 55.485 219.95 55.555 ;
    RECT 219.74 55.845 219.95 55.915 ;
    RECT 219.74 56.205 219.95 56.275 ;
    RECT 356.32 55.485 356.53 55.555 ;
    RECT 356.32 55.845 356.53 55.915 ;
    RECT 356.32 56.205 356.53 56.275 ;
    RECT 355.86 55.485 356.07 55.555 ;
    RECT 355.86 55.845 356.07 55.915 ;
    RECT 355.86 56.205 356.07 56.275 ;
    RECT 353.0 55.485 353.21 55.555 ;
    RECT 353.0 55.845 353.21 55.915 ;
    RECT 353.0 56.205 353.21 56.275 ;
    RECT 352.54 55.485 352.75 55.555 ;
    RECT 352.54 55.845 352.75 55.915 ;
    RECT 352.54 56.205 352.75 56.275 ;
    RECT 216.88 55.485 217.09 55.555 ;
    RECT 216.88 55.845 217.09 55.915 ;
    RECT 216.88 56.205 217.09 56.275 ;
    RECT 216.42 55.485 216.63 55.555 ;
    RECT 216.42 55.845 216.63 55.915 ;
    RECT 216.42 56.205 216.63 56.275 ;
    RECT 349.68 55.485 349.89 55.555 ;
    RECT 349.68 55.845 349.89 55.915 ;
    RECT 349.68 56.205 349.89 56.275 ;
    RECT 349.22 55.485 349.43 55.555 ;
    RECT 349.22 55.845 349.43 55.915 ;
    RECT 349.22 56.205 349.43 56.275 ;
    RECT 213.56 55.485 213.77 55.555 ;
    RECT 213.56 55.845 213.77 55.915 ;
    RECT 213.56 56.205 213.77 56.275 ;
    RECT 213.1 55.485 213.31 55.555 ;
    RECT 213.1 55.845 213.31 55.915 ;
    RECT 213.1 56.205 213.31 56.275 ;
    RECT 346.36 55.485 346.57 55.555 ;
    RECT 346.36 55.845 346.57 55.915 ;
    RECT 346.36 56.205 346.57 56.275 ;
    RECT 345.9 55.485 346.11 55.555 ;
    RECT 345.9 55.845 346.11 55.915 ;
    RECT 345.9 56.205 346.11 56.275 ;
    RECT 210.24 55.485 210.45 55.555 ;
    RECT 210.24 55.845 210.45 55.915 ;
    RECT 210.24 56.205 210.45 56.275 ;
    RECT 209.78 55.485 209.99 55.555 ;
    RECT 209.78 55.845 209.99 55.915 ;
    RECT 209.78 56.205 209.99 56.275 ;
    RECT 343.04 55.485 343.25 55.555 ;
    RECT 343.04 55.845 343.25 55.915 ;
    RECT 343.04 56.205 343.25 56.275 ;
    RECT 342.58 55.485 342.79 55.555 ;
    RECT 342.58 55.845 342.79 55.915 ;
    RECT 342.58 56.205 342.79 56.275 ;
    RECT 206.92 55.485 207.13 55.555 ;
    RECT 206.92 55.845 207.13 55.915 ;
    RECT 206.92 56.205 207.13 56.275 ;
    RECT 206.46 55.485 206.67 55.555 ;
    RECT 206.46 55.845 206.67 55.915 ;
    RECT 206.46 56.205 206.67 56.275 ;
    RECT 339.72 55.485 339.93 55.555 ;
    RECT 339.72 55.845 339.93 55.915 ;
    RECT 339.72 56.205 339.93 56.275 ;
    RECT 339.26 55.485 339.47 55.555 ;
    RECT 339.26 55.845 339.47 55.915 ;
    RECT 339.26 56.205 339.47 56.275 ;
    RECT 203.6 55.485 203.81 55.555 ;
    RECT 203.6 55.845 203.81 55.915 ;
    RECT 203.6 56.205 203.81 56.275 ;
    RECT 203.14 55.485 203.35 55.555 ;
    RECT 203.14 55.845 203.35 55.915 ;
    RECT 203.14 56.205 203.35 56.275 ;
    RECT 336.4 55.485 336.61 55.555 ;
    RECT 336.4 55.845 336.61 55.915 ;
    RECT 336.4 56.205 336.61 56.275 ;
    RECT 335.94 55.485 336.15 55.555 ;
    RECT 335.94 55.845 336.15 55.915 ;
    RECT 335.94 56.205 336.15 56.275 ;
    RECT 266.68 55.485 266.89 55.555 ;
    RECT 266.68 55.845 266.89 55.915 ;
    RECT 266.68 56.205 266.89 56.275 ;
    RECT 266.22 55.485 266.43 55.555 ;
    RECT 266.22 55.845 266.43 55.915 ;
    RECT 266.22 56.205 266.43 56.275 ;
    RECT 263.36 55.485 263.57 55.555 ;
    RECT 263.36 55.845 263.57 55.915 ;
    RECT 263.36 56.205 263.57 56.275 ;
    RECT 262.9 55.485 263.11 55.555 ;
    RECT 262.9 55.845 263.11 55.915 ;
    RECT 262.9 56.205 263.11 56.275 ;
    RECT 260.04 55.485 260.25 55.555 ;
    RECT 260.04 55.845 260.25 55.915 ;
    RECT 260.04 56.205 260.25 56.275 ;
    RECT 259.58 55.485 259.79 55.555 ;
    RECT 259.58 55.845 259.79 55.915 ;
    RECT 259.58 56.205 259.79 56.275 ;
    RECT 256.72 55.485 256.93 55.555 ;
    RECT 256.72 55.845 256.93 55.915 ;
    RECT 256.72 56.205 256.93 56.275 ;
    RECT 256.26 55.485 256.47 55.555 ;
    RECT 256.26 55.845 256.47 55.915 ;
    RECT 256.26 56.205 256.47 56.275 ;
    RECT 253.4 55.485 253.61 55.555 ;
    RECT 253.4 55.845 253.61 55.915 ;
    RECT 253.4 56.205 253.61 56.275 ;
    RECT 252.94 55.485 253.15 55.555 ;
    RECT 252.94 55.845 253.15 55.915 ;
    RECT 252.94 56.205 253.15 56.275 ;
    RECT 250.08 55.485 250.29 55.555 ;
    RECT 250.08 55.845 250.29 55.915 ;
    RECT 250.08 56.205 250.29 56.275 ;
    RECT 249.62 55.485 249.83 55.555 ;
    RECT 249.62 55.845 249.83 55.915 ;
    RECT 249.62 56.205 249.83 56.275 ;
    RECT 246.76 55.485 246.97 55.555 ;
    RECT 246.76 55.845 246.97 55.915 ;
    RECT 246.76 56.205 246.97 56.275 ;
    RECT 246.3 55.485 246.51 55.555 ;
    RECT 246.3 55.845 246.51 55.915 ;
    RECT 246.3 56.205 246.51 56.275 ;
    RECT 243.44 55.485 243.65 55.555 ;
    RECT 243.44 55.845 243.65 55.915 ;
    RECT 243.44 56.205 243.65 56.275 ;
    RECT 242.98 55.485 243.19 55.555 ;
    RECT 242.98 55.845 243.19 55.915 ;
    RECT 242.98 56.205 243.19 56.275 ;
    RECT 240.12 55.485 240.33 55.555 ;
    RECT 240.12 55.845 240.33 55.915 ;
    RECT 240.12 56.205 240.33 56.275 ;
    RECT 239.66 55.485 239.87 55.555 ;
    RECT 239.66 55.845 239.87 55.915 ;
    RECT 239.66 56.205 239.87 56.275 ;
    RECT 236.8 55.485 237.01 55.555 ;
    RECT 236.8 55.845 237.01 55.915 ;
    RECT 236.8 56.205 237.01 56.275 ;
    RECT 236.34 55.485 236.55 55.555 ;
    RECT 236.34 55.845 236.55 55.915 ;
    RECT 236.34 56.205 236.55 56.275 ;
    RECT 374.15 55.845 374.22 55.915 ;
    RECT 333.08 55.485 333.29 55.555 ;
    RECT 333.08 55.845 333.29 55.915 ;
    RECT 333.08 56.205 333.29 56.275 ;
    RECT 332.62 55.485 332.83 55.555 ;
    RECT 332.62 55.845 332.83 55.915 ;
    RECT 332.62 56.205 332.83 56.275 ;
    RECT 329.76 55.485 329.97 55.555 ;
    RECT 329.76 55.845 329.97 55.915 ;
    RECT 329.76 56.205 329.97 56.275 ;
    RECT 329.3 55.485 329.51 55.555 ;
    RECT 329.3 55.845 329.51 55.915 ;
    RECT 329.3 56.205 329.51 56.275 ;
    RECT 326.44 55.485 326.65 55.555 ;
    RECT 326.44 55.845 326.65 55.915 ;
    RECT 326.44 56.205 326.65 56.275 ;
    RECT 325.98 55.485 326.19 55.555 ;
    RECT 325.98 55.845 326.19 55.915 ;
    RECT 325.98 56.205 326.19 56.275 ;
    RECT 323.12 55.485 323.33 55.555 ;
    RECT 323.12 55.845 323.33 55.915 ;
    RECT 323.12 56.205 323.33 56.275 ;
    RECT 322.66 55.485 322.87 55.555 ;
    RECT 322.66 55.845 322.87 55.915 ;
    RECT 322.66 56.205 322.87 56.275 ;
    RECT 319.8 55.485 320.01 55.555 ;
    RECT 319.8 55.845 320.01 55.915 ;
    RECT 319.8 56.205 320.01 56.275 ;
    RECT 319.34 55.485 319.55 55.555 ;
    RECT 319.34 55.845 319.55 55.915 ;
    RECT 319.34 56.205 319.55 56.275 ;
    RECT 316.48 55.485 316.69 55.555 ;
    RECT 316.48 55.845 316.69 55.915 ;
    RECT 316.48 56.205 316.69 56.275 ;
    RECT 316.02 55.485 316.23 55.555 ;
    RECT 316.02 55.845 316.23 55.915 ;
    RECT 316.02 56.205 316.23 56.275 ;
    RECT 313.16 55.485 313.37 55.555 ;
    RECT 313.16 55.845 313.37 55.915 ;
    RECT 313.16 56.205 313.37 56.275 ;
    RECT 312.7 55.485 312.91 55.555 ;
    RECT 312.7 55.845 312.91 55.915 ;
    RECT 312.7 56.205 312.91 56.275 ;
    RECT 309.84 55.485 310.05 55.555 ;
    RECT 309.84 55.845 310.05 55.915 ;
    RECT 309.84 56.205 310.05 56.275 ;
    RECT 309.38 55.485 309.59 55.555 ;
    RECT 309.38 55.845 309.59 55.915 ;
    RECT 309.38 56.205 309.59 56.275 ;
    RECT 306.52 55.485 306.73 55.555 ;
    RECT 306.52 55.845 306.73 55.915 ;
    RECT 306.52 56.205 306.73 56.275 ;
    RECT 306.06 55.485 306.27 55.555 ;
    RECT 306.06 55.845 306.27 55.915 ;
    RECT 306.06 56.205 306.27 56.275 ;
    RECT 303.2 54.765 303.41 54.835 ;
    RECT 303.2 55.125 303.41 55.195 ;
    RECT 303.2 55.485 303.41 55.555 ;
    RECT 302.74 54.765 302.95 54.835 ;
    RECT 302.74 55.125 302.95 55.195 ;
    RECT 302.74 55.485 302.95 55.555 ;
    RECT 372.92 54.765 373.13 54.835 ;
    RECT 372.92 55.125 373.13 55.195 ;
    RECT 372.92 55.485 373.13 55.555 ;
    RECT 372.46 54.765 372.67 54.835 ;
    RECT 372.46 55.125 372.67 55.195 ;
    RECT 372.46 55.485 372.67 55.555 ;
    RECT 369.6 54.765 369.81 54.835 ;
    RECT 369.6 55.125 369.81 55.195 ;
    RECT 369.6 55.485 369.81 55.555 ;
    RECT 369.14 54.765 369.35 54.835 ;
    RECT 369.14 55.125 369.35 55.195 ;
    RECT 369.14 55.485 369.35 55.555 ;
    RECT 200.605 55.125 200.675 55.195 ;
    RECT 299.88 54.765 300.09 54.835 ;
    RECT 299.88 55.125 300.09 55.195 ;
    RECT 299.88 55.485 300.09 55.555 ;
    RECT 299.42 54.765 299.63 54.835 ;
    RECT 299.42 55.125 299.63 55.195 ;
    RECT 299.42 55.485 299.63 55.555 ;
    RECT 296.56 54.765 296.77 54.835 ;
    RECT 296.56 55.125 296.77 55.195 ;
    RECT 296.56 55.485 296.77 55.555 ;
    RECT 296.1 54.765 296.31 54.835 ;
    RECT 296.1 55.125 296.31 55.195 ;
    RECT 296.1 55.485 296.31 55.555 ;
    RECT 293.24 54.765 293.45 54.835 ;
    RECT 293.24 55.125 293.45 55.195 ;
    RECT 293.24 55.485 293.45 55.555 ;
    RECT 292.78 54.765 292.99 54.835 ;
    RECT 292.78 55.125 292.99 55.195 ;
    RECT 292.78 55.485 292.99 55.555 ;
    RECT 289.92 54.765 290.13 54.835 ;
    RECT 289.92 55.125 290.13 55.195 ;
    RECT 289.92 55.485 290.13 55.555 ;
    RECT 289.46 54.765 289.67 54.835 ;
    RECT 289.46 55.125 289.67 55.195 ;
    RECT 289.46 55.485 289.67 55.555 ;
    RECT 286.6 54.765 286.81 54.835 ;
    RECT 286.6 55.125 286.81 55.195 ;
    RECT 286.6 55.485 286.81 55.555 ;
    RECT 286.14 54.765 286.35 54.835 ;
    RECT 286.14 55.125 286.35 55.195 ;
    RECT 286.14 55.485 286.35 55.555 ;
    RECT 283.28 54.765 283.49 54.835 ;
    RECT 283.28 55.125 283.49 55.195 ;
    RECT 283.28 55.485 283.49 55.555 ;
    RECT 282.82 54.765 283.03 54.835 ;
    RECT 282.82 55.125 283.03 55.195 ;
    RECT 282.82 55.485 283.03 55.555 ;
    RECT 279.96 54.765 280.17 54.835 ;
    RECT 279.96 55.125 280.17 55.195 ;
    RECT 279.96 55.485 280.17 55.555 ;
    RECT 279.5 54.765 279.71 54.835 ;
    RECT 279.5 55.125 279.71 55.195 ;
    RECT 279.5 55.485 279.71 55.555 ;
    RECT 276.64 54.765 276.85 54.835 ;
    RECT 276.64 55.125 276.85 55.195 ;
    RECT 276.64 55.485 276.85 55.555 ;
    RECT 276.18 54.765 276.39 54.835 ;
    RECT 276.18 55.125 276.39 55.195 ;
    RECT 276.18 55.485 276.39 55.555 ;
    RECT 273.32 54.765 273.53 54.835 ;
    RECT 273.32 55.125 273.53 55.195 ;
    RECT 273.32 55.485 273.53 55.555 ;
    RECT 272.86 54.765 273.07 54.835 ;
    RECT 272.86 55.125 273.07 55.195 ;
    RECT 272.86 55.485 273.07 55.555 ;
    RECT 270.0 54.765 270.21 54.835 ;
    RECT 270.0 55.125 270.21 55.195 ;
    RECT 270.0 55.485 270.21 55.555 ;
    RECT 269.54 54.765 269.75 54.835 ;
    RECT 269.54 55.125 269.75 55.195 ;
    RECT 269.54 55.485 269.75 55.555 ;
    RECT 233.48 54.765 233.69 54.835 ;
    RECT 233.48 55.125 233.69 55.195 ;
    RECT 233.48 55.485 233.69 55.555 ;
    RECT 233.02 54.765 233.23 54.835 ;
    RECT 233.02 55.125 233.23 55.195 ;
    RECT 233.02 55.485 233.23 55.555 ;
    RECT 230.16 54.765 230.37 54.835 ;
    RECT 230.16 55.125 230.37 55.195 ;
    RECT 230.16 55.485 230.37 55.555 ;
    RECT 229.7 54.765 229.91 54.835 ;
    RECT 229.7 55.125 229.91 55.195 ;
    RECT 229.7 55.485 229.91 55.555 ;
    RECT 366.28 54.765 366.49 54.835 ;
    RECT 366.28 55.125 366.49 55.195 ;
    RECT 366.28 55.485 366.49 55.555 ;
    RECT 365.82 54.765 366.03 54.835 ;
    RECT 365.82 55.125 366.03 55.195 ;
    RECT 365.82 55.485 366.03 55.555 ;
    RECT 226.84 54.765 227.05 54.835 ;
    RECT 226.84 55.125 227.05 55.195 ;
    RECT 226.84 55.485 227.05 55.555 ;
    RECT 226.38 54.765 226.59 54.835 ;
    RECT 226.38 55.125 226.59 55.195 ;
    RECT 226.38 55.485 226.59 55.555 ;
    RECT 362.96 54.765 363.17 54.835 ;
    RECT 362.96 55.125 363.17 55.195 ;
    RECT 362.96 55.485 363.17 55.555 ;
    RECT 362.5 54.765 362.71 54.835 ;
    RECT 362.5 55.125 362.71 55.195 ;
    RECT 362.5 55.485 362.71 55.555 ;
    RECT 223.52 54.765 223.73 54.835 ;
    RECT 223.52 55.125 223.73 55.195 ;
    RECT 223.52 55.485 223.73 55.555 ;
    RECT 223.06 54.765 223.27 54.835 ;
    RECT 223.06 55.125 223.27 55.195 ;
    RECT 223.06 55.485 223.27 55.555 ;
    RECT 359.64 54.765 359.85 54.835 ;
    RECT 359.64 55.125 359.85 55.195 ;
    RECT 359.64 55.485 359.85 55.555 ;
    RECT 359.18 54.765 359.39 54.835 ;
    RECT 359.18 55.125 359.39 55.195 ;
    RECT 359.18 55.485 359.39 55.555 ;
    RECT 220.2 54.765 220.41 54.835 ;
    RECT 220.2 55.125 220.41 55.195 ;
    RECT 220.2 55.485 220.41 55.555 ;
    RECT 219.74 54.765 219.95 54.835 ;
    RECT 219.74 55.125 219.95 55.195 ;
    RECT 219.74 55.485 219.95 55.555 ;
    RECT 356.32 54.765 356.53 54.835 ;
    RECT 356.32 55.125 356.53 55.195 ;
    RECT 356.32 55.485 356.53 55.555 ;
    RECT 355.86 54.765 356.07 54.835 ;
    RECT 355.86 55.125 356.07 55.195 ;
    RECT 355.86 55.485 356.07 55.555 ;
    RECT 353.0 54.765 353.21 54.835 ;
    RECT 353.0 55.125 353.21 55.195 ;
    RECT 353.0 55.485 353.21 55.555 ;
    RECT 352.54 54.765 352.75 54.835 ;
    RECT 352.54 55.125 352.75 55.195 ;
    RECT 352.54 55.485 352.75 55.555 ;
    RECT 216.88 54.765 217.09 54.835 ;
    RECT 216.88 55.125 217.09 55.195 ;
    RECT 216.88 55.485 217.09 55.555 ;
    RECT 216.42 54.765 216.63 54.835 ;
    RECT 216.42 55.125 216.63 55.195 ;
    RECT 216.42 55.485 216.63 55.555 ;
    RECT 349.68 54.765 349.89 54.835 ;
    RECT 349.68 55.125 349.89 55.195 ;
    RECT 349.68 55.485 349.89 55.555 ;
    RECT 349.22 54.765 349.43 54.835 ;
    RECT 349.22 55.125 349.43 55.195 ;
    RECT 349.22 55.485 349.43 55.555 ;
    RECT 213.56 54.765 213.77 54.835 ;
    RECT 213.56 55.125 213.77 55.195 ;
    RECT 213.56 55.485 213.77 55.555 ;
    RECT 213.1 54.765 213.31 54.835 ;
    RECT 213.1 55.125 213.31 55.195 ;
    RECT 213.1 55.485 213.31 55.555 ;
    RECT 346.36 54.765 346.57 54.835 ;
    RECT 346.36 55.125 346.57 55.195 ;
    RECT 346.36 55.485 346.57 55.555 ;
    RECT 345.9 54.765 346.11 54.835 ;
    RECT 345.9 55.125 346.11 55.195 ;
    RECT 345.9 55.485 346.11 55.555 ;
    RECT 210.24 54.765 210.45 54.835 ;
    RECT 210.24 55.125 210.45 55.195 ;
    RECT 210.24 55.485 210.45 55.555 ;
    RECT 209.78 54.765 209.99 54.835 ;
    RECT 209.78 55.125 209.99 55.195 ;
    RECT 209.78 55.485 209.99 55.555 ;
    RECT 343.04 54.765 343.25 54.835 ;
    RECT 343.04 55.125 343.25 55.195 ;
    RECT 343.04 55.485 343.25 55.555 ;
    RECT 342.58 54.765 342.79 54.835 ;
    RECT 342.58 55.125 342.79 55.195 ;
    RECT 342.58 55.485 342.79 55.555 ;
    RECT 206.92 54.765 207.13 54.835 ;
    RECT 206.92 55.125 207.13 55.195 ;
    RECT 206.92 55.485 207.13 55.555 ;
    RECT 206.46 54.765 206.67 54.835 ;
    RECT 206.46 55.125 206.67 55.195 ;
    RECT 206.46 55.485 206.67 55.555 ;
    RECT 339.72 54.765 339.93 54.835 ;
    RECT 339.72 55.125 339.93 55.195 ;
    RECT 339.72 55.485 339.93 55.555 ;
    RECT 339.26 54.765 339.47 54.835 ;
    RECT 339.26 55.125 339.47 55.195 ;
    RECT 339.26 55.485 339.47 55.555 ;
    RECT 203.6 54.765 203.81 54.835 ;
    RECT 203.6 55.125 203.81 55.195 ;
    RECT 203.6 55.485 203.81 55.555 ;
    RECT 203.14 54.765 203.35 54.835 ;
    RECT 203.14 55.125 203.35 55.195 ;
    RECT 203.14 55.485 203.35 55.555 ;
    RECT 336.4 54.765 336.61 54.835 ;
    RECT 336.4 55.125 336.61 55.195 ;
    RECT 336.4 55.485 336.61 55.555 ;
    RECT 335.94 54.765 336.15 54.835 ;
    RECT 335.94 55.125 336.15 55.195 ;
    RECT 335.94 55.485 336.15 55.555 ;
    RECT 266.68 54.765 266.89 54.835 ;
    RECT 266.68 55.125 266.89 55.195 ;
    RECT 266.68 55.485 266.89 55.555 ;
    RECT 266.22 54.765 266.43 54.835 ;
    RECT 266.22 55.125 266.43 55.195 ;
    RECT 266.22 55.485 266.43 55.555 ;
    RECT 263.36 54.765 263.57 54.835 ;
    RECT 263.36 55.125 263.57 55.195 ;
    RECT 263.36 55.485 263.57 55.555 ;
    RECT 262.9 54.765 263.11 54.835 ;
    RECT 262.9 55.125 263.11 55.195 ;
    RECT 262.9 55.485 263.11 55.555 ;
    RECT 260.04 54.765 260.25 54.835 ;
    RECT 260.04 55.125 260.25 55.195 ;
    RECT 260.04 55.485 260.25 55.555 ;
    RECT 259.58 54.765 259.79 54.835 ;
    RECT 259.58 55.125 259.79 55.195 ;
    RECT 259.58 55.485 259.79 55.555 ;
    RECT 256.72 54.765 256.93 54.835 ;
    RECT 256.72 55.125 256.93 55.195 ;
    RECT 256.72 55.485 256.93 55.555 ;
    RECT 256.26 54.765 256.47 54.835 ;
    RECT 256.26 55.125 256.47 55.195 ;
    RECT 256.26 55.485 256.47 55.555 ;
    RECT 253.4 54.765 253.61 54.835 ;
    RECT 253.4 55.125 253.61 55.195 ;
    RECT 253.4 55.485 253.61 55.555 ;
    RECT 252.94 54.765 253.15 54.835 ;
    RECT 252.94 55.125 253.15 55.195 ;
    RECT 252.94 55.485 253.15 55.555 ;
    RECT 250.08 54.765 250.29 54.835 ;
    RECT 250.08 55.125 250.29 55.195 ;
    RECT 250.08 55.485 250.29 55.555 ;
    RECT 249.62 54.765 249.83 54.835 ;
    RECT 249.62 55.125 249.83 55.195 ;
    RECT 249.62 55.485 249.83 55.555 ;
    RECT 246.76 54.765 246.97 54.835 ;
    RECT 246.76 55.125 246.97 55.195 ;
    RECT 246.76 55.485 246.97 55.555 ;
    RECT 246.3 54.765 246.51 54.835 ;
    RECT 246.3 55.125 246.51 55.195 ;
    RECT 246.3 55.485 246.51 55.555 ;
    RECT 243.44 54.765 243.65 54.835 ;
    RECT 243.44 55.125 243.65 55.195 ;
    RECT 243.44 55.485 243.65 55.555 ;
    RECT 242.98 54.765 243.19 54.835 ;
    RECT 242.98 55.125 243.19 55.195 ;
    RECT 242.98 55.485 243.19 55.555 ;
    RECT 240.12 54.765 240.33 54.835 ;
    RECT 240.12 55.125 240.33 55.195 ;
    RECT 240.12 55.485 240.33 55.555 ;
    RECT 239.66 54.765 239.87 54.835 ;
    RECT 239.66 55.125 239.87 55.195 ;
    RECT 239.66 55.485 239.87 55.555 ;
    RECT 236.8 54.765 237.01 54.835 ;
    RECT 236.8 55.125 237.01 55.195 ;
    RECT 236.8 55.485 237.01 55.555 ;
    RECT 236.34 54.765 236.55 54.835 ;
    RECT 236.34 55.125 236.55 55.195 ;
    RECT 236.34 55.485 236.55 55.555 ;
    RECT 374.15 55.125 374.22 55.195 ;
    RECT 333.08 54.765 333.29 54.835 ;
    RECT 333.08 55.125 333.29 55.195 ;
    RECT 333.08 55.485 333.29 55.555 ;
    RECT 332.62 54.765 332.83 54.835 ;
    RECT 332.62 55.125 332.83 55.195 ;
    RECT 332.62 55.485 332.83 55.555 ;
    RECT 329.76 54.765 329.97 54.835 ;
    RECT 329.76 55.125 329.97 55.195 ;
    RECT 329.76 55.485 329.97 55.555 ;
    RECT 329.3 54.765 329.51 54.835 ;
    RECT 329.3 55.125 329.51 55.195 ;
    RECT 329.3 55.485 329.51 55.555 ;
    RECT 326.44 54.765 326.65 54.835 ;
    RECT 326.44 55.125 326.65 55.195 ;
    RECT 326.44 55.485 326.65 55.555 ;
    RECT 325.98 54.765 326.19 54.835 ;
    RECT 325.98 55.125 326.19 55.195 ;
    RECT 325.98 55.485 326.19 55.555 ;
    RECT 323.12 54.765 323.33 54.835 ;
    RECT 323.12 55.125 323.33 55.195 ;
    RECT 323.12 55.485 323.33 55.555 ;
    RECT 322.66 54.765 322.87 54.835 ;
    RECT 322.66 55.125 322.87 55.195 ;
    RECT 322.66 55.485 322.87 55.555 ;
    RECT 319.8 54.765 320.01 54.835 ;
    RECT 319.8 55.125 320.01 55.195 ;
    RECT 319.8 55.485 320.01 55.555 ;
    RECT 319.34 54.765 319.55 54.835 ;
    RECT 319.34 55.125 319.55 55.195 ;
    RECT 319.34 55.485 319.55 55.555 ;
    RECT 316.48 54.765 316.69 54.835 ;
    RECT 316.48 55.125 316.69 55.195 ;
    RECT 316.48 55.485 316.69 55.555 ;
    RECT 316.02 54.765 316.23 54.835 ;
    RECT 316.02 55.125 316.23 55.195 ;
    RECT 316.02 55.485 316.23 55.555 ;
    RECT 313.16 54.765 313.37 54.835 ;
    RECT 313.16 55.125 313.37 55.195 ;
    RECT 313.16 55.485 313.37 55.555 ;
    RECT 312.7 54.765 312.91 54.835 ;
    RECT 312.7 55.125 312.91 55.195 ;
    RECT 312.7 55.485 312.91 55.555 ;
    RECT 309.84 54.765 310.05 54.835 ;
    RECT 309.84 55.125 310.05 55.195 ;
    RECT 309.84 55.485 310.05 55.555 ;
    RECT 309.38 54.765 309.59 54.835 ;
    RECT 309.38 55.125 309.59 55.195 ;
    RECT 309.38 55.485 309.59 55.555 ;
    RECT 306.52 54.765 306.73 54.835 ;
    RECT 306.52 55.125 306.73 55.195 ;
    RECT 306.52 55.485 306.73 55.555 ;
    RECT 306.06 54.765 306.27 54.835 ;
    RECT 306.06 55.125 306.27 55.195 ;
    RECT 306.06 55.485 306.27 55.555 ;
    RECT 303.2 54.045 303.41 54.115 ;
    RECT 303.2 54.405 303.41 54.475 ;
    RECT 303.2 54.765 303.41 54.835 ;
    RECT 302.74 54.045 302.95 54.115 ;
    RECT 302.74 54.405 302.95 54.475 ;
    RECT 302.74 54.765 302.95 54.835 ;
    RECT 372.92 54.045 373.13 54.115 ;
    RECT 372.92 54.405 373.13 54.475 ;
    RECT 372.92 54.765 373.13 54.835 ;
    RECT 372.46 54.045 372.67 54.115 ;
    RECT 372.46 54.405 372.67 54.475 ;
    RECT 372.46 54.765 372.67 54.835 ;
    RECT 369.6 54.045 369.81 54.115 ;
    RECT 369.6 54.405 369.81 54.475 ;
    RECT 369.6 54.765 369.81 54.835 ;
    RECT 369.14 54.045 369.35 54.115 ;
    RECT 369.14 54.405 369.35 54.475 ;
    RECT 369.14 54.765 369.35 54.835 ;
    RECT 200.605 54.405 200.675 54.475 ;
    RECT 299.88 54.045 300.09 54.115 ;
    RECT 299.88 54.405 300.09 54.475 ;
    RECT 299.88 54.765 300.09 54.835 ;
    RECT 299.42 54.045 299.63 54.115 ;
    RECT 299.42 54.405 299.63 54.475 ;
    RECT 299.42 54.765 299.63 54.835 ;
    RECT 296.56 54.045 296.77 54.115 ;
    RECT 296.56 54.405 296.77 54.475 ;
    RECT 296.56 54.765 296.77 54.835 ;
    RECT 296.1 54.045 296.31 54.115 ;
    RECT 296.1 54.405 296.31 54.475 ;
    RECT 296.1 54.765 296.31 54.835 ;
    RECT 293.24 54.045 293.45 54.115 ;
    RECT 293.24 54.405 293.45 54.475 ;
    RECT 293.24 54.765 293.45 54.835 ;
    RECT 292.78 54.045 292.99 54.115 ;
    RECT 292.78 54.405 292.99 54.475 ;
    RECT 292.78 54.765 292.99 54.835 ;
    RECT 289.92 54.045 290.13 54.115 ;
    RECT 289.92 54.405 290.13 54.475 ;
    RECT 289.92 54.765 290.13 54.835 ;
    RECT 289.46 54.045 289.67 54.115 ;
    RECT 289.46 54.405 289.67 54.475 ;
    RECT 289.46 54.765 289.67 54.835 ;
    RECT 286.6 54.045 286.81 54.115 ;
    RECT 286.6 54.405 286.81 54.475 ;
    RECT 286.6 54.765 286.81 54.835 ;
    RECT 286.14 54.045 286.35 54.115 ;
    RECT 286.14 54.405 286.35 54.475 ;
    RECT 286.14 54.765 286.35 54.835 ;
    RECT 283.28 54.045 283.49 54.115 ;
    RECT 283.28 54.405 283.49 54.475 ;
    RECT 283.28 54.765 283.49 54.835 ;
    RECT 282.82 54.045 283.03 54.115 ;
    RECT 282.82 54.405 283.03 54.475 ;
    RECT 282.82 54.765 283.03 54.835 ;
    RECT 279.96 54.045 280.17 54.115 ;
    RECT 279.96 54.405 280.17 54.475 ;
    RECT 279.96 54.765 280.17 54.835 ;
    RECT 279.5 54.045 279.71 54.115 ;
    RECT 279.5 54.405 279.71 54.475 ;
    RECT 279.5 54.765 279.71 54.835 ;
    RECT 276.64 54.045 276.85 54.115 ;
    RECT 276.64 54.405 276.85 54.475 ;
    RECT 276.64 54.765 276.85 54.835 ;
    RECT 276.18 54.045 276.39 54.115 ;
    RECT 276.18 54.405 276.39 54.475 ;
    RECT 276.18 54.765 276.39 54.835 ;
    RECT 273.32 54.045 273.53 54.115 ;
    RECT 273.32 54.405 273.53 54.475 ;
    RECT 273.32 54.765 273.53 54.835 ;
    RECT 272.86 54.045 273.07 54.115 ;
    RECT 272.86 54.405 273.07 54.475 ;
    RECT 272.86 54.765 273.07 54.835 ;
    RECT 270.0 54.045 270.21 54.115 ;
    RECT 270.0 54.405 270.21 54.475 ;
    RECT 270.0 54.765 270.21 54.835 ;
    RECT 269.54 54.045 269.75 54.115 ;
    RECT 269.54 54.405 269.75 54.475 ;
    RECT 269.54 54.765 269.75 54.835 ;
    RECT 233.48 54.045 233.69 54.115 ;
    RECT 233.48 54.405 233.69 54.475 ;
    RECT 233.48 54.765 233.69 54.835 ;
    RECT 233.02 54.045 233.23 54.115 ;
    RECT 233.02 54.405 233.23 54.475 ;
    RECT 233.02 54.765 233.23 54.835 ;
    RECT 230.16 54.045 230.37 54.115 ;
    RECT 230.16 54.405 230.37 54.475 ;
    RECT 230.16 54.765 230.37 54.835 ;
    RECT 229.7 54.045 229.91 54.115 ;
    RECT 229.7 54.405 229.91 54.475 ;
    RECT 229.7 54.765 229.91 54.835 ;
    RECT 366.28 54.045 366.49 54.115 ;
    RECT 366.28 54.405 366.49 54.475 ;
    RECT 366.28 54.765 366.49 54.835 ;
    RECT 365.82 54.045 366.03 54.115 ;
    RECT 365.82 54.405 366.03 54.475 ;
    RECT 365.82 54.765 366.03 54.835 ;
    RECT 226.84 54.045 227.05 54.115 ;
    RECT 226.84 54.405 227.05 54.475 ;
    RECT 226.84 54.765 227.05 54.835 ;
    RECT 226.38 54.045 226.59 54.115 ;
    RECT 226.38 54.405 226.59 54.475 ;
    RECT 226.38 54.765 226.59 54.835 ;
    RECT 362.96 54.045 363.17 54.115 ;
    RECT 362.96 54.405 363.17 54.475 ;
    RECT 362.96 54.765 363.17 54.835 ;
    RECT 362.5 54.045 362.71 54.115 ;
    RECT 362.5 54.405 362.71 54.475 ;
    RECT 362.5 54.765 362.71 54.835 ;
    RECT 223.52 54.045 223.73 54.115 ;
    RECT 223.52 54.405 223.73 54.475 ;
    RECT 223.52 54.765 223.73 54.835 ;
    RECT 223.06 54.045 223.27 54.115 ;
    RECT 223.06 54.405 223.27 54.475 ;
    RECT 223.06 54.765 223.27 54.835 ;
    RECT 359.64 54.045 359.85 54.115 ;
    RECT 359.64 54.405 359.85 54.475 ;
    RECT 359.64 54.765 359.85 54.835 ;
    RECT 359.18 54.045 359.39 54.115 ;
    RECT 359.18 54.405 359.39 54.475 ;
    RECT 359.18 54.765 359.39 54.835 ;
    RECT 220.2 54.045 220.41 54.115 ;
    RECT 220.2 54.405 220.41 54.475 ;
    RECT 220.2 54.765 220.41 54.835 ;
    RECT 219.74 54.045 219.95 54.115 ;
    RECT 219.74 54.405 219.95 54.475 ;
    RECT 219.74 54.765 219.95 54.835 ;
    RECT 356.32 54.045 356.53 54.115 ;
    RECT 356.32 54.405 356.53 54.475 ;
    RECT 356.32 54.765 356.53 54.835 ;
    RECT 355.86 54.045 356.07 54.115 ;
    RECT 355.86 54.405 356.07 54.475 ;
    RECT 355.86 54.765 356.07 54.835 ;
    RECT 353.0 54.045 353.21 54.115 ;
    RECT 353.0 54.405 353.21 54.475 ;
    RECT 353.0 54.765 353.21 54.835 ;
    RECT 352.54 54.045 352.75 54.115 ;
    RECT 352.54 54.405 352.75 54.475 ;
    RECT 352.54 54.765 352.75 54.835 ;
    RECT 216.88 54.045 217.09 54.115 ;
    RECT 216.88 54.405 217.09 54.475 ;
    RECT 216.88 54.765 217.09 54.835 ;
    RECT 216.42 54.045 216.63 54.115 ;
    RECT 216.42 54.405 216.63 54.475 ;
    RECT 216.42 54.765 216.63 54.835 ;
    RECT 349.68 54.045 349.89 54.115 ;
    RECT 349.68 54.405 349.89 54.475 ;
    RECT 349.68 54.765 349.89 54.835 ;
    RECT 349.22 54.045 349.43 54.115 ;
    RECT 349.22 54.405 349.43 54.475 ;
    RECT 349.22 54.765 349.43 54.835 ;
    RECT 213.56 54.045 213.77 54.115 ;
    RECT 213.56 54.405 213.77 54.475 ;
    RECT 213.56 54.765 213.77 54.835 ;
    RECT 213.1 54.045 213.31 54.115 ;
    RECT 213.1 54.405 213.31 54.475 ;
    RECT 213.1 54.765 213.31 54.835 ;
    RECT 346.36 54.045 346.57 54.115 ;
    RECT 346.36 54.405 346.57 54.475 ;
    RECT 346.36 54.765 346.57 54.835 ;
    RECT 345.9 54.045 346.11 54.115 ;
    RECT 345.9 54.405 346.11 54.475 ;
    RECT 345.9 54.765 346.11 54.835 ;
    RECT 210.24 54.045 210.45 54.115 ;
    RECT 210.24 54.405 210.45 54.475 ;
    RECT 210.24 54.765 210.45 54.835 ;
    RECT 209.78 54.045 209.99 54.115 ;
    RECT 209.78 54.405 209.99 54.475 ;
    RECT 209.78 54.765 209.99 54.835 ;
    RECT 343.04 54.045 343.25 54.115 ;
    RECT 343.04 54.405 343.25 54.475 ;
    RECT 343.04 54.765 343.25 54.835 ;
    RECT 342.58 54.045 342.79 54.115 ;
    RECT 342.58 54.405 342.79 54.475 ;
    RECT 342.58 54.765 342.79 54.835 ;
    RECT 206.92 54.045 207.13 54.115 ;
    RECT 206.92 54.405 207.13 54.475 ;
    RECT 206.92 54.765 207.13 54.835 ;
    RECT 206.46 54.045 206.67 54.115 ;
    RECT 206.46 54.405 206.67 54.475 ;
    RECT 206.46 54.765 206.67 54.835 ;
    RECT 339.72 54.045 339.93 54.115 ;
    RECT 339.72 54.405 339.93 54.475 ;
    RECT 339.72 54.765 339.93 54.835 ;
    RECT 339.26 54.045 339.47 54.115 ;
    RECT 339.26 54.405 339.47 54.475 ;
    RECT 339.26 54.765 339.47 54.835 ;
    RECT 203.6 54.045 203.81 54.115 ;
    RECT 203.6 54.405 203.81 54.475 ;
    RECT 203.6 54.765 203.81 54.835 ;
    RECT 203.14 54.045 203.35 54.115 ;
    RECT 203.14 54.405 203.35 54.475 ;
    RECT 203.14 54.765 203.35 54.835 ;
    RECT 336.4 54.045 336.61 54.115 ;
    RECT 336.4 54.405 336.61 54.475 ;
    RECT 336.4 54.765 336.61 54.835 ;
    RECT 335.94 54.045 336.15 54.115 ;
    RECT 335.94 54.405 336.15 54.475 ;
    RECT 335.94 54.765 336.15 54.835 ;
    RECT 266.68 54.045 266.89 54.115 ;
    RECT 266.68 54.405 266.89 54.475 ;
    RECT 266.68 54.765 266.89 54.835 ;
    RECT 266.22 54.045 266.43 54.115 ;
    RECT 266.22 54.405 266.43 54.475 ;
    RECT 266.22 54.765 266.43 54.835 ;
    RECT 263.36 54.045 263.57 54.115 ;
    RECT 263.36 54.405 263.57 54.475 ;
    RECT 263.36 54.765 263.57 54.835 ;
    RECT 262.9 54.045 263.11 54.115 ;
    RECT 262.9 54.405 263.11 54.475 ;
    RECT 262.9 54.765 263.11 54.835 ;
    RECT 260.04 54.045 260.25 54.115 ;
    RECT 260.04 54.405 260.25 54.475 ;
    RECT 260.04 54.765 260.25 54.835 ;
    RECT 259.58 54.045 259.79 54.115 ;
    RECT 259.58 54.405 259.79 54.475 ;
    RECT 259.58 54.765 259.79 54.835 ;
    RECT 256.72 54.045 256.93 54.115 ;
    RECT 256.72 54.405 256.93 54.475 ;
    RECT 256.72 54.765 256.93 54.835 ;
    RECT 256.26 54.045 256.47 54.115 ;
    RECT 256.26 54.405 256.47 54.475 ;
    RECT 256.26 54.765 256.47 54.835 ;
    RECT 253.4 54.045 253.61 54.115 ;
    RECT 253.4 54.405 253.61 54.475 ;
    RECT 253.4 54.765 253.61 54.835 ;
    RECT 252.94 54.045 253.15 54.115 ;
    RECT 252.94 54.405 253.15 54.475 ;
    RECT 252.94 54.765 253.15 54.835 ;
    RECT 250.08 54.045 250.29 54.115 ;
    RECT 250.08 54.405 250.29 54.475 ;
    RECT 250.08 54.765 250.29 54.835 ;
    RECT 249.62 54.045 249.83 54.115 ;
    RECT 249.62 54.405 249.83 54.475 ;
    RECT 249.62 54.765 249.83 54.835 ;
    RECT 246.76 54.045 246.97 54.115 ;
    RECT 246.76 54.405 246.97 54.475 ;
    RECT 246.76 54.765 246.97 54.835 ;
    RECT 246.3 54.045 246.51 54.115 ;
    RECT 246.3 54.405 246.51 54.475 ;
    RECT 246.3 54.765 246.51 54.835 ;
    RECT 243.44 54.045 243.65 54.115 ;
    RECT 243.44 54.405 243.65 54.475 ;
    RECT 243.44 54.765 243.65 54.835 ;
    RECT 242.98 54.045 243.19 54.115 ;
    RECT 242.98 54.405 243.19 54.475 ;
    RECT 242.98 54.765 243.19 54.835 ;
    RECT 240.12 54.045 240.33 54.115 ;
    RECT 240.12 54.405 240.33 54.475 ;
    RECT 240.12 54.765 240.33 54.835 ;
    RECT 239.66 54.045 239.87 54.115 ;
    RECT 239.66 54.405 239.87 54.475 ;
    RECT 239.66 54.765 239.87 54.835 ;
    RECT 236.8 54.045 237.01 54.115 ;
    RECT 236.8 54.405 237.01 54.475 ;
    RECT 236.8 54.765 237.01 54.835 ;
    RECT 236.34 54.045 236.55 54.115 ;
    RECT 236.34 54.405 236.55 54.475 ;
    RECT 236.34 54.765 236.55 54.835 ;
    RECT 374.15 54.405 374.22 54.475 ;
    RECT 333.08 54.045 333.29 54.115 ;
    RECT 333.08 54.405 333.29 54.475 ;
    RECT 333.08 54.765 333.29 54.835 ;
    RECT 332.62 54.045 332.83 54.115 ;
    RECT 332.62 54.405 332.83 54.475 ;
    RECT 332.62 54.765 332.83 54.835 ;
    RECT 329.76 54.045 329.97 54.115 ;
    RECT 329.76 54.405 329.97 54.475 ;
    RECT 329.76 54.765 329.97 54.835 ;
    RECT 329.3 54.045 329.51 54.115 ;
    RECT 329.3 54.405 329.51 54.475 ;
    RECT 329.3 54.765 329.51 54.835 ;
    RECT 326.44 54.045 326.65 54.115 ;
    RECT 326.44 54.405 326.65 54.475 ;
    RECT 326.44 54.765 326.65 54.835 ;
    RECT 325.98 54.045 326.19 54.115 ;
    RECT 325.98 54.405 326.19 54.475 ;
    RECT 325.98 54.765 326.19 54.835 ;
    RECT 323.12 54.045 323.33 54.115 ;
    RECT 323.12 54.405 323.33 54.475 ;
    RECT 323.12 54.765 323.33 54.835 ;
    RECT 322.66 54.045 322.87 54.115 ;
    RECT 322.66 54.405 322.87 54.475 ;
    RECT 322.66 54.765 322.87 54.835 ;
    RECT 319.8 54.045 320.01 54.115 ;
    RECT 319.8 54.405 320.01 54.475 ;
    RECT 319.8 54.765 320.01 54.835 ;
    RECT 319.34 54.045 319.55 54.115 ;
    RECT 319.34 54.405 319.55 54.475 ;
    RECT 319.34 54.765 319.55 54.835 ;
    RECT 316.48 54.045 316.69 54.115 ;
    RECT 316.48 54.405 316.69 54.475 ;
    RECT 316.48 54.765 316.69 54.835 ;
    RECT 316.02 54.045 316.23 54.115 ;
    RECT 316.02 54.405 316.23 54.475 ;
    RECT 316.02 54.765 316.23 54.835 ;
    RECT 313.16 54.045 313.37 54.115 ;
    RECT 313.16 54.405 313.37 54.475 ;
    RECT 313.16 54.765 313.37 54.835 ;
    RECT 312.7 54.045 312.91 54.115 ;
    RECT 312.7 54.405 312.91 54.475 ;
    RECT 312.7 54.765 312.91 54.835 ;
    RECT 309.84 54.045 310.05 54.115 ;
    RECT 309.84 54.405 310.05 54.475 ;
    RECT 309.84 54.765 310.05 54.835 ;
    RECT 309.38 54.045 309.59 54.115 ;
    RECT 309.38 54.405 309.59 54.475 ;
    RECT 309.38 54.765 309.59 54.835 ;
    RECT 306.52 54.045 306.73 54.115 ;
    RECT 306.52 54.405 306.73 54.475 ;
    RECT 306.52 54.765 306.73 54.835 ;
    RECT 306.06 54.045 306.27 54.115 ;
    RECT 306.06 54.405 306.27 54.475 ;
    RECT 306.06 54.765 306.27 54.835 ;
    RECT 303.2 53.325 303.41 53.395 ;
    RECT 303.2 53.685 303.41 53.755 ;
    RECT 303.2 54.045 303.41 54.115 ;
    RECT 302.74 53.325 302.95 53.395 ;
    RECT 302.74 53.685 302.95 53.755 ;
    RECT 302.74 54.045 302.95 54.115 ;
    RECT 372.92 53.325 373.13 53.395 ;
    RECT 372.92 53.685 373.13 53.755 ;
    RECT 372.92 54.045 373.13 54.115 ;
    RECT 372.46 53.325 372.67 53.395 ;
    RECT 372.46 53.685 372.67 53.755 ;
    RECT 372.46 54.045 372.67 54.115 ;
    RECT 369.6 53.325 369.81 53.395 ;
    RECT 369.6 53.685 369.81 53.755 ;
    RECT 369.6 54.045 369.81 54.115 ;
    RECT 369.14 53.325 369.35 53.395 ;
    RECT 369.14 53.685 369.35 53.755 ;
    RECT 369.14 54.045 369.35 54.115 ;
    RECT 200.605 53.685 200.675 53.755 ;
    RECT 299.88 53.325 300.09 53.395 ;
    RECT 299.88 53.685 300.09 53.755 ;
    RECT 299.88 54.045 300.09 54.115 ;
    RECT 299.42 53.325 299.63 53.395 ;
    RECT 299.42 53.685 299.63 53.755 ;
    RECT 299.42 54.045 299.63 54.115 ;
    RECT 296.56 53.325 296.77 53.395 ;
    RECT 296.56 53.685 296.77 53.755 ;
    RECT 296.56 54.045 296.77 54.115 ;
    RECT 296.1 53.325 296.31 53.395 ;
    RECT 296.1 53.685 296.31 53.755 ;
    RECT 296.1 54.045 296.31 54.115 ;
    RECT 293.24 53.325 293.45 53.395 ;
    RECT 293.24 53.685 293.45 53.755 ;
    RECT 293.24 54.045 293.45 54.115 ;
    RECT 292.78 53.325 292.99 53.395 ;
    RECT 292.78 53.685 292.99 53.755 ;
    RECT 292.78 54.045 292.99 54.115 ;
    RECT 289.92 53.325 290.13 53.395 ;
    RECT 289.92 53.685 290.13 53.755 ;
    RECT 289.92 54.045 290.13 54.115 ;
    RECT 289.46 53.325 289.67 53.395 ;
    RECT 289.46 53.685 289.67 53.755 ;
    RECT 289.46 54.045 289.67 54.115 ;
    RECT 286.6 53.325 286.81 53.395 ;
    RECT 286.6 53.685 286.81 53.755 ;
    RECT 286.6 54.045 286.81 54.115 ;
    RECT 286.14 53.325 286.35 53.395 ;
    RECT 286.14 53.685 286.35 53.755 ;
    RECT 286.14 54.045 286.35 54.115 ;
    RECT 283.28 53.325 283.49 53.395 ;
    RECT 283.28 53.685 283.49 53.755 ;
    RECT 283.28 54.045 283.49 54.115 ;
    RECT 282.82 53.325 283.03 53.395 ;
    RECT 282.82 53.685 283.03 53.755 ;
    RECT 282.82 54.045 283.03 54.115 ;
    RECT 279.96 53.325 280.17 53.395 ;
    RECT 279.96 53.685 280.17 53.755 ;
    RECT 279.96 54.045 280.17 54.115 ;
    RECT 279.5 53.325 279.71 53.395 ;
    RECT 279.5 53.685 279.71 53.755 ;
    RECT 279.5 54.045 279.71 54.115 ;
    RECT 276.64 53.325 276.85 53.395 ;
    RECT 276.64 53.685 276.85 53.755 ;
    RECT 276.64 54.045 276.85 54.115 ;
    RECT 276.18 53.325 276.39 53.395 ;
    RECT 276.18 53.685 276.39 53.755 ;
    RECT 276.18 54.045 276.39 54.115 ;
    RECT 273.32 53.325 273.53 53.395 ;
    RECT 273.32 53.685 273.53 53.755 ;
    RECT 273.32 54.045 273.53 54.115 ;
    RECT 272.86 53.325 273.07 53.395 ;
    RECT 272.86 53.685 273.07 53.755 ;
    RECT 272.86 54.045 273.07 54.115 ;
    RECT 270.0 53.325 270.21 53.395 ;
    RECT 270.0 53.685 270.21 53.755 ;
    RECT 270.0 54.045 270.21 54.115 ;
    RECT 269.54 53.325 269.75 53.395 ;
    RECT 269.54 53.685 269.75 53.755 ;
    RECT 269.54 54.045 269.75 54.115 ;
    RECT 233.48 53.325 233.69 53.395 ;
    RECT 233.48 53.685 233.69 53.755 ;
    RECT 233.48 54.045 233.69 54.115 ;
    RECT 233.02 53.325 233.23 53.395 ;
    RECT 233.02 53.685 233.23 53.755 ;
    RECT 233.02 54.045 233.23 54.115 ;
    RECT 230.16 53.325 230.37 53.395 ;
    RECT 230.16 53.685 230.37 53.755 ;
    RECT 230.16 54.045 230.37 54.115 ;
    RECT 229.7 53.325 229.91 53.395 ;
    RECT 229.7 53.685 229.91 53.755 ;
    RECT 229.7 54.045 229.91 54.115 ;
    RECT 366.28 53.325 366.49 53.395 ;
    RECT 366.28 53.685 366.49 53.755 ;
    RECT 366.28 54.045 366.49 54.115 ;
    RECT 365.82 53.325 366.03 53.395 ;
    RECT 365.82 53.685 366.03 53.755 ;
    RECT 365.82 54.045 366.03 54.115 ;
    RECT 226.84 53.325 227.05 53.395 ;
    RECT 226.84 53.685 227.05 53.755 ;
    RECT 226.84 54.045 227.05 54.115 ;
    RECT 226.38 53.325 226.59 53.395 ;
    RECT 226.38 53.685 226.59 53.755 ;
    RECT 226.38 54.045 226.59 54.115 ;
    RECT 362.96 53.325 363.17 53.395 ;
    RECT 362.96 53.685 363.17 53.755 ;
    RECT 362.96 54.045 363.17 54.115 ;
    RECT 362.5 53.325 362.71 53.395 ;
    RECT 362.5 53.685 362.71 53.755 ;
    RECT 362.5 54.045 362.71 54.115 ;
    RECT 223.52 53.325 223.73 53.395 ;
    RECT 223.52 53.685 223.73 53.755 ;
    RECT 223.52 54.045 223.73 54.115 ;
    RECT 223.06 53.325 223.27 53.395 ;
    RECT 223.06 53.685 223.27 53.755 ;
    RECT 223.06 54.045 223.27 54.115 ;
    RECT 359.64 53.325 359.85 53.395 ;
    RECT 359.64 53.685 359.85 53.755 ;
    RECT 359.64 54.045 359.85 54.115 ;
    RECT 359.18 53.325 359.39 53.395 ;
    RECT 359.18 53.685 359.39 53.755 ;
    RECT 359.18 54.045 359.39 54.115 ;
    RECT 220.2 53.325 220.41 53.395 ;
    RECT 220.2 53.685 220.41 53.755 ;
    RECT 220.2 54.045 220.41 54.115 ;
    RECT 219.74 53.325 219.95 53.395 ;
    RECT 219.74 53.685 219.95 53.755 ;
    RECT 219.74 54.045 219.95 54.115 ;
    RECT 356.32 53.325 356.53 53.395 ;
    RECT 356.32 53.685 356.53 53.755 ;
    RECT 356.32 54.045 356.53 54.115 ;
    RECT 355.86 53.325 356.07 53.395 ;
    RECT 355.86 53.685 356.07 53.755 ;
    RECT 355.86 54.045 356.07 54.115 ;
    RECT 353.0 53.325 353.21 53.395 ;
    RECT 353.0 53.685 353.21 53.755 ;
    RECT 353.0 54.045 353.21 54.115 ;
    RECT 352.54 53.325 352.75 53.395 ;
    RECT 352.54 53.685 352.75 53.755 ;
    RECT 352.54 54.045 352.75 54.115 ;
    RECT 216.88 53.325 217.09 53.395 ;
    RECT 216.88 53.685 217.09 53.755 ;
    RECT 216.88 54.045 217.09 54.115 ;
    RECT 216.42 53.325 216.63 53.395 ;
    RECT 216.42 53.685 216.63 53.755 ;
    RECT 216.42 54.045 216.63 54.115 ;
    RECT 349.68 53.325 349.89 53.395 ;
    RECT 349.68 53.685 349.89 53.755 ;
    RECT 349.68 54.045 349.89 54.115 ;
    RECT 349.22 53.325 349.43 53.395 ;
    RECT 349.22 53.685 349.43 53.755 ;
    RECT 349.22 54.045 349.43 54.115 ;
    RECT 213.56 53.325 213.77 53.395 ;
    RECT 213.56 53.685 213.77 53.755 ;
    RECT 213.56 54.045 213.77 54.115 ;
    RECT 213.1 53.325 213.31 53.395 ;
    RECT 213.1 53.685 213.31 53.755 ;
    RECT 213.1 54.045 213.31 54.115 ;
    RECT 346.36 53.325 346.57 53.395 ;
    RECT 346.36 53.685 346.57 53.755 ;
    RECT 346.36 54.045 346.57 54.115 ;
    RECT 345.9 53.325 346.11 53.395 ;
    RECT 345.9 53.685 346.11 53.755 ;
    RECT 345.9 54.045 346.11 54.115 ;
    RECT 210.24 53.325 210.45 53.395 ;
    RECT 210.24 53.685 210.45 53.755 ;
    RECT 210.24 54.045 210.45 54.115 ;
    RECT 209.78 53.325 209.99 53.395 ;
    RECT 209.78 53.685 209.99 53.755 ;
    RECT 209.78 54.045 209.99 54.115 ;
    RECT 343.04 53.325 343.25 53.395 ;
    RECT 343.04 53.685 343.25 53.755 ;
    RECT 343.04 54.045 343.25 54.115 ;
    RECT 342.58 53.325 342.79 53.395 ;
    RECT 342.58 53.685 342.79 53.755 ;
    RECT 342.58 54.045 342.79 54.115 ;
    RECT 206.92 53.325 207.13 53.395 ;
    RECT 206.92 53.685 207.13 53.755 ;
    RECT 206.92 54.045 207.13 54.115 ;
    RECT 206.46 53.325 206.67 53.395 ;
    RECT 206.46 53.685 206.67 53.755 ;
    RECT 206.46 54.045 206.67 54.115 ;
    RECT 339.72 53.325 339.93 53.395 ;
    RECT 339.72 53.685 339.93 53.755 ;
    RECT 339.72 54.045 339.93 54.115 ;
    RECT 339.26 53.325 339.47 53.395 ;
    RECT 339.26 53.685 339.47 53.755 ;
    RECT 339.26 54.045 339.47 54.115 ;
    RECT 203.6 53.325 203.81 53.395 ;
    RECT 203.6 53.685 203.81 53.755 ;
    RECT 203.6 54.045 203.81 54.115 ;
    RECT 203.14 53.325 203.35 53.395 ;
    RECT 203.14 53.685 203.35 53.755 ;
    RECT 203.14 54.045 203.35 54.115 ;
    RECT 336.4 53.325 336.61 53.395 ;
    RECT 336.4 53.685 336.61 53.755 ;
    RECT 336.4 54.045 336.61 54.115 ;
    RECT 335.94 53.325 336.15 53.395 ;
    RECT 335.94 53.685 336.15 53.755 ;
    RECT 335.94 54.045 336.15 54.115 ;
    RECT 266.68 53.325 266.89 53.395 ;
    RECT 266.68 53.685 266.89 53.755 ;
    RECT 266.68 54.045 266.89 54.115 ;
    RECT 266.22 53.325 266.43 53.395 ;
    RECT 266.22 53.685 266.43 53.755 ;
    RECT 266.22 54.045 266.43 54.115 ;
    RECT 263.36 53.325 263.57 53.395 ;
    RECT 263.36 53.685 263.57 53.755 ;
    RECT 263.36 54.045 263.57 54.115 ;
    RECT 262.9 53.325 263.11 53.395 ;
    RECT 262.9 53.685 263.11 53.755 ;
    RECT 262.9 54.045 263.11 54.115 ;
    RECT 260.04 53.325 260.25 53.395 ;
    RECT 260.04 53.685 260.25 53.755 ;
    RECT 260.04 54.045 260.25 54.115 ;
    RECT 259.58 53.325 259.79 53.395 ;
    RECT 259.58 53.685 259.79 53.755 ;
    RECT 259.58 54.045 259.79 54.115 ;
    RECT 256.72 53.325 256.93 53.395 ;
    RECT 256.72 53.685 256.93 53.755 ;
    RECT 256.72 54.045 256.93 54.115 ;
    RECT 256.26 53.325 256.47 53.395 ;
    RECT 256.26 53.685 256.47 53.755 ;
    RECT 256.26 54.045 256.47 54.115 ;
    RECT 253.4 53.325 253.61 53.395 ;
    RECT 253.4 53.685 253.61 53.755 ;
    RECT 253.4 54.045 253.61 54.115 ;
    RECT 252.94 53.325 253.15 53.395 ;
    RECT 252.94 53.685 253.15 53.755 ;
    RECT 252.94 54.045 253.15 54.115 ;
    RECT 250.08 53.325 250.29 53.395 ;
    RECT 250.08 53.685 250.29 53.755 ;
    RECT 250.08 54.045 250.29 54.115 ;
    RECT 249.62 53.325 249.83 53.395 ;
    RECT 249.62 53.685 249.83 53.755 ;
    RECT 249.62 54.045 249.83 54.115 ;
    RECT 246.76 53.325 246.97 53.395 ;
    RECT 246.76 53.685 246.97 53.755 ;
    RECT 246.76 54.045 246.97 54.115 ;
    RECT 246.3 53.325 246.51 53.395 ;
    RECT 246.3 53.685 246.51 53.755 ;
    RECT 246.3 54.045 246.51 54.115 ;
    RECT 243.44 53.325 243.65 53.395 ;
    RECT 243.44 53.685 243.65 53.755 ;
    RECT 243.44 54.045 243.65 54.115 ;
    RECT 242.98 53.325 243.19 53.395 ;
    RECT 242.98 53.685 243.19 53.755 ;
    RECT 242.98 54.045 243.19 54.115 ;
    RECT 240.12 53.325 240.33 53.395 ;
    RECT 240.12 53.685 240.33 53.755 ;
    RECT 240.12 54.045 240.33 54.115 ;
    RECT 239.66 53.325 239.87 53.395 ;
    RECT 239.66 53.685 239.87 53.755 ;
    RECT 239.66 54.045 239.87 54.115 ;
    RECT 236.8 53.325 237.01 53.395 ;
    RECT 236.8 53.685 237.01 53.755 ;
    RECT 236.8 54.045 237.01 54.115 ;
    RECT 236.34 53.325 236.55 53.395 ;
    RECT 236.34 53.685 236.55 53.755 ;
    RECT 236.34 54.045 236.55 54.115 ;
    RECT 374.15 53.685 374.22 53.755 ;
    RECT 333.08 53.325 333.29 53.395 ;
    RECT 333.08 53.685 333.29 53.755 ;
    RECT 333.08 54.045 333.29 54.115 ;
    RECT 332.62 53.325 332.83 53.395 ;
    RECT 332.62 53.685 332.83 53.755 ;
    RECT 332.62 54.045 332.83 54.115 ;
    RECT 329.76 53.325 329.97 53.395 ;
    RECT 329.76 53.685 329.97 53.755 ;
    RECT 329.76 54.045 329.97 54.115 ;
    RECT 329.3 53.325 329.51 53.395 ;
    RECT 329.3 53.685 329.51 53.755 ;
    RECT 329.3 54.045 329.51 54.115 ;
    RECT 326.44 53.325 326.65 53.395 ;
    RECT 326.44 53.685 326.65 53.755 ;
    RECT 326.44 54.045 326.65 54.115 ;
    RECT 325.98 53.325 326.19 53.395 ;
    RECT 325.98 53.685 326.19 53.755 ;
    RECT 325.98 54.045 326.19 54.115 ;
    RECT 323.12 53.325 323.33 53.395 ;
    RECT 323.12 53.685 323.33 53.755 ;
    RECT 323.12 54.045 323.33 54.115 ;
    RECT 322.66 53.325 322.87 53.395 ;
    RECT 322.66 53.685 322.87 53.755 ;
    RECT 322.66 54.045 322.87 54.115 ;
    RECT 319.8 53.325 320.01 53.395 ;
    RECT 319.8 53.685 320.01 53.755 ;
    RECT 319.8 54.045 320.01 54.115 ;
    RECT 319.34 53.325 319.55 53.395 ;
    RECT 319.34 53.685 319.55 53.755 ;
    RECT 319.34 54.045 319.55 54.115 ;
    RECT 316.48 53.325 316.69 53.395 ;
    RECT 316.48 53.685 316.69 53.755 ;
    RECT 316.48 54.045 316.69 54.115 ;
    RECT 316.02 53.325 316.23 53.395 ;
    RECT 316.02 53.685 316.23 53.755 ;
    RECT 316.02 54.045 316.23 54.115 ;
    RECT 313.16 53.325 313.37 53.395 ;
    RECT 313.16 53.685 313.37 53.755 ;
    RECT 313.16 54.045 313.37 54.115 ;
    RECT 312.7 53.325 312.91 53.395 ;
    RECT 312.7 53.685 312.91 53.755 ;
    RECT 312.7 54.045 312.91 54.115 ;
    RECT 309.84 53.325 310.05 53.395 ;
    RECT 309.84 53.685 310.05 53.755 ;
    RECT 309.84 54.045 310.05 54.115 ;
    RECT 309.38 53.325 309.59 53.395 ;
    RECT 309.38 53.685 309.59 53.755 ;
    RECT 309.38 54.045 309.59 54.115 ;
    RECT 306.52 53.325 306.73 53.395 ;
    RECT 306.52 53.685 306.73 53.755 ;
    RECT 306.52 54.045 306.73 54.115 ;
    RECT 306.06 53.325 306.27 53.395 ;
    RECT 306.06 53.685 306.27 53.755 ;
    RECT 306.06 54.045 306.27 54.115 ;
    RECT 303.2 52.605 303.41 52.675 ;
    RECT 303.2 52.965 303.41 53.035 ;
    RECT 303.2 53.325 303.41 53.395 ;
    RECT 302.74 52.605 302.95 52.675 ;
    RECT 302.74 52.965 302.95 53.035 ;
    RECT 302.74 53.325 302.95 53.395 ;
    RECT 372.92 52.605 373.13 52.675 ;
    RECT 372.92 52.965 373.13 53.035 ;
    RECT 372.92 53.325 373.13 53.395 ;
    RECT 372.46 52.605 372.67 52.675 ;
    RECT 372.46 52.965 372.67 53.035 ;
    RECT 372.46 53.325 372.67 53.395 ;
    RECT 369.6 52.605 369.81 52.675 ;
    RECT 369.6 52.965 369.81 53.035 ;
    RECT 369.6 53.325 369.81 53.395 ;
    RECT 369.14 52.605 369.35 52.675 ;
    RECT 369.14 52.965 369.35 53.035 ;
    RECT 369.14 53.325 369.35 53.395 ;
    RECT 200.605 52.965 200.675 53.035 ;
    RECT 299.88 52.605 300.09 52.675 ;
    RECT 299.88 52.965 300.09 53.035 ;
    RECT 299.88 53.325 300.09 53.395 ;
    RECT 299.42 52.605 299.63 52.675 ;
    RECT 299.42 52.965 299.63 53.035 ;
    RECT 299.42 53.325 299.63 53.395 ;
    RECT 296.56 52.605 296.77 52.675 ;
    RECT 296.56 52.965 296.77 53.035 ;
    RECT 296.56 53.325 296.77 53.395 ;
    RECT 296.1 52.605 296.31 52.675 ;
    RECT 296.1 52.965 296.31 53.035 ;
    RECT 296.1 53.325 296.31 53.395 ;
    RECT 293.24 52.605 293.45 52.675 ;
    RECT 293.24 52.965 293.45 53.035 ;
    RECT 293.24 53.325 293.45 53.395 ;
    RECT 292.78 52.605 292.99 52.675 ;
    RECT 292.78 52.965 292.99 53.035 ;
    RECT 292.78 53.325 292.99 53.395 ;
    RECT 289.92 52.605 290.13 52.675 ;
    RECT 289.92 52.965 290.13 53.035 ;
    RECT 289.92 53.325 290.13 53.395 ;
    RECT 289.46 52.605 289.67 52.675 ;
    RECT 289.46 52.965 289.67 53.035 ;
    RECT 289.46 53.325 289.67 53.395 ;
    RECT 286.6 52.605 286.81 52.675 ;
    RECT 286.6 52.965 286.81 53.035 ;
    RECT 286.6 53.325 286.81 53.395 ;
    RECT 286.14 52.605 286.35 52.675 ;
    RECT 286.14 52.965 286.35 53.035 ;
    RECT 286.14 53.325 286.35 53.395 ;
    RECT 283.28 52.605 283.49 52.675 ;
    RECT 283.28 52.965 283.49 53.035 ;
    RECT 283.28 53.325 283.49 53.395 ;
    RECT 282.82 52.605 283.03 52.675 ;
    RECT 282.82 52.965 283.03 53.035 ;
    RECT 282.82 53.325 283.03 53.395 ;
    RECT 279.96 52.605 280.17 52.675 ;
    RECT 279.96 52.965 280.17 53.035 ;
    RECT 279.96 53.325 280.17 53.395 ;
    RECT 279.5 52.605 279.71 52.675 ;
    RECT 279.5 52.965 279.71 53.035 ;
    RECT 279.5 53.325 279.71 53.395 ;
    RECT 276.64 52.605 276.85 52.675 ;
    RECT 276.64 52.965 276.85 53.035 ;
    RECT 276.64 53.325 276.85 53.395 ;
    RECT 276.18 52.605 276.39 52.675 ;
    RECT 276.18 52.965 276.39 53.035 ;
    RECT 276.18 53.325 276.39 53.395 ;
    RECT 273.32 52.605 273.53 52.675 ;
    RECT 273.32 52.965 273.53 53.035 ;
    RECT 273.32 53.325 273.53 53.395 ;
    RECT 272.86 52.605 273.07 52.675 ;
    RECT 272.86 52.965 273.07 53.035 ;
    RECT 272.86 53.325 273.07 53.395 ;
    RECT 270.0 52.605 270.21 52.675 ;
    RECT 270.0 52.965 270.21 53.035 ;
    RECT 270.0 53.325 270.21 53.395 ;
    RECT 269.54 52.605 269.75 52.675 ;
    RECT 269.54 52.965 269.75 53.035 ;
    RECT 269.54 53.325 269.75 53.395 ;
    RECT 233.48 52.605 233.69 52.675 ;
    RECT 233.48 52.965 233.69 53.035 ;
    RECT 233.48 53.325 233.69 53.395 ;
    RECT 233.02 52.605 233.23 52.675 ;
    RECT 233.02 52.965 233.23 53.035 ;
    RECT 233.02 53.325 233.23 53.395 ;
    RECT 230.16 52.605 230.37 52.675 ;
    RECT 230.16 52.965 230.37 53.035 ;
    RECT 230.16 53.325 230.37 53.395 ;
    RECT 229.7 52.605 229.91 52.675 ;
    RECT 229.7 52.965 229.91 53.035 ;
    RECT 229.7 53.325 229.91 53.395 ;
    RECT 366.28 52.605 366.49 52.675 ;
    RECT 366.28 52.965 366.49 53.035 ;
    RECT 366.28 53.325 366.49 53.395 ;
    RECT 365.82 52.605 366.03 52.675 ;
    RECT 365.82 52.965 366.03 53.035 ;
    RECT 365.82 53.325 366.03 53.395 ;
    RECT 226.84 52.605 227.05 52.675 ;
    RECT 226.84 52.965 227.05 53.035 ;
    RECT 226.84 53.325 227.05 53.395 ;
    RECT 226.38 52.605 226.59 52.675 ;
    RECT 226.38 52.965 226.59 53.035 ;
    RECT 226.38 53.325 226.59 53.395 ;
    RECT 362.96 52.605 363.17 52.675 ;
    RECT 362.96 52.965 363.17 53.035 ;
    RECT 362.96 53.325 363.17 53.395 ;
    RECT 362.5 52.605 362.71 52.675 ;
    RECT 362.5 52.965 362.71 53.035 ;
    RECT 362.5 53.325 362.71 53.395 ;
    RECT 223.52 52.605 223.73 52.675 ;
    RECT 223.52 52.965 223.73 53.035 ;
    RECT 223.52 53.325 223.73 53.395 ;
    RECT 223.06 52.605 223.27 52.675 ;
    RECT 223.06 52.965 223.27 53.035 ;
    RECT 223.06 53.325 223.27 53.395 ;
    RECT 359.64 52.605 359.85 52.675 ;
    RECT 359.64 52.965 359.85 53.035 ;
    RECT 359.64 53.325 359.85 53.395 ;
    RECT 359.18 52.605 359.39 52.675 ;
    RECT 359.18 52.965 359.39 53.035 ;
    RECT 359.18 53.325 359.39 53.395 ;
    RECT 220.2 52.605 220.41 52.675 ;
    RECT 220.2 52.965 220.41 53.035 ;
    RECT 220.2 53.325 220.41 53.395 ;
    RECT 219.74 52.605 219.95 52.675 ;
    RECT 219.74 52.965 219.95 53.035 ;
    RECT 219.74 53.325 219.95 53.395 ;
    RECT 356.32 52.605 356.53 52.675 ;
    RECT 356.32 52.965 356.53 53.035 ;
    RECT 356.32 53.325 356.53 53.395 ;
    RECT 355.86 52.605 356.07 52.675 ;
    RECT 355.86 52.965 356.07 53.035 ;
    RECT 355.86 53.325 356.07 53.395 ;
    RECT 353.0 52.605 353.21 52.675 ;
    RECT 353.0 52.965 353.21 53.035 ;
    RECT 353.0 53.325 353.21 53.395 ;
    RECT 352.54 52.605 352.75 52.675 ;
    RECT 352.54 52.965 352.75 53.035 ;
    RECT 352.54 53.325 352.75 53.395 ;
    RECT 216.88 52.605 217.09 52.675 ;
    RECT 216.88 52.965 217.09 53.035 ;
    RECT 216.88 53.325 217.09 53.395 ;
    RECT 216.42 52.605 216.63 52.675 ;
    RECT 216.42 52.965 216.63 53.035 ;
    RECT 216.42 53.325 216.63 53.395 ;
    RECT 349.68 52.605 349.89 52.675 ;
    RECT 349.68 52.965 349.89 53.035 ;
    RECT 349.68 53.325 349.89 53.395 ;
    RECT 349.22 52.605 349.43 52.675 ;
    RECT 349.22 52.965 349.43 53.035 ;
    RECT 349.22 53.325 349.43 53.395 ;
    RECT 213.56 52.605 213.77 52.675 ;
    RECT 213.56 52.965 213.77 53.035 ;
    RECT 213.56 53.325 213.77 53.395 ;
    RECT 213.1 52.605 213.31 52.675 ;
    RECT 213.1 52.965 213.31 53.035 ;
    RECT 213.1 53.325 213.31 53.395 ;
    RECT 346.36 52.605 346.57 52.675 ;
    RECT 346.36 52.965 346.57 53.035 ;
    RECT 346.36 53.325 346.57 53.395 ;
    RECT 345.9 52.605 346.11 52.675 ;
    RECT 345.9 52.965 346.11 53.035 ;
    RECT 345.9 53.325 346.11 53.395 ;
    RECT 210.24 52.605 210.45 52.675 ;
    RECT 210.24 52.965 210.45 53.035 ;
    RECT 210.24 53.325 210.45 53.395 ;
    RECT 209.78 52.605 209.99 52.675 ;
    RECT 209.78 52.965 209.99 53.035 ;
    RECT 209.78 53.325 209.99 53.395 ;
    RECT 343.04 52.605 343.25 52.675 ;
    RECT 343.04 52.965 343.25 53.035 ;
    RECT 343.04 53.325 343.25 53.395 ;
    RECT 342.58 52.605 342.79 52.675 ;
    RECT 342.58 52.965 342.79 53.035 ;
    RECT 342.58 53.325 342.79 53.395 ;
    RECT 206.92 52.605 207.13 52.675 ;
    RECT 206.92 52.965 207.13 53.035 ;
    RECT 206.92 53.325 207.13 53.395 ;
    RECT 206.46 52.605 206.67 52.675 ;
    RECT 206.46 52.965 206.67 53.035 ;
    RECT 206.46 53.325 206.67 53.395 ;
    RECT 339.72 52.605 339.93 52.675 ;
    RECT 339.72 52.965 339.93 53.035 ;
    RECT 339.72 53.325 339.93 53.395 ;
    RECT 339.26 52.605 339.47 52.675 ;
    RECT 339.26 52.965 339.47 53.035 ;
    RECT 339.26 53.325 339.47 53.395 ;
    RECT 203.6 52.605 203.81 52.675 ;
    RECT 203.6 52.965 203.81 53.035 ;
    RECT 203.6 53.325 203.81 53.395 ;
    RECT 203.14 52.605 203.35 52.675 ;
    RECT 203.14 52.965 203.35 53.035 ;
    RECT 203.14 53.325 203.35 53.395 ;
    RECT 336.4 52.605 336.61 52.675 ;
    RECT 336.4 52.965 336.61 53.035 ;
    RECT 336.4 53.325 336.61 53.395 ;
    RECT 335.94 52.605 336.15 52.675 ;
    RECT 335.94 52.965 336.15 53.035 ;
    RECT 335.94 53.325 336.15 53.395 ;
    RECT 266.68 52.605 266.89 52.675 ;
    RECT 266.68 52.965 266.89 53.035 ;
    RECT 266.68 53.325 266.89 53.395 ;
    RECT 266.22 52.605 266.43 52.675 ;
    RECT 266.22 52.965 266.43 53.035 ;
    RECT 266.22 53.325 266.43 53.395 ;
    RECT 263.36 52.605 263.57 52.675 ;
    RECT 263.36 52.965 263.57 53.035 ;
    RECT 263.36 53.325 263.57 53.395 ;
    RECT 262.9 52.605 263.11 52.675 ;
    RECT 262.9 52.965 263.11 53.035 ;
    RECT 262.9 53.325 263.11 53.395 ;
    RECT 260.04 52.605 260.25 52.675 ;
    RECT 260.04 52.965 260.25 53.035 ;
    RECT 260.04 53.325 260.25 53.395 ;
    RECT 259.58 52.605 259.79 52.675 ;
    RECT 259.58 52.965 259.79 53.035 ;
    RECT 259.58 53.325 259.79 53.395 ;
    RECT 256.72 52.605 256.93 52.675 ;
    RECT 256.72 52.965 256.93 53.035 ;
    RECT 256.72 53.325 256.93 53.395 ;
    RECT 256.26 52.605 256.47 52.675 ;
    RECT 256.26 52.965 256.47 53.035 ;
    RECT 256.26 53.325 256.47 53.395 ;
    RECT 253.4 52.605 253.61 52.675 ;
    RECT 253.4 52.965 253.61 53.035 ;
    RECT 253.4 53.325 253.61 53.395 ;
    RECT 252.94 52.605 253.15 52.675 ;
    RECT 252.94 52.965 253.15 53.035 ;
    RECT 252.94 53.325 253.15 53.395 ;
    RECT 250.08 52.605 250.29 52.675 ;
    RECT 250.08 52.965 250.29 53.035 ;
    RECT 250.08 53.325 250.29 53.395 ;
    RECT 249.62 52.605 249.83 52.675 ;
    RECT 249.62 52.965 249.83 53.035 ;
    RECT 249.62 53.325 249.83 53.395 ;
    RECT 246.76 52.605 246.97 52.675 ;
    RECT 246.76 52.965 246.97 53.035 ;
    RECT 246.76 53.325 246.97 53.395 ;
    RECT 246.3 52.605 246.51 52.675 ;
    RECT 246.3 52.965 246.51 53.035 ;
    RECT 246.3 53.325 246.51 53.395 ;
    RECT 243.44 52.605 243.65 52.675 ;
    RECT 243.44 52.965 243.65 53.035 ;
    RECT 243.44 53.325 243.65 53.395 ;
    RECT 242.98 52.605 243.19 52.675 ;
    RECT 242.98 52.965 243.19 53.035 ;
    RECT 242.98 53.325 243.19 53.395 ;
    RECT 240.12 52.605 240.33 52.675 ;
    RECT 240.12 52.965 240.33 53.035 ;
    RECT 240.12 53.325 240.33 53.395 ;
    RECT 239.66 52.605 239.87 52.675 ;
    RECT 239.66 52.965 239.87 53.035 ;
    RECT 239.66 53.325 239.87 53.395 ;
    RECT 236.8 52.605 237.01 52.675 ;
    RECT 236.8 52.965 237.01 53.035 ;
    RECT 236.8 53.325 237.01 53.395 ;
    RECT 236.34 52.605 236.55 52.675 ;
    RECT 236.34 52.965 236.55 53.035 ;
    RECT 236.34 53.325 236.55 53.395 ;
    RECT 374.15 52.965 374.22 53.035 ;
    RECT 333.08 52.605 333.29 52.675 ;
    RECT 333.08 52.965 333.29 53.035 ;
    RECT 333.08 53.325 333.29 53.395 ;
    RECT 332.62 52.605 332.83 52.675 ;
    RECT 332.62 52.965 332.83 53.035 ;
    RECT 332.62 53.325 332.83 53.395 ;
    RECT 329.76 52.605 329.97 52.675 ;
    RECT 329.76 52.965 329.97 53.035 ;
    RECT 329.76 53.325 329.97 53.395 ;
    RECT 329.3 52.605 329.51 52.675 ;
    RECT 329.3 52.965 329.51 53.035 ;
    RECT 329.3 53.325 329.51 53.395 ;
    RECT 326.44 52.605 326.65 52.675 ;
    RECT 326.44 52.965 326.65 53.035 ;
    RECT 326.44 53.325 326.65 53.395 ;
    RECT 325.98 52.605 326.19 52.675 ;
    RECT 325.98 52.965 326.19 53.035 ;
    RECT 325.98 53.325 326.19 53.395 ;
    RECT 323.12 52.605 323.33 52.675 ;
    RECT 323.12 52.965 323.33 53.035 ;
    RECT 323.12 53.325 323.33 53.395 ;
    RECT 322.66 52.605 322.87 52.675 ;
    RECT 322.66 52.965 322.87 53.035 ;
    RECT 322.66 53.325 322.87 53.395 ;
    RECT 319.8 52.605 320.01 52.675 ;
    RECT 319.8 52.965 320.01 53.035 ;
    RECT 319.8 53.325 320.01 53.395 ;
    RECT 319.34 52.605 319.55 52.675 ;
    RECT 319.34 52.965 319.55 53.035 ;
    RECT 319.34 53.325 319.55 53.395 ;
    RECT 316.48 52.605 316.69 52.675 ;
    RECT 316.48 52.965 316.69 53.035 ;
    RECT 316.48 53.325 316.69 53.395 ;
    RECT 316.02 52.605 316.23 52.675 ;
    RECT 316.02 52.965 316.23 53.035 ;
    RECT 316.02 53.325 316.23 53.395 ;
    RECT 313.16 52.605 313.37 52.675 ;
    RECT 313.16 52.965 313.37 53.035 ;
    RECT 313.16 53.325 313.37 53.395 ;
    RECT 312.7 52.605 312.91 52.675 ;
    RECT 312.7 52.965 312.91 53.035 ;
    RECT 312.7 53.325 312.91 53.395 ;
    RECT 309.84 52.605 310.05 52.675 ;
    RECT 309.84 52.965 310.05 53.035 ;
    RECT 309.84 53.325 310.05 53.395 ;
    RECT 309.38 52.605 309.59 52.675 ;
    RECT 309.38 52.965 309.59 53.035 ;
    RECT 309.38 53.325 309.59 53.395 ;
    RECT 306.52 52.605 306.73 52.675 ;
    RECT 306.52 52.965 306.73 53.035 ;
    RECT 306.52 53.325 306.73 53.395 ;
    RECT 306.06 52.605 306.27 52.675 ;
    RECT 306.06 52.965 306.27 53.035 ;
    RECT 306.06 53.325 306.27 53.395 ;
    RECT 303.2 51.885 303.41 51.955 ;
    RECT 303.2 52.245 303.41 52.315 ;
    RECT 303.2 52.605 303.41 52.675 ;
    RECT 302.74 51.885 302.95 51.955 ;
    RECT 302.74 52.245 302.95 52.315 ;
    RECT 302.74 52.605 302.95 52.675 ;
    RECT 372.92 51.885 373.13 51.955 ;
    RECT 372.92 52.245 373.13 52.315 ;
    RECT 372.92 52.605 373.13 52.675 ;
    RECT 372.46 51.885 372.67 51.955 ;
    RECT 372.46 52.245 372.67 52.315 ;
    RECT 372.46 52.605 372.67 52.675 ;
    RECT 369.6 51.885 369.81 51.955 ;
    RECT 369.6 52.245 369.81 52.315 ;
    RECT 369.6 52.605 369.81 52.675 ;
    RECT 369.14 51.885 369.35 51.955 ;
    RECT 369.14 52.245 369.35 52.315 ;
    RECT 369.14 52.605 369.35 52.675 ;
    RECT 200.605 52.245 200.675 52.315 ;
    RECT 299.88 51.885 300.09 51.955 ;
    RECT 299.88 52.245 300.09 52.315 ;
    RECT 299.88 52.605 300.09 52.675 ;
    RECT 299.42 51.885 299.63 51.955 ;
    RECT 299.42 52.245 299.63 52.315 ;
    RECT 299.42 52.605 299.63 52.675 ;
    RECT 296.56 51.885 296.77 51.955 ;
    RECT 296.56 52.245 296.77 52.315 ;
    RECT 296.56 52.605 296.77 52.675 ;
    RECT 296.1 51.885 296.31 51.955 ;
    RECT 296.1 52.245 296.31 52.315 ;
    RECT 296.1 52.605 296.31 52.675 ;
    RECT 293.24 51.885 293.45 51.955 ;
    RECT 293.24 52.245 293.45 52.315 ;
    RECT 293.24 52.605 293.45 52.675 ;
    RECT 292.78 51.885 292.99 51.955 ;
    RECT 292.78 52.245 292.99 52.315 ;
    RECT 292.78 52.605 292.99 52.675 ;
    RECT 289.92 51.885 290.13 51.955 ;
    RECT 289.92 52.245 290.13 52.315 ;
    RECT 289.92 52.605 290.13 52.675 ;
    RECT 289.46 51.885 289.67 51.955 ;
    RECT 289.46 52.245 289.67 52.315 ;
    RECT 289.46 52.605 289.67 52.675 ;
    RECT 286.6 51.885 286.81 51.955 ;
    RECT 286.6 52.245 286.81 52.315 ;
    RECT 286.6 52.605 286.81 52.675 ;
    RECT 286.14 51.885 286.35 51.955 ;
    RECT 286.14 52.245 286.35 52.315 ;
    RECT 286.14 52.605 286.35 52.675 ;
    RECT 283.28 51.885 283.49 51.955 ;
    RECT 283.28 52.245 283.49 52.315 ;
    RECT 283.28 52.605 283.49 52.675 ;
    RECT 282.82 51.885 283.03 51.955 ;
    RECT 282.82 52.245 283.03 52.315 ;
    RECT 282.82 52.605 283.03 52.675 ;
    RECT 279.96 51.885 280.17 51.955 ;
    RECT 279.96 52.245 280.17 52.315 ;
    RECT 279.96 52.605 280.17 52.675 ;
    RECT 279.5 51.885 279.71 51.955 ;
    RECT 279.5 52.245 279.71 52.315 ;
    RECT 279.5 52.605 279.71 52.675 ;
    RECT 276.64 51.885 276.85 51.955 ;
    RECT 276.64 52.245 276.85 52.315 ;
    RECT 276.64 52.605 276.85 52.675 ;
    RECT 276.18 51.885 276.39 51.955 ;
    RECT 276.18 52.245 276.39 52.315 ;
    RECT 276.18 52.605 276.39 52.675 ;
    RECT 273.32 51.885 273.53 51.955 ;
    RECT 273.32 52.245 273.53 52.315 ;
    RECT 273.32 52.605 273.53 52.675 ;
    RECT 272.86 51.885 273.07 51.955 ;
    RECT 272.86 52.245 273.07 52.315 ;
    RECT 272.86 52.605 273.07 52.675 ;
    RECT 270.0 51.885 270.21 51.955 ;
    RECT 270.0 52.245 270.21 52.315 ;
    RECT 270.0 52.605 270.21 52.675 ;
    RECT 269.54 51.885 269.75 51.955 ;
    RECT 269.54 52.245 269.75 52.315 ;
    RECT 269.54 52.605 269.75 52.675 ;
    RECT 233.48 51.885 233.69 51.955 ;
    RECT 233.48 52.245 233.69 52.315 ;
    RECT 233.48 52.605 233.69 52.675 ;
    RECT 233.02 51.885 233.23 51.955 ;
    RECT 233.02 52.245 233.23 52.315 ;
    RECT 233.02 52.605 233.23 52.675 ;
    RECT 230.16 51.885 230.37 51.955 ;
    RECT 230.16 52.245 230.37 52.315 ;
    RECT 230.16 52.605 230.37 52.675 ;
    RECT 229.7 51.885 229.91 51.955 ;
    RECT 229.7 52.245 229.91 52.315 ;
    RECT 229.7 52.605 229.91 52.675 ;
    RECT 366.28 51.885 366.49 51.955 ;
    RECT 366.28 52.245 366.49 52.315 ;
    RECT 366.28 52.605 366.49 52.675 ;
    RECT 365.82 51.885 366.03 51.955 ;
    RECT 365.82 52.245 366.03 52.315 ;
    RECT 365.82 52.605 366.03 52.675 ;
    RECT 226.84 51.885 227.05 51.955 ;
    RECT 226.84 52.245 227.05 52.315 ;
    RECT 226.84 52.605 227.05 52.675 ;
    RECT 226.38 51.885 226.59 51.955 ;
    RECT 226.38 52.245 226.59 52.315 ;
    RECT 226.38 52.605 226.59 52.675 ;
    RECT 362.96 51.885 363.17 51.955 ;
    RECT 362.96 52.245 363.17 52.315 ;
    RECT 362.96 52.605 363.17 52.675 ;
    RECT 362.5 51.885 362.71 51.955 ;
    RECT 362.5 52.245 362.71 52.315 ;
    RECT 362.5 52.605 362.71 52.675 ;
    RECT 223.52 51.885 223.73 51.955 ;
    RECT 223.52 52.245 223.73 52.315 ;
    RECT 223.52 52.605 223.73 52.675 ;
    RECT 223.06 51.885 223.27 51.955 ;
    RECT 223.06 52.245 223.27 52.315 ;
    RECT 223.06 52.605 223.27 52.675 ;
    RECT 359.64 51.885 359.85 51.955 ;
    RECT 359.64 52.245 359.85 52.315 ;
    RECT 359.64 52.605 359.85 52.675 ;
    RECT 359.18 51.885 359.39 51.955 ;
    RECT 359.18 52.245 359.39 52.315 ;
    RECT 359.18 52.605 359.39 52.675 ;
    RECT 220.2 51.885 220.41 51.955 ;
    RECT 220.2 52.245 220.41 52.315 ;
    RECT 220.2 52.605 220.41 52.675 ;
    RECT 219.74 51.885 219.95 51.955 ;
    RECT 219.74 52.245 219.95 52.315 ;
    RECT 219.74 52.605 219.95 52.675 ;
    RECT 356.32 51.885 356.53 51.955 ;
    RECT 356.32 52.245 356.53 52.315 ;
    RECT 356.32 52.605 356.53 52.675 ;
    RECT 355.86 51.885 356.07 51.955 ;
    RECT 355.86 52.245 356.07 52.315 ;
    RECT 355.86 52.605 356.07 52.675 ;
    RECT 353.0 51.885 353.21 51.955 ;
    RECT 353.0 52.245 353.21 52.315 ;
    RECT 353.0 52.605 353.21 52.675 ;
    RECT 352.54 51.885 352.75 51.955 ;
    RECT 352.54 52.245 352.75 52.315 ;
    RECT 352.54 52.605 352.75 52.675 ;
    RECT 216.88 51.885 217.09 51.955 ;
    RECT 216.88 52.245 217.09 52.315 ;
    RECT 216.88 52.605 217.09 52.675 ;
    RECT 216.42 51.885 216.63 51.955 ;
    RECT 216.42 52.245 216.63 52.315 ;
    RECT 216.42 52.605 216.63 52.675 ;
    RECT 349.68 51.885 349.89 51.955 ;
    RECT 349.68 52.245 349.89 52.315 ;
    RECT 349.68 52.605 349.89 52.675 ;
    RECT 349.22 51.885 349.43 51.955 ;
    RECT 349.22 52.245 349.43 52.315 ;
    RECT 349.22 52.605 349.43 52.675 ;
    RECT 213.56 51.885 213.77 51.955 ;
    RECT 213.56 52.245 213.77 52.315 ;
    RECT 213.56 52.605 213.77 52.675 ;
    RECT 213.1 51.885 213.31 51.955 ;
    RECT 213.1 52.245 213.31 52.315 ;
    RECT 213.1 52.605 213.31 52.675 ;
    RECT 346.36 51.885 346.57 51.955 ;
    RECT 346.36 52.245 346.57 52.315 ;
    RECT 346.36 52.605 346.57 52.675 ;
    RECT 345.9 51.885 346.11 51.955 ;
    RECT 345.9 52.245 346.11 52.315 ;
    RECT 345.9 52.605 346.11 52.675 ;
    RECT 210.24 51.885 210.45 51.955 ;
    RECT 210.24 52.245 210.45 52.315 ;
    RECT 210.24 52.605 210.45 52.675 ;
    RECT 209.78 51.885 209.99 51.955 ;
    RECT 209.78 52.245 209.99 52.315 ;
    RECT 209.78 52.605 209.99 52.675 ;
    RECT 343.04 51.885 343.25 51.955 ;
    RECT 343.04 52.245 343.25 52.315 ;
    RECT 343.04 52.605 343.25 52.675 ;
    RECT 342.58 51.885 342.79 51.955 ;
    RECT 342.58 52.245 342.79 52.315 ;
    RECT 342.58 52.605 342.79 52.675 ;
    RECT 206.92 51.885 207.13 51.955 ;
    RECT 206.92 52.245 207.13 52.315 ;
    RECT 206.92 52.605 207.13 52.675 ;
    RECT 206.46 51.885 206.67 51.955 ;
    RECT 206.46 52.245 206.67 52.315 ;
    RECT 206.46 52.605 206.67 52.675 ;
    RECT 339.72 51.885 339.93 51.955 ;
    RECT 339.72 52.245 339.93 52.315 ;
    RECT 339.72 52.605 339.93 52.675 ;
    RECT 339.26 51.885 339.47 51.955 ;
    RECT 339.26 52.245 339.47 52.315 ;
    RECT 339.26 52.605 339.47 52.675 ;
    RECT 203.6 51.885 203.81 51.955 ;
    RECT 203.6 52.245 203.81 52.315 ;
    RECT 203.6 52.605 203.81 52.675 ;
    RECT 203.14 51.885 203.35 51.955 ;
    RECT 203.14 52.245 203.35 52.315 ;
    RECT 203.14 52.605 203.35 52.675 ;
    RECT 336.4 51.885 336.61 51.955 ;
    RECT 336.4 52.245 336.61 52.315 ;
    RECT 336.4 52.605 336.61 52.675 ;
    RECT 335.94 51.885 336.15 51.955 ;
    RECT 335.94 52.245 336.15 52.315 ;
    RECT 335.94 52.605 336.15 52.675 ;
    RECT 266.68 51.885 266.89 51.955 ;
    RECT 266.68 52.245 266.89 52.315 ;
    RECT 266.68 52.605 266.89 52.675 ;
    RECT 266.22 51.885 266.43 51.955 ;
    RECT 266.22 52.245 266.43 52.315 ;
    RECT 266.22 52.605 266.43 52.675 ;
    RECT 263.36 51.885 263.57 51.955 ;
    RECT 263.36 52.245 263.57 52.315 ;
    RECT 263.36 52.605 263.57 52.675 ;
    RECT 262.9 51.885 263.11 51.955 ;
    RECT 262.9 52.245 263.11 52.315 ;
    RECT 262.9 52.605 263.11 52.675 ;
    RECT 260.04 51.885 260.25 51.955 ;
    RECT 260.04 52.245 260.25 52.315 ;
    RECT 260.04 52.605 260.25 52.675 ;
    RECT 259.58 51.885 259.79 51.955 ;
    RECT 259.58 52.245 259.79 52.315 ;
    RECT 259.58 52.605 259.79 52.675 ;
    RECT 256.72 51.885 256.93 51.955 ;
    RECT 256.72 52.245 256.93 52.315 ;
    RECT 256.72 52.605 256.93 52.675 ;
    RECT 256.26 51.885 256.47 51.955 ;
    RECT 256.26 52.245 256.47 52.315 ;
    RECT 256.26 52.605 256.47 52.675 ;
    RECT 253.4 51.885 253.61 51.955 ;
    RECT 253.4 52.245 253.61 52.315 ;
    RECT 253.4 52.605 253.61 52.675 ;
    RECT 252.94 51.885 253.15 51.955 ;
    RECT 252.94 52.245 253.15 52.315 ;
    RECT 252.94 52.605 253.15 52.675 ;
    RECT 250.08 51.885 250.29 51.955 ;
    RECT 250.08 52.245 250.29 52.315 ;
    RECT 250.08 52.605 250.29 52.675 ;
    RECT 249.62 51.885 249.83 51.955 ;
    RECT 249.62 52.245 249.83 52.315 ;
    RECT 249.62 52.605 249.83 52.675 ;
    RECT 246.76 51.885 246.97 51.955 ;
    RECT 246.76 52.245 246.97 52.315 ;
    RECT 246.76 52.605 246.97 52.675 ;
    RECT 246.3 51.885 246.51 51.955 ;
    RECT 246.3 52.245 246.51 52.315 ;
    RECT 246.3 52.605 246.51 52.675 ;
    RECT 243.44 51.885 243.65 51.955 ;
    RECT 243.44 52.245 243.65 52.315 ;
    RECT 243.44 52.605 243.65 52.675 ;
    RECT 242.98 51.885 243.19 51.955 ;
    RECT 242.98 52.245 243.19 52.315 ;
    RECT 242.98 52.605 243.19 52.675 ;
    RECT 240.12 51.885 240.33 51.955 ;
    RECT 240.12 52.245 240.33 52.315 ;
    RECT 240.12 52.605 240.33 52.675 ;
    RECT 239.66 51.885 239.87 51.955 ;
    RECT 239.66 52.245 239.87 52.315 ;
    RECT 239.66 52.605 239.87 52.675 ;
    RECT 236.8 51.885 237.01 51.955 ;
    RECT 236.8 52.245 237.01 52.315 ;
    RECT 236.8 52.605 237.01 52.675 ;
    RECT 236.34 51.885 236.55 51.955 ;
    RECT 236.34 52.245 236.55 52.315 ;
    RECT 236.34 52.605 236.55 52.675 ;
    RECT 374.15 52.245 374.22 52.315 ;
    RECT 333.08 51.885 333.29 51.955 ;
    RECT 333.08 52.245 333.29 52.315 ;
    RECT 333.08 52.605 333.29 52.675 ;
    RECT 332.62 51.885 332.83 51.955 ;
    RECT 332.62 52.245 332.83 52.315 ;
    RECT 332.62 52.605 332.83 52.675 ;
    RECT 329.76 51.885 329.97 51.955 ;
    RECT 329.76 52.245 329.97 52.315 ;
    RECT 329.76 52.605 329.97 52.675 ;
    RECT 329.3 51.885 329.51 51.955 ;
    RECT 329.3 52.245 329.51 52.315 ;
    RECT 329.3 52.605 329.51 52.675 ;
    RECT 326.44 51.885 326.65 51.955 ;
    RECT 326.44 52.245 326.65 52.315 ;
    RECT 326.44 52.605 326.65 52.675 ;
    RECT 325.98 51.885 326.19 51.955 ;
    RECT 325.98 52.245 326.19 52.315 ;
    RECT 325.98 52.605 326.19 52.675 ;
    RECT 323.12 51.885 323.33 51.955 ;
    RECT 323.12 52.245 323.33 52.315 ;
    RECT 323.12 52.605 323.33 52.675 ;
    RECT 322.66 51.885 322.87 51.955 ;
    RECT 322.66 52.245 322.87 52.315 ;
    RECT 322.66 52.605 322.87 52.675 ;
    RECT 319.8 51.885 320.01 51.955 ;
    RECT 319.8 52.245 320.01 52.315 ;
    RECT 319.8 52.605 320.01 52.675 ;
    RECT 319.34 51.885 319.55 51.955 ;
    RECT 319.34 52.245 319.55 52.315 ;
    RECT 319.34 52.605 319.55 52.675 ;
    RECT 316.48 51.885 316.69 51.955 ;
    RECT 316.48 52.245 316.69 52.315 ;
    RECT 316.48 52.605 316.69 52.675 ;
    RECT 316.02 51.885 316.23 51.955 ;
    RECT 316.02 52.245 316.23 52.315 ;
    RECT 316.02 52.605 316.23 52.675 ;
    RECT 313.16 51.885 313.37 51.955 ;
    RECT 313.16 52.245 313.37 52.315 ;
    RECT 313.16 52.605 313.37 52.675 ;
    RECT 312.7 51.885 312.91 51.955 ;
    RECT 312.7 52.245 312.91 52.315 ;
    RECT 312.7 52.605 312.91 52.675 ;
    RECT 309.84 51.885 310.05 51.955 ;
    RECT 309.84 52.245 310.05 52.315 ;
    RECT 309.84 52.605 310.05 52.675 ;
    RECT 309.38 51.885 309.59 51.955 ;
    RECT 309.38 52.245 309.59 52.315 ;
    RECT 309.38 52.605 309.59 52.675 ;
    RECT 306.52 51.885 306.73 51.955 ;
    RECT 306.52 52.245 306.73 52.315 ;
    RECT 306.52 52.605 306.73 52.675 ;
    RECT 306.06 51.885 306.27 51.955 ;
    RECT 306.06 52.245 306.27 52.315 ;
    RECT 306.06 52.605 306.27 52.675 ;
    RECT 303.2 51.165 303.41 51.235 ;
    RECT 303.2 51.525 303.41 51.595 ;
    RECT 303.2 51.885 303.41 51.955 ;
    RECT 302.74 51.165 302.95 51.235 ;
    RECT 302.74 51.525 302.95 51.595 ;
    RECT 302.74 51.885 302.95 51.955 ;
    RECT 372.92 51.165 373.13 51.235 ;
    RECT 372.92 51.525 373.13 51.595 ;
    RECT 372.92 51.885 373.13 51.955 ;
    RECT 372.46 51.165 372.67 51.235 ;
    RECT 372.46 51.525 372.67 51.595 ;
    RECT 372.46 51.885 372.67 51.955 ;
    RECT 369.6 51.165 369.81 51.235 ;
    RECT 369.6 51.525 369.81 51.595 ;
    RECT 369.6 51.885 369.81 51.955 ;
    RECT 369.14 51.165 369.35 51.235 ;
    RECT 369.14 51.525 369.35 51.595 ;
    RECT 369.14 51.885 369.35 51.955 ;
    RECT 200.605 51.525 200.675 51.595 ;
    RECT 299.88 51.165 300.09 51.235 ;
    RECT 299.88 51.525 300.09 51.595 ;
    RECT 299.88 51.885 300.09 51.955 ;
    RECT 299.42 51.165 299.63 51.235 ;
    RECT 299.42 51.525 299.63 51.595 ;
    RECT 299.42 51.885 299.63 51.955 ;
    RECT 296.56 51.165 296.77 51.235 ;
    RECT 296.56 51.525 296.77 51.595 ;
    RECT 296.56 51.885 296.77 51.955 ;
    RECT 296.1 51.165 296.31 51.235 ;
    RECT 296.1 51.525 296.31 51.595 ;
    RECT 296.1 51.885 296.31 51.955 ;
    RECT 293.24 51.165 293.45 51.235 ;
    RECT 293.24 51.525 293.45 51.595 ;
    RECT 293.24 51.885 293.45 51.955 ;
    RECT 292.78 51.165 292.99 51.235 ;
    RECT 292.78 51.525 292.99 51.595 ;
    RECT 292.78 51.885 292.99 51.955 ;
    RECT 289.92 51.165 290.13 51.235 ;
    RECT 289.92 51.525 290.13 51.595 ;
    RECT 289.92 51.885 290.13 51.955 ;
    RECT 289.46 51.165 289.67 51.235 ;
    RECT 289.46 51.525 289.67 51.595 ;
    RECT 289.46 51.885 289.67 51.955 ;
    RECT 286.6 51.165 286.81 51.235 ;
    RECT 286.6 51.525 286.81 51.595 ;
    RECT 286.6 51.885 286.81 51.955 ;
    RECT 286.14 51.165 286.35 51.235 ;
    RECT 286.14 51.525 286.35 51.595 ;
    RECT 286.14 51.885 286.35 51.955 ;
    RECT 283.28 51.165 283.49 51.235 ;
    RECT 283.28 51.525 283.49 51.595 ;
    RECT 283.28 51.885 283.49 51.955 ;
    RECT 282.82 51.165 283.03 51.235 ;
    RECT 282.82 51.525 283.03 51.595 ;
    RECT 282.82 51.885 283.03 51.955 ;
    RECT 279.96 51.165 280.17 51.235 ;
    RECT 279.96 51.525 280.17 51.595 ;
    RECT 279.96 51.885 280.17 51.955 ;
    RECT 279.5 51.165 279.71 51.235 ;
    RECT 279.5 51.525 279.71 51.595 ;
    RECT 279.5 51.885 279.71 51.955 ;
    RECT 276.64 51.165 276.85 51.235 ;
    RECT 276.64 51.525 276.85 51.595 ;
    RECT 276.64 51.885 276.85 51.955 ;
    RECT 276.18 51.165 276.39 51.235 ;
    RECT 276.18 51.525 276.39 51.595 ;
    RECT 276.18 51.885 276.39 51.955 ;
    RECT 273.32 51.165 273.53 51.235 ;
    RECT 273.32 51.525 273.53 51.595 ;
    RECT 273.32 51.885 273.53 51.955 ;
    RECT 272.86 51.165 273.07 51.235 ;
    RECT 272.86 51.525 273.07 51.595 ;
    RECT 272.86 51.885 273.07 51.955 ;
    RECT 270.0 51.165 270.21 51.235 ;
    RECT 270.0 51.525 270.21 51.595 ;
    RECT 270.0 51.885 270.21 51.955 ;
    RECT 269.54 51.165 269.75 51.235 ;
    RECT 269.54 51.525 269.75 51.595 ;
    RECT 269.54 51.885 269.75 51.955 ;
    RECT 233.48 51.165 233.69 51.235 ;
    RECT 233.48 51.525 233.69 51.595 ;
    RECT 233.48 51.885 233.69 51.955 ;
    RECT 233.02 51.165 233.23 51.235 ;
    RECT 233.02 51.525 233.23 51.595 ;
    RECT 233.02 51.885 233.23 51.955 ;
    RECT 230.16 51.165 230.37 51.235 ;
    RECT 230.16 51.525 230.37 51.595 ;
    RECT 230.16 51.885 230.37 51.955 ;
    RECT 229.7 51.165 229.91 51.235 ;
    RECT 229.7 51.525 229.91 51.595 ;
    RECT 229.7 51.885 229.91 51.955 ;
    RECT 366.28 51.165 366.49 51.235 ;
    RECT 366.28 51.525 366.49 51.595 ;
    RECT 366.28 51.885 366.49 51.955 ;
    RECT 365.82 51.165 366.03 51.235 ;
    RECT 365.82 51.525 366.03 51.595 ;
    RECT 365.82 51.885 366.03 51.955 ;
    RECT 226.84 51.165 227.05 51.235 ;
    RECT 226.84 51.525 227.05 51.595 ;
    RECT 226.84 51.885 227.05 51.955 ;
    RECT 226.38 51.165 226.59 51.235 ;
    RECT 226.38 51.525 226.59 51.595 ;
    RECT 226.38 51.885 226.59 51.955 ;
    RECT 362.96 51.165 363.17 51.235 ;
    RECT 362.96 51.525 363.17 51.595 ;
    RECT 362.96 51.885 363.17 51.955 ;
    RECT 362.5 51.165 362.71 51.235 ;
    RECT 362.5 51.525 362.71 51.595 ;
    RECT 362.5 51.885 362.71 51.955 ;
    RECT 223.52 51.165 223.73 51.235 ;
    RECT 223.52 51.525 223.73 51.595 ;
    RECT 223.52 51.885 223.73 51.955 ;
    RECT 223.06 51.165 223.27 51.235 ;
    RECT 223.06 51.525 223.27 51.595 ;
    RECT 223.06 51.885 223.27 51.955 ;
    RECT 359.64 51.165 359.85 51.235 ;
    RECT 359.64 51.525 359.85 51.595 ;
    RECT 359.64 51.885 359.85 51.955 ;
    RECT 359.18 51.165 359.39 51.235 ;
    RECT 359.18 51.525 359.39 51.595 ;
    RECT 359.18 51.885 359.39 51.955 ;
    RECT 220.2 51.165 220.41 51.235 ;
    RECT 220.2 51.525 220.41 51.595 ;
    RECT 220.2 51.885 220.41 51.955 ;
    RECT 219.74 51.165 219.95 51.235 ;
    RECT 219.74 51.525 219.95 51.595 ;
    RECT 219.74 51.885 219.95 51.955 ;
    RECT 356.32 51.165 356.53 51.235 ;
    RECT 356.32 51.525 356.53 51.595 ;
    RECT 356.32 51.885 356.53 51.955 ;
    RECT 355.86 51.165 356.07 51.235 ;
    RECT 355.86 51.525 356.07 51.595 ;
    RECT 355.86 51.885 356.07 51.955 ;
    RECT 353.0 51.165 353.21 51.235 ;
    RECT 353.0 51.525 353.21 51.595 ;
    RECT 353.0 51.885 353.21 51.955 ;
    RECT 352.54 51.165 352.75 51.235 ;
    RECT 352.54 51.525 352.75 51.595 ;
    RECT 352.54 51.885 352.75 51.955 ;
    RECT 216.88 51.165 217.09 51.235 ;
    RECT 216.88 51.525 217.09 51.595 ;
    RECT 216.88 51.885 217.09 51.955 ;
    RECT 216.42 51.165 216.63 51.235 ;
    RECT 216.42 51.525 216.63 51.595 ;
    RECT 216.42 51.885 216.63 51.955 ;
    RECT 349.68 51.165 349.89 51.235 ;
    RECT 349.68 51.525 349.89 51.595 ;
    RECT 349.68 51.885 349.89 51.955 ;
    RECT 349.22 51.165 349.43 51.235 ;
    RECT 349.22 51.525 349.43 51.595 ;
    RECT 349.22 51.885 349.43 51.955 ;
    RECT 213.56 51.165 213.77 51.235 ;
    RECT 213.56 51.525 213.77 51.595 ;
    RECT 213.56 51.885 213.77 51.955 ;
    RECT 213.1 51.165 213.31 51.235 ;
    RECT 213.1 51.525 213.31 51.595 ;
    RECT 213.1 51.885 213.31 51.955 ;
    RECT 346.36 51.165 346.57 51.235 ;
    RECT 346.36 51.525 346.57 51.595 ;
    RECT 346.36 51.885 346.57 51.955 ;
    RECT 345.9 51.165 346.11 51.235 ;
    RECT 345.9 51.525 346.11 51.595 ;
    RECT 345.9 51.885 346.11 51.955 ;
    RECT 210.24 51.165 210.45 51.235 ;
    RECT 210.24 51.525 210.45 51.595 ;
    RECT 210.24 51.885 210.45 51.955 ;
    RECT 209.78 51.165 209.99 51.235 ;
    RECT 209.78 51.525 209.99 51.595 ;
    RECT 209.78 51.885 209.99 51.955 ;
    RECT 343.04 51.165 343.25 51.235 ;
    RECT 343.04 51.525 343.25 51.595 ;
    RECT 343.04 51.885 343.25 51.955 ;
    RECT 342.58 51.165 342.79 51.235 ;
    RECT 342.58 51.525 342.79 51.595 ;
    RECT 342.58 51.885 342.79 51.955 ;
    RECT 206.92 51.165 207.13 51.235 ;
    RECT 206.92 51.525 207.13 51.595 ;
    RECT 206.92 51.885 207.13 51.955 ;
    RECT 206.46 51.165 206.67 51.235 ;
    RECT 206.46 51.525 206.67 51.595 ;
    RECT 206.46 51.885 206.67 51.955 ;
    RECT 339.72 51.165 339.93 51.235 ;
    RECT 339.72 51.525 339.93 51.595 ;
    RECT 339.72 51.885 339.93 51.955 ;
    RECT 339.26 51.165 339.47 51.235 ;
    RECT 339.26 51.525 339.47 51.595 ;
    RECT 339.26 51.885 339.47 51.955 ;
    RECT 203.6 51.165 203.81 51.235 ;
    RECT 203.6 51.525 203.81 51.595 ;
    RECT 203.6 51.885 203.81 51.955 ;
    RECT 203.14 51.165 203.35 51.235 ;
    RECT 203.14 51.525 203.35 51.595 ;
    RECT 203.14 51.885 203.35 51.955 ;
    RECT 336.4 51.165 336.61 51.235 ;
    RECT 336.4 51.525 336.61 51.595 ;
    RECT 336.4 51.885 336.61 51.955 ;
    RECT 335.94 51.165 336.15 51.235 ;
    RECT 335.94 51.525 336.15 51.595 ;
    RECT 335.94 51.885 336.15 51.955 ;
    RECT 266.68 51.165 266.89 51.235 ;
    RECT 266.68 51.525 266.89 51.595 ;
    RECT 266.68 51.885 266.89 51.955 ;
    RECT 266.22 51.165 266.43 51.235 ;
    RECT 266.22 51.525 266.43 51.595 ;
    RECT 266.22 51.885 266.43 51.955 ;
    RECT 263.36 51.165 263.57 51.235 ;
    RECT 263.36 51.525 263.57 51.595 ;
    RECT 263.36 51.885 263.57 51.955 ;
    RECT 262.9 51.165 263.11 51.235 ;
    RECT 262.9 51.525 263.11 51.595 ;
    RECT 262.9 51.885 263.11 51.955 ;
    RECT 260.04 51.165 260.25 51.235 ;
    RECT 260.04 51.525 260.25 51.595 ;
    RECT 260.04 51.885 260.25 51.955 ;
    RECT 259.58 51.165 259.79 51.235 ;
    RECT 259.58 51.525 259.79 51.595 ;
    RECT 259.58 51.885 259.79 51.955 ;
    RECT 256.72 51.165 256.93 51.235 ;
    RECT 256.72 51.525 256.93 51.595 ;
    RECT 256.72 51.885 256.93 51.955 ;
    RECT 256.26 51.165 256.47 51.235 ;
    RECT 256.26 51.525 256.47 51.595 ;
    RECT 256.26 51.885 256.47 51.955 ;
    RECT 253.4 51.165 253.61 51.235 ;
    RECT 253.4 51.525 253.61 51.595 ;
    RECT 253.4 51.885 253.61 51.955 ;
    RECT 252.94 51.165 253.15 51.235 ;
    RECT 252.94 51.525 253.15 51.595 ;
    RECT 252.94 51.885 253.15 51.955 ;
    RECT 250.08 51.165 250.29 51.235 ;
    RECT 250.08 51.525 250.29 51.595 ;
    RECT 250.08 51.885 250.29 51.955 ;
    RECT 249.62 51.165 249.83 51.235 ;
    RECT 249.62 51.525 249.83 51.595 ;
    RECT 249.62 51.885 249.83 51.955 ;
    RECT 246.76 51.165 246.97 51.235 ;
    RECT 246.76 51.525 246.97 51.595 ;
    RECT 246.76 51.885 246.97 51.955 ;
    RECT 246.3 51.165 246.51 51.235 ;
    RECT 246.3 51.525 246.51 51.595 ;
    RECT 246.3 51.885 246.51 51.955 ;
    RECT 243.44 51.165 243.65 51.235 ;
    RECT 243.44 51.525 243.65 51.595 ;
    RECT 243.44 51.885 243.65 51.955 ;
    RECT 242.98 51.165 243.19 51.235 ;
    RECT 242.98 51.525 243.19 51.595 ;
    RECT 242.98 51.885 243.19 51.955 ;
    RECT 240.12 51.165 240.33 51.235 ;
    RECT 240.12 51.525 240.33 51.595 ;
    RECT 240.12 51.885 240.33 51.955 ;
    RECT 239.66 51.165 239.87 51.235 ;
    RECT 239.66 51.525 239.87 51.595 ;
    RECT 239.66 51.885 239.87 51.955 ;
    RECT 236.8 51.165 237.01 51.235 ;
    RECT 236.8 51.525 237.01 51.595 ;
    RECT 236.8 51.885 237.01 51.955 ;
    RECT 236.34 51.165 236.55 51.235 ;
    RECT 236.34 51.525 236.55 51.595 ;
    RECT 236.34 51.885 236.55 51.955 ;
    RECT 374.15 51.525 374.22 51.595 ;
    RECT 333.08 51.165 333.29 51.235 ;
    RECT 333.08 51.525 333.29 51.595 ;
    RECT 333.08 51.885 333.29 51.955 ;
    RECT 332.62 51.165 332.83 51.235 ;
    RECT 332.62 51.525 332.83 51.595 ;
    RECT 332.62 51.885 332.83 51.955 ;
    RECT 329.76 51.165 329.97 51.235 ;
    RECT 329.76 51.525 329.97 51.595 ;
    RECT 329.76 51.885 329.97 51.955 ;
    RECT 329.3 51.165 329.51 51.235 ;
    RECT 329.3 51.525 329.51 51.595 ;
    RECT 329.3 51.885 329.51 51.955 ;
    RECT 326.44 51.165 326.65 51.235 ;
    RECT 326.44 51.525 326.65 51.595 ;
    RECT 326.44 51.885 326.65 51.955 ;
    RECT 325.98 51.165 326.19 51.235 ;
    RECT 325.98 51.525 326.19 51.595 ;
    RECT 325.98 51.885 326.19 51.955 ;
    RECT 323.12 51.165 323.33 51.235 ;
    RECT 323.12 51.525 323.33 51.595 ;
    RECT 323.12 51.885 323.33 51.955 ;
    RECT 322.66 51.165 322.87 51.235 ;
    RECT 322.66 51.525 322.87 51.595 ;
    RECT 322.66 51.885 322.87 51.955 ;
    RECT 319.8 51.165 320.01 51.235 ;
    RECT 319.8 51.525 320.01 51.595 ;
    RECT 319.8 51.885 320.01 51.955 ;
    RECT 319.34 51.165 319.55 51.235 ;
    RECT 319.34 51.525 319.55 51.595 ;
    RECT 319.34 51.885 319.55 51.955 ;
    RECT 316.48 51.165 316.69 51.235 ;
    RECT 316.48 51.525 316.69 51.595 ;
    RECT 316.48 51.885 316.69 51.955 ;
    RECT 316.02 51.165 316.23 51.235 ;
    RECT 316.02 51.525 316.23 51.595 ;
    RECT 316.02 51.885 316.23 51.955 ;
    RECT 313.16 51.165 313.37 51.235 ;
    RECT 313.16 51.525 313.37 51.595 ;
    RECT 313.16 51.885 313.37 51.955 ;
    RECT 312.7 51.165 312.91 51.235 ;
    RECT 312.7 51.525 312.91 51.595 ;
    RECT 312.7 51.885 312.91 51.955 ;
    RECT 309.84 51.165 310.05 51.235 ;
    RECT 309.84 51.525 310.05 51.595 ;
    RECT 309.84 51.885 310.05 51.955 ;
    RECT 309.38 51.165 309.59 51.235 ;
    RECT 309.38 51.525 309.59 51.595 ;
    RECT 309.38 51.885 309.59 51.955 ;
    RECT 306.52 51.165 306.73 51.235 ;
    RECT 306.52 51.525 306.73 51.595 ;
    RECT 306.52 51.885 306.73 51.955 ;
    RECT 306.06 51.165 306.27 51.235 ;
    RECT 306.06 51.525 306.27 51.595 ;
    RECT 306.06 51.885 306.27 51.955 ;
    RECT 303.2 50.445 303.41 50.515 ;
    RECT 303.2 50.805 303.41 50.875 ;
    RECT 303.2 51.165 303.41 51.235 ;
    RECT 302.74 50.445 302.95 50.515 ;
    RECT 302.74 50.805 302.95 50.875 ;
    RECT 302.74 51.165 302.95 51.235 ;
    RECT 372.92 50.445 373.13 50.515 ;
    RECT 372.92 50.805 373.13 50.875 ;
    RECT 372.92 51.165 373.13 51.235 ;
    RECT 372.46 50.445 372.67 50.515 ;
    RECT 372.46 50.805 372.67 50.875 ;
    RECT 372.46 51.165 372.67 51.235 ;
    RECT 369.6 50.445 369.81 50.515 ;
    RECT 369.6 50.805 369.81 50.875 ;
    RECT 369.6 51.165 369.81 51.235 ;
    RECT 369.14 50.445 369.35 50.515 ;
    RECT 369.14 50.805 369.35 50.875 ;
    RECT 369.14 51.165 369.35 51.235 ;
    RECT 200.605 50.805 200.675 50.875 ;
    RECT 299.88 50.445 300.09 50.515 ;
    RECT 299.88 50.805 300.09 50.875 ;
    RECT 299.88 51.165 300.09 51.235 ;
    RECT 299.42 50.445 299.63 50.515 ;
    RECT 299.42 50.805 299.63 50.875 ;
    RECT 299.42 51.165 299.63 51.235 ;
    RECT 296.56 50.445 296.77 50.515 ;
    RECT 296.56 50.805 296.77 50.875 ;
    RECT 296.56 51.165 296.77 51.235 ;
    RECT 296.1 50.445 296.31 50.515 ;
    RECT 296.1 50.805 296.31 50.875 ;
    RECT 296.1 51.165 296.31 51.235 ;
    RECT 293.24 50.445 293.45 50.515 ;
    RECT 293.24 50.805 293.45 50.875 ;
    RECT 293.24 51.165 293.45 51.235 ;
    RECT 292.78 50.445 292.99 50.515 ;
    RECT 292.78 50.805 292.99 50.875 ;
    RECT 292.78 51.165 292.99 51.235 ;
    RECT 289.92 50.445 290.13 50.515 ;
    RECT 289.92 50.805 290.13 50.875 ;
    RECT 289.92 51.165 290.13 51.235 ;
    RECT 289.46 50.445 289.67 50.515 ;
    RECT 289.46 50.805 289.67 50.875 ;
    RECT 289.46 51.165 289.67 51.235 ;
    RECT 286.6 50.445 286.81 50.515 ;
    RECT 286.6 50.805 286.81 50.875 ;
    RECT 286.6 51.165 286.81 51.235 ;
    RECT 286.14 50.445 286.35 50.515 ;
    RECT 286.14 50.805 286.35 50.875 ;
    RECT 286.14 51.165 286.35 51.235 ;
    RECT 283.28 50.445 283.49 50.515 ;
    RECT 283.28 50.805 283.49 50.875 ;
    RECT 283.28 51.165 283.49 51.235 ;
    RECT 282.82 50.445 283.03 50.515 ;
    RECT 282.82 50.805 283.03 50.875 ;
    RECT 282.82 51.165 283.03 51.235 ;
    RECT 279.96 50.445 280.17 50.515 ;
    RECT 279.96 50.805 280.17 50.875 ;
    RECT 279.96 51.165 280.17 51.235 ;
    RECT 279.5 50.445 279.71 50.515 ;
    RECT 279.5 50.805 279.71 50.875 ;
    RECT 279.5 51.165 279.71 51.235 ;
    RECT 276.64 50.445 276.85 50.515 ;
    RECT 276.64 50.805 276.85 50.875 ;
    RECT 276.64 51.165 276.85 51.235 ;
    RECT 276.18 50.445 276.39 50.515 ;
    RECT 276.18 50.805 276.39 50.875 ;
    RECT 276.18 51.165 276.39 51.235 ;
    RECT 273.32 50.445 273.53 50.515 ;
    RECT 273.32 50.805 273.53 50.875 ;
    RECT 273.32 51.165 273.53 51.235 ;
    RECT 272.86 50.445 273.07 50.515 ;
    RECT 272.86 50.805 273.07 50.875 ;
    RECT 272.86 51.165 273.07 51.235 ;
    RECT 270.0 50.445 270.21 50.515 ;
    RECT 270.0 50.805 270.21 50.875 ;
    RECT 270.0 51.165 270.21 51.235 ;
    RECT 269.54 50.445 269.75 50.515 ;
    RECT 269.54 50.805 269.75 50.875 ;
    RECT 269.54 51.165 269.75 51.235 ;
    RECT 233.48 50.445 233.69 50.515 ;
    RECT 233.48 50.805 233.69 50.875 ;
    RECT 233.48 51.165 233.69 51.235 ;
    RECT 233.02 50.445 233.23 50.515 ;
    RECT 233.02 50.805 233.23 50.875 ;
    RECT 233.02 51.165 233.23 51.235 ;
    RECT 230.16 50.445 230.37 50.515 ;
    RECT 230.16 50.805 230.37 50.875 ;
    RECT 230.16 51.165 230.37 51.235 ;
    RECT 229.7 50.445 229.91 50.515 ;
    RECT 229.7 50.805 229.91 50.875 ;
    RECT 229.7 51.165 229.91 51.235 ;
    RECT 366.28 50.445 366.49 50.515 ;
    RECT 366.28 50.805 366.49 50.875 ;
    RECT 366.28 51.165 366.49 51.235 ;
    RECT 365.82 50.445 366.03 50.515 ;
    RECT 365.82 50.805 366.03 50.875 ;
    RECT 365.82 51.165 366.03 51.235 ;
    RECT 226.84 50.445 227.05 50.515 ;
    RECT 226.84 50.805 227.05 50.875 ;
    RECT 226.84 51.165 227.05 51.235 ;
    RECT 226.38 50.445 226.59 50.515 ;
    RECT 226.38 50.805 226.59 50.875 ;
    RECT 226.38 51.165 226.59 51.235 ;
    RECT 362.96 50.445 363.17 50.515 ;
    RECT 362.96 50.805 363.17 50.875 ;
    RECT 362.96 51.165 363.17 51.235 ;
    RECT 362.5 50.445 362.71 50.515 ;
    RECT 362.5 50.805 362.71 50.875 ;
    RECT 362.5 51.165 362.71 51.235 ;
    RECT 223.52 50.445 223.73 50.515 ;
    RECT 223.52 50.805 223.73 50.875 ;
    RECT 223.52 51.165 223.73 51.235 ;
    RECT 223.06 50.445 223.27 50.515 ;
    RECT 223.06 50.805 223.27 50.875 ;
    RECT 223.06 51.165 223.27 51.235 ;
    RECT 359.64 50.445 359.85 50.515 ;
    RECT 359.64 50.805 359.85 50.875 ;
    RECT 359.64 51.165 359.85 51.235 ;
    RECT 359.18 50.445 359.39 50.515 ;
    RECT 359.18 50.805 359.39 50.875 ;
    RECT 359.18 51.165 359.39 51.235 ;
    RECT 220.2 50.445 220.41 50.515 ;
    RECT 220.2 50.805 220.41 50.875 ;
    RECT 220.2 51.165 220.41 51.235 ;
    RECT 219.74 50.445 219.95 50.515 ;
    RECT 219.74 50.805 219.95 50.875 ;
    RECT 219.74 51.165 219.95 51.235 ;
    RECT 356.32 50.445 356.53 50.515 ;
    RECT 356.32 50.805 356.53 50.875 ;
    RECT 356.32 51.165 356.53 51.235 ;
    RECT 355.86 50.445 356.07 50.515 ;
    RECT 355.86 50.805 356.07 50.875 ;
    RECT 355.86 51.165 356.07 51.235 ;
    RECT 353.0 50.445 353.21 50.515 ;
    RECT 353.0 50.805 353.21 50.875 ;
    RECT 353.0 51.165 353.21 51.235 ;
    RECT 352.54 50.445 352.75 50.515 ;
    RECT 352.54 50.805 352.75 50.875 ;
    RECT 352.54 51.165 352.75 51.235 ;
    RECT 216.88 50.445 217.09 50.515 ;
    RECT 216.88 50.805 217.09 50.875 ;
    RECT 216.88 51.165 217.09 51.235 ;
    RECT 216.42 50.445 216.63 50.515 ;
    RECT 216.42 50.805 216.63 50.875 ;
    RECT 216.42 51.165 216.63 51.235 ;
    RECT 349.68 50.445 349.89 50.515 ;
    RECT 349.68 50.805 349.89 50.875 ;
    RECT 349.68 51.165 349.89 51.235 ;
    RECT 349.22 50.445 349.43 50.515 ;
    RECT 349.22 50.805 349.43 50.875 ;
    RECT 349.22 51.165 349.43 51.235 ;
    RECT 213.56 50.445 213.77 50.515 ;
    RECT 213.56 50.805 213.77 50.875 ;
    RECT 213.56 51.165 213.77 51.235 ;
    RECT 213.1 50.445 213.31 50.515 ;
    RECT 213.1 50.805 213.31 50.875 ;
    RECT 213.1 51.165 213.31 51.235 ;
    RECT 346.36 50.445 346.57 50.515 ;
    RECT 346.36 50.805 346.57 50.875 ;
    RECT 346.36 51.165 346.57 51.235 ;
    RECT 345.9 50.445 346.11 50.515 ;
    RECT 345.9 50.805 346.11 50.875 ;
    RECT 345.9 51.165 346.11 51.235 ;
    RECT 210.24 50.445 210.45 50.515 ;
    RECT 210.24 50.805 210.45 50.875 ;
    RECT 210.24 51.165 210.45 51.235 ;
    RECT 209.78 50.445 209.99 50.515 ;
    RECT 209.78 50.805 209.99 50.875 ;
    RECT 209.78 51.165 209.99 51.235 ;
    RECT 343.04 50.445 343.25 50.515 ;
    RECT 343.04 50.805 343.25 50.875 ;
    RECT 343.04 51.165 343.25 51.235 ;
    RECT 342.58 50.445 342.79 50.515 ;
    RECT 342.58 50.805 342.79 50.875 ;
    RECT 342.58 51.165 342.79 51.235 ;
    RECT 206.92 50.445 207.13 50.515 ;
    RECT 206.92 50.805 207.13 50.875 ;
    RECT 206.92 51.165 207.13 51.235 ;
    RECT 206.46 50.445 206.67 50.515 ;
    RECT 206.46 50.805 206.67 50.875 ;
    RECT 206.46 51.165 206.67 51.235 ;
    RECT 339.72 50.445 339.93 50.515 ;
    RECT 339.72 50.805 339.93 50.875 ;
    RECT 339.72 51.165 339.93 51.235 ;
    RECT 339.26 50.445 339.47 50.515 ;
    RECT 339.26 50.805 339.47 50.875 ;
    RECT 339.26 51.165 339.47 51.235 ;
    RECT 203.6 50.445 203.81 50.515 ;
    RECT 203.6 50.805 203.81 50.875 ;
    RECT 203.6 51.165 203.81 51.235 ;
    RECT 203.14 50.445 203.35 50.515 ;
    RECT 203.14 50.805 203.35 50.875 ;
    RECT 203.14 51.165 203.35 51.235 ;
    RECT 336.4 50.445 336.61 50.515 ;
    RECT 336.4 50.805 336.61 50.875 ;
    RECT 336.4 51.165 336.61 51.235 ;
    RECT 335.94 50.445 336.15 50.515 ;
    RECT 335.94 50.805 336.15 50.875 ;
    RECT 335.94 51.165 336.15 51.235 ;
    RECT 266.68 50.445 266.89 50.515 ;
    RECT 266.68 50.805 266.89 50.875 ;
    RECT 266.68 51.165 266.89 51.235 ;
    RECT 266.22 50.445 266.43 50.515 ;
    RECT 266.22 50.805 266.43 50.875 ;
    RECT 266.22 51.165 266.43 51.235 ;
    RECT 263.36 50.445 263.57 50.515 ;
    RECT 263.36 50.805 263.57 50.875 ;
    RECT 263.36 51.165 263.57 51.235 ;
    RECT 262.9 50.445 263.11 50.515 ;
    RECT 262.9 50.805 263.11 50.875 ;
    RECT 262.9 51.165 263.11 51.235 ;
    RECT 260.04 50.445 260.25 50.515 ;
    RECT 260.04 50.805 260.25 50.875 ;
    RECT 260.04 51.165 260.25 51.235 ;
    RECT 259.58 50.445 259.79 50.515 ;
    RECT 259.58 50.805 259.79 50.875 ;
    RECT 259.58 51.165 259.79 51.235 ;
    RECT 256.72 50.445 256.93 50.515 ;
    RECT 256.72 50.805 256.93 50.875 ;
    RECT 256.72 51.165 256.93 51.235 ;
    RECT 256.26 50.445 256.47 50.515 ;
    RECT 256.26 50.805 256.47 50.875 ;
    RECT 256.26 51.165 256.47 51.235 ;
    RECT 253.4 50.445 253.61 50.515 ;
    RECT 253.4 50.805 253.61 50.875 ;
    RECT 253.4 51.165 253.61 51.235 ;
    RECT 252.94 50.445 253.15 50.515 ;
    RECT 252.94 50.805 253.15 50.875 ;
    RECT 252.94 51.165 253.15 51.235 ;
    RECT 250.08 50.445 250.29 50.515 ;
    RECT 250.08 50.805 250.29 50.875 ;
    RECT 250.08 51.165 250.29 51.235 ;
    RECT 249.62 50.445 249.83 50.515 ;
    RECT 249.62 50.805 249.83 50.875 ;
    RECT 249.62 51.165 249.83 51.235 ;
    RECT 246.76 50.445 246.97 50.515 ;
    RECT 246.76 50.805 246.97 50.875 ;
    RECT 246.76 51.165 246.97 51.235 ;
    RECT 246.3 50.445 246.51 50.515 ;
    RECT 246.3 50.805 246.51 50.875 ;
    RECT 246.3 51.165 246.51 51.235 ;
    RECT 243.44 50.445 243.65 50.515 ;
    RECT 243.44 50.805 243.65 50.875 ;
    RECT 243.44 51.165 243.65 51.235 ;
    RECT 242.98 50.445 243.19 50.515 ;
    RECT 242.98 50.805 243.19 50.875 ;
    RECT 242.98 51.165 243.19 51.235 ;
    RECT 240.12 50.445 240.33 50.515 ;
    RECT 240.12 50.805 240.33 50.875 ;
    RECT 240.12 51.165 240.33 51.235 ;
    RECT 239.66 50.445 239.87 50.515 ;
    RECT 239.66 50.805 239.87 50.875 ;
    RECT 239.66 51.165 239.87 51.235 ;
    RECT 236.8 50.445 237.01 50.515 ;
    RECT 236.8 50.805 237.01 50.875 ;
    RECT 236.8 51.165 237.01 51.235 ;
    RECT 236.34 50.445 236.55 50.515 ;
    RECT 236.34 50.805 236.55 50.875 ;
    RECT 236.34 51.165 236.55 51.235 ;
    RECT 374.15 50.805 374.22 50.875 ;
    RECT 333.08 50.445 333.29 50.515 ;
    RECT 333.08 50.805 333.29 50.875 ;
    RECT 333.08 51.165 333.29 51.235 ;
    RECT 332.62 50.445 332.83 50.515 ;
    RECT 332.62 50.805 332.83 50.875 ;
    RECT 332.62 51.165 332.83 51.235 ;
    RECT 329.76 50.445 329.97 50.515 ;
    RECT 329.76 50.805 329.97 50.875 ;
    RECT 329.76 51.165 329.97 51.235 ;
    RECT 329.3 50.445 329.51 50.515 ;
    RECT 329.3 50.805 329.51 50.875 ;
    RECT 329.3 51.165 329.51 51.235 ;
    RECT 326.44 50.445 326.65 50.515 ;
    RECT 326.44 50.805 326.65 50.875 ;
    RECT 326.44 51.165 326.65 51.235 ;
    RECT 325.98 50.445 326.19 50.515 ;
    RECT 325.98 50.805 326.19 50.875 ;
    RECT 325.98 51.165 326.19 51.235 ;
    RECT 323.12 50.445 323.33 50.515 ;
    RECT 323.12 50.805 323.33 50.875 ;
    RECT 323.12 51.165 323.33 51.235 ;
    RECT 322.66 50.445 322.87 50.515 ;
    RECT 322.66 50.805 322.87 50.875 ;
    RECT 322.66 51.165 322.87 51.235 ;
    RECT 319.8 50.445 320.01 50.515 ;
    RECT 319.8 50.805 320.01 50.875 ;
    RECT 319.8 51.165 320.01 51.235 ;
    RECT 319.34 50.445 319.55 50.515 ;
    RECT 319.34 50.805 319.55 50.875 ;
    RECT 319.34 51.165 319.55 51.235 ;
    RECT 316.48 50.445 316.69 50.515 ;
    RECT 316.48 50.805 316.69 50.875 ;
    RECT 316.48 51.165 316.69 51.235 ;
    RECT 316.02 50.445 316.23 50.515 ;
    RECT 316.02 50.805 316.23 50.875 ;
    RECT 316.02 51.165 316.23 51.235 ;
    RECT 313.16 50.445 313.37 50.515 ;
    RECT 313.16 50.805 313.37 50.875 ;
    RECT 313.16 51.165 313.37 51.235 ;
    RECT 312.7 50.445 312.91 50.515 ;
    RECT 312.7 50.805 312.91 50.875 ;
    RECT 312.7 51.165 312.91 51.235 ;
    RECT 309.84 50.445 310.05 50.515 ;
    RECT 309.84 50.805 310.05 50.875 ;
    RECT 309.84 51.165 310.05 51.235 ;
    RECT 309.38 50.445 309.59 50.515 ;
    RECT 309.38 50.805 309.59 50.875 ;
    RECT 309.38 51.165 309.59 51.235 ;
    RECT 306.52 50.445 306.73 50.515 ;
    RECT 306.52 50.805 306.73 50.875 ;
    RECT 306.52 51.165 306.73 51.235 ;
    RECT 306.06 50.445 306.27 50.515 ;
    RECT 306.06 50.805 306.27 50.875 ;
    RECT 306.06 51.165 306.27 51.235 ;
    RECT 303.2 11.565 303.41 11.635 ;
    RECT 303.2 11.925 303.41 11.995 ;
    RECT 303.2 12.285 303.41 12.355 ;
    RECT 302.74 11.565 302.95 11.635 ;
    RECT 302.74 11.925 302.95 11.995 ;
    RECT 302.74 12.285 302.95 12.355 ;
    RECT 369.6 11.565 369.81 11.635 ;
    RECT 369.6 11.925 369.81 11.995 ;
    RECT 369.6 12.285 369.81 12.355 ;
    RECT 369.14 11.565 369.35 11.635 ;
    RECT 369.14 11.925 369.35 11.995 ;
    RECT 369.14 12.285 369.35 12.355 ;
    RECT 299.88 11.565 300.09 11.635 ;
    RECT 299.88 11.925 300.09 11.995 ;
    RECT 299.88 12.285 300.09 12.355 ;
    RECT 299.42 11.565 299.63 11.635 ;
    RECT 299.42 11.925 299.63 11.995 ;
    RECT 299.42 12.285 299.63 12.355 ;
    RECT 296.56 11.565 296.77 11.635 ;
    RECT 296.56 11.925 296.77 11.995 ;
    RECT 296.56 12.285 296.77 12.355 ;
    RECT 296.1 11.565 296.31 11.635 ;
    RECT 296.1 11.925 296.31 11.995 ;
    RECT 296.1 12.285 296.31 12.355 ;
    RECT 293.24 11.565 293.45 11.635 ;
    RECT 293.24 11.925 293.45 11.995 ;
    RECT 293.24 12.285 293.45 12.355 ;
    RECT 292.78 11.565 292.99 11.635 ;
    RECT 292.78 11.925 292.99 11.995 ;
    RECT 292.78 12.285 292.99 12.355 ;
    RECT 289.92 11.565 290.13 11.635 ;
    RECT 289.92 11.925 290.13 11.995 ;
    RECT 289.92 12.285 290.13 12.355 ;
    RECT 289.46 11.565 289.67 11.635 ;
    RECT 289.46 11.925 289.67 11.995 ;
    RECT 289.46 12.285 289.67 12.355 ;
    RECT 286.6 11.565 286.81 11.635 ;
    RECT 286.6 11.925 286.81 11.995 ;
    RECT 286.6 12.285 286.81 12.355 ;
    RECT 286.14 11.565 286.35 11.635 ;
    RECT 286.14 11.925 286.35 11.995 ;
    RECT 286.14 12.285 286.35 12.355 ;
    RECT 283.28 11.565 283.49 11.635 ;
    RECT 283.28 11.925 283.49 11.995 ;
    RECT 283.28 12.285 283.49 12.355 ;
    RECT 282.82 11.565 283.03 11.635 ;
    RECT 282.82 11.925 283.03 11.995 ;
    RECT 282.82 12.285 283.03 12.355 ;
    RECT 279.96 11.565 280.17 11.635 ;
    RECT 279.96 11.925 280.17 11.995 ;
    RECT 279.96 12.285 280.17 12.355 ;
    RECT 279.5 11.565 279.71 11.635 ;
    RECT 279.5 11.925 279.71 11.995 ;
    RECT 279.5 12.285 279.71 12.355 ;
    RECT 276.64 11.565 276.85 11.635 ;
    RECT 276.64 11.925 276.85 11.995 ;
    RECT 276.64 12.285 276.85 12.355 ;
    RECT 276.18 11.565 276.39 11.635 ;
    RECT 276.18 11.925 276.39 11.995 ;
    RECT 276.18 12.285 276.39 12.355 ;
    RECT 273.32 11.565 273.53 11.635 ;
    RECT 273.32 11.925 273.53 11.995 ;
    RECT 273.32 12.285 273.53 12.355 ;
    RECT 272.86 11.565 273.07 11.635 ;
    RECT 272.86 11.925 273.07 11.995 ;
    RECT 272.86 12.285 273.07 12.355 ;
    RECT 270.0 11.565 270.21 11.635 ;
    RECT 270.0 11.925 270.21 11.995 ;
    RECT 270.0 12.285 270.21 12.355 ;
    RECT 269.54 11.565 269.75 11.635 ;
    RECT 269.54 11.925 269.75 11.995 ;
    RECT 269.54 12.285 269.75 12.355 ;
    RECT 233.48 11.565 233.69 11.635 ;
    RECT 233.48 11.925 233.69 11.995 ;
    RECT 233.48 12.285 233.69 12.355 ;
    RECT 233.02 11.565 233.23 11.635 ;
    RECT 233.02 11.925 233.23 11.995 ;
    RECT 233.02 12.285 233.23 12.355 ;
    RECT 230.16 11.565 230.37 11.635 ;
    RECT 230.16 11.925 230.37 11.995 ;
    RECT 230.16 12.285 230.37 12.355 ;
    RECT 229.7 11.565 229.91 11.635 ;
    RECT 229.7 11.925 229.91 11.995 ;
    RECT 229.7 12.285 229.91 12.355 ;
    RECT 366.28 11.565 366.49 11.635 ;
    RECT 366.28 11.925 366.49 11.995 ;
    RECT 366.28 12.285 366.49 12.355 ;
    RECT 365.82 11.565 366.03 11.635 ;
    RECT 365.82 11.925 366.03 11.995 ;
    RECT 365.82 12.285 366.03 12.355 ;
    RECT 226.84 11.565 227.05 11.635 ;
    RECT 226.84 11.925 227.05 11.995 ;
    RECT 226.84 12.285 227.05 12.355 ;
    RECT 226.38 11.565 226.59 11.635 ;
    RECT 226.38 11.925 226.59 11.995 ;
    RECT 226.38 12.285 226.59 12.355 ;
    RECT 362.96 11.565 363.17 11.635 ;
    RECT 362.96 11.925 363.17 11.995 ;
    RECT 362.96 12.285 363.17 12.355 ;
    RECT 362.5 11.565 362.71 11.635 ;
    RECT 362.5 11.925 362.71 11.995 ;
    RECT 362.5 12.285 362.71 12.355 ;
    RECT 223.52 11.565 223.73 11.635 ;
    RECT 223.52 11.925 223.73 11.995 ;
    RECT 223.52 12.285 223.73 12.355 ;
    RECT 223.06 11.565 223.27 11.635 ;
    RECT 223.06 11.925 223.27 11.995 ;
    RECT 223.06 12.285 223.27 12.355 ;
    RECT 359.64 11.565 359.85 11.635 ;
    RECT 359.64 11.925 359.85 11.995 ;
    RECT 359.64 12.285 359.85 12.355 ;
    RECT 359.18 11.565 359.39 11.635 ;
    RECT 359.18 11.925 359.39 11.995 ;
    RECT 359.18 12.285 359.39 12.355 ;
    RECT 200.605 11.925 200.675 11.995 ;
    RECT 220.2 11.565 220.41 11.635 ;
    RECT 220.2 11.925 220.41 11.995 ;
    RECT 220.2 12.285 220.41 12.355 ;
    RECT 219.74 11.565 219.95 11.635 ;
    RECT 219.74 11.925 219.95 11.995 ;
    RECT 219.74 12.285 219.95 12.355 ;
    RECT 356.32 11.565 356.53 11.635 ;
    RECT 356.32 11.925 356.53 11.995 ;
    RECT 356.32 12.285 356.53 12.355 ;
    RECT 355.86 11.565 356.07 11.635 ;
    RECT 355.86 11.925 356.07 11.995 ;
    RECT 355.86 12.285 356.07 12.355 ;
    RECT 353.0 11.565 353.21 11.635 ;
    RECT 353.0 11.925 353.21 11.995 ;
    RECT 353.0 12.285 353.21 12.355 ;
    RECT 352.54 11.565 352.75 11.635 ;
    RECT 352.54 11.925 352.75 11.995 ;
    RECT 352.54 12.285 352.75 12.355 ;
    RECT 216.88 11.565 217.09 11.635 ;
    RECT 216.88 11.925 217.09 11.995 ;
    RECT 216.88 12.285 217.09 12.355 ;
    RECT 216.42 11.565 216.63 11.635 ;
    RECT 216.42 11.925 216.63 11.995 ;
    RECT 216.42 12.285 216.63 12.355 ;
    RECT 349.68 11.565 349.89 11.635 ;
    RECT 349.68 11.925 349.89 11.995 ;
    RECT 349.68 12.285 349.89 12.355 ;
    RECT 349.22 11.565 349.43 11.635 ;
    RECT 349.22 11.925 349.43 11.995 ;
    RECT 349.22 12.285 349.43 12.355 ;
    RECT 213.56 11.565 213.77 11.635 ;
    RECT 213.56 11.925 213.77 11.995 ;
    RECT 213.56 12.285 213.77 12.355 ;
    RECT 213.1 11.565 213.31 11.635 ;
    RECT 213.1 11.925 213.31 11.995 ;
    RECT 213.1 12.285 213.31 12.355 ;
    RECT 346.36 11.565 346.57 11.635 ;
    RECT 346.36 11.925 346.57 11.995 ;
    RECT 346.36 12.285 346.57 12.355 ;
    RECT 345.9 11.565 346.11 11.635 ;
    RECT 345.9 11.925 346.11 11.995 ;
    RECT 345.9 12.285 346.11 12.355 ;
    RECT 210.24 11.565 210.45 11.635 ;
    RECT 210.24 11.925 210.45 11.995 ;
    RECT 210.24 12.285 210.45 12.355 ;
    RECT 209.78 11.565 209.99 11.635 ;
    RECT 209.78 11.925 209.99 11.995 ;
    RECT 209.78 12.285 209.99 12.355 ;
    RECT 343.04 11.565 343.25 11.635 ;
    RECT 343.04 11.925 343.25 11.995 ;
    RECT 343.04 12.285 343.25 12.355 ;
    RECT 342.58 11.565 342.79 11.635 ;
    RECT 342.58 11.925 342.79 11.995 ;
    RECT 342.58 12.285 342.79 12.355 ;
    RECT 206.92 11.565 207.13 11.635 ;
    RECT 206.92 11.925 207.13 11.995 ;
    RECT 206.92 12.285 207.13 12.355 ;
    RECT 206.46 11.565 206.67 11.635 ;
    RECT 206.46 11.925 206.67 11.995 ;
    RECT 206.46 12.285 206.67 12.355 ;
    RECT 339.72 11.565 339.93 11.635 ;
    RECT 339.72 11.925 339.93 11.995 ;
    RECT 339.72 12.285 339.93 12.355 ;
    RECT 339.26 11.565 339.47 11.635 ;
    RECT 339.26 11.925 339.47 11.995 ;
    RECT 339.26 12.285 339.47 12.355 ;
    RECT 336.4 11.565 336.61 11.635 ;
    RECT 336.4 11.925 336.61 11.995 ;
    RECT 336.4 12.285 336.61 12.355 ;
    RECT 335.94 11.565 336.15 11.635 ;
    RECT 335.94 11.925 336.15 11.995 ;
    RECT 335.94 12.285 336.15 12.355 ;
    RECT 266.68 11.565 266.89 11.635 ;
    RECT 266.68 11.925 266.89 11.995 ;
    RECT 266.68 12.285 266.89 12.355 ;
    RECT 266.22 11.565 266.43 11.635 ;
    RECT 266.22 11.925 266.43 11.995 ;
    RECT 266.22 12.285 266.43 12.355 ;
    RECT 263.36 11.565 263.57 11.635 ;
    RECT 263.36 11.925 263.57 11.995 ;
    RECT 263.36 12.285 263.57 12.355 ;
    RECT 262.9 11.565 263.11 11.635 ;
    RECT 262.9 11.925 263.11 11.995 ;
    RECT 262.9 12.285 263.11 12.355 ;
    RECT 372.92 11.565 373.13 11.635 ;
    RECT 372.92 11.925 373.13 11.995 ;
    RECT 372.92 12.285 373.13 12.355 ;
    RECT 372.46 11.565 372.67 11.635 ;
    RECT 372.46 11.925 372.67 11.995 ;
    RECT 372.46 12.285 372.67 12.355 ;
    RECT 260.04 11.565 260.25 11.635 ;
    RECT 260.04 11.925 260.25 11.995 ;
    RECT 260.04 12.285 260.25 12.355 ;
    RECT 259.58 11.565 259.79 11.635 ;
    RECT 259.58 11.925 259.79 11.995 ;
    RECT 259.58 12.285 259.79 12.355 ;
    RECT 256.72 11.565 256.93 11.635 ;
    RECT 256.72 11.925 256.93 11.995 ;
    RECT 256.72 12.285 256.93 12.355 ;
    RECT 256.26 11.565 256.47 11.635 ;
    RECT 256.26 11.925 256.47 11.995 ;
    RECT 256.26 12.285 256.47 12.355 ;
    RECT 253.4 11.565 253.61 11.635 ;
    RECT 253.4 11.925 253.61 11.995 ;
    RECT 253.4 12.285 253.61 12.355 ;
    RECT 252.94 11.565 253.15 11.635 ;
    RECT 252.94 11.925 253.15 11.995 ;
    RECT 252.94 12.285 253.15 12.355 ;
    RECT 250.08 11.565 250.29 11.635 ;
    RECT 250.08 11.925 250.29 11.995 ;
    RECT 250.08 12.285 250.29 12.355 ;
    RECT 249.62 11.565 249.83 11.635 ;
    RECT 249.62 11.925 249.83 11.995 ;
    RECT 249.62 12.285 249.83 12.355 ;
    RECT 246.76 11.565 246.97 11.635 ;
    RECT 246.76 11.925 246.97 11.995 ;
    RECT 246.76 12.285 246.97 12.355 ;
    RECT 246.3 11.565 246.51 11.635 ;
    RECT 246.3 11.925 246.51 11.995 ;
    RECT 246.3 12.285 246.51 12.355 ;
    RECT 243.44 11.565 243.65 11.635 ;
    RECT 243.44 11.925 243.65 11.995 ;
    RECT 243.44 12.285 243.65 12.355 ;
    RECT 242.98 11.565 243.19 11.635 ;
    RECT 242.98 11.925 243.19 11.995 ;
    RECT 242.98 12.285 243.19 12.355 ;
    RECT 203.6 11.565 203.81 11.635 ;
    RECT 203.6 11.925 203.81 11.995 ;
    RECT 203.6 12.285 203.81 12.355 ;
    RECT 203.14 11.565 203.35 11.635 ;
    RECT 203.14 11.925 203.35 11.995 ;
    RECT 203.14 12.285 203.35 12.355 ;
    RECT 240.12 11.565 240.33 11.635 ;
    RECT 240.12 11.925 240.33 11.995 ;
    RECT 240.12 12.285 240.33 12.355 ;
    RECT 239.66 11.565 239.87 11.635 ;
    RECT 239.66 11.925 239.87 11.995 ;
    RECT 239.66 12.285 239.87 12.355 ;
    RECT 236.8 11.565 237.01 11.635 ;
    RECT 236.8 11.925 237.01 11.995 ;
    RECT 236.8 12.285 237.01 12.355 ;
    RECT 236.34 11.565 236.55 11.635 ;
    RECT 236.34 11.925 236.55 11.995 ;
    RECT 236.34 12.285 236.55 12.355 ;
    RECT 333.08 11.565 333.29 11.635 ;
    RECT 333.08 11.925 333.29 11.995 ;
    RECT 333.08 12.285 333.29 12.355 ;
    RECT 332.62 11.565 332.83 11.635 ;
    RECT 332.62 11.925 332.83 11.995 ;
    RECT 332.62 12.285 332.83 12.355 ;
    RECT 329.76 11.565 329.97 11.635 ;
    RECT 329.76 11.925 329.97 11.995 ;
    RECT 329.76 12.285 329.97 12.355 ;
    RECT 329.3 11.565 329.51 11.635 ;
    RECT 329.3 11.925 329.51 11.995 ;
    RECT 329.3 12.285 329.51 12.355 ;
    RECT 326.44 11.565 326.65 11.635 ;
    RECT 326.44 11.925 326.65 11.995 ;
    RECT 326.44 12.285 326.65 12.355 ;
    RECT 325.98 11.565 326.19 11.635 ;
    RECT 325.98 11.925 326.19 11.995 ;
    RECT 325.98 12.285 326.19 12.355 ;
    RECT 374.15 11.925 374.22 11.995 ;
    RECT 323.12 11.565 323.33 11.635 ;
    RECT 323.12 11.925 323.33 11.995 ;
    RECT 323.12 12.285 323.33 12.355 ;
    RECT 322.66 11.565 322.87 11.635 ;
    RECT 322.66 11.925 322.87 11.995 ;
    RECT 322.66 12.285 322.87 12.355 ;
    RECT 319.8 11.565 320.01 11.635 ;
    RECT 319.8 11.925 320.01 11.995 ;
    RECT 319.8 12.285 320.01 12.355 ;
    RECT 319.34 11.565 319.55 11.635 ;
    RECT 319.34 11.925 319.55 11.995 ;
    RECT 319.34 12.285 319.55 12.355 ;
    RECT 316.48 11.565 316.69 11.635 ;
    RECT 316.48 11.925 316.69 11.995 ;
    RECT 316.48 12.285 316.69 12.355 ;
    RECT 316.02 11.565 316.23 11.635 ;
    RECT 316.02 11.925 316.23 11.995 ;
    RECT 316.02 12.285 316.23 12.355 ;
    RECT 313.16 11.565 313.37 11.635 ;
    RECT 313.16 11.925 313.37 11.995 ;
    RECT 313.16 12.285 313.37 12.355 ;
    RECT 312.7 11.565 312.91 11.635 ;
    RECT 312.7 11.925 312.91 11.995 ;
    RECT 312.7 12.285 312.91 12.355 ;
    RECT 309.84 11.565 310.05 11.635 ;
    RECT 309.84 11.925 310.05 11.995 ;
    RECT 309.84 12.285 310.05 12.355 ;
    RECT 309.38 11.565 309.59 11.635 ;
    RECT 309.38 11.925 309.59 11.995 ;
    RECT 309.38 12.285 309.59 12.355 ;
    RECT 306.52 11.565 306.73 11.635 ;
    RECT 306.52 11.925 306.73 11.995 ;
    RECT 306.52 12.285 306.73 12.355 ;
    RECT 306.06 11.565 306.27 11.635 ;
    RECT 306.06 11.925 306.27 11.995 ;
    RECT 306.06 12.285 306.27 12.355 ;
    RECT 303.2 49.725 303.41 49.795 ;
    RECT 303.2 50.085 303.41 50.155 ;
    RECT 303.2 50.445 303.41 50.515 ;
    RECT 302.74 49.725 302.95 49.795 ;
    RECT 302.74 50.085 302.95 50.155 ;
    RECT 302.74 50.445 302.95 50.515 ;
    RECT 372.92 49.725 373.13 49.795 ;
    RECT 372.92 50.085 373.13 50.155 ;
    RECT 372.92 50.445 373.13 50.515 ;
    RECT 372.46 49.725 372.67 49.795 ;
    RECT 372.46 50.085 372.67 50.155 ;
    RECT 372.46 50.445 372.67 50.515 ;
    RECT 369.6 49.725 369.81 49.795 ;
    RECT 369.6 50.085 369.81 50.155 ;
    RECT 369.6 50.445 369.81 50.515 ;
    RECT 369.14 49.725 369.35 49.795 ;
    RECT 369.14 50.085 369.35 50.155 ;
    RECT 369.14 50.445 369.35 50.515 ;
    RECT 200.605 50.085 200.675 50.155 ;
    RECT 299.88 49.725 300.09 49.795 ;
    RECT 299.88 50.085 300.09 50.155 ;
    RECT 299.88 50.445 300.09 50.515 ;
    RECT 299.42 49.725 299.63 49.795 ;
    RECT 299.42 50.085 299.63 50.155 ;
    RECT 299.42 50.445 299.63 50.515 ;
    RECT 296.56 49.725 296.77 49.795 ;
    RECT 296.56 50.085 296.77 50.155 ;
    RECT 296.56 50.445 296.77 50.515 ;
    RECT 296.1 49.725 296.31 49.795 ;
    RECT 296.1 50.085 296.31 50.155 ;
    RECT 296.1 50.445 296.31 50.515 ;
    RECT 293.24 49.725 293.45 49.795 ;
    RECT 293.24 50.085 293.45 50.155 ;
    RECT 293.24 50.445 293.45 50.515 ;
    RECT 292.78 49.725 292.99 49.795 ;
    RECT 292.78 50.085 292.99 50.155 ;
    RECT 292.78 50.445 292.99 50.515 ;
    RECT 289.92 49.725 290.13 49.795 ;
    RECT 289.92 50.085 290.13 50.155 ;
    RECT 289.92 50.445 290.13 50.515 ;
    RECT 289.46 49.725 289.67 49.795 ;
    RECT 289.46 50.085 289.67 50.155 ;
    RECT 289.46 50.445 289.67 50.515 ;
    RECT 286.6 49.725 286.81 49.795 ;
    RECT 286.6 50.085 286.81 50.155 ;
    RECT 286.6 50.445 286.81 50.515 ;
    RECT 286.14 49.725 286.35 49.795 ;
    RECT 286.14 50.085 286.35 50.155 ;
    RECT 286.14 50.445 286.35 50.515 ;
    RECT 283.28 49.725 283.49 49.795 ;
    RECT 283.28 50.085 283.49 50.155 ;
    RECT 283.28 50.445 283.49 50.515 ;
    RECT 282.82 49.725 283.03 49.795 ;
    RECT 282.82 50.085 283.03 50.155 ;
    RECT 282.82 50.445 283.03 50.515 ;
    RECT 279.96 49.725 280.17 49.795 ;
    RECT 279.96 50.085 280.17 50.155 ;
    RECT 279.96 50.445 280.17 50.515 ;
    RECT 279.5 49.725 279.71 49.795 ;
    RECT 279.5 50.085 279.71 50.155 ;
    RECT 279.5 50.445 279.71 50.515 ;
    RECT 276.64 49.725 276.85 49.795 ;
    RECT 276.64 50.085 276.85 50.155 ;
    RECT 276.64 50.445 276.85 50.515 ;
    RECT 276.18 49.725 276.39 49.795 ;
    RECT 276.18 50.085 276.39 50.155 ;
    RECT 276.18 50.445 276.39 50.515 ;
    RECT 273.32 49.725 273.53 49.795 ;
    RECT 273.32 50.085 273.53 50.155 ;
    RECT 273.32 50.445 273.53 50.515 ;
    RECT 272.86 49.725 273.07 49.795 ;
    RECT 272.86 50.085 273.07 50.155 ;
    RECT 272.86 50.445 273.07 50.515 ;
    RECT 270.0 49.725 270.21 49.795 ;
    RECT 270.0 50.085 270.21 50.155 ;
    RECT 270.0 50.445 270.21 50.515 ;
    RECT 269.54 49.725 269.75 49.795 ;
    RECT 269.54 50.085 269.75 50.155 ;
    RECT 269.54 50.445 269.75 50.515 ;
    RECT 233.48 49.725 233.69 49.795 ;
    RECT 233.48 50.085 233.69 50.155 ;
    RECT 233.48 50.445 233.69 50.515 ;
    RECT 233.02 49.725 233.23 49.795 ;
    RECT 233.02 50.085 233.23 50.155 ;
    RECT 233.02 50.445 233.23 50.515 ;
    RECT 230.16 49.725 230.37 49.795 ;
    RECT 230.16 50.085 230.37 50.155 ;
    RECT 230.16 50.445 230.37 50.515 ;
    RECT 229.7 49.725 229.91 49.795 ;
    RECT 229.7 50.085 229.91 50.155 ;
    RECT 229.7 50.445 229.91 50.515 ;
    RECT 366.28 49.725 366.49 49.795 ;
    RECT 366.28 50.085 366.49 50.155 ;
    RECT 366.28 50.445 366.49 50.515 ;
    RECT 365.82 49.725 366.03 49.795 ;
    RECT 365.82 50.085 366.03 50.155 ;
    RECT 365.82 50.445 366.03 50.515 ;
    RECT 226.84 49.725 227.05 49.795 ;
    RECT 226.84 50.085 227.05 50.155 ;
    RECT 226.84 50.445 227.05 50.515 ;
    RECT 226.38 49.725 226.59 49.795 ;
    RECT 226.38 50.085 226.59 50.155 ;
    RECT 226.38 50.445 226.59 50.515 ;
    RECT 362.96 49.725 363.17 49.795 ;
    RECT 362.96 50.085 363.17 50.155 ;
    RECT 362.96 50.445 363.17 50.515 ;
    RECT 362.5 49.725 362.71 49.795 ;
    RECT 362.5 50.085 362.71 50.155 ;
    RECT 362.5 50.445 362.71 50.515 ;
    RECT 223.52 49.725 223.73 49.795 ;
    RECT 223.52 50.085 223.73 50.155 ;
    RECT 223.52 50.445 223.73 50.515 ;
    RECT 223.06 49.725 223.27 49.795 ;
    RECT 223.06 50.085 223.27 50.155 ;
    RECT 223.06 50.445 223.27 50.515 ;
    RECT 359.64 49.725 359.85 49.795 ;
    RECT 359.64 50.085 359.85 50.155 ;
    RECT 359.64 50.445 359.85 50.515 ;
    RECT 359.18 49.725 359.39 49.795 ;
    RECT 359.18 50.085 359.39 50.155 ;
    RECT 359.18 50.445 359.39 50.515 ;
    RECT 220.2 49.725 220.41 49.795 ;
    RECT 220.2 50.085 220.41 50.155 ;
    RECT 220.2 50.445 220.41 50.515 ;
    RECT 219.74 49.725 219.95 49.795 ;
    RECT 219.74 50.085 219.95 50.155 ;
    RECT 219.74 50.445 219.95 50.515 ;
    RECT 356.32 49.725 356.53 49.795 ;
    RECT 356.32 50.085 356.53 50.155 ;
    RECT 356.32 50.445 356.53 50.515 ;
    RECT 355.86 49.725 356.07 49.795 ;
    RECT 355.86 50.085 356.07 50.155 ;
    RECT 355.86 50.445 356.07 50.515 ;
    RECT 353.0 49.725 353.21 49.795 ;
    RECT 353.0 50.085 353.21 50.155 ;
    RECT 353.0 50.445 353.21 50.515 ;
    RECT 352.54 49.725 352.75 49.795 ;
    RECT 352.54 50.085 352.75 50.155 ;
    RECT 352.54 50.445 352.75 50.515 ;
    RECT 216.88 49.725 217.09 49.795 ;
    RECT 216.88 50.085 217.09 50.155 ;
    RECT 216.88 50.445 217.09 50.515 ;
    RECT 216.42 49.725 216.63 49.795 ;
    RECT 216.42 50.085 216.63 50.155 ;
    RECT 216.42 50.445 216.63 50.515 ;
    RECT 349.68 49.725 349.89 49.795 ;
    RECT 349.68 50.085 349.89 50.155 ;
    RECT 349.68 50.445 349.89 50.515 ;
    RECT 349.22 49.725 349.43 49.795 ;
    RECT 349.22 50.085 349.43 50.155 ;
    RECT 349.22 50.445 349.43 50.515 ;
    RECT 213.56 49.725 213.77 49.795 ;
    RECT 213.56 50.085 213.77 50.155 ;
    RECT 213.56 50.445 213.77 50.515 ;
    RECT 213.1 49.725 213.31 49.795 ;
    RECT 213.1 50.085 213.31 50.155 ;
    RECT 213.1 50.445 213.31 50.515 ;
    RECT 346.36 49.725 346.57 49.795 ;
    RECT 346.36 50.085 346.57 50.155 ;
    RECT 346.36 50.445 346.57 50.515 ;
    RECT 345.9 49.725 346.11 49.795 ;
    RECT 345.9 50.085 346.11 50.155 ;
    RECT 345.9 50.445 346.11 50.515 ;
    RECT 210.24 49.725 210.45 49.795 ;
    RECT 210.24 50.085 210.45 50.155 ;
    RECT 210.24 50.445 210.45 50.515 ;
    RECT 209.78 49.725 209.99 49.795 ;
    RECT 209.78 50.085 209.99 50.155 ;
    RECT 209.78 50.445 209.99 50.515 ;
    RECT 343.04 49.725 343.25 49.795 ;
    RECT 343.04 50.085 343.25 50.155 ;
    RECT 343.04 50.445 343.25 50.515 ;
    RECT 342.58 49.725 342.79 49.795 ;
    RECT 342.58 50.085 342.79 50.155 ;
    RECT 342.58 50.445 342.79 50.515 ;
    RECT 206.92 49.725 207.13 49.795 ;
    RECT 206.92 50.085 207.13 50.155 ;
    RECT 206.92 50.445 207.13 50.515 ;
    RECT 206.46 49.725 206.67 49.795 ;
    RECT 206.46 50.085 206.67 50.155 ;
    RECT 206.46 50.445 206.67 50.515 ;
    RECT 339.72 49.725 339.93 49.795 ;
    RECT 339.72 50.085 339.93 50.155 ;
    RECT 339.72 50.445 339.93 50.515 ;
    RECT 339.26 49.725 339.47 49.795 ;
    RECT 339.26 50.085 339.47 50.155 ;
    RECT 339.26 50.445 339.47 50.515 ;
    RECT 203.6 49.725 203.81 49.795 ;
    RECT 203.6 50.085 203.81 50.155 ;
    RECT 203.6 50.445 203.81 50.515 ;
    RECT 203.14 49.725 203.35 49.795 ;
    RECT 203.14 50.085 203.35 50.155 ;
    RECT 203.14 50.445 203.35 50.515 ;
    RECT 336.4 49.725 336.61 49.795 ;
    RECT 336.4 50.085 336.61 50.155 ;
    RECT 336.4 50.445 336.61 50.515 ;
    RECT 335.94 49.725 336.15 49.795 ;
    RECT 335.94 50.085 336.15 50.155 ;
    RECT 335.94 50.445 336.15 50.515 ;
    RECT 266.68 49.725 266.89 49.795 ;
    RECT 266.68 50.085 266.89 50.155 ;
    RECT 266.68 50.445 266.89 50.515 ;
    RECT 266.22 49.725 266.43 49.795 ;
    RECT 266.22 50.085 266.43 50.155 ;
    RECT 266.22 50.445 266.43 50.515 ;
    RECT 263.36 49.725 263.57 49.795 ;
    RECT 263.36 50.085 263.57 50.155 ;
    RECT 263.36 50.445 263.57 50.515 ;
    RECT 262.9 49.725 263.11 49.795 ;
    RECT 262.9 50.085 263.11 50.155 ;
    RECT 262.9 50.445 263.11 50.515 ;
    RECT 260.04 49.725 260.25 49.795 ;
    RECT 260.04 50.085 260.25 50.155 ;
    RECT 260.04 50.445 260.25 50.515 ;
    RECT 259.58 49.725 259.79 49.795 ;
    RECT 259.58 50.085 259.79 50.155 ;
    RECT 259.58 50.445 259.79 50.515 ;
    RECT 256.72 49.725 256.93 49.795 ;
    RECT 256.72 50.085 256.93 50.155 ;
    RECT 256.72 50.445 256.93 50.515 ;
    RECT 256.26 49.725 256.47 49.795 ;
    RECT 256.26 50.085 256.47 50.155 ;
    RECT 256.26 50.445 256.47 50.515 ;
    RECT 253.4 49.725 253.61 49.795 ;
    RECT 253.4 50.085 253.61 50.155 ;
    RECT 253.4 50.445 253.61 50.515 ;
    RECT 252.94 49.725 253.15 49.795 ;
    RECT 252.94 50.085 253.15 50.155 ;
    RECT 252.94 50.445 253.15 50.515 ;
    RECT 250.08 49.725 250.29 49.795 ;
    RECT 250.08 50.085 250.29 50.155 ;
    RECT 250.08 50.445 250.29 50.515 ;
    RECT 249.62 49.725 249.83 49.795 ;
    RECT 249.62 50.085 249.83 50.155 ;
    RECT 249.62 50.445 249.83 50.515 ;
    RECT 246.76 49.725 246.97 49.795 ;
    RECT 246.76 50.085 246.97 50.155 ;
    RECT 246.76 50.445 246.97 50.515 ;
    RECT 246.3 49.725 246.51 49.795 ;
    RECT 246.3 50.085 246.51 50.155 ;
    RECT 246.3 50.445 246.51 50.515 ;
    RECT 243.44 49.725 243.65 49.795 ;
    RECT 243.44 50.085 243.65 50.155 ;
    RECT 243.44 50.445 243.65 50.515 ;
    RECT 242.98 49.725 243.19 49.795 ;
    RECT 242.98 50.085 243.19 50.155 ;
    RECT 242.98 50.445 243.19 50.515 ;
    RECT 240.12 49.725 240.33 49.795 ;
    RECT 240.12 50.085 240.33 50.155 ;
    RECT 240.12 50.445 240.33 50.515 ;
    RECT 239.66 49.725 239.87 49.795 ;
    RECT 239.66 50.085 239.87 50.155 ;
    RECT 239.66 50.445 239.87 50.515 ;
    RECT 236.8 49.725 237.01 49.795 ;
    RECT 236.8 50.085 237.01 50.155 ;
    RECT 236.8 50.445 237.01 50.515 ;
    RECT 236.34 49.725 236.55 49.795 ;
    RECT 236.34 50.085 236.55 50.155 ;
    RECT 236.34 50.445 236.55 50.515 ;
    RECT 374.15 50.085 374.22 50.155 ;
    RECT 333.08 49.725 333.29 49.795 ;
    RECT 333.08 50.085 333.29 50.155 ;
    RECT 333.08 50.445 333.29 50.515 ;
    RECT 332.62 49.725 332.83 49.795 ;
    RECT 332.62 50.085 332.83 50.155 ;
    RECT 332.62 50.445 332.83 50.515 ;
    RECT 329.76 49.725 329.97 49.795 ;
    RECT 329.76 50.085 329.97 50.155 ;
    RECT 329.76 50.445 329.97 50.515 ;
    RECT 329.3 49.725 329.51 49.795 ;
    RECT 329.3 50.085 329.51 50.155 ;
    RECT 329.3 50.445 329.51 50.515 ;
    RECT 326.44 49.725 326.65 49.795 ;
    RECT 326.44 50.085 326.65 50.155 ;
    RECT 326.44 50.445 326.65 50.515 ;
    RECT 325.98 49.725 326.19 49.795 ;
    RECT 325.98 50.085 326.19 50.155 ;
    RECT 325.98 50.445 326.19 50.515 ;
    RECT 323.12 49.725 323.33 49.795 ;
    RECT 323.12 50.085 323.33 50.155 ;
    RECT 323.12 50.445 323.33 50.515 ;
    RECT 322.66 49.725 322.87 49.795 ;
    RECT 322.66 50.085 322.87 50.155 ;
    RECT 322.66 50.445 322.87 50.515 ;
    RECT 319.8 49.725 320.01 49.795 ;
    RECT 319.8 50.085 320.01 50.155 ;
    RECT 319.8 50.445 320.01 50.515 ;
    RECT 319.34 49.725 319.55 49.795 ;
    RECT 319.34 50.085 319.55 50.155 ;
    RECT 319.34 50.445 319.55 50.515 ;
    RECT 316.48 49.725 316.69 49.795 ;
    RECT 316.48 50.085 316.69 50.155 ;
    RECT 316.48 50.445 316.69 50.515 ;
    RECT 316.02 49.725 316.23 49.795 ;
    RECT 316.02 50.085 316.23 50.155 ;
    RECT 316.02 50.445 316.23 50.515 ;
    RECT 313.16 49.725 313.37 49.795 ;
    RECT 313.16 50.085 313.37 50.155 ;
    RECT 313.16 50.445 313.37 50.515 ;
    RECT 312.7 49.725 312.91 49.795 ;
    RECT 312.7 50.085 312.91 50.155 ;
    RECT 312.7 50.445 312.91 50.515 ;
    RECT 309.84 49.725 310.05 49.795 ;
    RECT 309.84 50.085 310.05 50.155 ;
    RECT 309.84 50.445 310.05 50.515 ;
    RECT 309.38 49.725 309.59 49.795 ;
    RECT 309.38 50.085 309.59 50.155 ;
    RECT 309.38 50.445 309.59 50.515 ;
    RECT 306.52 49.725 306.73 49.795 ;
    RECT 306.52 50.085 306.73 50.155 ;
    RECT 306.52 50.445 306.73 50.515 ;
    RECT 306.06 49.725 306.27 49.795 ;
    RECT 306.06 50.085 306.27 50.155 ;
    RECT 306.06 50.445 306.27 50.515 ;
    RECT 303.2 49.005 303.41 49.075 ;
    RECT 303.2 49.365 303.41 49.435 ;
    RECT 303.2 49.725 303.41 49.795 ;
    RECT 302.74 49.005 302.95 49.075 ;
    RECT 302.74 49.365 302.95 49.435 ;
    RECT 302.74 49.725 302.95 49.795 ;
    RECT 372.92 49.005 373.13 49.075 ;
    RECT 372.92 49.365 373.13 49.435 ;
    RECT 372.92 49.725 373.13 49.795 ;
    RECT 372.46 49.005 372.67 49.075 ;
    RECT 372.46 49.365 372.67 49.435 ;
    RECT 372.46 49.725 372.67 49.795 ;
    RECT 369.6 49.005 369.81 49.075 ;
    RECT 369.6 49.365 369.81 49.435 ;
    RECT 369.6 49.725 369.81 49.795 ;
    RECT 369.14 49.005 369.35 49.075 ;
    RECT 369.14 49.365 369.35 49.435 ;
    RECT 369.14 49.725 369.35 49.795 ;
    RECT 200.605 49.365 200.675 49.435 ;
    RECT 299.88 49.005 300.09 49.075 ;
    RECT 299.88 49.365 300.09 49.435 ;
    RECT 299.88 49.725 300.09 49.795 ;
    RECT 299.42 49.005 299.63 49.075 ;
    RECT 299.42 49.365 299.63 49.435 ;
    RECT 299.42 49.725 299.63 49.795 ;
    RECT 296.56 49.005 296.77 49.075 ;
    RECT 296.56 49.365 296.77 49.435 ;
    RECT 296.56 49.725 296.77 49.795 ;
    RECT 296.1 49.005 296.31 49.075 ;
    RECT 296.1 49.365 296.31 49.435 ;
    RECT 296.1 49.725 296.31 49.795 ;
    RECT 293.24 49.005 293.45 49.075 ;
    RECT 293.24 49.365 293.45 49.435 ;
    RECT 293.24 49.725 293.45 49.795 ;
    RECT 292.78 49.005 292.99 49.075 ;
    RECT 292.78 49.365 292.99 49.435 ;
    RECT 292.78 49.725 292.99 49.795 ;
    RECT 289.92 49.005 290.13 49.075 ;
    RECT 289.92 49.365 290.13 49.435 ;
    RECT 289.92 49.725 290.13 49.795 ;
    RECT 289.46 49.005 289.67 49.075 ;
    RECT 289.46 49.365 289.67 49.435 ;
    RECT 289.46 49.725 289.67 49.795 ;
    RECT 286.6 49.005 286.81 49.075 ;
    RECT 286.6 49.365 286.81 49.435 ;
    RECT 286.6 49.725 286.81 49.795 ;
    RECT 286.14 49.005 286.35 49.075 ;
    RECT 286.14 49.365 286.35 49.435 ;
    RECT 286.14 49.725 286.35 49.795 ;
    RECT 283.28 49.005 283.49 49.075 ;
    RECT 283.28 49.365 283.49 49.435 ;
    RECT 283.28 49.725 283.49 49.795 ;
    RECT 282.82 49.005 283.03 49.075 ;
    RECT 282.82 49.365 283.03 49.435 ;
    RECT 282.82 49.725 283.03 49.795 ;
    RECT 279.96 49.005 280.17 49.075 ;
    RECT 279.96 49.365 280.17 49.435 ;
    RECT 279.96 49.725 280.17 49.795 ;
    RECT 279.5 49.005 279.71 49.075 ;
    RECT 279.5 49.365 279.71 49.435 ;
    RECT 279.5 49.725 279.71 49.795 ;
    RECT 276.64 49.005 276.85 49.075 ;
    RECT 276.64 49.365 276.85 49.435 ;
    RECT 276.64 49.725 276.85 49.795 ;
    RECT 276.18 49.005 276.39 49.075 ;
    RECT 276.18 49.365 276.39 49.435 ;
    RECT 276.18 49.725 276.39 49.795 ;
    RECT 273.32 49.005 273.53 49.075 ;
    RECT 273.32 49.365 273.53 49.435 ;
    RECT 273.32 49.725 273.53 49.795 ;
    RECT 272.86 49.005 273.07 49.075 ;
    RECT 272.86 49.365 273.07 49.435 ;
    RECT 272.86 49.725 273.07 49.795 ;
    RECT 270.0 49.005 270.21 49.075 ;
    RECT 270.0 49.365 270.21 49.435 ;
    RECT 270.0 49.725 270.21 49.795 ;
    RECT 269.54 49.005 269.75 49.075 ;
    RECT 269.54 49.365 269.75 49.435 ;
    RECT 269.54 49.725 269.75 49.795 ;
    RECT 233.48 49.005 233.69 49.075 ;
    RECT 233.48 49.365 233.69 49.435 ;
    RECT 233.48 49.725 233.69 49.795 ;
    RECT 233.02 49.005 233.23 49.075 ;
    RECT 233.02 49.365 233.23 49.435 ;
    RECT 233.02 49.725 233.23 49.795 ;
    RECT 230.16 49.005 230.37 49.075 ;
    RECT 230.16 49.365 230.37 49.435 ;
    RECT 230.16 49.725 230.37 49.795 ;
    RECT 229.7 49.005 229.91 49.075 ;
    RECT 229.7 49.365 229.91 49.435 ;
    RECT 229.7 49.725 229.91 49.795 ;
    RECT 366.28 49.005 366.49 49.075 ;
    RECT 366.28 49.365 366.49 49.435 ;
    RECT 366.28 49.725 366.49 49.795 ;
    RECT 365.82 49.005 366.03 49.075 ;
    RECT 365.82 49.365 366.03 49.435 ;
    RECT 365.82 49.725 366.03 49.795 ;
    RECT 226.84 49.005 227.05 49.075 ;
    RECT 226.84 49.365 227.05 49.435 ;
    RECT 226.84 49.725 227.05 49.795 ;
    RECT 226.38 49.005 226.59 49.075 ;
    RECT 226.38 49.365 226.59 49.435 ;
    RECT 226.38 49.725 226.59 49.795 ;
    RECT 362.96 49.005 363.17 49.075 ;
    RECT 362.96 49.365 363.17 49.435 ;
    RECT 362.96 49.725 363.17 49.795 ;
    RECT 362.5 49.005 362.71 49.075 ;
    RECT 362.5 49.365 362.71 49.435 ;
    RECT 362.5 49.725 362.71 49.795 ;
    RECT 223.52 49.005 223.73 49.075 ;
    RECT 223.52 49.365 223.73 49.435 ;
    RECT 223.52 49.725 223.73 49.795 ;
    RECT 223.06 49.005 223.27 49.075 ;
    RECT 223.06 49.365 223.27 49.435 ;
    RECT 223.06 49.725 223.27 49.795 ;
    RECT 359.64 49.005 359.85 49.075 ;
    RECT 359.64 49.365 359.85 49.435 ;
    RECT 359.64 49.725 359.85 49.795 ;
    RECT 359.18 49.005 359.39 49.075 ;
    RECT 359.18 49.365 359.39 49.435 ;
    RECT 359.18 49.725 359.39 49.795 ;
    RECT 220.2 49.005 220.41 49.075 ;
    RECT 220.2 49.365 220.41 49.435 ;
    RECT 220.2 49.725 220.41 49.795 ;
    RECT 219.74 49.005 219.95 49.075 ;
    RECT 219.74 49.365 219.95 49.435 ;
    RECT 219.74 49.725 219.95 49.795 ;
    RECT 356.32 49.005 356.53 49.075 ;
    RECT 356.32 49.365 356.53 49.435 ;
    RECT 356.32 49.725 356.53 49.795 ;
    RECT 355.86 49.005 356.07 49.075 ;
    RECT 355.86 49.365 356.07 49.435 ;
    RECT 355.86 49.725 356.07 49.795 ;
    RECT 353.0 49.005 353.21 49.075 ;
    RECT 353.0 49.365 353.21 49.435 ;
    RECT 353.0 49.725 353.21 49.795 ;
    RECT 352.54 49.005 352.75 49.075 ;
    RECT 352.54 49.365 352.75 49.435 ;
    RECT 352.54 49.725 352.75 49.795 ;
    RECT 216.88 49.005 217.09 49.075 ;
    RECT 216.88 49.365 217.09 49.435 ;
    RECT 216.88 49.725 217.09 49.795 ;
    RECT 216.42 49.005 216.63 49.075 ;
    RECT 216.42 49.365 216.63 49.435 ;
    RECT 216.42 49.725 216.63 49.795 ;
    RECT 349.68 49.005 349.89 49.075 ;
    RECT 349.68 49.365 349.89 49.435 ;
    RECT 349.68 49.725 349.89 49.795 ;
    RECT 349.22 49.005 349.43 49.075 ;
    RECT 349.22 49.365 349.43 49.435 ;
    RECT 349.22 49.725 349.43 49.795 ;
    RECT 213.56 49.005 213.77 49.075 ;
    RECT 213.56 49.365 213.77 49.435 ;
    RECT 213.56 49.725 213.77 49.795 ;
    RECT 213.1 49.005 213.31 49.075 ;
    RECT 213.1 49.365 213.31 49.435 ;
    RECT 213.1 49.725 213.31 49.795 ;
    RECT 346.36 49.005 346.57 49.075 ;
    RECT 346.36 49.365 346.57 49.435 ;
    RECT 346.36 49.725 346.57 49.795 ;
    RECT 345.9 49.005 346.11 49.075 ;
    RECT 345.9 49.365 346.11 49.435 ;
    RECT 345.9 49.725 346.11 49.795 ;
    RECT 210.24 49.005 210.45 49.075 ;
    RECT 210.24 49.365 210.45 49.435 ;
    RECT 210.24 49.725 210.45 49.795 ;
    RECT 209.78 49.005 209.99 49.075 ;
    RECT 209.78 49.365 209.99 49.435 ;
    RECT 209.78 49.725 209.99 49.795 ;
    RECT 343.04 49.005 343.25 49.075 ;
    RECT 343.04 49.365 343.25 49.435 ;
    RECT 343.04 49.725 343.25 49.795 ;
    RECT 342.58 49.005 342.79 49.075 ;
    RECT 342.58 49.365 342.79 49.435 ;
    RECT 342.58 49.725 342.79 49.795 ;
    RECT 206.92 49.005 207.13 49.075 ;
    RECT 206.92 49.365 207.13 49.435 ;
    RECT 206.92 49.725 207.13 49.795 ;
    RECT 206.46 49.005 206.67 49.075 ;
    RECT 206.46 49.365 206.67 49.435 ;
    RECT 206.46 49.725 206.67 49.795 ;
    RECT 339.72 49.005 339.93 49.075 ;
    RECT 339.72 49.365 339.93 49.435 ;
    RECT 339.72 49.725 339.93 49.795 ;
    RECT 339.26 49.005 339.47 49.075 ;
    RECT 339.26 49.365 339.47 49.435 ;
    RECT 339.26 49.725 339.47 49.795 ;
    RECT 203.6 49.005 203.81 49.075 ;
    RECT 203.6 49.365 203.81 49.435 ;
    RECT 203.6 49.725 203.81 49.795 ;
    RECT 203.14 49.005 203.35 49.075 ;
    RECT 203.14 49.365 203.35 49.435 ;
    RECT 203.14 49.725 203.35 49.795 ;
    RECT 336.4 49.005 336.61 49.075 ;
    RECT 336.4 49.365 336.61 49.435 ;
    RECT 336.4 49.725 336.61 49.795 ;
    RECT 335.94 49.005 336.15 49.075 ;
    RECT 335.94 49.365 336.15 49.435 ;
    RECT 335.94 49.725 336.15 49.795 ;
    RECT 266.68 49.005 266.89 49.075 ;
    RECT 266.68 49.365 266.89 49.435 ;
    RECT 266.68 49.725 266.89 49.795 ;
    RECT 266.22 49.005 266.43 49.075 ;
    RECT 266.22 49.365 266.43 49.435 ;
    RECT 266.22 49.725 266.43 49.795 ;
    RECT 263.36 49.005 263.57 49.075 ;
    RECT 263.36 49.365 263.57 49.435 ;
    RECT 263.36 49.725 263.57 49.795 ;
    RECT 262.9 49.005 263.11 49.075 ;
    RECT 262.9 49.365 263.11 49.435 ;
    RECT 262.9 49.725 263.11 49.795 ;
    RECT 260.04 49.005 260.25 49.075 ;
    RECT 260.04 49.365 260.25 49.435 ;
    RECT 260.04 49.725 260.25 49.795 ;
    RECT 259.58 49.005 259.79 49.075 ;
    RECT 259.58 49.365 259.79 49.435 ;
    RECT 259.58 49.725 259.79 49.795 ;
    RECT 256.72 49.005 256.93 49.075 ;
    RECT 256.72 49.365 256.93 49.435 ;
    RECT 256.72 49.725 256.93 49.795 ;
    RECT 256.26 49.005 256.47 49.075 ;
    RECT 256.26 49.365 256.47 49.435 ;
    RECT 256.26 49.725 256.47 49.795 ;
    RECT 253.4 49.005 253.61 49.075 ;
    RECT 253.4 49.365 253.61 49.435 ;
    RECT 253.4 49.725 253.61 49.795 ;
    RECT 252.94 49.005 253.15 49.075 ;
    RECT 252.94 49.365 253.15 49.435 ;
    RECT 252.94 49.725 253.15 49.795 ;
    RECT 250.08 49.005 250.29 49.075 ;
    RECT 250.08 49.365 250.29 49.435 ;
    RECT 250.08 49.725 250.29 49.795 ;
    RECT 249.62 49.005 249.83 49.075 ;
    RECT 249.62 49.365 249.83 49.435 ;
    RECT 249.62 49.725 249.83 49.795 ;
    RECT 246.76 49.005 246.97 49.075 ;
    RECT 246.76 49.365 246.97 49.435 ;
    RECT 246.76 49.725 246.97 49.795 ;
    RECT 246.3 49.005 246.51 49.075 ;
    RECT 246.3 49.365 246.51 49.435 ;
    RECT 246.3 49.725 246.51 49.795 ;
    RECT 243.44 49.005 243.65 49.075 ;
    RECT 243.44 49.365 243.65 49.435 ;
    RECT 243.44 49.725 243.65 49.795 ;
    RECT 242.98 49.005 243.19 49.075 ;
    RECT 242.98 49.365 243.19 49.435 ;
    RECT 242.98 49.725 243.19 49.795 ;
    RECT 240.12 49.005 240.33 49.075 ;
    RECT 240.12 49.365 240.33 49.435 ;
    RECT 240.12 49.725 240.33 49.795 ;
    RECT 239.66 49.005 239.87 49.075 ;
    RECT 239.66 49.365 239.87 49.435 ;
    RECT 239.66 49.725 239.87 49.795 ;
    RECT 236.8 49.005 237.01 49.075 ;
    RECT 236.8 49.365 237.01 49.435 ;
    RECT 236.8 49.725 237.01 49.795 ;
    RECT 236.34 49.005 236.55 49.075 ;
    RECT 236.34 49.365 236.55 49.435 ;
    RECT 236.34 49.725 236.55 49.795 ;
    RECT 374.15 49.365 374.22 49.435 ;
    RECT 333.08 49.005 333.29 49.075 ;
    RECT 333.08 49.365 333.29 49.435 ;
    RECT 333.08 49.725 333.29 49.795 ;
    RECT 332.62 49.005 332.83 49.075 ;
    RECT 332.62 49.365 332.83 49.435 ;
    RECT 332.62 49.725 332.83 49.795 ;
    RECT 329.76 49.005 329.97 49.075 ;
    RECT 329.76 49.365 329.97 49.435 ;
    RECT 329.76 49.725 329.97 49.795 ;
    RECT 329.3 49.005 329.51 49.075 ;
    RECT 329.3 49.365 329.51 49.435 ;
    RECT 329.3 49.725 329.51 49.795 ;
    RECT 326.44 49.005 326.65 49.075 ;
    RECT 326.44 49.365 326.65 49.435 ;
    RECT 326.44 49.725 326.65 49.795 ;
    RECT 325.98 49.005 326.19 49.075 ;
    RECT 325.98 49.365 326.19 49.435 ;
    RECT 325.98 49.725 326.19 49.795 ;
    RECT 323.12 49.005 323.33 49.075 ;
    RECT 323.12 49.365 323.33 49.435 ;
    RECT 323.12 49.725 323.33 49.795 ;
    RECT 322.66 49.005 322.87 49.075 ;
    RECT 322.66 49.365 322.87 49.435 ;
    RECT 322.66 49.725 322.87 49.795 ;
    RECT 319.8 49.005 320.01 49.075 ;
    RECT 319.8 49.365 320.01 49.435 ;
    RECT 319.8 49.725 320.01 49.795 ;
    RECT 319.34 49.005 319.55 49.075 ;
    RECT 319.34 49.365 319.55 49.435 ;
    RECT 319.34 49.725 319.55 49.795 ;
    RECT 316.48 49.005 316.69 49.075 ;
    RECT 316.48 49.365 316.69 49.435 ;
    RECT 316.48 49.725 316.69 49.795 ;
    RECT 316.02 49.005 316.23 49.075 ;
    RECT 316.02 49.365 316.23 49.435 ;
    RECT 316.02 49.725 316.23 49.795 ;
    RECT 313.16 49.005 313.37 49.075 ;
    RECT 313.16 49.365 313.37 49.435 ;
    RECT 313.16 49.725 313.37 49.795 ;
    RECT 312.7 49.005 312.91 49.075 ;
    RECT 312.7 49.365 312.91 49.435 ;
    RECT 312.7 49.725 312.91 49.795 ;
    RECT 309.84 49.005 310.05 49.075 ;
    RECT 309.84 49.365 310.05 49.435 ;
    RECT 309.84 49.725 310.05 49.795 ;
    RECT 309.38 49.005 309.59 49.075 ;
    RECT 309.38 49.365 309.59 49.435 ;
    RECT 309.38 49.725 309.59 49.795 ;
    RECT 306.52 49.005 306.73 49.075 ;
    RECT 306.52 49.365 306.73 49.435 ;
    RECT 306.52 49.725 306.73 49.795 ;
    RECT 306.06 49.005 306.27 49.075 ;
    RECT 306.06 49.365 306.27 49.435 ;
    RECT 306.06 49.725 306.27 49.795 ;
    RECT 303.2 48.285 303.41 48.355 ;
    RECT 303.2 48.645 303.41 48.715 ;
    RECT 303.2 49.005 303.41 49.075 ;
    RECT 302.74 48.285 302.95 48.355 ;
    RECT 302.74 48.645 302.95 48.715 ;
    RECT 302.74 49.005 302.95 49.075 ;
    RECT 372.92 48.285 373.13 48.355 ;
    RECT 372.92 48.645 373.13 48.715 ;
    RECT 372.92 49.005 373.13 49.075 ;
    RECT 372.46 48.285 372.67 48.355 ;
    RECT 372.46 48.645 372.67 48.715 ;
    RECT 372.46 49.005 372.67 49.075 ;
    RECT 369.6 48.285 369.81 48.355 ;
    RECT 369.6 48.645 369.81 48.715 ;
    RECT 369.6 49.005 369.81 49.075 ;
    RECT 369.14 48.285 369.35 48.355 ;
    RECT 369.14 48.645 369.35 48.715 ;
    RECT 369.14 49.005 369.35 49.075 ;
    RECT 200.605 48.645 200.675 48.715 ;
    RECT 299.88 48.285 300.09 48.355 ;
    RECT 299.88 48.645 300.09 48.715 ;
    RECT 299.88 49.005 300.09 49.075 ;
    RECT 299.42 48.285 299.63 48.355 ;
    RECT 299.42 48.645 299.63 48.715 ;
    RECT 299.42 49.005 299.63 49.075 ;
    RECT 296.56 48.285 296.77 48.355 ;
    RECT 296.56 48.645 296.77 48.715 ;
    RECT 296.56 49.005 296.77 49.075 ;
    RECT 296.1 48.285 296.31 48.355 ;
    RECT 296.1 48.645 296.31 48.715 ;
    RECT 296.1 49.005 296.31 49.075 ;
    RECT 293.24 48.285 293.45 48.355 ;
    RECT 293.24 48.645 293.45 48.715 ;
    RECT 293.24 49.005 293.45 49.075 ;
    RECT 292.78 48.285 292.99 48.355 ;
    RECT 292.78 48.645 292.99 48.715 ;
    RECT 292.78 49.005 292.99 49.075 ;
    RECT 289.92 48.285 290.13 48.355 ;
    RECT 289.92 48.645 290.13 48.715 ;
    RECT 289.92 49.005 290.13 49.075 ;
    RECT 289.46 48.285 289.67 48.355 ;
    RECT 289.46 48.645 289.67 48.715 ;
    RECT 289.46 49.005 289.67 49.075 ;
    RECT 286.6 48.285 286.81 48.355 ;
    RECT 286.6 48.645 286.81 48.715 ;
    RECT 286.6 49.005 286.81 49.075 ;
    RECT 286.14 48.285 286.35 48.355 ;
    RECT 286.14 48.645 286.35 48.715 ;
    RECT 286.14 49.005 286.35 49.075 ;
    RECT 283.28 48.285 283.49 48.355 ;
    RECT 283.28 48.645 283.49 48.715 ;
    RECT 283.28 49.005 283.49 49.075 ;
    RECT 282.82 48.285 283.03 48.355 ;
    RECT 282.82 48.645 283.03 48.715 ;
    RECT 282.82 49.005 283.03 49.075 ;
    RECT 279.96 48.285 280.17 48.355 ;
    RECT 279.96 48.645 280.17 48.715 ;
    RECT 279.96 49.005 280.17 49.075 ;
    RECT 279.5 48.285 279.71 48.355 ;
    RECT 279.5 48.645 279.71 48.715 ;
    RECT 279.5 49.005 279.71 49.075 ;
    RECT 276.64 48.285 276.85 48.355 ;
    RECT 276.64 48.645 276.85 48.715 ;
    RECT 276.64 49.005 276.85 49.075 ;
    RECT 276.18 48.285 276.39 48.355 ;
    RECT 276.18 48.645 276.39 48.715 ;
    RECT 276.18 49.005 276.39 49.075 ;
    RECT 273.32 48.285 273.53 48.355 ;
    RECT 273.32 48.645 273.53 48.715 ;
    RECT 273.32 49.005 273.53 49.075 ;
    RECT 272.86 48.285 273.07 48.355 ;
    RECT 272.86 48.645 273.07 48.715 ;
    RECT 272.86 49.005 273.07 49.075 ;
    RECT 270.0 48.285 270.21 48.355 ;
    RECT 270.0 48.645 270.21 48.715 ;
    RECT 270.0 49.005 270.21 49.075 ;
    RECT 269.54 48.285 269.75 48.355 ;
    RECT 269.54 48.645 269.75 48.715 ;
    RECT 269.54 49.005 269.75 49.075 ;
    RECT 233.48 48.285 233.69 48.355 ;
    RECT 233.48 48.645 233.69 48.715 ;
    RECT 233.48 49.005 233.69 49.075 ;
    RECT 233.02 48.285 233.23 48.355 ;
    RECT 233.02 48.645 233.23 48.715 ;
    RECT 233.02 49.005 233.23 49.075 ;
    RECT 230.16 48.285 230.37 48.355 ;
    RECT 230.16 48.645 230.37 48.715 ;
    RECT 230.16 49.005 230.37 49.075 ;
    RECT 229.7 48.285 229.91 48.355 ;
    RECT 229.7 48.645 229.91 48.715 ;
    RECT 229.7 49.005 229.91 49.075 ;
    RECT 366.28 48.285 366.49 48.355 ;
    RECT 366.28 48.645 366.49 48.715 ;
    RECT 366.28 49.005 366.49 49.075 ;
    RECT 365.82 48.285 366.03 48.355 ;
    RECT 365.82 48.645 366.03 48.715 ;
    RECT 365.82 49.005 366.03 49.075 ;
    RECT 226.84 48.285 227.05 48.355 ;
    RECT 226.84 48.645 227.05 48.715 ;
    RECT 226.84 49.005 227.05 49.075 ;
    RECT 226.38 48.285 226.59 48.355 ;
    RECT 226.38 48.645 226.59 48.715 ;
    RECT 226.38 49.005 226.59 49.075 ;
    RECT 362.96 48.285 363.17 48.355 ;
    RECT 362.96 48.645 363.17 48.715 ;
    RECT 362.96 49.005 363.17 49.075 ;
    RECT 362.5 48.285 362.71 48.355 ;
    RECT 362.5 48.645 362.71 48.715 ;
    RECT 362.5 49.005 362.71 49.075 ;
    RECT 223.52 48.285 223.73 48.355 ;
    RECT 223.52 48.645 223.73 48.715 ;
    RECT 223.52 49.005 223.73 49.075 ;
    RECT 223.06 48.285 223.27 48.355 ;
    RECT 223.06 48.645 223.27 48.715 ;
    RECT 223.06 49.005 223.27 49.075 ;
    RECT 359.64 48.285 359.85 48.355 ;
    RECT 359.64 48.645 359.85 48.715 ;
    RECT 359.64 49.005 359.85 49.075 ;
    RECT 359.18 48.285 359.39 48.355 ;
    RECT 359.18 48.645 359.39 48.715 ;
    RECT 359.18 49.005 359.39 49.075 ;
    RECT 220.2 48.285 220.41 48.355 ;
    RECT 220.2 48.645 220.41 48.715 ;
    RECT 220.2 49.005 220.41 49.075 ;
    RECT 219.74 48.285 219.95 48.355 ;
    RECT 219.74 48.645 219.95 48.715 ;
    RECT 219.74 49.005 219.95 49.075 ;
    RECT 356.32 48.285 356.53 48.355 ;
    RECT 356.32 48.645 356.53 48.715 ;
    RECT 356.32 49.005 356.53 49.075 ;
    RECT 355.86 48.285 356.07 48.355 ;
    RECT 355.86 48.645 356.07 48.715 ;
    RECT 355.86 49.005 356.07 49.075 ;
    RECT 353.0 48.285 353.21 48.355 ;
    RECT 353.0 48.645 353.21 48.715 ;
    RECT 353.0 49.005 353.21 49.075 ;
    RECT 352.54 48.285 352.75 48.355 ;
    RECT 352.54 48.645 352.75 48.715 ;
    RECT 352.54 49.005 352.75 49.075 ;
    RECT 216.88 48.285 217.09 48.355 ;
    RECT 216.88 48.645 217.09 48.715 ;
    RECT 216.88 49.005 217.09 49.075 ;
    RECT 216.42 48.285 216.63 48.355 ;
    RECT 216.42 48.645 216.63 48.715 ;
    RECT 216.42 49.005 216.63 49.075 ;
    RECT 349.68 48.285 349.89 48.355 ;
    RECT 349.68 48.645 349.89 48.715 ;
    RECT 349.68 49.005 349.89 49.075 ;
    RECT 349.22 48.285 349.43 48.355 ;
    RECT 349.22 48.645 349.43 48.715 ;
    RECT 349.22 49.005 349.43 49.075 ;
    RECT 213.56 48.285 213.77 48.355 ;
    RECT 213.56 48.645 213.77 48.715 ;
    RECT 213.56 49.005 213.77 49.075 ;
    RECT 213.1 48.285 213.31 48.355 ;
    RECT 213.1 48.645 213.31 48.715 ;
    RECT 213.1 49.005 213.31 49.075 ;
    RECT 346.36 48.285 346.57 48.355 ;
    RECT 346.36 48.645 346.57 48.715 ;
    RECT 346.36 49.005 346.57 49.075 ;
    RECT 345.9 48.285 346.11 48.355 ;
    RECT 345.9 48.645 346.11 48.715 ;
    RECT 345.9 49.005 346.11 49.075 ;
    RECT 210.24 48.285 210.45 48.355 ;
    RECT 210.24 48.645 210.45 48.715 ;
    RECT 210.24 49.005 210.45 49.075 ;
    RECT 209.78 48.285 209.99 48.355 ;
    RECT 209.78 48.645 209.99 48.715 ;
    RECT 209.78 49.005 209.99 49.075 ;
    RECT 343.04 48.285 343.25 48.355 ;
    RECT 343.04 48.645 343.25 48.715 ;
    RECT 343.04 49.005 343.25 49.075 ;
    RECT 342.58 48.285 342.79 48.355 ;
    RECT 342.58 48.645 342.79 48.715 ;
    RECT 342.58 49.005 342.79 49.075 ;
    RECT 206.92 48.285 207.13 48.355 ;
    RECT 206.92 48.645 207.13 48.715 ;
    RECT 206.92 49.005 207.13 49.075 ;
    RECT 206.46 48.285 206.67 48.355 ;
    RECT 206.46 48.645 206.67 48.715 ;
    RECT 206.46 49.005 206.67 49.075 ;
    RECT 339.72 48.285 339.93 48.355 ;
    RECT 339.72 48.645 339.93 48.715 ;
    RECT 339.72 49.005 339.93 49.075 ;
    RECT 339.26 48.285 339.47 48.355 ;
    RECT 339.26 48.645 339.47 48.715 ;
    RECT 339.26 49.005 339.47 49.075 ;
    RECT 203.6 48.285 203.81 48.355 ;
    RECT 203.6 48.645 203.81 48.715 ;
    RECT 203.6 49.005 203.81 49.075 ;
    RECT 203.14 48.285 203.35 48.355 ;
    RECT 203.14 48.645 203.35 48.715 ;
    RECT 203.14 49.005 203.35 49.075 ;
    RECT 336.4 48.285 336.61 48.355 ;
    RECT 336.4 48.645 336.61 48.715 ;
    RECT 336.4 49.005 336.61 49.075 ;
    RECT 335.94 48.285 336.15 48.355 ;
    RECT 335.94 48.645 336.15 48.715 ;
    RECT 335.94 49.005 336.15 49.075 ;
    RECT 266.68 48.285 266.89 48.355 ;
    RECT 266.68 48.645 266.89 48.715 ;
    RECT 266.68 49.005 266.89 49.075 ;
    RECT 266.22 48.285 266.43 48.355 ;
    RECT 266.22 48.645 266.43 48.715 ;
    RECT 266.22 49.005 266.43 49.075 ;
    RECT 263.36 48.285 263.57 48.355 ;
    RECT 263.36 48.645 263.57 48.715 ;
    RECT 263.36 49.005 263.57 49.075 ;
    RECT 262.9 48.285 263.11 48.355 ;
    RECT 262.9 48.645 263.11 48.715 ;
    RECT 262.9 49.005 263.11 49.075 ;
    RECT 260.04 48.285 260.25 48.355 ;
    RECT 260.04 48.645 260.25 48.715 ;
    RECT 260.04 49.005 260.25 49.075 ;
    RECT 259.58 48.285 259.79 48.355 ;
    RECT 259.58 48.645 259.79 48.715 ;
    RECT 259.58 49.005 259.79 49.075 ;
    RECT 256.72 48.285 256.93 48.355 ;
    RECT 256.72 48.645 256.93 48.715 ;
    RECT 256.72 49.005 256.93 49.075 ;
    RECT 256.26 48.285 256.47 48.355 ;
    RECT 256.26 48.645 256.47 48.715 ;
    RECT 256.26 49.005 256.47 49.075 ;
    RECT 253.4 48.285 253.61 48.355 ;
    RECT 253.4 48.645 253.61 48.715 ;
    RECT 253.4 49.005 253.61 49.075 ;
    RECT 252.94 48.285 253.15 48.355 ;
    RECT 252.94 48.645 253.15 48.715 ;
    RECT 252.94 49.005 253.15 49.075 ;
    RECT 250.08 48.285 250.29 48.355 ;
    RECT 250.08 48.645 250.29 48.715 ;
    RECT 250.08 49.005 250.29 49.075 ;
    RECT 249.62 48.285 249.83 48.355 ;
    RECT 249.62 48.645 249.83 48.715 ;
    RECT 249.62 49.005 249.83 49.075 ;
    RECT 246.76 48.285 246.97 48.355 ;
    RECT 246.76 48.645 246.97 48.715 ;
    RECT 246.76 49.005 246.97 49.075 ;
    RECT 246.3 48.285 246.51 48.355 ;
    RECT 246.3 48.645 246.51 48.715 ;
    RECT 246.3 49.005 246.51 49.075 ;
    RECT 243.44 48.285 243.65 48.355 ;
    RECT 243.44 48.645 243.65 48.715 ;
    RECT 243.44 49.005 243.65 49.075 ;
    RECT 242.98 48.285 243.19 48.355 ;
    RECT 242.98 48.645 243.19 48.715 ;
    RECT 242.98 49.005 243.19 49.075 ;
    RECT 240.12 48.285 240.33 48.355 ;
    RECT 240.12 48.645 240.33 48.715 ;
    RECT 240.12 49.005 240.33 49.075 ;
    RECT 239.66 48.285 239.87 48.355 ;
    RECT 239.66 48.645 239.87 48.715 ;
    RECT 239.66 49.005 239.87 49.075 ;
    RECT 236.8 48.285 237.01 48.355 ;
    RECT 236.8 48.645 237.01 48.715 ;
    RECT 236.8 49.005 237.01 49.075 ;
    RECT 236.34 48.285 236.55 48.355 ;
    RECT 236.34 48.645 236.55 48.715 ;
    RECT 236.34 49.005 236.55 49.075 ;
    RECT 374.15 48.645 374.22 48.715 ;
    RECT 333.08 48.285 333.29 48.355 ;
    RECT 333.08 48.645 333.29 48.715 ;
    RECT 333.08 49.005 333.29 49.075 ;
    RECT 332.62 48.285 332.83 48.355 ;
    RECT 332.62 48.645 332.83 48.715 ;
    RECT 332.62 49.005 332.83 49.075 ;
    RECT 329.76 48.285 329.97 48.355 ;
    RECT 329.76 48.645 329.97 48.715 ;
    RECT 329.76 49.005 329.97 49.075 ;
    RECT 329.3 48.285 329.51 48.355 ;
    RECT 329.3 48.645 329.51 48.715 ;
    RECT 329.3 49.005 329.51 49.075 ;
    RECT 326.44 48.285 326.65 48.355 ;
    RECT 326.44 48.645 326.65 48.715 ;
    RECT 326.44 49.005 326.65 49.075 ;
    RECT 325.98 48.285 326.19 48.355 ;
    RECT 325.98 48.645 326.19 48.715 ;
    RECT 325.98 49.005 326.19 49.075 ;
    RECT 323.12 48.285 323.33 48.355 ;
    RECT 323.12 48.645 323.33 48.715 ;
    RECT 323.12 49.005 323.33 49.075 ;
    RECT 322.66 48.285 322.87 48.355 ;
    RECT 322.66 48.645 322.87 48.715 ;
    RECT 322.66 49.005 322.87 49.075 ;
    RECT 319.8 48.285 320.01 48.355 ;
    RECT 319.8 48.645 320.01 48.715 ;
    RECT 319.8 49.005 320.01 49.075 ;
    RECT 319.34 48.285 319.55 48.355 ;
    RECT 319.34 48.645 319.55 48.715 ;
    RECT 319.34 49.005 319.55 49.075 ;
    RECT 316.48 48.285 316.69 48.355 ;
    RECT 316.48 48.645 316.69 48.715 ;
    RECT 316.48 49.005 316.69 49.075 ;
    RECT 316.02 48.285 316.23 48.355 ;
    RECT 316.02 48.645 316.23 48.715 ;
    RECT 316.02 49.005 316.23 49.075 ;
    RECT 313.16 48.285 313.37 48.355 ;
    RECT 313.16 48.645 313.37 48.715 ;
    RECT 313.16 49.005 313.37 49.075 ;
    RECT 312.7 48.285 312.91 48.355 ;
    RECT 312.7 48.645 312.91 48.715 ;
    RECT 312.7 49.005 312.91 49.075 ;
    RECT 309.84 48.285 310.05 48.355 ;
    RECT 309.84 48.645 310.05 48.715 ;
    RECT 309.84 49.005 310.05 49.075 ;
    RECT 309.38 48.285 309.59 48.355 ;
    RECT 309.38 48.645 309.59 48.715 ;
    RECT 309.38 49.005 309.59 49.075 ;
    RECT 306.52 48.285 306.73 48.355 ;
    RECT 306.52 48.645 306.73 48.715 ;
    RECT 306.52 49.005 306.73 49.075 ;
    RECT 306.06 48.285 306.27 48.355 ;
    RECT 306.06 48.645 306.27 48.715 ;
    RECT 306.06 49.005 306.27 49.075 ;
    RECT 303.2 47.565 303.41 47.635 ;
    RECT 303.2 47.925 303.41 47.995 ;
    RECT 303.2 48.285 303.41 48.355 ;
    RECT 302.74 47.565 302.95 47.635 ;
    RECT 302.74 47.925 302.95 47.995 ;
    RECT 302.74 48.285 302.95 48.355 ;
    RECT 372.92 47.565 373.13 47.635 ;
    RECT 372.92 47.925 373.13 47.995 ;
    RECT 372.92 48.285 373.13 48.355 ;
    RECT 372.46 47.565 372.67 47.635 ;
    RECT 372.46 47.925 372.67 47.995 ;
    RECT 372.46 48.285 372.67 48.355 ;
    RECT 369.6 47.565 369.81 47.635 ;
    RECT 369.6 47.925 369.81 47.995 ;
    RECT 369.6 48.285 369.81 48.355 ;
    RECT 369.14 47.565 369.35 47.635 ;
    RECT 369.14 47.925 369.35 47.995 ;
    RECT 369.14 48.285 369.35 48.355 ;
    RECT 200.605 47.925 200.675 47.995 ;
    RECT 299.88 47.565 300.09 47.635 ;
    RECT 299.88 47.925 300.09 47.995 ;
    RECT 299.88 48.285 300.09 48.355 ;
    RECT 299.42 47.565 299.63 47.635 ;
    RECT 299.42 47.925 299.63 47.995 ;
    RECT 299.42 48.285 299.63 48.355 ;
    RECT 296.56 47.565 296.77 47.635 ;
    RECT 296.56 47.925 296.77 47.995 ;
    RECT 296.56 48.285 296.77 48.355 ;
    RECT 296.1 47.565 296.31 47.635 ;
    RECT 296.1 47.925 296.31 47.995 ;
    RECT 296.1 48.285 296.31 48.355 ;
    RECT 293.24 47.565 293.45 47.635 ;
    RECT 293.24 47.925 293.45 47.995 ;
    RECT 293.24 48.285 293.45 48.355 ;
    RECT 292.78 47.565 292.99 47.635 ;
    RECT 292.78 47.925 292.99 47.995 ;
    RECT 292.78 48.285 292.99 48.355 ;
    RECT 289.92 47.565 290.13 47.635 ;
    RECT 289.92 47.925 290.13 47.995 ;
    RECT 289.92 48.285 290.13 48.355 ;
    RECT 289.46 47.565 289.67 47.635 ;
    RECT 289.46 47.925 289.67 47.995 ;
    RECT 289.46 48.285 289.67 48.355 ;
    RECT 286.6 47.565 286.81 47.635 ;
    RECT 286.6 47.925 286.81 47.995 ;
    RECT 286.6 48.285 286.81 48.355 ;
    RECT 286.14 47.565 286.35 47.635 ;
    RECT 286.14 47.925 286.35 47.995 ;
    RECT 286.14 48.285 286.35 48.355 ;
    RECT 283.28 47.565 283.49 47.635 ;
    RECT 283.28 47.925 283.49 47.995 ;
    RECT 283.28 48.285 283.49 48.355 ;
    RECT 282.82 47.565 283.03 47.635 ;
    RECT 282.82 47.925 283.03 47.995 ;
    RECT 282.82 48.285 283.03 48.355 ;
    RECT 279.96 47.565 280.17 47.635 ;
    RECT 279.96 47.925 280.17 47.995 ;
    RECT 279.96 48.285 280.17 48.355 ;
    RECT 279.5 47.565 279.71 47.635 ;
    RECT 279.5 47.925 279.71 47.995 ;
    RECT 279.5 48.285 279.71 48.355 ;
    RECT 276.64 47.565 276.85 47.635 ;
    RECT 276.64 47.925 276.85 47.995 ;
    RECT 276.64 48.285 276.85 48.355 ;
    RECT 276.18 47.565 276.39 47.635 ;
    RECT 276.18 47.925 276.39 47.995 ;
    RECT 276.18 48.285 276.39 48.355 ;
    RECT 273.32 47.565 273.53 47.635 ;
    RECT 273.32 47.925 273.53 47.995 ;
    RECT 273.32 48.285 273.53 48.355 ;
    RECT 272.86 47.565 273.07 47.635 ;
    RECT 272.86 47.925 273.07 47.995 ;
    RECT 272.86 48.285 273.07 48.355 ;
    RECT 270.0 47.565 270.21 47.635 ;
    RECT 270.0 47.925 270.21 47.995 ;
    RECT 270.0 48.285 270.21 48.355 ;
    RECT 269.54 47.565 269.75 47.635 ;
    RECT 269.54 47.925 269.75 47.995 ;
    RECT 269.54 48.285 269.75 48.355 ;
    RECT 233.48 47.565 233.69 47.635 ;
    RECT 233.48 47.925 233.69 47.995 ;
    RECT 233.48 48.285 233.69 48.355 ;
    RECT 233.02 47.565 233.23 47.635 ;
    RECT 233.02 47.925 233.23 47.995 ;
    RECT 233.02 48.285 233.23 48.355 ;
    RECT 230.16 47.565 230.37 47.635 ;
    RECT 230.16 47.925 230.37 47.995 ;
    RECT 230.16 48.285 230.37 48.355 ;
    RECT 229.7 47.565 229.91 47.635 ;
    RECT 229.7 47.925 229.91 47.995 ;
    RECT 229.7 48.285 229.91 48.355 ;
    RECT 366.28 47.565 366.49 47.635 ;
    RECT 366.28 47.925 366.49 47.995 ;
    RECT 366.28 48.285 366.49 48.355 ;
    RECT 365.82 47.565 366.03 47.635 ;
    RECT 365.82 47.925 366.03 47.995 ;
    RECT 365.82 48.285 366.03 48.355 ;
    RECT 226.84 47.565 227.05 47.635 ;
    RECT 226.84 47.925 227.05 47.995 ;
    RECT 226.84 48.285 227.05 48.355 ;
    RECT 226.38 47.565 226.59 47.635 ;
    RECT 226.38 47.925 226.59 47.995 ;
    RECT 226.38 48.285 226.59 48.355 ;
    RECT 362.96 47.565 363.17 47.635 ;
    RECT 362.96 47.925 363.17 47.995 ;
    RECT 362.96 48.285 363.17 48.355 ;
    RECT 362.5 47.565 362.71 47.635 ;
    RECT 362.5 47.925 362.71 47.995 ;
    RECT 362.5 48.285 362.71 48.355 ;
    RECT 223.52 47.565 223.73 47.635 ;
    RECT 223.52 47.925 223.73 47.995 ;
    RECT 223.52 48.285 223.73 48.355 ;
    RECT 223.06 47.565 223.27 47.635 ;
    RECT 223.06 47.925 223.27 47.995 ;
    RECT 223.06 48.285 223.27 48.355 ;
    RECT 359.64 47.565 359.85 47.635 ;
    RECT 359.64 47.925 359.85 47.995 ;
    RECT 359.64 48.285 359.85 48.355 ;
    RECT 359.18 47.565 359.39 47.635 ;
    RECT 359.18 47.925 359.39 47.995 ;
    RECT 359.18 48.285 359.39 48.355 ;
    RECT 220.2 47.565 220.41 47.635 ;
    RECT 220.2 47.925 220.41 47.995 ;
    RECT 220.2 48.285 220.41 48.355 ;
    RECT 219.74 47.565 219.95 47.635 ;
    RECT 219.74 47.925 219.95 47.995 ;
    RECT 219.74 48.285 219.95 48.355 ;
    RECT 356.32 47.565 356.53 47.635 ;
    RECT 356.32 47.925 356.53 47.995 ;
    RECT 356.32 48.285 356.53 48.355 ;
    RECT 355.86 47.565 356.07 47.635 ;
    RECT 355.86 47.925 356.07 47.995 ;
    RECT 355.86 48.285 356.07 48.355 ;
    RECT 353.0 47.565 353.21 47.635 ;
    RECT 353.0 47.925 353.21 47.995 ;
    RECT 353.0 48.285 353.21 48.355 ;
    RECT 352.54 47.565 352.75 47.635 ;
    RECT 352.54 47.925 352.75 47.995 ;
    RECT 352.54 48.285 352.75 48.355 ;
    RECT 216.88 47.565 217.09 47.635 ;
    RECT 216.88 47.925 217.09 47.995 ;
    RECT 216.88 48.285 217.09 48.355 ;
    RECT 216.42 47.565 216.63 47.635 ;
    RECT 216.42 47.925 216.63 47.995 ;
    RECT 216.42 48.285 216.63 48.355 ;
    RECT 349.68 47.565 349.89 47.635 ;
    RECT 349.68 47.925 349.89 47.995 ;
    RECT 349.68 48.285 349.89 48.355 ;
    RECT 349.22 47.565 349.43 47.635 ;
    RECT 349.22 47.925 349.43 47.995 ;
    RECT 349.22 48.285 349.43 48.355 ;
    RECT 213.56 47.565 213.77 47.635 ;
    RECT 213.56 47.925 213.77 47.995 ;
    RECT 213.56 48.285 213.77 48.355 ;
    RECT 213.1 47.565 213.31 47.635 ;
    RECT 213.1 47.925 213.31 47.995 ;
    RECT 213.1 48.285 213.31 48.355 ;
    RECT 346.36 47.565 346.57 47.635 ;
    RECT 346.36 47.925 346.57 47.995 ;
    RECT 346.36 48.285 346.57 48.355 ;
    RECT 345.9 47.565 346.11 47.635 ;
    RECT 345.9 47.925 346.11 47.995 ;
    RECT 345.9 48.285 346.11 48.355 ;
    RECT 210.24 47.565 210.45 47.635 ;
    RECT 210.24 47.925 210.45 47.995 ;
    RECT 210.24 48.285 210.45 48.355 ;
    RECT 209.78 47.565 209.99 47.635 ;
    RECT 209.78 47.925 209.99 47.995 ;
    RECT 209.78 48.285 209.99 48.355 ;
    RECT 343.04 47.565 343.25 47.635 ;
    RECT 343.04 47.925 343.25 47.995 ;
    RECT 343.04 48.285 343.25 48.355 ;
    RECT 342.58 47.565 342.79 47.635 ;
    RECT 342.58 47.925 342.79 47.995 ;
    RECT 342.58 48.285 342.79 48.355 ;
    RECT 206.92 47.565 207.13 47.635 ;
    RECT 206.92 47.925 207.13 47.995 ;
    RECT 206.92 48.285 207.13 48.355 ;
    RECT 206.46 47.565 206.67 47.635 ;
    RECT 206.46 47.925 206.67 47.995 ;
    RECT 206.46 48.285 206.67 48.355 ;
    RECT 339.72 47.565 339.93 47.635 ;
    RECT 339.72 47.925 339.93 47.995 ;
    RECT 339.72 48.285 339.93 48.355 ;
    RECT 339.26 47.565 339.47 47.635 ;
    RECT 339.26 47.925 339.47 47.995 ;
    RECT 339.26 48.285 339.47 48.355 ;
    RECT 203.6 47.565 203.81 47.635 ;
    RECT 203.6 47.925 203.81 47.995 ;
    RECT 203.6 48.285 203.81 48.355 ;
    RECT 203.14 47.565 203.35 47.635 ;
    RECT 203.14 47.925 203.35 47.995 ;
    RECT 203.14 48.285 203.35 48.355 ;
    RECT 336.4 47.565 336.61 47.635 ;
    RECT 336.4 47.925 336.61 47.995 ;
    RECT 336.4 48.285 336.61 48.355 ;
    RECT 335.94 47.565 336.15 47.635 ;
    RECT 335.94 47.925 336.15 47.995 ;
    RECT 335.94 48.285 336.15 48.355 ;
    RECT 266.68 47.565 266.89 47.635 ;
    RECT 266.68 47.925 266.89 47.995 ;
    RECT 266.68 48.285 266.89 48.355 ;
    RECT 266.22 47.565 266.43 47.635 ;
    RECT 266.22 47.925 266.43 47.995 ;
    RECT 266.22 48.285 266.43 48.355 ;
    RECT 263.36 47.565 263.57 47.635 ;
    RECT 263.36 47.925 263.57 47.995 ;
    RECT 263.36 48.285 263.57 48.355 ;
    RECT 262.9 47.565 263.11 47.635 ;
    RECT 262.9 47.925 263.11 47.995 ;
    RECT 262.9 48.285 263.11 48.355 ;
    RECT 260.04 47.565 260.25 47.635 ;
    RECT 260.04 47.925 260.25 47.995 ;
    RECT 260.04 48.285 260.25 48.355 ;
    RECT 259.58 47.565 259.79 47.635 ;
    RECT 259.58 47.925 259.79 47.995 ;
    RECT 259.58 48.285 259.79 48.355 ;
    RECT 256.72 47.565 256.93 47.635 ;
    RECT 256.72 47.925 256.93 47.995 ;
    RECT 256.72 48.285 256.93 48.355 ;
    RECT 256.26 47.565 256.47 47.635 ;
    RECT 256.26 47.925 256.47 47.995 ;
    RECT 256.26 48.285 256.47 48.355 ;
    RECT 253.4 47.565 253.61 47.635 ;
    RECT 253.4 47.925 253.61 47.995 ;
    RECT 253.4 48.285 253.61 48.355 ;
    RECT 252.94 47.565 253.15 47.635 ;
    RECT 252.94 47.925 253.15 47.995 ;
    RECT 252.94 48.285 253.15 48.355 ;
    RECT 250.08 47.565 250.29 47.635 ;
    RECT 250.08 47.925 250.29 47.995 ;
    RECT 250.08 48.285 250.29 48.355 ;
    RECT 249.62 47.565 249.83 47.635 ;
    RECT 249.62 47.925 249.83 47.995 ;
    RECT 249.62 48.285 249.83 48.355 ;
    RECT 246.76 47.565 246.97 47.635 ;
    RECT 246.76 47.925 246.97 47.995 ;
    RECT 246.76 48.285 246.97 48.355 ;
    RECT 246.3 47.565 246.51 47.635 ;
    RECT 246.3 47.925 246.51 47.995 ;
    RECT 246.3 48.285 246.51 48.355 ;
    RECT 243.44 47.565 243.65 47.635 ;
    RECT 243.44 47.925 243.65 47.995 ;
    RECT 243.44 48.285 243.65 48.355 ;
    RECT 242.98 47.565 243.19 47.635 ;
    RECT 242.98 47.925 243.19 47.995 ;
    RECT 242.98 48.285 243.19 48.355 ;
    RECT 240.12 47.565 240.33 47.635 ;
    RECT 240.12 47.925 240.33 47.995 ;
    RECT 240.12 48.285 240.33 48.355 ;
    RECT 239.66 47.565 239.87 47.635 ;
    RECT 239.66 47.925 239.87 47.995 ;
    RECT 239.66 48.285 239.87 48.355 ;
    RECT 236.8 47.565 237.01 47.635 ;
    RECT 236.8 47.925 237.01 47.995 ;
    RECT 236.8 48.285 237.01 48.355 ;
    RECT 236.34 47.565 236.55 47.635 ;
    RECT 236.34 47.925 236.55 47.995 ;
    RECT 236.34 48.285 236.55 48.355 ;
    RECT 374.15 47.925 374.22 47.995 ;
    RECT 333.08 47.565 333.29 47.635 ;
    RECT 333.08 47.925 333.29 47.995 ;
    RECT 333.08 48.285 333.29 48.355 ;
    RECT 332.62 47.565 332.83 47.635 ;
    RECT 332.62 47.925 332.83 47.995 ;
    RECT 332.62 48.285 332.83 48.355 ;
    RECT 329.76 47.565 329.97 47.635 ;
    RECT 329.76 47.925 329.97 47.995 ;
    RECT 329.76 48.285 329.97 48.355 ;
    RECT 329.3 47.565 329.51 47.635 ;
    RECT 329.3 47.925 329.51 47.995 ;
    RECT 329.3 48.285 329.51 48.355 ;
    RECT 326.44 47.565 326.65 47.635 ;
    RECT 326.44 47.925 326.65 47.995 ;
    RECT 326.44 48.285 326.65 48.355 ;
    RECT 325.98 47.565 326.19 47.635 ;
    RECT 325.98 47.925 326.19 47.995 ;
    RECT 325.98 48.285 326.19 48.355 ;
    RECT 323.12 47.565 323.33 47.635 ;
    RECT 323.12 47.925 323.33 47.995 ;
    RECT 323.12 48.285 323.33 48.355 ;
    RECT 322.66 47.565 322.87 47.635 ;
    RECT 322.66 47.925 322.87 47.995 ;
    RECT 322.66 48.285 322.87 48.355 ;
    RECT 319.8 47.565 320.01 47.635 ;
    RECT 319.8 47.925 320.01 47.995 ;
    RECT 319.8 48.285 320.01 48.355 ;
    RECT 319.34 47.565 319.55 47.635 ;
    RECT 319.34 47.925 319.55 47.995 ;
    RECT 319.34 48.285 319.55 48.355 ;
    RECT 316.48 47.565 316.69 47.635 ;
    RECT 316.48 47.925 316.69 47.995 ;
    RECT 316.48 48.285 316.69 48.355 ;
    RECT 316.02 47.565 316.23 47.635 ;
    RECT 316.02 47.925 316.23 47.995 ;
    RECT 316.02 48.285 316.23 48.355 ;
    RECT 313.16 47.565 313.37 47.635 ;
    RECT 313.16 47.925 313.37 47.995 ;
    RECT 313.16 48.285 313.37 48.355 ;
    RECT 312.7 47.565 312.91 47.635 ;
    RECT 312.7 47.925 312.91 47.995 ;
    RECT 312.7 48.285 312.91 48.355 ;
    RECT 309.84 47.565 310.05 47.635 ;
    RECT 309.84 47.925 310.05 47.995 ;
    RECT 309.84 48.285 310.05 48.355 ;
    RECT 309.38 47.565 309.59 47.635 ;
    RECT 309.38 47.925 309.59 47.995 ;
    RECT 309.38 48.285 309.59 48.355 ;
    RECT 306.52 47.565 306.73 47.635 ;
    RECT 306.52 47.925 306.73 47.995 ;
    RECT 306.52 48.285 306.73 48.355 ;
    RECT 306.06 47.565 306.27 47.635 ;
    RECT 306.06 47.925 306.27 47.995 ;
    RECT 306.06 48.285 306.27 48.355 ;
    RECT 303.2 46.845 303.41 46.915 ;
    RECT 303.2 47.205 303.41 47.275 ;
    RECT 303.2 47.565 303.41 47.635 ;
    RECT 302.74 46.845 302.95 46.915 ;
    RECT 302.74 47.205 302.95 47.275 ;
    RECT 302.74 47.565 302.95 47.635 ;
    RECT 372.92 46.845 373.13 46.915 ;
    RECT 372.92 47.205 373.13 47.275 ;
    RECT 372.92 47.565 373.13 47.635 ;
    RECT 372.46 46.845 372.67 46.915 ;
    RECT 372.46 47.205 372.67 47.275 ;
    RECT 372.46 47.565 372.67 47.635 ;
    RECT 369.6 46.845 369.81 46.915 ;
    RECT 369.6 47.205 369.81 47.275 ;
    RECT 369.6 47.565 369.81 47.635 ;
    RECT 369.14 46.845 369.35 46.915 ;
    RECT 369.14 47.205 369.35 47.275 ;
    RECT 369.14 47.565 369.35 47.635 ;
    RECT 200.605 47.205 200.675 47.275 ;
    RECT 299.88 46.845 300.09 46.915 ;
    RECT 299.88 47.205 300.09 47.275 ;
    RECT 299.88 47.565 300.09 47.635 ;
    RECT 299.42 46.845 299.63 46.915 ;
    RECT 299.42 47.205 299.63 47.275 ;
    RECT 299.42 47.565 299.63 47.635 ;
    RECT 296.56 46.845 296.77 46.915 ;
    RECT 296.56 47.205 296.77 47.275 ;
    RECT 296.56 47.565 296.77 47.635 ;
    RECT 296.1 46.845 296.31 46.915 ;
    RECT 296.1 47.205 296.31 47.275 ;
    RECT 296.1 47.565 296.31 47.635 ;
    RECT 293.24 46.845 293.45 46.915 ;
    RECT 293.24 47.205 293.45 47.275 ;
    RECT 293.24 47.565 293.45 47.635 ;
    RECT 292.78 46.845 292.99 46.915 ;
    RECT 292.78 47.205 292.99 47.275 ;
    RECT 292.78 47.565 292.99 47.635 ;
    RECT 289.92 46.845 290.13 46.915 ;
    RECT 289.92 47.205 290.13 47.275 ;
    RECT 289.92 47.565 290.13 47.635 ;
    RECT 289.46 46.845 289.67 46.915 ;
    RECT 289.46 47.205 289.67 47.275 ;
    RECT 289.46 47.565 289.67 47.635 ;
    RECT 286.6 46.845 286.81 46.915 ;
    RECT 286.6 47.205 286.81 47.275 ;
    RECT 286.6 47.565 286.81 47.635 ;
    RECT 286.14 46.845 286.35 46.915 ;
    RECT 286.14 47.205 286.35 47.275 ;
    RECT 286.14 47.565 286.35 47.635 ;
    RECT 283.28 46.845 283.49 46.915 ;
    RECT 283.28 47.205 283.49 47.275 ;
    RECT 283.28 47.565 283.49 47.635 ;
    RECT 282.82 46.845 283.03 46.915 ;
    RECT 282.82 47.205 283.03 47.275 ;
    RECT 282.82 47.565 283.03 47.635 ;
    RECT 279.96 46.845 280.17 46.915 ;
    RECT 279.96 47.205 280.17 47.275 ;
    RECT 279.96 47.565 280.17 47.635 ;
    RECT 279.5 46.845 279.71 46.915 ;
    RECT 279.5 47.205 279.71 47.275 ;
    RECT 279.5 47.565 279.71 47.635 ;
    RECT 276.64 46.845 276.85 46.915 ;
    RECT 276.64 47.205 276.85 47.275 ;
    RECT 276.64 47.565 276.85 47.635 ;
    RECT 276.18 46.845 276.39 46.915 ;
    RECT 276.18 47.205 276.39 47.275 ;
    RECT 276.18 47.565 276.39 47.635 ;
    RECT 273.32 46.845 273.53 46.915 ;
    RECT 273.32 47.205 273.53 47.275 ;
    RECT 273.32 47.565 273.53 47.635 ;
    RECT 272.86 46.845 273.07 46.915 ;
    RECT 272.86 47.205 273.07 47.275 ;
    RECT 272.86 47.565 273.07 47.635 ;
    RECT 270.0 46.845 270.21 46.915 ;
    RECT 270.0 47.205 270.21 47.275 ;
    RECT 270.0 47.565 270.21 47.635 ;
    RECT 269.54 46.845 269.75 46.915 ;
    RECT 269.54 47.205 269.75 47.275 ;
    RECT 269.54 47.565 269.75 47.635 ;
    RECT 233.48 46.845 233.69 46.915 ;
    RECT 233.48 47.205 233.69 47.275 ;
    RECT 233.48 47.565 233.69 47.635 ;
    RECT 233.02 46.845 233.23 46.915 ;
    RECT 233.02 47.205 233.23 47.275 ;
    RECT 233.02 47.565 233.23 47.635 ;
    RECT 230.16 46.845 230.37 46.915 ;
    RECT 230.16 47.205 230.37 47.275 ;
    RECT 230.16 47.565 230.37 47.635 ;
    RECT 229.7 46.845 229.91 46.915 ;
    RECT 229.7 47.205 229.91 47.275 ;
    RECT 229.7 47.565 229.91 47.635 ;
    RECT 366.28 46.845 366.49 46.915 ;
    RECT 366.28 47.205 366.49 47.275 ;
    RECT 366.28 47.565 366.49 47.635 ;
    RECT 365.82 46.845 366.03 46.915 ;
    RECT 365.82 47.205 366.03 47.275 ;
    RECT 365.82 47.565 366.03 47.635 ;
    RECT 226.84 46.845 227.05 46.915 ;
    RECT 226.84 47.205 227.05 47.275 ;
    RECT 226.84 47.565 227.05 47.635 ;
    RECT 226.38 46.845 226.59 46.915 ;
    RECT 226.38 47.205 226.59 47.275 ;
    RECT 226.38 47.565 226.59 47.635 ;
    RECT 362.96 46.845 363.17 46.915 ;
    RECT 362.96 47.205 363.17 47.275 ;
    RECT 362.96 47.565 363.17 47.635 ;
    RECT 362.5 46.845 362.71 46.915 ;
    RECT 362.5 47.205 362.71 47.275 ;
    RECT 362.5 47.565 362.71 47.635 ;
    RECT 223.52 46.845 223.73 46.915 ;
    RECT 223.52 47.205 223.73 47.275 ;
    RECT 223.52 47.565 223.73 47.635 ;
    RECT 223.06 46.845 223.27 46.915 ;
    RECT 223.06 47.205 223.27 47.275 ;
    RECT 223.06 47.565 223.27 47.635 ;
    RECT 359.64 46.845 359.85 46.915 ;
    RECT 359.64 47.205 359.85 47.275 ;
    RECT 359.64 47.565 359.85 47.635 ;
    RECT 359.18 46.845 359.39 46.915 ;
    RECT 359.18 47.205 359.39 47.275 ;
    RECT 359.18 47.565 359.39 47.635 ;
    RECT 220.2 46.845 220.41 46.915 ;
    RECT 220.2 47.205 220.41 47.275 ;
    RECT 220.2 47.565 220.41 47.635 ;
    RECT 219.74 46.845 219.95 46.915 ;
    RECT 219.74 47.205 219.95 47.275 ;
    RECT 219.74 47.565 219.95 47.635 ;
    RECT 356.32 46.845 356.53 46.915 ;
    RECT 356.32 47.205 356.53 47.275 ;
    RECT 356.32 47.565 356.53 47.635 ;
    RECT 355.86 46.845 356.07 46.915 ;
    RECT 355.86 47.205 356.07 47.275 ;
    RECT 355.86 47.565 356.07 47.635 ;
    RECT 353.0 46.845 353.21 46.915 ;
    RECT 353.0 47.205 353.21 47.275 ;
    RECT 353.0 47.565 353.21 47.635 ;
    RECT 352.54 46.845 352.75 46.915 ;
    RECT 352.54 47.205 352.75 47.275 ;
    RECT 352.54 47.565 352.75 47.635 ;
    RECT 216.88 46.845 217.09 46.915 ;
    RECT 216.88 47.205 217.09 47.275 ;
    RECT 216.88 47.565 217.09 47.635 ;
    RECT 216.42 46.845 216.63 46.915 ;
    RECT 216.42 47.205 216.63 47.275 ;
    RECT 216.42 47.565 216.63 47.635 ;
    RECT 349.68 46.845 349.89 46.915 ;
    RECT 349.68 47.205 349.89 47.275 ;
    RECT 349.68 47.565 349.89 47.635 ;
    RECT 349.22 46.845 349.43 46.915 ;
    RECT 349.22 47.205 349.43 47.275 ;
    RECT 349.22 47.565 349.43 47.635 ;
    RECT 213.56 46.845 213.77 46.915 ;
    RECT 213.56 47.205 213.77 47.275 ;
    RECT 213.56 47.565 213.77 47.635 ;
    RECT 213.1 46.845 213.31 46.915 ;
    RECT 213.1 47.205 213.31 47.275 ;
    RECT 213.1 47.565 213.31 47.635 ;
    RECT 346.36 46.845 346.57 46.915 ;
    RECT 346.36 47.205 346.57 47.275 ;
    RECT 346.36 47.565 346.57 47.635 ;
    RECT 345.9 46.845 346.11 46.915 ;
    RECT 345.9 47.205 346.11 47.275 ;
    RECT 345.9 47.565 346.11 47.635 ;
    RECT 210.24 46.845 210.45 46.915 ;
    RECT 210.24 47.205 210.45 47.275 ;
    RECT 210.24 47.565 210.45 47.635 ;
    RECT 209.78 46.845 209.99 46.915 ;
    RECT 209.78 47.205 209.99 47.275 ;
    RECT 209.78 47.565 209.99 47.635 ;
    RECT 343.04 46.845 343.25 46.915 ;
    RECT 343.04 47.205 343.25 47.275 ;
    RECT 343.04 47.565 343.25 47.635 ;
    RECT 342.58 46.845 342.79 46.915 ;
    RECT 342.58 47.205 342.79 47.275 ;
    RECT 342.58 47.565 342.79 47.635 ;
    RECT 206.92 46.845 207.13 46.915 ;
    RECT 206.92 47.205 207.13 47.275 ;
    RECT 206.92 47.565 207.13 47.635 ;
    RECT 206.46 46.845 206.67 46.915 ;
    RECT 206.46 47.205 206.67 47.275 ;
    RECT 206.46 47.565 206.67 47.635 ;
    RECT 339.72 46.845 339.93 46.915 ;
    RECT 339.72 47.205 339.93 47.275 ;
    RECT 339.72 47.565 339.93 47.635 ;
    RECT 339.26 46.845 339.47 46.915 ;
    RECT 339.26 47.205 339.47 47.275 ;
    RECT 339.26 47.565 339.47 47.635 ;
    RECT 203.6 46.845 203.81 46.915 ;
    RECT 203.6 47.205 203.81 47.275 ;
    RECT 203.6 47.565 203.81 47.635 ;
    RECT 203.14 46.845 203.35 46.915 ;
    RECT 203.14 47.205 203.35 47.275 ;
    RECT 203.14 47.565 203.35 47.635 ;
    RECT 336.4 46.845 336.61 46.915 ;
    RECT 336.4 47.205 336.61 47.275 ;
    RECT 336.4 47.565 336.61 47.635 ;
    RECT 335.94 46.845 336.15 46.915 ;
    RECT 335.94 47.205 336.15 47.275 ;
    RECT 335.94 47.565 336.15 47.635 ;
    RECT 266.68 46.845 266.89 46.915 ;
    RECT 266.68 47.205 266.89 47.275 ;
    RECT 266.68 47.565 266.89 47.635 ;
    RECT 266.22 46.845 266.43 46.915 ;
    RECT 266.22 47.205 266.43 47.275 ;
    RECT 266.22 47.565 266.43 47.635 ;
    RECT 263.36 46.845 263.57 46.915 ;
    RECT 263.36 47.205 263.57 47.275 ;
    RECT 263.36 47.565 263.57 47.635 ;
    RECT 262.9 46.845 263.11 46.915 ;
    RECT 262.9 47.205 263.11 47.275 ;
    RECT 262.9 47.565 263.11 47.635 ;
    RECT 260.04 46.845 260.25 46.915 ;
    RECT 260.04 47.205 260.25 47.275 ;
    RECT 260.04 47.565 260.25 47.635 ;
    RECT 259.58 46.845 259.79 46.915 ;
    RECT 259.58 47.205 259.79 47.275 ;
    RECT 259.58 47.565 259.79 47.635 ;
    RECT 256.72 46.845 256.93 46.915 ;
    RECT 256.72 47.205 256.93 47.275 ;
    RECT 256.72 47.565 256.93 47.635 ;
    RECT 256.26 46.845 256.47 46.915 ;
    RECT 256.26 47.205 256.47 47.275 ;
    RECT 256.26 47.565 256.47 47.635 ;
    RECT 253.4 46.845 253.61 46.915 ;
    RECT 253.4 47.205 253.61 47.275 ;
    RECT 253.4 47.565 253.61 47.635 ;
    RECT 252.94 46.845 253.15 46.915 ;
    RECT 252.94 47.205 253.15 47.275 ;
    RECT 252.94 47.565 253.15 47.635 ;
    RECT 250.08 46.845 250.29 46.915 ;
    RECT 250.08 47.205 250.29 47.275 ;
    RECT 250.08 47.565 250.29 47.635 ;
    RECT 249.62 46.845 249.83 46.915 ;
    RECT 249.62 47.205 249.83 47.275 ;
    RECT 249.62 47.565 249.83 47.635 ;
    RECT 246.76 46.845 246.97 46.915 ;
    RECT 246.76 47.205 246.97 47.275 ;
    RECT 246.76 47.565 246.97 47.635 ;
    RECT 246.3 46.845 246.51 46.915 ;
    RECT 246.3 47.205 246.51 47.275 ;
    RECT 246.3 47.565 246.51 47.635 ;
    RECT 243.44 46.845 243.65 46.915 ;
    RECT 243.44 47.205 243.65 47.275 ;
    RECT 243.44 47.565 243.65 47.635 ;
    RECT 242.98 46.845 243.19 46.915 ;
    RECT 242.98 47.205 243.19 47.275 ;
    RECT 242.98 47.565 243.19 47.635 ;
    RECT 240.12 46.845 240.33 46.915 ;
    RECT 240.12 47.205 240.33 47.275 ;
    RECT 240.12 47.565 240.33 47.635 ;
    RECT 239.66 46.845 239.87 46.915 ;
    RECT 239.66 47.205 239.87 47.275 ;
    RECT 239.66 47.565 239.87 47.635 ;
    RECT 236.8 46.845 237.01 46.915 ;
    RECT 236.8 47.205 237.01 47.275 ;
    RECT 236.8 47.565 237.01 47.635 ;
    RECT 236.34 46.845 236.55 46.915 ;
    RECT 236.34 47.205 236.55 47.275 ;
    RECT 236.34 47.565 236.55 47.635 ;
    RECT 374.15 47.205 374.22 47.275 ;
    RECT 333.08 46.845 333.29 46.915 ;
    RECT 333.08 47.205 333.29 47.275 ;
    RECT 333.08 47.565 333.29 47.635 ;
    RECT 332.62 46.845 332.83 46.915 ;
    RECT 332.62 47.205 332.83 47.275 ;
    RECT 332.62 47.565 332.83 47.635 ;
    RECT 329.76 46.845 329.97 46.915 ;
    RECT 329.76 47.205 329.97 47.275 ;
    RECT 329.76 47.565 329.97 47.635 ;
    RECT 329.3 46.845 329.51 46.915 ;
    RECT 329.3 47.205 329.51 47.275 ;
    RECT 329.3 47.565 329.51 47.635 ;
    RECT 326.44 46.845 326.65 46.915 ;
    RECT 326.44 47.205 326.65 47.275 ;
    RECT 326.44 47.565 326.65 47.635 ;
    RECT 325.98 46.845 326.19 46.915 ;
    RECT 325.98 47.205 326.19 47.275 ;
    RECT 325.98 47.565 326.19 47.635 ;
    RECT 323.12 46.845 323.33 46.915 ;
    RECT 323.12 47.205 323.33 47.275 ;
    RECT 323.12 47.565 323.33 47.635 ;
    RECT 322.66 46.845 322.87 46.915 ;
    RECT 322.66 47.205 322.87 47.275 ;
    RECT 322.66 47.565 322.87 47.635 ;
    RECT 319.8 46.845 320.01 46.915 ;
    RECT 319.8 47.205 320.01 47.275 ;
    RECT 319.8 47.565 320.01 47.635 ;
    RECT 319.34 46.845 319.55 46.915 ;
    RECT 319.34 47.205 319.55 47.275 ;
    RECT 319.34 47.565 319.55 47.635 ;
    RECT 316.48 46.845 316.69 46.915 ;
    RECT 316.48 47.205 316.69 47.275 ;
    RECT 316.48 47.565 316.69 47.635 ;
    RECT 316.02 46.845 316.23 46.915 ;
    RECT 316.02 47.205 316.23 47.275 ;
    RECT 316.02 47.565 316.23 47.635 ;
    RECT 313.16 46.845 313.37 46.915 ;
    RECT 313.16 47.205 313.37 47.275 ;
    RECT 313.16 47.565 313.37 47.635 ;
    RECT 312.7 46.845 312.91 46.915 ;
    RECT 312.7 47.205 312.91 47.275 ;
    RECT 312.7 47.565 312.91 47.635 ;
    RECT 309.84 46.845 310.05 46.915 ;
    RECT 309.84 47.205 310.05 47.275 ;
    RECT 309.84 47.565 310.05 47.635 ;
    RECT 309.38 46.845 309.59 46.915 ;
    RECT 309.38 47.205 309.59 47.275 ;
    RECT 309.38 47.565 309.59 47.635 ;
    RECT 306.52 46.845 306.73 46.915 ;
    RECT 306.52 47.205 306.73 47.275 ;
    RECT 306.52 47.565 306.73 47.635 ;
    RECT 306.06 46.845 306.27 46.915 ;
    RECT 306.06 47.205 306.27 47.275 ;
    RECT 306.06 47.565 306.27 47.635 ;
    RECT 303.2 46.125 303.41 46.195 ;
    RECT 303.2 46.485 303.41 46.555 ;
    RECT 303.2 46.845 303.41 46.915 ;
    RECT 302.74 46.125 302.95 46.195 ;
    RECT 302.74 46.485 302.95 46.555 ;
    RECT 302.74 46.845 302.95 46.915 ;
    RECT 372.92 46.125 373.13 46.195 ;
    RECT 372.92 46.485 373.13 46.555 ;
    RECT 372.92 46.845 373.13 46.915 ;
    RECT 372.46 46.125 372.67 46.195 ;
    RECT 372.46 46.485 372.67 46.555 ;
    RECT 372.46 46.845 372.67 46.915 ;
    RECT 369.6 46.125 369.81 46.195 ;
    RECT 369.6 46.485 369.81 46.555 ;
    RECT 369.6 46.845 369.81 46.915 ;
    RECT 369.14 46.125 369.35 46.195 ;
    RECT 369.14 46.485 369.35 46.555 ;
    RECT 369.14 46.845 369.35 46.915 ;
    RECT 200.605 46.485 200.675 46.555 ;
    RECT 299.88 46.125 300.09 46.195 ;
    RECT 299.88 46.485 300.09 46.555 ;
    RECT 299.88 46.845 300.09 46.915 ;
    RECT 299.42 46.125 299.63 46.195 ;
    RECT 299.42 46.485 299.63 46.555 ;
    RECT 299.42 46.845 299.63 46.915 ;
    RECT 296.56 46.125 296.77 46.195 ;
    RECT 296.56 46.485 296.77 46.555 ;
    RECT 296.56 46.845 296.77 46.915 ;
    RECT 296.1 46.125 296.31 46.195 ;
    RECT 296.1 46.485 296.31 46.555 ;
    RECT 296.1 46.845 296.31 46.915 ;
    RECT 293.24 46.125 293.45 46.195 ;
    RECT 293.24 46.485 293.45 46.555 ;
    RECT 293.24 46.845 293.45 46.915 ;
    RECT 292.78 46.125 292.99 46.195 ;
    RECT 292.78 46.485 292.99 46.555 ;
    RECT 292.78 46.845 292.99 46.915 ;
    RECT 289.92 46.125 290.13 46.195 ;
    RECT 289.92 46.485 290.13 46.555 ;
    RECT 289.92 46.845 290.13 46.915 ;
    RECT 289.46 46.125 289.67 46.195 ;
    RECT 289.46 46.485 289.67 46.555 ;
    RECT 289.46 46.845 289.67 46.915 ;
    RECT 286.6 46.125 286.81 46.195 ;
    RECT 286.6 46.485 286.81 46.555 ;
    RECT 286.6 46.845 286.81 46.915 ;
    RECT 286.14 46.125 286.35 46.195 ;
    RECT 286.14 46.485 286.35 46.555 ;
    RECT 286.14 46.845 286.35 46.915 ;
    RECT 283.28 46.125 283.49 46.195 ;
    RECT 283.28 46.485 283.49 46.555 ;
    RECT 283.28 46.845 283.49 46.915 ;
    RECT 282.82 46.125 283.03 46.195 ;
    RECT 282.82 46.485 283.03 46.555 ;
    RECT 282.82 46.845 283.03 46.915 ;
    RECT 279.96 46.125 280.17 46.195 ;
    RECT 279.96 46.485 280.17 46.555 ;
    RECT 279.96 46.845 280.17 46.915 ;
    RECT 279.5 46.125 279.71 46.195 ;
    RECT 279.5 46.485 279.71 46.555 ;
    RECT 279.5 46.845 279.71 46.915 ;
    RECT 276.64 46.125 276.85 46.195 ;
    RECT 276.64 46.485 276.85 46.555 ;
    RECT 276.64 46.845 276.85 46.915 ;
    RECT 276.18 46.125 276.39 46.195 ;
    RECT 276.18 46.485 276.39 46.555 ;
    RECT 276.18 46.845 276.39 46.915 ;
    RECT 273.32 46.125 273.53 46.195 ;
    RECT 273.32 46.485 273.53 46.555 ;
    RECT 273.32 46.845 273.53 46.915 ;
    RECT 272.86 46.125 273.07 46.195 ;
    RECT 272.86 46.485 273.07 46.555 ;
    RECT 272.86 46.845 273.07 46.915 ;
    RECT 270.0 46.125 270.21 46.195 ;
    RECT 270.0 46.485 270.21 46.555 ;
    RECT 270.0 46.845 270.21 46.915 ;
    RECT 269.54 46.125 269.75 46.195 ;
    RECT 269.54 46.485 269.75 46.555 ;
    RECT 269.54 46.845 269.75 46.915 ;
    RECT 233.48 46.125 233.69 46.195 ;
    RECT 233.48 46.485 233.69 46.555 ;
    RECT 233.48 46.845 233.69 46.915 ;
    RECT 233.02 46.125 233.23 46.195 ;
    RECT 233.02 46.485 233.23 46.555 ;
    RECT 233.02 46.845 233.23 46.915 ;
    RECT 230.16 46.125 230.37 46.195 ;
    RECT 230.16 46.485 230.37 46.555 ;
    RECT 230.16 46.845 230.37 46.915 ;
    RECT 229.7 46.125 229.91 46.195 ;
    RECT 229.7 46.485 229.91 46.555 ;
    RECT 229.7 46.845 229.91 46.915 ;
    RECT 366.28 46.125 366.49 46.195 ;
    RECT 366.28 46.485 366.49 46.555 ;
    RECT 366.28 46.845 366.49 46.915 ;
    RECT 365.82 46.125 366.03 46.195 ;
    RECT 365.82 46.485 366.03 46.555 ;
    RECT 365.82 46.845 366.03 46.915 ;
    RECT 226.84 46.125 227.05 46.195 ;
    RECT 226.84 46.485 227.05 46.555 ;
    RECT 226.84 46.845 227.05 46.915 ;
    RECT 226.38 46.125 226.59 46.195 ;
    RECT 226.38 46.485 226.59 46.555 ;
    RECT 226.38 46.845 226.59 46.915 ;
    RECT 362.96 46.125 363.17 46.195 ;
    RECT 362.96 46.485 363.17 46.555 ;
    RECT 362.96 46.845 363.17 46.915 ;
    RECT 362.5 46.125 362.71 46.195 ;
    RECT 362.5 46.485 362.71 46.555 ;
    RECT 362.5 46.845 362.71 46.915 ;
    RECT 223.52 46.125 223.73 46.195 ;
    RECT 223.52 46.485 223.73 46.555 ;
    RECT 223.52 46.845 223.73 46.915 ;
    RECT 223.06 46.125 223.27 46.195 ;
    RECT 223.06 46.485 223.27 46.555 ;
    RECT 223.06 46.845 223.27 46.915 ;
    RECT 359.64 46.125 359.85 46.195 ;
    RECT 359.64 46.485 359.85 46.555 ;
    RECT 359.64 46.845 359.85 46.915 ;
    RECT 359.18 46.125 359.39 46.195 ;
    RECT 359.18 46.485 359.39 46.555 ;
    RECT 359.18 46.845 359.39 46.915 ;
    RECT 220.2 46.125 220.41 46.195 ;
    RECT 220.2 46.485 220.41 46.555 ;
    RECT 220.2 46.845 220.41 46.915 ;
    RECT 219.74 46.125 219.95 46.195 ;
    RECT 219.74 46.485 219.95 46.555 ;
    RECT 219.74 46.845 219.95 46.915 ;
    RECT 356.32 46.125 356.53 46.195 ;
    RECT 356.32 46.485 356.53 46.555 ;
    RECT 356.32 46.845 356.53 46.915 ;
    RECT 355.86 46.125 356.07 46.195 ;
    RECT 355.86 46.485 356.07 46.555 ;
    RECT 355.86 46.845 356.07 46.915 ;
    RECT 353.0 46.125 353.21 46.195 ;
    RECT 353.0 46.485 353.21 46.555 ;
    RECT 353.0 46.845 353.21 46.915 ;
    RECT 352.54 46.125 352.75 46.195 ;
    RECT 352.54 46.485 352.75 46.555 ;
    RECT 352.54 46.845 352.75 46.915 ;
    RECT 216.88 46.125 217.09 46.195 ;
    RECT 216.88 46.485 217.09 46.555 ;
    RECT 216.88 46.845 217.09 46.915 ;
    RECT 216.42 46.125 216.63 46.195 ;
    RECT 216.42 46.485 216.63 46.555 ;
    RECT 216.42 46.845 216.63 46.915 ;
    RECT 349.68 46.125 349.89 46.195 ;
    RECT 349.68 46.485 349.89 46.555 ;
    RECT 349.68 46.845 349.89 46.915 ;
    RECT 349.22 46.125 349.43 46.195 ;
    RECT 349.22 46.485 349.43 46.555 ;
    RECT 349.22 46.845 349.43 46.915 ;
    RECT 213.56 46.125 213.77 46.195 ;
    RECT 213.56 46.485 213.77 46.555 ;
    RECT 213.56 46.845 213.77 46.915 ;
    RECT 213.1 46.125 213.31 46.195 ;
    RECT 213.1 46.485 213.31 46.555 ;
    RECT 213.1 46.845 213.31 46.915 ;
    RECT 346.36 46.125 346.57 46.195 ;
    RECT 346.36 46.485 346.57 46.555 ;
    RECT 346.36 46.845 346.57 46.915 ;
    RECT 345.9 46.125 346.11 46.195 ;
    RECT 345.9 46.485 346.11 46.555 ;
    RECT 345.9 46.845 346.11 46.915 ;
    RECT 210.24 46.125 210.45 46.195 ;
    RECT 210.24 46.485 210.45 46.555 ;
    RECT 210.24 46.845 210.45 46.915 ;
    RECT 209.78 46.125 209.99 46.195 ;
    RECT 209.78 46.485 209.99 46.555 ;
    RECT 209.78 46.845 209.99 46.915 ;
    RECT 343.04 46.125 343.25 46.195 ;
    RECT 343.04 46.485 343.25 46.555 ;
    RECT 343.04 46.845 343.25 46.915 ;
    RECT 342.58 46.125 342.79 46.195 ;
    RECT 342.58 46.485 342.79 46.555 ;
    RECT 342.58 46.845 342.79 46.915 ;
    RECT 206.92 46.125 207.13 46.195 ;
    RECT 206.92 46.485 207.13 46.555 ;
    RECT 206.92 46.845 207.13 46.915 ;
    RECT 206.46 46.125 206.67 46.195 ;
    RECT 206.46 46.485 206.67 46.555 ;
    RECT 206.46 46.845 206.67 46.915 ;
    RECT 339.72 46.125 339.93 46.195 ;
    RECT 339.72 46.485 339.93 46.555 ;
    RECT 339.72 46.845 339.93 46.915 ;
    RECT 339.26 46.125 339.47 46.195 ;
    RECT 339.26 46.485 339.47 46.555 ;
    RECT 339.26 46.845 339.47 46.915 ;
    RECT 203.6 46.125 203.81 46.195 ;
    RECT 203.6 46.485 203.81 46.555 ;
    RECT 203.6 46.845 203.81 46.915 ;
    RECT 203.14 46.125 203.35 46.195 ;
    RECT 203.14 46.485 203.35 46.555 ;
    RECT 203.14 46.845 203.35 46.915 ;
    RECT 336.4 46.125 336.61 46.195 ;
    RECT 336.4 46.485 336.61 46.555 ;
    RECT 336.4 46.845 336.61 46.915 ;
    RECT 335.94 46.125 336.15 46.195 ;
    RECT 335.94 46.485 336.15 46.555 ;
    RECT 335.94 46.845 336.15 46.915 ;
    RECT 266.68 46.125 266.89 46.195 ;
    RECT 266.68 46.485 266.89 46.555 ;
    RECT 266.68 46.845 266.89 46.915 ;
    RECT 266.22 46.125 266.43 46.195 ;
    RECT 266.22 46.485 266.43 46.555 ;
    RECT 266.22 46.845 266.43 46.915 ;
    RECT 263.36 46.125 263.57 46.195 ;
    RECT 263.36 46.485 263.57 46.555 ;
    RECT 263.36 46.845 263.57 46.915 ;
    RECT 262.9 46.125 263.11 46.195 ;
    RECT 262.9 46.485 263.11 46.555 ;
    RECT 262.9 46.845 263.11 46.915 ;
    RECT 260.04 46.125 260.25 46.195 ;
    RECT 260.04 46.485 260.25 46.555 ;
    RECT 260.04 46.845 260.25 46.915 ;
    RECT 259.58 46.125 259.79 46.195 ;
    RECT 259.58 46.485 259.79 46.555 ;
    RECT 259.58 46.845 259.79 46.915 ;
    RECT 256.72 46.125 256.93 46.195 ;
    RECT 256.72 46.485 256.93 46.555 ;
    RECT 256.72 46.845 256.93 46.915 ;
    RECT 256.26 46.125 256.47 46.195 ;
    RECT 256.26 46.485 256.47 46.555 ;
    RECT 256.26 46.845 256.47 46.915 ;
    RECT 253.4 46.125 253.61 46.195 ;
    RECT 253.4 46.485 253.61 46.555 ;
    RECT 253.4 46.845 253.61 46.915 ;
    RECT 252.94 46.125 253.15 46.195 ;
    RECT 252.94 46.485 253.15 46.555 ;
    RECT 252.94 46.845 253.15 46.915 ;
    RECT 250.08 46.125 250.29 46.195 ;
    RECT 250.08 46.485 250.29 46.555 ;
    RECT 250.08 46.845 250.29 46.915 ;
    RECT 249.62 46.125 249.83 46.195 ;
    RECT 249.62 46.485 249.83 46.555 ;
    RECT 249.62 46.845 249.83 46.915 ;
    RECT 246.76 46.125 246.97 46.195 ;
    RECT 246.76 46.485 246.97 46.555 ;
    RECT 246.76 46.845 246.97 46.915 ;
    RECT 246.3 46.125 246.51 46.195 ;
    RECT 246.3 46.485 246.51 46.555 ;
    RECT 246.3 46.845 246.51 46.915 ;
    RECT 243.44 46.125 243.65 46.195 ;
    RECT 243.44 46.485 243.65 46.555 ;
    RECT 243.44 46.845 243.65 46.915 ;
    RECT 242.98 46.125 243.19 46.195 ;
    RECT 242.98 46.485 243.19 46.555 ;
    RECT 242.98 46.845 243.19 46.915 ;
    RECT 240.12 46.125 240.33 46.195 ;
    RECT 240.12 46.485 240.33 46.555 ;
    RECT 240.12 46.845 240.33 46.915 ;
    RECT 239.66 46.125 239.87 46.195 ;
    RECT 239.66 46.485 239.87 46.555 ;
    RECT 239.66 46.845 239.87 46.915 ;
    RECT 236.8 46.125 237.01 46.195 ;
    RECT 236.8 46.485 237.01 46.555 ;
    RECT 236.8 46.845 237.01 46.915 ;
    RECT 236.34 46.125 236.55 46.195 ;
    RECT 236.34 46.485 236.55 46.555 ;
    RECT 236.34 46.845 236.55 46.915 ;
    RECT 374.15 46.485 374.22 46.555 ;
    RECT 333.08 46.125 333.29 46.195 ;
    RECT 333.08 46.485 333.29 46.555 ;
    RECT 333.08 46.845 333.29 46.915 ;
    RECT 332.62 46.125 332.83 46.195 ;
    RECT 332.62 46.485 332.83 46.555 ;
    RECT 332.62 46.845 332.83 46.915 ;
    RECT 329.76 46.125 329.97 46.195 ;
    RECT 329.76 46.485 329.97 46.555 ;
    RECT 329.76 46.845 329.97 46.915 ;
    RECT 329.3 46.125 329.51 46.195 ;
    RECT 329.3 46.485 329.51 46.555 ;
    RECT 329.3 46.845 329.51 46.915 ;
    RECT 326.44 46.125 326.65 46.195 ;
    RECT 326.44 46.485 326.65 46.555 ;
    RECT 326.44 46.845 326.65 46.915 ;
    RECT 325.98 46.125 326.19 46.195 ;
    RECT 325.98 46.485 326.19 46.555 ;
    RECT 325.98 46.845 326.19 46.915 ;
    RECT 323.12 46.125 323.33 46.195 ;
    RECT 323.12 46.485 323.33 46.555 ;
    RECT 323.12 46.845 323.33 46.915 ;
    RECT 322.66 46.125 322.87 46.195 ;
    RECT 322.66 46.485 322.87 46.555 ;
    RECT 322.66 46.845 322.87 46.915 ;
    RECT 319.8 46.125 320.01 46.195 ;
    RECT 319.8 46.485 320.01 46.555 ;
    RECT 319.8 46.845 320.01 46.915 ;
    RECT 319.34 46.125 319.55 46.195 ;
    RECT 319.34 46.485 319.55 46.555 ;
    RECT 319.34 46.845 319.55 46.915 ;
    RECT 316.48 46.125 316.69 46.195 ;
    RECT 316.48 46.485 316.69 46.555 ;
    RECT 316.48 46.845 316.69 46.915 ;
    RECT 316.02 46.125 316.23 46.195 ;
    RECT 316.02 46.485 316.23 46.555 ;
    RECT 316.02 46.845 316.23 46.915 ;
    RECT 313.16 46.125 313.37 46.195 ;
    RECT 313.16 46.485 313.37 46.555 ;
    RECT 313.16 46.845 313.37 46.915 ;
    RECT 312.7 46.125 312.91 46.195 ;
    RECT 312.7 46.485 312.91 46.555 ;
    RECT 312.7 46.845 312.91 46.915 ;
    RECT 309.84 46.125 310.05 46.195 ;
    RECT 309.84 46.485 310.05 46.555 ;
    RECT 309.84 46.845 310.05 46.915 ;
    RECT 309.38 46.125 309.59 46.195 ;
    RECT 309.38 46.485 309.59 46.555 ;
    RECT 309.38 46.845 309.59 46.915 ;
    RECT 306.52 46.125 306.73 46.195 ;
    RECT 306.52 46.485 306.73 46.555 ;
    RECT 306.52 46.845 306.73 46.915 ;
    RECT 306.06 46.125 306.27 46.195 ;
    RECT 306.06 46.485 306.27 46.555 ;
    RECT 306.06 46.845 306.27 46.915 ;
    RECT 303.2 45.405 303.41 45.475 ;
    RECT 303.2 45.765 303.41 45.835 ;
    RECT 303.2 46.125 303.41 46.195 ;
    RECT 302.74 45.405 302.95 45.475 ;
    RECT 302.74 45.765 302.95 45.835 ;
    RECT 302.74 46.125 302.95 46.195 ;
    RECT 372.92 45.405 373.13 45.475 ;
    RECT 372.92 45.765 373.13 45.835 ;
    RECT 372.92 46.125 373.13 46.195 ;
    RECT 372.46 45.405 372.67 45.475 ;
    RECT 372.46 45.765 372.67 45.835 ;
    RECT 372.46 46.125 372.67 46.195 ;
    RECT 369.6 45.405 369.81 45.475 ;
    RECT 369.6 45.765 369.81 45.835 ;
    RECT 369.6 46.125 369.81 46.195 ;
    RECT 369.14 45.405 369.35 45.475 ;
    RECT 369.14 45.765 369.35 45.835 ;
    RECT 369.14 46.125 369.35 46.195 ;
    RECT 200.605 45.765 200.675 45.835 ;
    RECT 299.88 45.405 300.09 45.475 ;
    RECT 299.88 45.765 300.09 45.835 ;
    RECT 299.88 46.125 300.09 46.195 ;
    RECT 299.42 45.405 299.63 45.475 ;
    RECT 299.42 45.765 299.63 45.835 ;
    RECT 299.42 46.125 299.63 46.195 ;
    RECT 296.56 45.405 296.77 45.475 ;
    RECT 296.56 45.765 296.77 45.835 ;
    RECT 296.56 46.125 296.77 46.195 ;
    RECT 296.1 45.405 296.31 45.475 ;
    RECT 296.1 45.765 296.31 45.835 ;
    RECT 296.1 46.125 296.31 46.195 ;
    RECT 293.24 45.405 293.45 45.475 ;
    RECT 293.24 45.765 293.45 45.835 ;
    RECT 293.24 46.125 293.45 46.195 ;
    RECT 292.78 45.405 292.99 45.475 ;
    RECT 292.78 45.765 292.99 45.835 ;
    RECT 292.78 46.125 292.99 46.195 ;
    RECT 289.92 45.405 290.13 45.475 ;
    RECT 289.92 45.765 290.13 45.835 ;
    RECT 289.92 46.125 290.13 46.195 ;
    RECT 289.46 45.405 289.67 45.475 ;
    RECT 289.46 45.765 289.67 45.835 ;
    RECT 289.46 46.125 289.67 46.195 ;
    RECT 286.6 45.405 286.81 45.475 ;
    RECT 286.6 45.765 286.81 45.835 ;
    RECT 286.6 46.125 286.81 46.195 ;
    RECT 286.14 45.405 286.35 45.475 ;
    RECT 286.14 45.765 286.35 45.835 ;
    RECT 286.14 46.125 286.35 46.195 ;
    RECT 283.28 45.405 283.49 45.475 ;
    RECT 283.28 45.765 283.49 45.835 ;
    RECT 283.28 46.125 283.49 46.195 ;
    RECT 282.82 45.405 283.03 45.475 ;
    RECT 282.82 45.765 283.03 45.835 ;
    RECT 282.82 46.125 283.03 46.195 ;
    RECT 279.96 45.405 280.17 45.475 ;
    RECT 279.96 45.765 280.17 45.835 ;
    RECT 279.96 46.125 280.17 46.195 ;
    RECT 279.5 45.405 279.71 45.475 ;
    RECT 279.5 45.765 279.71 45.835 ;
    RECT 279.5 46.125 279.71 46.195 ;
    RECT 276.64 45.405 276.85 45.475 ;
    RECT 276.64 45.765 276.85 45.835 ;
    RECT 276.64 46.125 276.85 46.195 ;
    RECT 276.18 45.405 276.39 45.475 ;
    RECT 276.18 45.765 276.39 45.835 ;
    RECT 276.18 46.125 276.39 46.195 ;
    RECT 273.32 45.405 273.53 45.475 ;
    RECT 273.32 45.765 273.53 45.835 ;
    RECT 273.32 46.125 273.53 46.195 ;
    RECT 272.86 45.405 273.07 45.475 ;
    RECT 272.86 45.765 273.07 45.835 ;
    RECT 272.86 46.125 273.07 46.195 ;
    RECT 270.0 45.405 270.21 45.475 ;
    RECT 270.0 45.765 270.21 45.835 ;
    RECT 270.0 46.125 270.21 46.195 ;
    RECT 269.54 45.405 269.75 45.475 ;
    RECT 269.54 45.765 269.75 45.835 ;
    RECT 269.54 46.125 269.75 46.195 ;
    RECT 233.48 45.405 233.69 45.475 ;
    RECT 233.48 45.765 233.69 45.835 ;
    RECT 233.48 46.125 233.69 46.195 ;
    RECT 233.02 45.405 233.23 45.475 ;
    RECT 233.02 45.765 233.23 45.835 ;
    RECT 233.02 46.125 233.23 46.195 ;
    RECT 230.16 45.405 230.37 45.475 ;
    RECT 230.16 45.765 230.37 45.835 ;
    RECT 230.16 46.125 230.37 46.195 ;
    RECT 229.7 45.405 229.91 45.475 ;
    RECT 229.7 45.765 229.91 45.835 ;
    RECT 229.7 46.125 229.91 46.195 ;
    RECT 366.28 45.405 366.49 45.475 ;
    RECT 366.28 45.765 366.49 45.835 ;
    RECT 366.28 46.125 366.49 46.195 ;
    RECT 365.82 45.405 366.03 45.475 ;
    RECT 365.82 45.765 366.03 45.835 ;
    RECT 365.82 46.125 366.03 46.195 ;
    RECT 226.84 45.405 227.05 45.475 ;
    RECT 226.84 45.765 227.05 45.835 ;
    RECT 226.84 46.125 227.05 46.195 ;
    RECT 226.38 45.405 226.59 45.475 ;
    RECT 226.38 45.765 226.59 45.835 ;
    RECT 226.38 46.125 226.59 46.195 ;
    RECT 362.96 45.405 363.17 45.475 ;
    RECT 362.96 45.765 363.17 45.835 ;
    RECT 362.96 46.125 363.17 46.195 ;
    RECT 362.5 45.405 362.71 45.475 ;
    RECT 362.5 45.765 362.71 45.835 ;
    RECT 362.5 46.125 362.71 46.195 ;
    RECT 223.52 45.405 223.73 45.475 ;
    RECT 223.52 45.765 223.73 45.835 ;
    RECT 223.52 46.125 223.73 46.195 ;
    RECT 223.06 45.405 223.27 45.475 ;
    RECT 223.06 45.765 223.27 45.835 ;
    RECT 223.06 46.125 223.27 46.195 ;
    RECT 359.64 45.405 359.85 45.475 ;
    RECT 359.64 45.765 359.85 45.835 ;
    RECT 359.64 46.125 359.85 46.195 ;
    RECT 359.18 45.405 359.39 45.475 ;
    RECT 359.18 45.765 359.39 45.835 ;
    RECT 359.18 46.125 359.39 46.195 ;
    RECT 220.2 45.405 220.41 45.475 ;
    RECT 220.2 45.765 220.41 45.835 ;
    RECT 220.2 46.125 220.41 46.195 ;
    RECT 219.74 45.405 219.95 45.475 ;
    RECT 219.74 45.765 219.95 45.835 ;
    RECT 219.74 46.125 219.95 46.195 ;
    RECT 356.32 45.405 356.53 45.475 ;
    RECT 356.32 45.765 356.53 45.835 ;
    RECT 356.32 46.125 356.53 46.195 ;
    RECT 355.86 45.405 356.07 45.475 ;
    RECT 355.86 45.765 356.07 45.835 ;
    RECT 355.86 46.125 356.07 46.195 ;
    RECT 353.0 45.405 353.21 45.475 ;
    RECT 353.0 45.765 353.21 45.835 ;
    RECT 353.0 46.125 353.21 46.195 ;
    RECT 352.54 45.405 352.75 45.475 ;
    RECT 352.54 45.765 352.75 45.835 ;
    RECT 352.54 46.125 352.75 46.195 ;
    RECT 216.88 45.405 217.09 45.475 ;
    RECT 216.88 45.765 217.09 45.835 ;
    RECT 216.88 46.125 217.09 46.195 ;
    RECT 216.42 45.405 216.63 45.475 ;
    RECT 216.42 45.765 216.63 45.835 ;
    RECT 216.42 46.125 216.63 46.195 ;
    RECT 349.68 45.405 349.89 45.475 ;
    RECT 349.68 45.765 349.89 45.835 ;
    RECT 349.68 46.125 349.89 46.195 ;
    RECT 349.22 45.405 349.43 45.475 ;
    RECT 349.22 45.765 349.43 45.835 ;
    RECT 349.22 46.125 349.43 46.195 ;
    RECT 213.56 45.405 213.77 45.475 ;
    RECT 213.56 45.765 213.77 45.835 ;
    RECT 213.56 46.125 213.77 46.195 ;
    RECT 213.1 45.405 213.31 45.475 ;
    RECT 213.1 45.765 213.31 45.835 ;
    RECT 213.1 46.125 213.31 46.195 ;
    RECT 346.36 45.405 346.57 45.475 ;
    RECT 346.36 45.765 346.57 45.835 ;
    RECT 346.36 46.125 346.57 46.195 ;
    RECT 345.9 45.405 346.11 45.475 ;
    RECT 345.9 45.765 346.11 45.835 ;
    RECT 345.9 46.125 346.11 46.195 ;
    RECT 210.24 45.405 210.45 45.475 ;
    RECT 210.24 45.765 210.45 45.835 ;
    RECT 210.24 46.125 210.45 46.195 ;
    RECT 209.78 45.405 209.99 45.475 ;
    RECT 209.78 45.765 209.99 45.835 ;
    RECT 209.78 46.125 209.99 46.195 ;
    RECT 343.04 45.405 343.25 45.475 ;
    RECT 343.04 45.765 343.25 45.835 ;
    RECT 343.04 46.125 343.25 46.195 ;
    RECT 342.58 45.405 342.79 45.475 ;
    RECT 342.58 45.765 342.79 45.835 ;
    RECT 342.58 46.125 342.79 46.195 ;
    RECT 206.92 45.405 207.13 45.475 ;
    RECT 206.92 45.765 207.13 45.835 ;
    RECT 206.92 46.125 207.13 46.195 ;
    RECT 206.46 45.405 206.67 45.475 ;
    RECT 206.46 45.765 206.67 45.835 ;
    RECT 206.46 46.125 206.67 46.195 ;
    RECT 339.72 45.405 339.93 45.475 ;
    RECT 339.72 45.765 339.93 45.835 ;
    RECT 339.72 46.125 339.93 46.195 ;
    RECT 339.26 45.405 339.47 45.475 ;
    RECT 339.26 45.765 339.47 45.835 ;
    RECT 339.26 46.125 339.47 46.195 ;
    RECT 203.6 45.405 203.81 45.475 ;
    RECT 203.6 45.765 203.81 45.835 ;
    RECT 203.6 46.125 203.81 46.195 ;
    RECT 203.14 45.405 203.35 45.475 ;
    RECT 203.14 45.765 203.35 45.835 ;
    RECT 203.14 46.125 203.35 46.195 ;
    RECT 336.4 45.405 336.61 45.475 ;
    RECT 336.4 45.765 336.61 45.835 ;
    RECT 336.4 46.125 336.61 46.195 ;
    RECT 335.94 45.405 336.15 45.475 ;
    RECT 335.94 45.765 336.15 45.835 ;
    RECT 335.94 46.125 336.15 46.195 ;
    RECT 266.68 45.405 266.89 45.475 ;
    RECT 266.68 45.765 266.89 45.835 ;
    RECT 266.68 46.125 266.89 46.195 ;
    RECT 266.22 45.405 266.43 45.475 ;
    RECT 266.22 45.765 266.43 45.835 ;
    RECT 266.22 46.125 266.43 46.195 ;
    RECT 263.36 45.405 263.57 45.475 ;
    RECT 263.36 45.765 263.57 45.835 ;
    RECT 263.36 46.125 263.57 46.195 ;
    RECT 262.9 45.405 263.11 45.475 ;
    RECT 262.9 45.765 263.11 45.835 ;
    RECT 262.9 46.125 263.11 46.195 ;
    RECT 260.04 45.405 260.25 45.475 ;
    RECT 260.04 45.765 260.25 45.835 ;
    RECT 260.04 46.125 260.25 46.195 ;
    RECT 259.58 45.405 259.79 45.475 ;
    RECT 259.58 45.765 259.79 45.835 ;
    RECT 259.58 46.125 259.79 46.195 ;
    RECT 256.72 45.405 256.93 45.475 ;
    RECT 256.72 45.765 256.93 45.835 ;
    RECT 256.72 46.125 256.93 46.195 ;
    RECT 256.26 45.405 256.47 45.475 ;
    RECT 256.26 45.765 256.47 45.835 ;
    RECT 256.26 46.125 256.47 46.195 ;
    RECT 253.4 45.405 253.61 45.475 ;
    RECT 253.4 45.765 253.61 45.835 ;
    RECT 253.4 46.125 253.61 46.195 ;
    RECT 252.94 45.405 253.15 45.475 ;
    RECT 252.94 45.765 253.15 45.835 ;
    RECT 252.94 46.125 253.15 46.195 ;
    RECT 250.08 45.405 250.29 45.475 ;
    RECT 250.08 45.765 250.29 45.835 ;
    RECT 250.08 46.125 250.29 46.195 ;
    RECT 249.62 45.405 249.83 45.475 ;
    RECT 249.62 45.765 249.83 45.835 ;
    RECT 249.62 46.125 249.83 46.195 ;
    RECT 246.76 45.405 246.97 45.475 ;
    RECT 246.76 45.765 246.97 45.835 ;
    RECT 246.76 46.125 246.97 46.195 ;
    RECT 246.3 45.405 246.51 45.475 ;
    RECT 246.3 45.765 246.51 45.835 ;
    RECT 246.3 46.125 246.51 46.195 ;
    RECT 243.44 45.405 243.65 45.475 ;
    RECT 243.44 45.765 243.65 45.835 ;
    RECT 243.44 46.125 243.65 46.195 ;
    RECT 242.98 45.405 243.19 45.475 ;
    RECT 242.98 45.765 243.19 45.835 ;
    RECT 242.98 46.125 243.19 46.195 ;
    RECT 240.12 45.405 240.33 45.475 ;
    RECT 240.12 45.765 240.33 45.835 ;
    RECT 240.12 46.125 240.33 46.195 ;
    RECT 239.66 45.405 239.87 45.475 ;
    RECT 239.66 45.765 239.87 45.835 ;
    RECT 239.66 46.125 239.87 46.195 ;
    RECT 236.8 45.405 237.01 45.475 ;
    RECT 236.8 45.765 237.01 45.835 ;
    RECT 236.8 46.125 237.01 46.195 ;
    RECT 236.34 45.405 236.55 45.475 ;
    RECT 236.34 45.765 236.55 45.835 ;
    RECT 236.34 46.125 236.55 46.195 ;
    RECT 374.15 45.765 374.22 45.835 ;
    RECT 333.08 45.405 333.29 45.475 ;
    RECT 333.08 45.765 333.29 45.835 ;
    RECT 333.08 46.125 333.29 46.195 ;
    RECT 332.62 45.405 332.83 45.475 ;
    RECT 332.62 45.765 332.83 45.835 ;
    RECT 332.62 46.125 332.83 46.195 ;
    RECT 329.76 45.405 329.97 45.475 ;
    RECT 329.76 45.765 329.97 45.835 ;
    RECT 329.76 46.125 329.97 46.195 ;
    RECT 329.3 45.405 329.51 45.475 ;
    RECT 329.3 45.765 329.51 45.835 ;
    RECT 329.3 46.125 329.51 46.195 ;
    RECT 326.44 45.405 326.65 45.475 ;
    RECT 326.44 45.765 326.65 45.835 ;
    RECT 326.44 46.125 326.65 46.195 ;
    RECT 325.98 45.405 326.19 45.475 ;
    RECT 325.98 45.765 326.19 45.835 ;
    RECT 325.98 46.125 326.19 46.195 ;
    RECT 323.12 45.405 323.33 45.475 ;
    RECT 323.12 45.765 323.33 45.835 ;
    RECT 323.12 46.125 323.33 46.195 ;
    RECT 322.66 45.405 322.87 45.475 ;
    RECT 322.66 45.765 322.87 45.835 ;
    RECT 322.66 46.125 322.87 46.195 ;
    RECT 319.8 45.405 320.01 45.475 ;
    RECT 319.8 45.765 320.01 45.835 ;
    RECT 319.8 46.125 320.01 46.195 ;
    RECT 319.34 45.405 319.55 45.475 ;
    RECT 319.34 45.765 319.55 45.835 ;
    RECT 319.34 46.125 319.55 46.195 ;
    RECT 316.48 45.405 316.69 45.475 ;
    RECT 316.48 45.765 316.69 45.835 ;
    RECT 316.48 46.125 316.69 46.195 ;
    RECT 316.02 45.405 316.23 45.475 ;
    RECT 316.02 45.765 316.23 45.835 ;
    RECT 316.02 46.125 316.23 46.195 ;
    RECT 313.16 45.405 313.37 45.475 ;
    RECT 313.16 45.765 313.37 45.835 ;
    RECT 313.16 46.125 313.37 46.195 ;
    RECT 312.7 45.405 312.91 45.475 ;
    RECT 312.7 45.765 312.91 45.835 ;
    RECT 312.7 46.125 312.91 46.195 ;
    RECT 309.84 45.405 310.05 45.475 ;
    RECT 309.84 45.765 310.05 45.835 ;
    RECT 309.84 46.125 310.05 46.195 ;
    RECT 309.38 45.405 309.59 45.475 ;
    RECT 309.38 45.765 309.59 45.835 ;
    RECT 309.38 46.125 309.59 46.195 ;
    RECT 306.52 45.405 306.73 45.475 ;
    RECT 306.52 45.765 306.73 45.835 ;
    RECT 306.52 46.125 306.73 46.195 ;
    RECT 306.06 45.405 306.27 45.475 ;
    RECT 306.06 45.765 306.27 45.835 ;
    RECT 306.06 46.125 306.27 46.195 ;
    RECT 303.2 44.685 303.41 44.755 ;
    RECT 303.2 45.045 303.41 45.115 ;
    RECT 303.2 45.405 303.41 45.475 ;
    RECT 302.74 44.685 302.95 44.755 ;
    RECT 302.74 45.045 302.95 45.115 ;
    RECT 302.74 45.405 302.95 45.475 ;
    RECT 372.92 44.685 373.13 44.755 ;
    RECT 372.92 45.045 373.13 45.115 ;
    RECT 372.92 45.405 373.13 45.475 ;
    RECT 372.46 44.685 372.67 44.755 ;
    RECT 372.46 45.045 372.67 45.115 ;
    RECT 372.46 45.405 372.67 45.475 ;
    RECT 369.6 44.685 369.81 44.755 ;
    RECT 369.6 45.045 369.81 45.115 ;
    RECT 369.6 45.405 369.81 45.475 ;
    RECT 369.14 44.685 369.35 44.755 ;
    RECT 369.14 45.045 369.35 45.115 ;
    RECT 369.14 45.405 369.35 45.475 ;
    RECT 200.605 45.045 200.675 45.115 ;
    RECT 299.88 44.685 300.09 44.755 ;
    RECT 299.88 45.045 300.09 45.115 ;
    RECT 299.88 45.405 300.09 45.475 ;
    RECT 299.42 44.685 299.63 44.755 ;
    RECT 299.42 45.045 299.63 45.115 ;
    RECT 299.42 45.405 299.63 45.475 ;
    RECT 296.56 44.685 296.77 44.755 ;
    RECT 296.56 45.045 296.77 45.115 ;
    RECT 296.56 45.405 296.77 45.475 ;
    RECT 296.1 44.685 296.31 44.755 ;
    RECT 296.1 45.045 296.31 45.115 ;
    RECT 296.1 45.405 296.31 45.475 ;
    RECT 293.24 44.685 293.45 44.755 ;
    RECT 293.24 45.045 293.45 45.115 ;
    RECT 293.24 45.405 293.45 45.475 ;
    RECT 292.78 44.685 292.99 44.755 ;
    RECT 292.78 45.045 292.99 45.115 ;
    RECT 292.78 45.405 292.99 45.475 ;
    RECT 289.92 44.685 290.13 44.755 ;
    RECT 289.92 45.045 290.13 45.115 ;
    RECT 289.92 45.405 290.13 45.475 ;
    RECT 289.46 44.685 289.67 44.755 ;
    RECT 289.46 45.045 289.67 45.115 ;
    RECT 289.46 45.405 289.67 45.475 ;
    RECT 286.6 44.685 286.81 44.755 ;
    RECT 286.6 45.045 286.81 45.115 ;
    RECT 286.6 45.405 286.81 45.475 ;
    RECT 286.14 44.685 286.35 44.755 ;
    RECT 286.14 45.045 286.35 45.115 ;
    RECT 286.14 45.405 286.35 45.475 ;
    RECT 283.28 44.685 283.49 44.755 ;
    RECT 283.28 45.045 283.49 45.115 ;
    RECT 283.28 45.405 283.49 45.475 ;
    RECT 282.82 44.685 283.03 44.755 ;
    RECT 282.82 45.045 283.03 45.115 ;
    RECT 282.82 45.405 283.03 45.475 ;
    RECT 279.96 44.685 280.17 44.755 ;
    RECT 279.96 45.045 280.17 45.115 ;
    RECT 279.96 45.405 280.17 45.475 ;
    RECT 279.5 44.685 279.71 44.755 ;
    RECT 279.5 45.045 279.71 45.115 ;
    RECT 279.5 45.405 279.71 45.475 ;
    RECT 276.64 44.685 276.85 44.755 ;
    RECT 276.64 45.045 276.85 45.115 ;
    RECT 276.64 45.405 276.85 45.475 ;
    RECT 276.18 44.685 276.39 44.755 ;
    RECT 276.18 45.045 276.39 45.115 ;
    RECT 276.18 45.405 276.39 45.475 ;
    RECT 273.32 44.685 273.53 44.755 ;
    RECT 273.32 45.045 273.53 45.115 ;
    RECT 273.32 45.405 273.53 45.475 ;
    RECT 272.86 44.685 273.07 44.755 ;
    RECT 272.86 45.045 273.07 45.115 ;
    RECT 272.86 45.405 273.07 45.475 ;
    RECT 270.0 44.685 270.21 44.755 ;
    RECT 270.0 45.045 270.21 45.115 ;
    RECT 270.0 45.405 270.21 45.475 ;
    RECT 269.54 44.685 269.75 44.755 ;
    RECT 269.54 45.045 269.75 45.115 ;
    RECT 269.54 45.405 269.75 45.475 ;
    RECT 233.48 44.685 233.69 44.755 ;
    RECT 233.48 45.045 233.69 45.115 ;
    RECT 233.48 45.405 233.69 45.475 ;
    RECT 233.02 44.685 233.23 44.755 ;
    RECT 233.02 45.045 233.23 45.115 ;
    RECT 233.02 45.405 233.23 45.475 ;
    RECT 230.16 44.685 230.37 44.755 ;
    RECT 230.16 45.045 230.37 45.115 ;
    RECT 230.16 45.405 230.37 45.475 ;
    RECT 229.7 44.685 229.91 44.755 ;
    RECT 229.7 45.045 229.91 45.115 ;
    RECT 229.7 45.405 229.91 45.475 ;
    RECT 366.28 44.685 366.49 44.755 ;
    RECT 366.28 45.045 366.49 45.115 ;
    RECT 366.28 45.405 366.49 45.475 ;
    RECT 365.82 44.685 366.03 44.755 ;
    RECT 365.82 45.045 366.03 45.115 ;
    RECT 365.82 45.405 366.03 45.475 ;
    RECT 226.84 44.685 227.05 44.755 ;
    RECT 226.84 45.045 227.05 45.115 ;
    RECT 226.84 45.405 227.05 45.475 ;
    RECT 226.38 44.685 226.59 44.755 ;
    RECT 226.38 45.045 226.59 45.115 ;
    RECT 226.38 45.405 226.59 45.475 ;
    RECT 362.96 44.685 363.17 44.755 ;
    RECT 362.96 45.045 363.17 45.115 ;
    RECT 362.96 45.405 363.17 45.475 ;
    RECT 362.5 44.685 362.71 44.755 ;
    RECT 362.5 45.045 362.71 45.115 ;
    RECT 362.5 45.405 362.71 45.475 ;
    RECT 223.52 44.685 223.73 44.755 ;
    RECT 223.52 45.045 223.73 45.115 ;
    RECT 223.52 45.405 223.73 45.475 ;
    RECT 223.06 44.685 223.27 44.755 ;
    RECT 223.06 45.045 223.27 45.115 ;
    RECT 223.06 45.405 223.27 45.475 ;
    RECT 359.64 44.685 359.85 44.755 ;
    RECT 359.64 45.045 359.85 45.115 ;
    RECT 359.64 45.405 359.85 45.475 ;
    RECT 359.18 44.685 359.39 44.755 ;
    RECT 359.18 45.045 359.39 45.115 ;
    RECT 359.18 45.405 359.39 45.475 ;
    RECT 220.2 44.685 220.41 44.755 ;
    RECT 220.2 45.045 220.41 45.115 ;
    RECT 220.2 45.405 220.41 45.475 ;
    RECT 219.74 44.685 219.95 44.755 ;
    RECT 219.74 45.045 219.95 45.115 ;
    RECT 219.74 45.405 219.95 45.475 ;
    RECT 356.32 44.685 356.53 44.755 ;
    RECT 356.32 45.045 356.53 45.115 ;
    RECT 356.32 45.405 356.53 45.475 ;
    RECT 355.86 44.685 356.07 44.755 ;
    RECT 355.86 45.045 356.07 45.115 ;
    RECT 355.86 45.405 356.07 45.475 ;
    RECT 353.0 44.685 353.21 44.755 ;
    RECT 353.0 45.045 353.21 45.115 ;
    RECT 353.0 45.405 353.21 45.475 ;
    RECT 352.54 44.685 352.75 44.755 ;
    RECT 352.54 45.045 352.75 45.115 ;
    RECT 352.54 45.405 352.75 45.475 ;
    RECT 216.88 44.685 217.09 44.755 ;
    RECT 216.88 45.045 217.09 45.115 ;
    RECT 216.88 45.405 217.09 45.475 ;
    RECT 216.42 44.685 216.63 44.755 ;
    RECT 216.42 45.045 216.63 45.115 ;
    RECT 216.42 45.405 216.63 45.475 ;
    RECT 349.68 44.685 349.89 44.755 ;
    RECT 349.68 45.045 349.89 45.115 ;
    RECT 349.68 45.405 349.89 45.475 ;
    RECT 349.22 44.685 349.43 44.755 ;
    RECT 349.22 45.045 349.43 45.115 ;
    RECT 349.22 45.405 349.43 45.475 ;
    RECT 213.56 44.685 213.77 44.755 ;
    RECT 213.56 45.045 213.77 45.115 ;
    RECT 213.56 45.405 213.77 45.475 ;
    RECT 213.1 44.685 213.31 44.755 ;
    RECT 213.1 45.045 213.31 45.115 ;
    RECT 213.1 45.405 213.31 45.475 ;
    RECT 346.36 44.685 346.57 44.755 ;
    RECT 346.36 45.045 346.57 45.115 ;
    RECT 346.36 45.405 346.57 45.475 ;
    RECT 345.9 44.685 346.11 44.755 ;
    RECT 345.9 45.045 346.11 45.115 ;
    RECT 345.9 45.405 346.11 45.475 ;
    RECT 210.24 44.685 210.45 44.755 ;
    RECT 210.24 45.045 210.45 45.115 ;
    RECT 210.24 45.405 210.45 45.475 ;
    RECT 209.78 44.685 209.99 44.755 ;
    RECT 209.78 45.045 209.99 45.115 ;
    RECT 209.78 45.405 209.99 45.475 ;
    RECT 343.04 44.685 343.25 44.755 ;
    RECT 343.04 45.045 343.25 45.115 ;
    RECT 343.04 45.405 343.25 45.475 ;
    RECT 342.58 44.685 342.79 44.755 ;
    RECT 342.58 45.045 342.79 45.115 ;
    RECT 342.58 45.405 342.79 45.475 ;
    RECT 206.92 44.685 207.13 44.755 ;
    RECT 206.92 45.045 207.13 45.115 ;
    RECT 206.92 45.405 207.13 45.475 ;
    RECT 206.46 44.685 206.67 44.755 ;
    RECT 206.46 45.045 206.67 45.115 ;
    RECT 206.46 45.405 206.67 45.475 ;
    RECT 339.72 44.685 339.93 44.755 ;
    RECT 339.72 45.045 339.93 45.115 ;
    RECT 339.72 45.405 339.93 45.475 ;
    RECT 339.26 44.685 339.47 44.755 ;
    RECT 339.26 45.045 339.47 45.115 ;
    RECT 339.26 45.405 339.47 45.475 ;
    RECT 203.6 44.685 203.81 44.755 ;
    RECT 203.6 45.045 203.81 45.115 ;
    RECT 203.6 45.405 203.81 45.475 ;
    RECT 203.14 44.685 203.35 44.755 ;
    RECT 203.14 45.045 203.35 45.115 ;
    RECT 203.14 45.405 203.35 45.475 ;
    RECT 336.4 44.685 336.61 44.755 ;
    RECT 336.4 45.045 336.61 45.115 ;
    RECT 336.4 45.405 336.61 45.475 ;
    RECT 335.94 44.685 336.15 44.755 ;
    RECT 335.94 45.045 336.15 45.115 ;
    RECT 335.94 45.405 336.15 45.475 ;
    RECT 266.68 44.685 266.89 44.755 ;
    RECT 266.68 45.045 266.89 45.115 ;
    RECT 266.68 45.405 266.89 45.475 ;
    RECT 266.22 44.685 266.43 44.755 ;
    RECT 266.22 45.045 266.43 45.115 ;
    RECT 266.22 45.405 266.43 45.475 ;
    RECT 263.36 44.685 263.57 44.755 ;
    RECT 263.36 45.045 263.57 45.115 ;
    RECT 263.36 45.405 263.57 45.475 ;
    RECT 262.9 44.685 263.11 44.755 ;
    RECT 262.9 45.045 263.11 45.115 ;
    RECT 262.9 45.405 263.11 45.475 ;
    RECT 260.04 44.685 260.25 44.755 ;
    RECT 260.04 45.045 260.25 45.115 ;
    RECT 260.04 45.405 260.25 45.475 ;
    RECT 259.58 44.685 259.79 44.755 ;
    RECT 259.58 45.045 259.79 45.115 ;
    RECT 259.58 45.405 259.79 45.475 ;
    RECT 256.72 44.685 256.93 44.755 ;
    RECT 256.72 45.045 256.93 45.115 ;
    RECT 256.72 45.405 256.93 45.475 ;
    RECT 256.26 44.685 256.47 44.755 ;
    RECT 256.26 45.045 256.47 45.115 ;
    RECT 256.26 45.405 256.47 45.475 ;
    RECT 253.4 44.685 253.61 44.755 ;
    RECT 253.4 45.045 253.61 45.115 ;
    RECT 253.4 45.405 253.61 45.475 ;
    RECT 252.94 44.685 253.15 44.755 ;
    RECT 252.94 45.045 253.15 45.115 ;
    RECT 252.94 45.405 253.15 45.475 ;
    RECT 250.08 44.685 250.29 44.755 ;
    RECT 250.08 45.045 250.29 45.115 ;
    RECT 250.08 45.405 250.29 45.475 ;
    RECT 249.62 44.685 249.83 44.755 ;
    RECT 249.62 45.045 249.83 45.115 ;
    RECT 249.62 45.405 249.83 45.475 ;
    RECT 246.76 44.685 246.97 44.755 ;
    RECT 246.76 45.045 246.97 45.115 ;
    RECT 246.76 45.405 246.97 45.475 ;
    RECT 246.3 44.685 246.51 44.755 ;
    RECT 246.3 45.045 246.51 45.115 ;
    RECT 246.3 45.405 246.51 45.475 ;
    RECT 243.44 44.685 243.65 44.755 ;
    RECT 243.44 45.045 243.65 45.115 ;
    RECT 243.44 45.405 243.65 45.475 ;
    RECT 242.98 44.685 243.19 44.755 ;
    RECT 242.98 45.045 243.19 45.115 ;
    RECT 242.98 45.405 243.19 45.475 ;
    RECT 240.12 44.685 240.33 44.755 ;
    RECT 240.12 45.045 240.33 45.115 ;
    RECT 240.12 45.405 240.33 45.475 ;
    RECT 239.66 44.685 239.87 44.755 ;
    RECT 239.66 45.045 239.87 45.115 ;
    RECT 239.66 45.405 239.87 45.475 ;
    RECT 236.8 44.685 237.01 44.755 ;
    RECT 236.8 45.045 237.01 45.115 ;
    RECT 236.8 45.405 237.01 45.475 ;
    RECT 236.34 44.685 236.55 44.755 ;
    RECT 236.34 45.045 236.55 45.115 ;
    RECT 236.34 45.405 236.55 45.475 ;
    RECT 374.15 45.045 374.22 45.115 ;
    RECT 333.08 44.685 333.29 44.755 ;
    RECT 333.08 45.045 333.29 45.115 ;
    RECT 333.08 45.405 333.29 45.475 ;
    RECT 332.62 44.685 332.83 44.755 ;
    RECT 332.62 45.045 332.83 45.115 ;
    RECT 332.62 45.405 332.83 45.475 ;
    RECT 329.76 44.685 329.97 44.755 ;
    RECT 329.76 45.045 329.97 45.115 ;
    RECT 329.76 45.405 329.97 45.475 ;
    RECT 329.3 44.685 329.51 44.755 ;
    RECT 329.3 45.045 329.51 45.115 ;
    RECT 329.3 45.405 329.51 45.475 ;
    RECT 326.44 44.685 326.65 44.755 ;
    RECT 326.44 45.045 326.65 45.115 ;
    RECT 326.44 45.405 326.65 45.475 ;
    RECT 325.98 44.685 326.19 44.755 ;
    RECT 325.98 45.045 326.19 45.115 ;
    RECT 325.98 45.405 326.19 45.475 ;
    RECT 323.12 44.685 323.33 44.755 ;
    RECT 323.12 45.045 323.33 45.115 ;
    RECT 323.12 45.405 323.33 45.475 ;
    RECT 322.66 44.685 322.87 44.755 ;
    RECT 322.66 45.045 322.87 45.115 ;
    RECT 322.66 45.405 322.87 45.475 ;
    RECT 319.8 44.685 320.01 44.755 ;
    RECT 319.8 45.045 320.01 45.115 ;
    RECT 319.8 45.405 320.01 45.475 ;
    RECT 319.34 44.685 319.55 44.755 ;
    RECT 319.34 45.045 319.55 45.115 ;
    RECT 319.34 45.405 319.55 45.475 ;
    RECT 316.48 44.685 316.69 44.755 ;
    RECT 316.48 45.045 316.69 45.115 ;
    RECT 316.48 45.405 316.69 45.475 ;
    RECT 316.02 44.685 316.23 44.755 ;
    RECT 316.02 45.045 316.23 45.115 ;
    RECT 316.02 45.405 316.23 45.475 ;
    RECT 313.16 44.685 313.37 44.755 ;
    RECT 313.16 45.045 313.37 45.115 ;
    RECT 313.16 45.405 313.37 45.475 ;
    RECT 312.7 44.685 312.91 44.755 ;
    RECT 312.7 45.045 312.91 45.115 ;
    RECT 312.7 45.405 312.91 45.475 ;
    RECT 309.84 44.685 310.05 44.755 ;
    RECT 309.84 45.045 310.05 45.115 ;
    RECT 309.84 45.405 310.05 45.475 ;
    RECT 309.38 44.685 309.59 44.755 ;
    RECT 309.38 45.045 309.59 45.115 ;
    RECT 309.38 45.405 309.59 45.475 ;
    RECT 306.52 44.685 306.73 44.755 ;
    RECT 306.52 45.045 306.73 45.115 ;
    RECT 306.52 45.405 306.73 45.475 ;
    RECT 306.06 44.685 306.27 44.755 ;
    RECT 306.06 45.045 306.27 45.115 ;
    RECT 306.06 45.405 306.27 45.475 ;
    RECT 303.2 43.965 303.41 44.035 ;
    RECT 303.2 44.325 303.41 44.395 ;
    RECT 303.2 44.685 303.41 44.755 ;
    RECT 302.74 43.965 302.95 44.035 ;
    RECT 302.74 44.325 302.95 44.395 ;
    RECT 302.74 44.685 302.95 44.755 ;
    RECT 372.92 43.965 373.13 44.035 ;
    RECT 372.92 44.325 373.13 44.395 ;
    RECT 372.92 44.685 373.13 44.755 ;
    RECT 372.46 43.965 372.67 44.035 ;
    RECT 372.46 44.325 372.67 44.395 ;
    RECT 372.46 44.685 372.67 44.755 ;
    RECT 369.6 43.965 369.81 44.035 ;
    RECT 369.6 44.325 369.81 44.395 ;
    RECT 369.6 44.685 369.81 44.755 ;
    RECT 369.14 43.965 369.35 44.035 ;
    RECT 369.14 44.325 369.35 44.395 ;
    RECT 369.14 44.685 369.35 44.755 ;
    RECT 200.605 44.325 200.675 44.395 ;
    RECT 299.88 43.965 300.09 44.035 ;
    RECT 299.88 44.325 300.09 44.395 ;
    RECT 299.88 44.685 300.09 44.755 ;
    RECT 299.42 43.965 299.63 44.035 ;
    RECT 299.42 44.325 299.63 44.395 ;
    RECT 299.42 44.685 299.63 44.755 ;
    RECT 296.56 43.965 296.77 44.035 ;
    RECT 296.56 44.325 296.77 44.395 ;
    RECT 296.56 44.685 296.77 44.755 ;
    RECT 296.1 43.965 296.31 44.035 ;
    RECT 296.1 44.325 296.31 44.395 ;
    RECT 296.1 44.685 296.31 44.755 ;
    RECT 293.24 43.965 293.45 44.035 ;
    RECT 293.24 44.325 293.45 44.395 ;
    RECT 293.24 44.685 293.45 44.755 ;
    RECT 292.78 43.965 292.99 44.035 ;
    RECT 292.78 44.325 292.99 44.395 ;
    RECT 292.78 44.685 292.99 44.755 ;
    RECT 289.92 43.965 290.13 44.035 ;
    RECT 289.92 44.325 290.13 44.395 ;
    RECT 289.92 44.685 290.13 44.755 ;
    RECT 289.46 43.965 289.67 44.035 ;
    RECT 289.46 44.325 289.67 44.395 ;
    RECT 289.46 44.685 289.67 44.755 ;
    RECT 286.6 43.965 286.81 44.035 ;
    RECT 286.6 44.325 286.81 44.395 ;
    RECT 286.6 44.685 286.81 44.755 ;
    RECT 286.14 43.965 286.35 44.035 ;
    RECT 286.14 44.325 286.35 44.395 ;
    RECT 286.14 44.685 286.35 44.755 ;
    RECT 283.28 43.965 283.49 44.035 ;
    RECT 283.28 44.325 283.49 44.395 ;
    RECT 283.28 44.685 283.49 44.755 ;
    RECT 282.82 43.965 283.03 44.035 ;
    RECT 282.82 44.325 283.03 44.395 ;
    RECT 282.82 44.685 283.03 44.755 ;
    RECT 279.96 43.965 280.17 44.035 ;
    RECT 279.96 44.325 280.17 44.395 ;
    RECT 279.96 44.685 280.17 44.755 ;
    RECT 279.5 43.965 279.71 44.035 ;
    RECT 279.5 44.325 279.71 44.395 ;
    RECT 279.5 44.685 279.71 44.755 ;
    RECT 276.64 43.965 276.85 44.035 ;
    RECT 276.64 44.325 276.85 44.395 ;
    RECT 276.64 44.685 276.85 44.755 ;
    RECT 276.18 43.965 276.39 44.035 ;
    RECT 276.18 44.325 276.39 44.395 ;
    RECT 276.18 44.685 276.39 44.755 ;
    RECT 273.32 43.965 273.53 44.035 ;
    RECT 273.32 44.325 273.53 44.395 ;
    RECT 273.32 44.685 273.53 44.755 ;
    RECT 272.86 43.965 273.07 44.035 ;
    RECT 272.86 44.325 273.07 44.395 ;
    RECT 272.86 44.685 273.07 44.755 ;
    RECT 270.0 43.965 270.21 44.035 ;
    RECT 270.0 44.325 270.21 44.395 ;
    RECT 270.0 44.685 270.21 44.755 ;
    RECT 269.54 43.965 269.75 44.035 ;
    RECT 269.54 44.325 269.75 44.395 ;
    RECT 269.54 44.685 269.75 44.755 ;
    RECT 233.48 43.965 233.69 44.035 ;
    RECT 233.48 44.325 233.69 44.395 ;
    RECT 233.48 44.685 233.69 44.755 ;
    RECT 233.02 43.965 233.23 44.035 ;
    RECT 233.02 44.325 233.23 44.395 ;
    RECT 233.02 44.685 233.23 44.755 ;
    RECT 230.16 43.965 230.37 44.035 ;
    RECT 230.16 44.325 230.37 44.395 ;
    RECT 230.16 44.685 230.37 44.755 ;
    RECT 229.7 43.965 229.91 44.035 ;
    RECT 229.7 44.325 229.91 44.395 ;
    RECT 229.7 44.685 229.91 44.755 ;
    RECT 366.28 43.965 366.49 44.035 ;
    RECT 366.28 44.325 366.49 44.395 ;
    RECT 366.28 44.685 366.49 44.755 ;
    RECT 365.82 43.965 366.03 44.035 ;
    RECT 365.82 44.325 366.03 44.395 ;
    RECT 365.82 44.685 366.03 44.755 ;
    RECT 226.84 43.965 227.05 44.035 ;
    RECT 226.84 44.325 227.05 44.395 ;
    RECT 226.84 44.685 227.05 44.755 ;
    RECT 226.38 43.965 226.59 44.035 ;
    RECT 226.38 44.325 226.59 44.395 ;
    RECT 226.38 44.685 226.59 44.755 ;
    RECT 362.96 43.965 363.17 44.035 ;
    RECT 362.96 44.325 363.17 44.395 ;
    RECT 362.96 44.685 363.17 44.755 ;
    RECT 362.5 43.965 362.71 44.035 ;
    RECT 362.5 44.325 362.71 44.395 ;
    RECT 362.5 44.685 362.71 44.755 ;
    RECT 223.52 43.965 223.73 44.035 ;
    RECT 223.52 44.325 223.73 44.395 ;
    RECT 223.52 44.685 223.73 44.755 ;
    RECT 223.06 43.965 223.27 44.035 ;
    RECT 223.06 44.325 223.27 44.395 ;
    RECT 223.06 44.685 223.27 44.755 ;
    RECT 359.64 43.965 359.85 44.035 ;
    RECT 359.64 44.325 359.85 44.395 ;
    RECT 359.64 44.685 359.85 44.755 ;
    RECT 359.18 43.965 359.39 44.035 ;
    RECT 359.18 44.325 359.39 44.395 ;
    RECT 359.18 44.685 359.39 44.755 ;
    RECT 220.2 43.965 220.41 44.035 ;
    RECT 220.2 44.325 220.41 44.395 ;
    RECT 220.2 44.685 220.41 44.755 ;
    RECT 219.74 43.965 219.95 44.035 ;
    RECT 219.74 44.325 219.95 44.395 ;
    RECT 219.74 44.685 219.95 44.755 ;
    RECT 356.32 43.965 356.53 44.035 ;
    RECT 356.32 44.325 356.53 44.395 ;
    RECT 356.32 44.685 356.53 44.755 ;
    RECT 355.86 43.965 356.07 44.035 ;
    RECT 355.86 44.325 356.07 44.395 ;
    RECT 355.86 44.685 356.07 44.755 ;
    RECT 353.0 43.965 353.21 44.035 ;
    RECT 353.0 44.325 353.21 44.395 ;
    RECT 353.0 44.685 353.21 44.755 ;
    RECT 352.54 43.965 352.75 44.035 ;
    RECT 352.54 44.325 352.75 44.395 ;
    RECT 352.54 44.685 352.75 44.755 ;
    RECT 216.88 43.965 217.09 44.035 ;
    RECT 216.88 44.325 217.09 44.395 ;
    RECT 216.88 44.685 217.09 44.755 ;
    RECT 216.42 43.965 216.63 44.035 ;
    RECT 216.42 44.325 216.63 44.395 ;
    RECT 216.42 44.685 216.63 44.755 ;
    RECT 349.68 43.965 349.89 44.035 ;
    RECT 349.68 44.325 349.89 44.395 ;
    RECT 349.68 44.685 349.89 44.755 ;
    RECT 349.22 43.965 349.43 44.035 ;
    RECT 349.22 44.325 349.43 44.395 ;
    RECT 349.22 44.685 349.43 44.755 ;
    RECT 213.56 43.965 213.77 44.035 ;
    RECT 213.56 44.325 213.77 44.395 ;
    RECT 213.56 44.685 213.77 44.755 ;
    RECT 213.1 43.965 213.31 44.035 ;
    RECT 213.1 44.325 213.31 44.395 ;
    RECT 213.1 44.685 213.31 44.755 ;
    RECT 346.36 43.965 346.57 44.035 ;
    RECT 346.36 44.325 346.57 44.395 ;
    RECT 346.36 44.685 346.57 44.755 ;
    RECT 345.9 43.965 346.11 44.035 ;
    RECT 345.9 44.325 346.11 44.395 ;
    RECT 345.9 44.685 346.11 44.755 ;
    RECT 210.24 43.965 210.45 44.035 ;
    RECT 210.24 44.325 210.45 44.395 ;
    RECT 210.24 44.685 210.45 44.755 ;
    RECT 209.78 43.965 209.99 44.035 ;
    RECT 209.78 44.325 209.99 44.395 ;
    RECT 209.78 44.685 209.99 44.755 ;
    RECT 343.04 43.965 343.25 44.035 ;
    RECT 343.04 44.325 343.25 44.395 ;
    RECT 343.04 44.685 343.25 44.755 ;
    RECT 342.58 43.965 342.79 44.035 ;
    RECT 342.58 44.325 342.79 44.395 ;
    RECT 342.58 44.685 342.79 44.755 ;
    RECT 206.92 43.965 207.13 44.035 ;
    RECT 206.92 44.325 207.13 44.395 ;
    RECT 206.92 44.685 207.13 44.755 ;
    RECT 206.46 43.965 206.67 44.035 ;
    RECT 206.46 44.325 206.67 44.395 ;
    RECT 206.46 44.685 206.67 44.755 ;
    RECT 339.72 43.965 339.93 44.035 ;
    RECT 339.72 44.325 339.93 44.395 ;
    RECT 339.72 44.685 339.93 44.755 ;
    RECT 339.26 43.965 339.47 44.035 ;
    RECT 339.26 44.325 339.47 44.395 ;
    RECT 339.26 44.685 339.47 44.755 ;
    RECT 203.6 43.965 203.81 44.035 ;
    RECT 203.6 44.325 203.81 44.395 ;
    RECT 203.6 44.685 203.81 44.755 ;
    RECT 203.14 43.965 203.35 44.035 ;
    RECT 203.14 44.325 203.35 44.395 ;
    RECT 203.14 44.685 203.35 44.755 ;
    RECT 336.4 43.965 336.61 44.035 ;
    RECT 336.4 44.325 336.61 44.395 ;
    RECT 336.4 44.685 336.61 44.755 ;
    RECT 335.94 43.965 336.15 44.035 ;
    RECT 335.94 44.325 336.15 44.395 ;
    RECT 335.94 44.685 336.15 44.755 ;
    RECT 266.68 43.965 266.89 44.035 ;
    RECT 266.68 44.325 266.89 44.395 ;
    RECT 266.68 44.685 266.89 44.755 ;
    RECT 266.22 43.965 266.43 44.035 ;
    RECT 266.22 44.325 266.43 44.395 ;
    RECT 266.22 44.685 266.43 44.755 ;
    RECT 263.36 43.965 263.57 44.035 ;
    RECT 263.36 44.325 263.57 44.395 ;
    RECT 263.36 44.685 263.57 44.755 ;
    RECT 262.9 43.965 263.11 44.035 ;
    RECT 262.9 44.325 263.11 44.395 ;
    RECT 262.9 44.685 263.11 44.755 ;
    RECT 260.04 43.965 260.25 44.035 ;
    RECT 260.04 44.325 260.25 44.395 ;
    RECT 260.04 44.685 260.25 44.755 ;
    RECT 259.58 43.965 259.79 44.035 ;
    RECT 259.58 44.325 259.79 44.395 ;
    RECT 259.58 44.685 259.79 44.755 ;
    RECT 256.72 43.965 256.93 44.035 ;
    RECT 256.72 44.325 256.93 44.395 ;
    RECT 256.72 44.685 256.93 44.755 ;
    RECT 256.26 43.965 256.47 44.035 ;
    RECT 256.26 44.325 256.47 44.395 ;
    RECT 256.26 44.685 256.47 44.755 ;
    RECT 253.4 43.965 253.61 44.035 ;
    RECT 253.4 44.325 253.61 44.395 ;
    RECT 253.4 44.685 253.61 44.755 ;
    RECT 252.94 43.965 253.15 44.035 ;
    RECT 252.94 44.325 253.15 44.395 ;
    RECT 252.94 44.685 253.15 44.755 ;
    RECT 250.08 43.965 250.29 44.035 ;
    RECT 250.08 44.325 250.29 44.395 ;
    RECT 250.08 44.685 250.29 44.755 ;
    RECT 249.62 43.965 249.83 44.035 ;
    RECT 249.62 44.325 249.83 44.395 ;
    RECT 249.62 44.685 249.83 44.755 ;
    RECT 246.76 43.965 246.97 44.035 ;
    RECT 246.76 44.325 246.97 44.395 ;
    RECT 246.76 44.685 246.97 44.755 ;
    RECT 246.3 43.965 246.51 44.035 ;
    RECT 246.3 44.325 246.51 44.395 ;
    RECT 246.3 44.685 246.51 44.755 ;
    RECT 243.44 43.965 243.65 44.035 ;
    RECT 243.44 44.325 243.65 44.395 ;
    RECT 243.44 44.685 243.65 44.755 ;
    RECT 242.98 43.965 243.19 44.035 ;
    RECT 242.98 44.325 243.19 44.395 ;
    RECT 242.98 44.685 243.19 44.755 ;
    RECT 240.12 43.965 240.33 44.035 ;
    RECT 240.12 44.325 240.33 44.395 ;
    RECT 240.12 44.685 240.33 44.755 ;
    RECT 239.66 43.965 239.87 44.035 ;
    RECT 239.66 44.325 239.87 44.395 ;
    RECT 239.66 44.685 239.87 44.755 ;
    RECT 236.8 43.965 237.01 44.035 ;
    RECT 236.8 44.325 237.01 44.395 ;
    RECT 236.8 44.685 237.01 44.755 ;
    RECT 236.34 43.965 236.55 44.035 ;
    RECT 236.34 44.325 236.55 44.395 ;
    RECT 236.34 44.685 236.55 44.755 ;
    RECT 374.15 44.325 374.22 44.395 ;
    RECT 333.08 43.965 333.29 44.035 ;
    RECT 333.08 44.325 333.29 44.395 ;
    RECT 333.08 44.685 333.29 44.755 ;
    RECT 332.62 43.965 332.83 44.035 ;
    RECT 332.62 44.325 332.83 44.395 ;
    RECT 332.62 44.685 332.83 44.755 ;
    RECT 329.76 43.965 329.97 44.035 ;
    RECT 329.76 44.325 329.97 44.395 ;
    RECT 329.76 44.685 329.97 44.755 ;
    RECT 329.3 43.965 329.51 44.035 ;
    RECT 329.3 44.325 329.51 44.395 ;
    RECT 329.3 44.685 329.51 44.755 ;
    RECT 326.44 43.965 326.65 44.035 ;
    RECT 326.44 44.325 326.65 44.395 ;
    RECT 326.44 44.685 326.65 44.755 ;
    RECT 325.98 43.965 326.19 44.035 ;
    RECT 325.98 44.325 326.19 44.395 ;
    RECT 325.98 44.685 326.19 44.755 ;
    RECT 323.12 43.965 323.33 44.035 ;
    RECT 323.12 44.325 323.33 44.395 ;
    RECT 323.12 44.685 323.33 44.755 ;
    RECT 322.66 43.965 322.87 44.035 ;
    RECT 322.66 44.325 322.87 44.395 ;
    RECT 322.66 44.685 322.87 44.755 ;
    RECT 319.8 43.965 320.01 44.035 ;
    RECT 319.8 44.325 320.01 44.395 ;
    RECT 319.8 44.685 320.01 44.755 ;
    RECT 319.34 43.965 319.55 44.035 ;
    RECT 319.34 44.325 319.55 44.395 ;
    RECT 319.34 44.685 319.55 44.755 ;
    RECT 316.48 43.965 316.69 44.035 ;
    RECT 316.48 44.325 316.69 44.395 ;
    RECT 316.48 44.685 316.69 44.755 ;
    RECT 316.02 43.965 316.23 44.035 ;
    RECT 316.02 44.325 316.23 44.395 ;
    RECT 316.02 44.685 316.23 44.755 ;
    RECT 313.16 43.965 313.37 44.035 ;
    RECT 313.16 44.325 313.37 44.395 ;
    RECT 313.16 44.685 313.37 44.755 ;
    RECT 312.7 43.965 312.91 44.035 ;
    RECT 312.7 44.325 312.91 44.395 ;
    RECT 312.7 44.685 312.91 44.755 ;
    RECT 309.84 43.965 310.05 44.035 ;
    RECT 309.84 44.325 310.05 44.395 ;
    RECT 309.84 44.685 310.05 44.755 ;
    RECT 309.38 43.965 309.59 44.035 ;
    RECT 309.38 44.325 309.59 44.395 ;
    RECT 309.38 44.685 309.59 44.755 ;
    RECT 306.52 43.965 306.73 44.035 ;
    RECT 306.52 44.325 306.73 44.395 ;
    RECT 306.52 44.685 306.73 44.755 ;
    RECT 306.06 43.965 306.27 44.035 ;
    RECT 306.06 44.325 306.27 44.395 ;
    RECT 306.06 44.685 306.27 44.755 ;
    RECT 303.2 43.245 303.41 43.315 ;
    RECT 303.2 43.605 303.41 43.675 ;
    RECT 303.2 43.965 303.41 44.035 ;
    RECT 302.74 43.245 302.95 43.315 ;
    RECT 302.74 43.605 302.95 43.675 ;
    RECT 302.74 43.965 302.95 44.035 ;
    RECT 372.92 43.245 373.13 43.315 ;
    RECT 372.92 43.605 373.13 43.675 ;
    RECT 372.92 43.965 373.13 44.035 ;
    RECT 372.46 43.245 372.67 43.315 ;
    RECT 372.46 43.605 372.67 43.675 ;
    RECT 372.46 43.965 372.67 44.035 ;
    RECT 369.6 43.245 369.81 43.315 ;
    RECT 369.6 43.605 369.81 43.675 ;
    RECT 369.6 43.965 369.81 44.035 ;
    RECT 369.14 43.245 369.35 43.315 ;
    RECT 369.14 43.605 369.35 43.675 ;
    RECT 369.14 43.965 369.35 44.035 ;
    RECT 200.605 43.605 200.675 43.675 ;
    RECT 299.88 43.245 300.09 43.315 ;
    RECT 299.88 43.605 300.09 43.675 ;
    RECT 299.88 43.965 300.09 44.035 ;
    RECT 299.42 43.245 299.63 43.315 ;
    RECT 299.42 43.605 299.63 43.675 ;
    RECT 299.42 43.965 299.63 44.035 ;
    RECT 296.56 43.245 296.77 43.315 ;
    RECT 296.56 43.605 296.77 43.675 ;
    RECT 296.56 43.965 296.77 44.035 ;
    RECT 296.1 43.245 296.31 43.315 ;
    RECT 296.1 43.605 296.31 43.675 ;
    RECT 296.1 43.965 296.31 44.035 ;
    RECT 293.24 43.245 293.45 43.315 ;
    RECT 293.24 43.605 293.45 43.675 ;
    RECT 293.24 43.965 293.45 44.035 ;
    RECT 292.78 43.245 292.99 43.315 ;
    RECT 292.78 43.605 292.99 43.675 ;
    RECT 292.78 43.965 292.99 44.035 ;
    RECT 289.92 43.245 290.13 43.315 ;
    RECT 289.92 43.605 290.13 43.675 ;
    RECT 289.92 43.965 290.13 44.035 ;
    RECT 289.46 43.245 289.67 43.315 ;
    RECT 289.46 43.605 289.67 43.675 ;
    RECT 289.46 43.965 289.67 44.035 ;
    RECT 286.6 43.245 286.81 43.315 ;
    RECT 286.6 43.605 286.81 43.675 ;
    RECT 286.6 43.965 286.81 44.035 ;
    RECT 286.14 43.245 286.35 43.315 ;
    RECT 286.14 43.605 286.35 43.675 ;
    RECT 286.14 43.965 286.35 44.035 ;
    RECT 283.28 43.245 283.49 43.315 ;
    RECT 283.28 43.605 283.49 43.675 ;
    RECT 283.28 43.965 283.49 44.035 ;
    RECT 282.82 43.245 283.03 43.315 ;
    RECT 282.82 43.605 283.03 43.675 ;
    RECT 282.82 43.965 283.03 44.035 ;
    RECT 279.96 43.245 280.17 43.315 ;
    RECT 279.96 43.605 280.17 43.675 ;
    RECT 279.96 43.965 280.17 44.035 ;
    RECT 279.5 43.245 279.71 43.315 ;
    RECT 279.5 43.605 279.71 43.675 ;
    RECT 279.5 43.965 279.71 44.035 ;
    RECT 276.64 43.245 276.85 43.315 ;
    RECT 276.64 43.605 276.85 43.675 ;
    RECT 276.64 43.965 276.85 44.035 ;
    RECT 276.18 43.245 276.39 43.315 ;
    RECT 276.18 43.605 276.39 43.675 ;
    RECT 276.18 43.965 276.39 44.035 ;
    RECT 273.32 43.245 273.53 43.315 ;
    RECT 273.32 43.605 273.53 43.675 ;
    RECT 273.32 43.965 273.53 44.035 ;
    RECT 272.86 43.245 273.07 43.315 ;
    RECT 272.86 43.605 273.07 43.675 ;
    RECT 272.86 43.965 273.07 44.035 ;
    RECT 270.0 43.245 270.21 43.315 ;
    RECT 270.0 43.605 270.21 43.675 ;
    RECT 270.0 43.965 270.21 44.035 ;
    RECT 269.54 43.245 269.75 43.315 ;
    RECT 269.54 43.605 269.75 43.675 ;
    RECT 269.54 43.965 269.75 44.035 ;
    RECT 233.48 43.245 233.69 43.315 ;
    RECT 233.48 43.605 233.69 43.675 ;
    RECT 233.48 43.965 233.69 44.035 ;
    RECT 233.02 43.245 233.23 43.315 ;
    RECT 233.02 43.605 233.23 43.675 ;
    RECT 233.02 43.965 233.23 44.035 ;
    RECT 230.16 43.245 230.37 43.315 ;
    RECT 230.16 43.605 230.37 43.675 ;
    RECT 230.16 43.965 230.37 44.035 ;
    RECT 229.7 43.245 229.91 43.315 ;
    RECT 229.7 43.605 229.91 43.675 ;
    RECT 229.7 43.965 229.91 44.035 ;
    RECT 366.28 43.245 366.49 43.315 ;
    RECT 366.28 43.605 366.49 43.675 ;
    RECT 366.28 43.965 366.49 44.035 ;
    RECT 365.82 43.245 366.03 43.315 ;
    RECT 365.82 43.605 366.03 43.675 ;
    RECT 365.82 43.965 366.03 44.035 ;
    RECT 226.84 43.245 227.05 43.315 ;
    RECT 226.84 43.605 227.05 43.675 ;
    RECT 226.84 43.965 227.05 44.035 ;
    RECT 226.38 43.245 226.59 43.315 ;
    RECT 226.38 43.605 226.59 43.675 ;
    RECT 226.38 43.965 226.59 44.035 ;
    RECT 362.96 43.245 363.17 43.315 ;
    RECT 362.96 43.605 363.17 43.675 ;
    RECT 362.96 43.965 363.17 44.035 ;
    RECT 362.5 43.245 362.71 43.315 ;
    RECT 362.5 43.605 362.71 43.675 ;
    RECT 362.5 43.965 362.71 44.035 ;
    RECT 223.52 43.245 223.73 43.315 ;
    RECT 223.52 43.605 223.73 43.675 ;
    RECT 223.52 43.965 223.73 44.035 ;
    RECT 223.06 43.245 223.27 43.315 ;
    RECT 223.06 43.605 223.27 43.675 ;
    RECT 223.06 43.965 223.27 44.035 ;
    RECT 359.64 43.245 359.85 43.315 ;
    RECT 359.64 43.605 359.85 43.675 ;
    RECT 359.64 43.965 359.85 44.035 ;
    RECT 359.18 43.245 359.39 43.315 ;
    RECT 359.18 43.605 359.39 43.675 ;
    RECT 359.18 43.965 359.39 44.035 ;
    RECT 220.2 43.245 220.41 43.315 ;
    RECT 220.2 43.605 220.41 43.675 ;
    RECT 220.2 43.965 220.41 44.035 ;
    RECT 219.74 43.245 219.95 43.315 ;
    RECT 219.74 43.605 219.95 43.675 ;
    RECT 219.74 43.965 219.95 44.035 ;
    RECT 356.32 43.245 356.53 43.315 ;
    RECT 356.32 43.605 356.53 43.675 ;
    RECT 356.32 43.965 356.53 44.035 ;
    RECT 355.86 43.245 356.07 43.315 ;
    RECT 355.86 43.605 356.07 43.675 ;
    RECT 355.86 43.965 356.07 44.035 ;
    RECT 353.0 43.245 353.21 43.315 ;
    RECT 353.0 43.605 353.21 43.675 ;
    RECT 353.0 43.965 353.21 44.035 ;
    RECT 352.54 43.245 352.75 43.315 ;
    RECT 352.54 43.605 352.75 43.675 ;
    RECT 352.54 43.965 352.75 44.035 ;
    RECT 216.88 43.245 217.09 43.315 ;
    RECT 216.88 43.605 217.09 43.675 ;
    RECT 216.88 43.965 217.09 44.035 ;
    RECT 216.42 43.245 216.63 43.315 ;
    RECT 216.42 43.605 216.63 43.675 ;
    RECT 216.42 43.965 216.63 44.035 ;
    RECT 349.68 43.245 349.89 43.315 ;
    RECT 349.68 43.605 349.89 43.675 ;
    RECT 349.68 43.965 349.89 44.035 ;
    RECT 349.22 43.245 349.43 43.315 ;
    RECT 349.22 43.605 349.43 43.675 ;
    RECT 349.22 43.965 349.43 44.035 ;
    RECT 213.56 43.245 213.77 43.315 ;
    RECT 213.56 43.605 213.77 43.675 ;
    RECT 213.56 43.965 213.77 44.035 ;
    RECT 213.1 43.245 213.31 43.315 ;
    RECT 213.1 43.605 213.31 43.675 ;
    RECT 213.1 43.965 213.31 44.035 ;
    RECT 346.36 43.245 346.57 43.315 ;
    RECT 346.36 43.605 346.57 43.675 ;
    RECT 346.36 43.965 346.57 44.035 ;
    RECT 345.9 43.245 346.11 43.315 ;
    RECT 345.9 43.605 346.11 43.675 ;
    RECT 345.9 43.965 346.11 44.035 ;
    RECT 210.24 43.245 210.45 43.315 ;
    RECT 210.24 43.605 210.45 43.675 ;
    RECT 210.24 43.965 210.45 44.035 ;
    RECT 209.78 43.245 209.99 43.315 ;
    RECT 209.78 43.605 209.99 43.675 ;
    RECT 209.78 43.965 209.99 44.035 ;
    RECT 343.04 43.245 343.25 43.315 ;
    RECT 343.04 43.605 343.25 43.675 ;
    RECT 343.04 43.965 343.25 44.035 ;
    RECT 342.58 43.245 342.79 43.315 ;
    RECT 342.58 43.605 342.79 43.675 ;
    RECT 342.58 43.965 342.79 44.035 ;
    RECT 206.92 43.245 207.13 43.315 ;
    RECT 206.92 43.605 207.13 43.675 ;
    RECT 206.92 43.965 207.13 44.035 ;
    RECT 206.46 43.245 206.67 43.315 ;
    RECT 206.46 43.605 206.67 43.675 ;
    RECT 206.46 43.965 206.67 44.035 ;
    RECT 339.72 43.245 339.93 43.315 ;
    RECT 339.72 43.605 339.93 43.675 ;
    RECT 339.72 43.965 339.93 44.035 ;
    RECT 339.26 43.245 339.47 43.315 ;
    RECT 339.26 43.605 339.47 43.675 ;
    RECT 339.26 43.965 339.47 44.035 ;
    RECT 203.6 43.245 203.81 43.315 ;
    RECT 203.6 43.605 203.81 43.675 ;
    RECT 203.6 43.965 203.81 44.035 ;
    RECT 203.14 43.245 203.35 43.315 ;
    RECT 203.14 43.605 203.35 43.675 ;
    RECT 203.14 43.965 203.35 44.035 ;
    RECT 336.4 43.245 336.61 43.315 ;
    RECT 336.4 43.605 336.61 43.675 ;
    RECT 336.4 43.965 336.61 44.035 ;
    RECT 335.94 43.245 336.15 43.315 ;
    RECT 335.94 43.605 336.15 43.675 ;
    RECT 335.94 43.965 336.15 44.035 ;
    RECT 266.68 43.245 266.89 43.315 ;
    RECT 266.68 43.605 266.89 43.675 ;
    RECT 266.68 43.965 266.89 44.035 ;
    RECT 266.22 43.245 266.43 43.315 ;
    RECT 266.22 43.605 266.43 43.675 ;
    RECT 266.22 43.965 266.43 44.035 ;
    RECT 263.36 43.245 263.57 43.315 ;
    RECT 263.36 43.605 263.57 43.675 ;
    RECT 263.36 43.965 263.57 44.035 ;
    RECT 262.9 43.245 263.11 43.315 ;
    RECT 262.9 43.605 263.11 43.675 ;
    RECT 262.9 43.965 263.11 44.035 ;
    RECT 260.04 43.245 260.25 43.315 ;
    RECT 260.04 43.605 260.25 43.675 ;
    RECT 260.04 43.965 260.25 44.035 ;
    RECT 259.58 43.245 259.79 43.315 ;
    RECT 259.58 43.605 259.79 43.675 ;
    RECT 259.58 43.965 259.79 44.035 ;
    RECT 256.72 43.245 256.93 43.315 ;
    RECT 256.72 43.605 256.93 43.675 ;
    RECT 256.72 43.965 256.93 44.035 ;
    RECT 256.26 43.245 256.47 43.315 ;
    RECT 256.26 43.605 256.47 43.675 ;
    RECT 256.26 43.965 256.47 44.035 ;
    RECT 253.4 43.245 253.61 43.315 ;
    RECT 253.4 43.605 253.61 43.675 ;
    RECT 253.4 43.965 253.61 44.035 ;
    RECT 252.94 43.245 253.15 43.315 ;
    RECT 252.94 43.605 253.15 43.675 ;
    RECT 252.94 43.965 253.15 44.035 ;
    RECT 250.08 43.245 250.29 43.315 ;
    RECT 250.08 43.605 250.29 43.675 ;
    RECT 250.08 43.965 250.29 44.035 ;
    RECT 249.62 43.245 249.83 43.315 ;
    RECT 249.62 43.605 249.83 43.675 ;
    RECT 249.62 43.965 249.83 44.035 ;
    RECT 246.76 43.245 246.97 43.315 ;
    RECT 246.76 43.605 246.97 43.675 ;
    RECT 246.76 43.965 246.97 44.035 ;
    RECT 246.3 43.245 246.51 43.315 ;
    RECT 246.3 43.605 246.51 43.675 ;
    RECT 246.3 43.965 246.51 44.035 ;
    RECT 243.44 43.245 243.65 43.315 ;
    RECT 243.44 43.605 243.65 43.675 ;
    RECT 243.44 43.965 243.65 44.035 ;
    RECT 242.98 43.245 243.19 43.315 ;
    RECT 242.98 43.605 243.19 43.675 ;
    RECT 242.98 43.965 243.19 44.035 ;
    RECT 240.12 43.245 240.33 43.315 ;
    RECT 240.12 43.605 240.33 43.675 ;
    RECT 240.12 43.965 240.33 44.035 ;
    RECT 239.66 43.245 239.87 43.315 ;
    RECT 239.66 43.605 239.87 43.675 ;
    RECT 239.66 43.965 239.87 44.035 ;
    RECT 236.8 43.245 237.01 43.315 ;
    RECT 236.8 43.605 237.01 43.675 ;
    RECT 236.8 43.965 237.01 44.035 ;
    RECT 236.34 43.245 236.55 43.315 ;
    RECT 236.34 43.605 236.55 43.675 ;
    RECT 236.34 43.965 236.55 44.035 ;
    RECT 374.15 43.605 374.22 43.675 ;
    RECT 333.08 43.245 333.29 43.315 ;
    RECT 333.08 43.605 333.29 43.675 ;
    RECT 333.08 43.965 333.29 44.035 ;
    RECT 332.62 43.245 332.83 43.315 ;
    RECT 332.62 43.605 332.83 43.675 ;
    RECT 332.62 43.965 332.83 44.035 ;
    RECT 329.76 43.245 329.97 43.315 ;
    RECT 329.76 43.605 329.97 43.675 ;
    RECT 329.76 43.965 329.97 44.035 ;
    RECT 329.3 43.245 329.51 43.315 ;
    RECT 329.3 43.605 329.51 43.675 ;
    RECT 329.3 43.965 329.51 44.035 ;
    RECT 326.44 43.245 326.65 43.315 ;
    RECT 326.44 43.605 326.65 43.675 ;
    RECT 326.44 43.965 326.65 44.035 ;
    RECT 325.98 43.245 326.19 43.315 ;
    RECT 325.98 43.605 326.19 43.675 ;
    RECT 325.98 43.965 326.19 44.035 ;
    RECT 323.12 43.245 323.33 43.315 ;
    RECT 323.12 43.605 323.33 43.675 ;
    RECT 323.12 43.965 323.33 44.035 ;
    RECT 322.66 43.245 322.87 43.315 ;
    RECT 322.66 43.605 322.87 43.675 ;
    RECT 322.66 43.965 322.87 44.035 ;
    RECT 319.8 43.245 320.01 43.315 ;
    RECT 319.8 43.605 320.01 43.675 ;
    RECT 319.8 43.965 320.01 44.035 ;
    RECT 319.34 43.245 319.55 43.315 ;
    RECT 319.34 43.605 319.55 43.675 ;
    RECT 319.34 43.965 319.55 44.035 ;
    RECT 316.48 43.245 316.69 43.315 ;
    RECT 316.48 43.605 316.69 43.675 ;
    RECT 316.48 43.965 316.69 44.035 ;
    RECT 316.02 43.245 316.23 43.315 ;
    RECT 316.02 43.605 316.23 43.675 ;
    RECT 316.02 43.965 316.23 44.035 ;
    RECT 313.16 43.245 313.37 43.315 ;
    RECT 313.16 43.605 313.37 43.675 ;
    RECT 313.16 43.965 313.37 44.035 ;
    RECT 312.7 43.245 312.91 43.315 ;
    RECT 312.7 43.605 312.91 43.675 ;
    RECT 312.7 43.965 312.91 44.035 ;
    RECT 309.84 43.245 310.05 43.315 ;
    RECT 309.84 43.605 310.05 43.675 ;
    RECT 309.84 43.965 310.05 44.035 ;
    RECT 309.38 43.245 309.59 43.315 ;
    RECT 309.38 43.605 309.59 43.675 ;
    RECT 309.38 43.965 309.59 44.035 ;
    RECT 306.52 43.245 306.73 43.315 ;
    RECT 306.52 43.605 306.73 43.675 ;
    RECT 306.52 43.965 306.73 44.035 ;
    RECT 306.06 43.245 306.27 43.315 ;
    RECT 306.06 43.605 306.27 43.675 ;
    RECT 306.06 43.965 306.27 44.035 ;
    RECT 303.2 42.525 303.41 42.595 ;
    RECT 303.2 42.885 303.41 42.955 ;
    RECT 303.2 43.245 303.41 43.315 ;
    RECT 302.74 42.525 302.95 42.595 ;
    RECT 302.74 42.885 302.95 42.955 ;
    RECT 302.74 43.245 302.95 43.315 ;
    RECT 372.92 42.525 373.13 42.595 ;
    RECT 372.92 42.885 373.13 42.955 ;
    RECT 372.92 43.245 373.13 43.315 ;
    RECT 372.46 42.525 372.67 42.595 ;
    RECT 372.46 42.885 372.67 42.955 ;
    RECT 372.46 43.245 372.67 43.315 ;
    RECT 369.6 42.525 369.81 42.595 ;
    RECT 369.6 42.885 369.81 42.955 ;
    RECT 369.6 43.245 369.81 43.315 ;
    RECT 369.14 42.525 369.35 42.595 ;
    RECT 369.14 42.885 369.35 42.955 ;
    RECT 369.14 43.245 369.35 43.315 ;
    RECT 200.605 42.885 200.675 42.955 ;
    RECT 299.88 42.525 300.09 42.595 ;
    RECT 299.88 42.885 300.09 42.955 ;
    RECT 299.88 43.245 300.09 43.315 ;
    RECT 299.42 42.525 299.63 42.595 ;
    RECT 299.42 42.885 299.63 42.955 ;
    RECT 299.42 43.245 299.63 43.315 ;
    RECT 296.56 42.525 296.77 42.595 ;
    RECT 296.56 42.885 296.77 42.955 ;
    RECT 296.56 43.245 296.77 43.315 ;
    RECT 296.1 42.525 296.31 42.595 ;
    RECT 296.1 42.885 296.31 42.955 ;
    RECT 296.1 43.245 296.31 43.315 ;
    RECT 293.24 42.525 293.45 42.595 ;
    RECT 293.24 42.885 293.45 42.955 ;
    RECT 293.24 43.245 293.45 43.315 ;
    RECT 292.78 42.525 292.99 42.595 ;
    RECT 292.78 42.885 292.99 42.955 ;
    RECT 292.78 43.245 292.99 43.315 ;
    RECT 289.92 42.525 290.13 42.595 ;
    RECT 289.92 42.885 290.13 42.955 ;
    RECT 289.92 43.245 290.13 43.315 ;
    RECT 289.46 42.525 289.67 42.595 ;
    RECT 289.46 42.885 289.67 42.955 ;
    RECT 289.46 43.245 289.67 43.315 ;
    RECT 286.6 42.525 286.81 42.595 ;
    RECT 286.6 42.885 286.81 42.955 ;
    RECT 286.6 43.245 286.81 43.315 ;
    RECT 286.14 42.525 286.35 42.595 ;
    RECT 286.14 42.885 286.35 42.955 ;
    RECT 286.14 43.245 286.35 43.315 ;
    RECT 283.28 42.525 283.49 42.595 ;
    RECT 283.28 42.885 283.49 42.955 ;
    RECT 283.28 43.245 283.49 43.315 ;
    RECT 282.82 42.525 283.03 42.595 ;
    RECT 282.82 42.885 283.03 42.955 ;
    RECT 282.82 43.245 283.03 43.315 ;
    RECT 279.96 42.525 280.17 42.595 ;
    RECT 279.96 42.885 280.17 42.955 ;
    RECT 279.96 43.245 280.17 43.315 ;
    RECT 279.5 42.525 279.71 42.595 ;
    RECT 279.5 42.885 279.71 42.955 ;
    RECT 279.5 43.245 279.71 43.315 ;
    RECT 276.64 42.525 276.85 42.595 ;
    RECT 276.64 42.885 276.85 42.955 ;
    RECT 276.64 43.245 276.85 43.315 ;
    RECT 276.18 42.525 276.39 42.595 ;
    RECT 276.18 42.885 276.39 42.955 ;
    RECT 276.18 43.245 276.39 43.315 ;
    RECT 273.32 42.525 273.53 42.595 ;
    RECT 273.32 42.885 273.53 42.955 ;
    RECT 273.32 43.245 273.53 43.315 ;
    RECT 272.86 42.525 273.07 42.595 ;
    RECT 272.86 42.885 273.07 42.955 ;
    RECT 272.86 43.245 273.07 43.315 ;
    RECT 270.0 42.525 270.21 42.595 ;
    RECT 270.0 42.885 270.21 42.955 ;
    RECT 270.0 43.245 270.21 43.315 ;
    RECT 269.54 42.525 269.75 42.595 ;
    RECT 269.54 42.885 269.75 42.955 ;
    RECT 269.54 43.245 269.75 43.315 ;
    RECT 233.48 42.525 233.69 42.595 ;
    RECT 233.48 42.885 233.69 42.955 ;
    RECT 233.48 43.245 233.69 43.315 ;
    RECT 233.02 42.525 233.23 42.595 ;
    RECT 233.02 42.885 233.23 42.955 ;
    RECT 233.02 43.245 233.23 43.315 ;
    RECT 230.16 42.525 230.37 42.595 ;
    RECT 230.16 42.885 230.37 42.955 ;
    RECT 230.16 43.245 230.37 43.315 ;
    RECT 229.7 42.525 229.91 42.595 ;
    RECT 229.7 42.885 229.91 42.955 ;
    RECT 229.7 43.245 229.91 43.315 ;
    RECT 366.28 42.525 366.49 42.595 ;
    RECT 366.28 42.885 366.49 42.955 ;
    RECT 366.28 43.245 366.49 43.315 ;
    RECT 365.82 42.525 366.03 42.595 ;
    RECT 365.82 42.885 366.03 42.955 ;
    RECT 365.82 43.245 366.03 43.315 ;
    RECT 226.84 42.525 227.05 42.595 ;
    RECT 226.84 42.885 227.05 42.955 ;
    RECT 226.84 43.245 227.05 43.315 ;
    RECT 226.38 42.525 226.59 42.595 ;
    RECT 226.38 42.885 226.59 42.955 ;
    RECT 226.38 43.245 226.59 43.315 ;
    RECT 362.96 42.525 363.17 42.595 ;
    RECT 362.96 42.885 363.17 42.955 ;
    RECT 362.96 43.245 363.17 43.315 ;
    RECT 362.5 42.525 362.71 42.595 ;
    RECT 362.5 42.885 362.71 42.955 ;
    RECT 362.5 43.245 362.71 43.315 ;
    RECT 223.52 42.525 223.73 42.595 ;
    RECT 223.52 42.885 223.73 42.955 ;
    RECT 223.52 43.245 223.73 43.315 ;
    RECT 223.06 42.525 223.27 42.595 ;
    RECT 223.06 42.885 223.27 42.955 ;
    RECT 223.06 43.245 223.27 43.315 ;
    RECT 359.64 42.525 359.85 42.595 ;
    RECT 359.64 42.885 359.85 42.955 ;
    RECT 359.64 43.245 359.85 43.315 ;
    RECT 359.18 42.525 359.39 42.595 ;
    RECT 359.18 42.885 359.39 42.955 ;
    RECT 359.18 43.245 359.39 43.315 ;
    RECT 220.2 42.525 220.41 42.595 ;
    RECT 220.2 42.885 220.41 42.955 ;
    RECT 220.2 43.245 220.41 43.315 ;
    RECT 219.74 42.525 219.95 42.595 ;
    RECT 219.74 42.885 219.95 42.955 ;
    RECT 219.74 43.245 219.95 43.315 ;
    RECT 356.32 42.525 356.53 42.595 ;
    RECT 356.32 42.885 356.53 42.955 ;
    RECT 356.32 43.245 356.53 43.315 ;
    RECT 355.86 42.525 356.07 42.595 ;
    RECT 355.86 42.885 356.07 42.955 ;
    RECT 355.86 43.245 356.07 43.315 ;
    RECT 353.0 42.525 353.21 42.595 ;
    RECT 353.0 42.885 353.21 42.955 ;
    RECT 353.0 43.245 353.21 43.315 ;
    RECT 352.54 42.525 352.75 42.595 ;
    RECT 352.54 42.885 352.75 42.955 ;
    RECT 352.54 43.245 352.75 43.315 ;
    RECT 216.88 42.525 217.09 42.595 ;
    RECT 216.88 42.885 217.09 42.955 ;
    RECT 216.88 43.245 217.09 43.315 ;
    RECT 216.42 42.525 216.63 42.595 ;
    RECT 216.42 42.885 216.63 42.955 ;
    RECT 216.42 43.245 216.63 43.315 ;
    RECT 349.68 42.525 349.89 42.595 ;
    RECT 349.68 42.885 349.89 42.955 ;
    RECT 349.68 43.245 349.89 43.315 ;
    RECT 349.22 42.525 349.43 42.595 ;
    RECT 349.22 42.885 349.43 42.955 ;
    RECT 349.22 43.245 349.43 43.315 ;
    RECT 213.56 42.525 213.77 42.595 ;
    RECT 213.56 42.885 213.77 42.955 ;
    RECT 213.56 43.245 213.77 43.315 ;
    RECT 213.1 42.525 213.31 42.595 ;
    RECT 213.1 42.885 213.31 42.955 ;
    RECT 213.1 43.245 213.31 43.315 ;
    RECT 346.36 42.525 346.57 42.595 ;
    RECT 346.36 42.885 346.57 42.955 ;
    RECT 346.36 43.245 346.57 43.315 ;
    RECT 345.9 42.525 346.11 42.595 ;
    RECT 345.9 42.885 346.11 42.955 ;
    RECT 345.9 43.245 346.11 43.315 ;
    RECT 210.24 42.525 210.45 42.595 ;
    RECT 210.24 42.885 210.45 42.955 ;
    RECT 210.24 43.245 210.45 43.315 ;
    RECT 209.78 42.525 209.99 42.595 ;
    RECT 209.78 42.885 209.99 42.955 ;
    RECT 209.78 43.245 209.99 43.315 ;
    RECT 343.04 42.525 343.25 42.595 ;
    RECT 343.04 42.885 343.25 42.955 ;
    RECT 343.04 43.245 343.25 43.315 ;
    RECT 342.58 42.525 342.79 42.595 ;
    RECT 342.58 42.885 342.79 42.955 ;
    RECT 342.58 43.245 342.79 43.315 ;
    RECT 206.92 42.525 207.13 42.595 ;
    RECT 206.92 42.885 207.13 42.955 ;
    RECT 206.92 43.245 207.13 43.315 ;
    RECT 206.46 42.525 206.67 42.595 ;
    RECT 206.46 42.885 206.67 42.955 ;
    RECT 206.46 43.245 206.67 43.315 ;
    RECT 339.72 42.525 339.93 42.595 ;
    RECT 339.72 42.885 339.93 42.955 ;
    RECT 339.72 43.245 339.93 43.315 ;
    RECT 339.26 42.525 339.47 42.595 ;
    RECT 339.26 42.885 339.47 42.955 ;
    RECT 339.26 43.245 339.47 43.315 ;
    RECT 203.6 42.525 203.81 42.595 ;
    RECT 203.6 42.885 203.81 42.955 ;
    RECT 203.6 43.245 203.81 43.315 ;
    RECT 203.14 42.525 203.35 42.595 ;
    RECT 203.14 42.885 203.35 42.955 ;
    RECT 203.14 43.245 203.35 43.315 ;
    RECT 336.4 42.525 336.61 42.595 ;
    RECT 336.4 42.885 336.61 42.955 ;
    RECT 336.4 43.245 336.61 43.315 ;
    RECT 335.94 42.525 336.15 42.595 ;
    RECT 335.94 42.885 336.15 42.955 ;
    RECT 335.94 43.245 336.15 43.315 ;
    RECT 266.68 42.525 266.89 42.595 ;
    RECT 266.68 42.885 266.89 42.955 ;
    RECT 266.68 43.245 266.89 43.315 ;
    RECT 266.22 42.525 266.43 42.595 ;
    RECT 266.22 42.885 266.43 42.955 ;
    RECT 266.22 43.245 266.43 43.315 ;
    RECT 263.36 42.525 263.57 42.595 ;
    RECT 263.36 42.885 263.57 42.955 ;
    RECT 263.36 43.245 263.57 43.315 ;
    RECT 262.9 42.525 263.11 42.595 ;
    RECT 262.9 42.885 263.11 42.955 ;
    RECT 262.9 43.245 263.11 43.315 ;
    RECT 260.04 42.525 260.25 42.595 ;
    RECT 260.04 42.885 260.25 42.955 ;
    RECT 260.04 43.245 260.25 43.315 ;
    RECT 259.58 42.525 259.79 42.595 ;
    RECT 259.58 42.885 259.79 42.955 ;
    RECT 259.58 43.245 259.79 43.315 ;
    RECT 256.72 42.525 256.93 42.595 ;
    RECT 256.72 42.885 256.93 42.955 ;
    RECT 256.72 43.245 256.93 43.315 ;
    RECT 256.26 42.525 256.47 42.595 ;
    RECT 256.26 42.885 256.47 42.955 ;
    RECT 256.26 43.245 256.47 43.315 ;
    RECT 253.4 42.525 253.61 42.595 ;
    RECT 253.4 42.885 253.61 42.955 ;
    RECT 253.4 43.245 253.61 43.315 ;
    RECT 252.94 42.525 253.15 42.595 ;
    RECT 252.94 42.885 253.15 42.955 ;
    RECT 252.94 43.245 253.15 43.315 ;
    RECT 250.08 42.525 250.29 42.595 ;
    RECT 250.08 42.885 250.29 42.955 ;
    RECT 250.08 43.245 250.29 43.315 ;
    RECT 249.62 42.525 249.83 42.595 ;
    RECT 249.62 42.885 249.83 42.955 ;
    RECT 249.62 43.245 249.83 43.315 ;
    RECT 246.76 42.525 246.97 42.595 ;
    RECT 246.76 42.885 246.97 42.955 ;
    RECT 246.76 43.245 246.97 43.315 ;
    RECT 246.3 42.525 246.51 42.595 ;
    RECT 246.3 42.885 246.51 42.955 ;
    RECT 246.3 43.245 246.51 43.315 ;
    RECT 243.44 42.525 243.65 42.595 ;
    RECT 243.44 42.885 243.65 42.955 ;
    RECT 243.44 43.245 243.65 43.315 ;
    RECT 242.98 42.525 243.19 42.595 ;
    RECT 242.98 42.885 243.19 42.955 ;
    RECT 242.98 43.245 243.19 43.315 ;
    RECT 240.12 42.525 240.33 42.595 ;
    RECT 240.12 42.885 240.33 42.955 ;
    RECT 240.12 43.245 240.33 43.315 ;
    RECT 239.66 42.525 239.87 42.595 ;
    RECT 239.66 42.885 239.87 42.955 ;
    RECT 239.66 43.245 239.87 43.315 ;
    RECT 236.8 42.525 237.01 42.595 ;
    RECT 236.8 42.885 237.01 42.955 ;
    RECT 236.8 43.245 237.01 43.315 ;
    RECT 236.34 42.525 236.55 42.595 ;
    RECT 236.34 42.885 236.55 42.955 ;
    RECT 236.34 43.245 236.55 43.315 ;
    RECT 374.15 42.885 374.22 42.955 ;
    RECT 333.08 42.525 333.29 42.595 ;
    RECT 333.08 42.885 333.29 42.955 ;
    RECT 333.08 43.245 333.29 43.315 ;
    RECT 332.62 42.525 332.83 42.595 ;
    RECT 332.62 42.885 332.83 42.955 ;
    RECT 332.62 43.245 332.83 43.315 ;
    RECT 329.76 42.525 329.97 42.595 ;
    RECT 329.76 42.885 329.97 42.955 ;
    RECT 329.76 43.245 329.97 43.315 ;
    RECT 329.3 42.525 329.51 42.595 ;
    RECT 329.3 42.885 329.51 42.955 ;
    RECT 329.3 43.245 329.51 43.315 ;
    RECT 326.44 42.525 326.65 42.595 ;
    RECT 326.44 42.885 326.65 42.955 ;
    RECT 326.44 43.245 326.65 43.315 ;
    RECT 325.98 42.525 326.19 42.595 ;
    RECT 325.98 42.885 326.19 42.955 ;
    RECT 325.98 43.245 326.19 43.315 ;
    RECT 323.12 42.525 323.33 42.595 ;
    RECT 323.12 42.885 323.33 42.955 ;
    RECT 323.12 43.245 323.33 43.315 ;
    RECT 322.66 42.525 322.87 42.595 ;
    RECT 322.66 42.885 322.87 42.955 ;
    RECT 322.66 43.245 322.87 43.315 ;
    RECT 319.8 42.525 320.01 42.595 ;
    RECT 319.8 42.885 320.01 42.955 ;
    RECT 319.8 43.245 320.01 43.315 ;
    RECT 319.34 42.525 319.55 42.595 ;
    RECT 319.34 42.885 319.55 42.955 ;
    RECT 319.34 43.245 319.55 43.315 ;
    RECT 316.48 42.525 316.69 42.595 ;
    RECT 316.48 42.885 316.69 42.955 ;
    RECT 316.48 43.245 316.69 43.315 ;
    RECT 316.02 42.525 316.23 42.595 ;
    RECT 316.02 42.885 316.23 42.955 ;
    RECT 316.02 43.245 316.23 43.315 ;
    RECT 313.16 42.525 313.37 42.595 ;
    RECT 313.16 42.885 313.37 42.955 ;
    RECT 313.16 43.245 313.37 43.315 ;
    RECT 312.7 42.525 312.91 42.595 ;
    RECT 312.7 42.885 312.91 42.955 ;
    RECT 312.7 43.245 312.91 43.315 ;
    RECT 309.84 42.525 310.05 42.595 ;
    RECT 309.84 42.885 310.05 42.955 ;
    RECT 309.84 43.245 310.05 43.315 ;
    RECT 309.38 42.525 309.59 42.595 ;
    RECT 309.38 42.885 309.59 42.955 ;
    RECT 309.38 43.245 309.59 43.315 ;
    RECT 306.52 42.525 306.73 42.595 ;
    RECT 306.52 42.885 306.73 42.955 ;
    RECT 306.52 43.245 306.73 43.315 ;
    RECT 306.06 42.525 306.27 42.595 ;
    RECT 306.06 42.885 306.27 42.955 ;
    RECT 306.06 43.245 306.27 43.315 ;
    RECT 303.2 41.805 303.41 41.875 ;
    RECT 303.2 42.165 303.41 42.235 ;
    RECT 303.2 42.525 303.41 42.595 ;
    RECT 302.74 41.805 302.95 41.875 ;
    RECT 302.74 42.165 302.95 42.235 ;
    RECT 302.74 42.525 302.95 42.595 ;
    RECT 372.92 41.805 373.13 41.875 ;
    RECT 372.92 42.165 373.13 42.235 ;
    RECT 372.92 42.525 373.13 42.595 ;
    RECT 372.46 41.805 372.67 41.875 ;
    RECT 372.46 42.165 372.67 42.235 ;
    RECT 372.46 42.525 372.67 42.595 ;
    RECT 369.6 41.805 369.81 41.875 ;
    RECT 369.6 42.165 369.81 42.235 ;
    RECT 369.6 42.525 369.81 42.595 ;
    RECT 369.14 41.805 369.35 41.875 ;
    RECT 369.14 42.165 369.35 42.235 ;
    RECT 369.14 42.525 369.35 42.595 ;
    RECT 200.605 42.165 200.675 42.235 ;
    RECT 299.88 41.805 300.09 41.875 ;
    RECT 299.88 42.165 300.09 42.235 ;
    RECT 299.88 42.525 300.09 42.595 ;
    RECT 299.42 41.805 299.63 41.875 ;
    RECT 299.42 42.165 299.63 42.235 ;
    RECT 299.42 42.525 299.63 42.595 ;
    RECT 296.56 41.805 296.77 41.875 ;
    RECT 296.56 42.165 296.77 42.235 ;
    RECT 296.56 42.525 296.77 42.595 ;
    RECT 296.1 41.805 296.31 41.875 ;
    RECT 296.1 42.165 296.31 42.235 ;
    RECT 296.1 42.525 296.31 42.595 ;
    RECT 293.24 41.805 293.45 41.875 ;
    RECT 293.24 42.165 293.45 42.235 ;
    RECT 293.24 42.525 293.45 42.595 ;
    RECT 292.78 41.805 292.99 41.875 ;
    RECT 292.78 42.165 292.99 42.235 ;
    RECT 292.78 42.525 292.99 42.595 ;
    RECT 289.92 41.805 290.13 41.875 ;
    RECT 289.92 42.165 290.13 42.235 ;
    RECT 289.92 42.525 290.13 42.595 ;
    RECT 289.46 41.805 289.67 41.875 ;
    RECT 289.46 42.165 289.67 42.235 ;
    RECT 289.46 42.525 289.67 42.595 ;
    RECT 286.6 41.805 286.81 41.875 ;
    RECT 286.6 42.165 286.81 42.235 ;
    RECT 286.6 42.525 286.81 42.595 ;
    RECT 286.14 41.805 286.35 41.875 ;
    RECT 286.14 42.165 286.35 42.235 ;
    RECT 286.14 42.525 286.35 42.595 ;
    RECT 283.28 41.805 283.49 41.875 ;
    RECT 283.28 42.165 283.49 42.235 ;
    RECT 283.28 42.525 283.49 42.595 ;
    RECT 282.82 41.805 283.03 41.875 ;
    RECT 282.82 42.165 283.03 42.235 ;
    RECT 282.82 42.525 283.03 42.595 ;
    RECT 279.96 41.805 280.17 41.875 ;
    RECT 279.96 42.165 280.17 42.235 ;
    RECT 279.96 42.525 280.17 42.595 ;
    RECT 279.5 41.805 279.71 41.875 ;
    RECT 279.5 42.165 279.71 42.235 ;
    RECT 279.5 42.525 279.71 42.595 ;
    RECT 276.64 41.805 276.85 41.875 ;
    RECT 276.64 42.165 276.85 42.235 ;
    RECT 276.64 42.525 276.85 42.595 ;
    RECT 276.18 41.805 276.39 41.875 ;
    RECT 276.18 42.165 276.39 42.235 ;
    RECT 276.18 42.525 276.39 42.595 ;
    RECT 273.32 41.805 273.53 41.875 ;
    RECT 273.32 42.165 273.53 42.235 ;
    RECT 273.32 42.525 273.53 42.595 ;
    RECT 272.86 41.805 273.07 41.875 ;
    RECT 272.86 42.165 273.07 42.235 ;
    RECT 272.86 42.525 273.07 42.595 ;
    RECT 270.0 41.805 270.21 41.875 ;
    RECT 270.0 42.165 270.21 42.235 ;
    RECT 270.0 42.525 270.21 42.595 ;
    RECT 269.54 41.805 269.75 41.875 ;
    RECT 269.54 42.165 269.75 42.235 ;
    RECT 269.54 42.525 269.75 42.595 ;
    RECT 233.48 41.805 233.69 41.875 ;
    RECT 233.48 42.165 233.69 42.235 ;
    RECT 233.48 42.525 233.69 42.595 ;
    RECT 233.02 41.805 233.23 41.875 ;
    RECT 233.02 42.165 233.23 42.235 ;
    RECT 233.02 42.525 233.23 42.595 ;
    RECT 230.16 41.805 230.37 41.875 ;
    RECT 230.16 42.165 230.37 42.235 ;
    RECT 230.16 42.525 230.37 42.595 ;
    RECT 229.7 41.805 229.91 41.875 ;
    RECT 229.7 42.165 229.91 42.235 ;
    RECT 229.7 42.525 229.91 42.595 ;
    RECT 366.28 41.805 366.49 41.875 ;
    RECT 366.28 42.165 366.49 42.235 ;
    RECT 366.28 42.525 366.49 42.595 ;
    RECT 365.82 41.805 366.03 41.875 ;
    RECT 365.82 42.165 366.03 42.235 ;
    RECT 365.82 42.525 366.03 42.595 ;
    RECT 226.84 41.805 227.05 41.875 ;
    RECT 226.84 42.165 227.05 42.235 ;
    RECT 226.84 42.525 227.05 42.595 ;
    RECT 226.38 41.805 226.59 41.875 ;
    RECT 226.38 42.165 226.59 42.235 ;
    RECT 226.38 42.525 226.59 42.595 ;
    RECT 362.96 41.805 363.17 41.875 ;
    RECT 362.96 42.165 363.17 42.235 ;
    RECT 362.96 42.525 363.17 42.595 ;
    RECT 362.5 41.805 362.71 41.875 ;
    RECT 362.5 42.165 362.71 42.235 ;
    RECT 362.5 42.525 362.71 42.595 ;
    RECT 223.52 41.805 223.73 41.875 ;
    RECT 223.52 42.165 223.73 42.235 ;
    RECT 223.52 42.525 223.73 42.595 ;
    RECT 223.06 41.805 223.27 41.875 ;
    RECT 223.06 42.165 223.27 42.235 ;
    RECT 223.06 42.525 223.27 42.595 ;
    RECT 359.64 41.805 359.85 41.875 ;
    RECT 359.64 42.165 359.85 42.235 ;
    RECT 359.64 42.525 359.85 42.595 ;
    RECT 359.18 41.805 359.39 41.875 ;
    RECT 359.18 42.165 359.39 42.235 ;
    RECT 359.18 42.525 359.39 42.595 ;
    RECT 220.2 41.805 220.41 41.875 ;
    RECT 220.2 42.165 220.41 42.235 ;
    RECT 220.2 42.525 220.41 42.595 ;
    RECT 219.74 41.805 219.95 41.875 ;
    RECT 219.74 42.165 219.95 42.235 ;
    RECT 219.74 42.525 219.95 42.595 ;
    RECT 356.32 41.805 356.53 41.875 ;
    RECT 356.32 42.165 356.53 42.235 ;
    RECT 356.32 42.525 356.53 42.595 ;
    RECT 355.86 41.805 356.07 41.875 ;
    RECT 355.86 42.165 356.07 42.235 ;
    RECT 355.86 42.525 356.07 42.595 ;
    RECT 353.0 41.805 353.21 41.875 ;
    RECT 353.0 42.165 353.21 42.235 ;
    RECT 353.0 42.525 353.21 42.595 ;
    RECT 352.54 41.805 352.75 41.875 ;
    RECT 352.54 42.165 352.75 42.235 ;
    RECT 352.54 42.525 352.75 42.595 ;
    RECT 216.88 41.805 217.09 41.875 ;
    RECT 216.88 42.165 217.09 42.235 ;
    RECT 216.88 42.525 217.09 42.595 ;
    RECT 216.42 41.805 216.63 41.875 ;
    RECT 216.42 42.165 216.63 42.235 ;
    RECT 216.42 42.525 216.63 42.595 ;
    RECT 349.68 41.805 349.89 41.875 ;
    RECT 349.68 42.165 349.89 42.235 ;
    RECT 349.68 42.525 349.89 42.595 ;
    RECT 349.22 41.805 349.43 41.875 ;
    RECT 349.22 42.165 349.43 42.235 ;
    RECT 349.22 42.525 349.43 42.595 ;
    RECT 213.56 41.805 213.77 41.875 ;
    RECT 213.56 42.165 213.77 42.235 ;
    RECT 213.56 42.525 213.77 42.595 ;
    RECT 213.1 41.805 213.31 41.875 ;
    RECT 213.1 42.165 213.31 42.235 ;
    RECT 213.1 42.525 213.31 42.595 ;
    RECT 346.36 41.805 346.57 41.875 ;
    RECT 346.36 42.165 346.57 42.235 ;
    RECT 346.36 42.525 346.57 42.595 ;
    RECT 345.9 41.805 346.11 41.875 ;
    RECT 345.9 42.165 346.11 42.235 ;
    RECT 345.9 42.525 346.11 42.595 ;
    RECT 210.24 41.805 210.45 41.875 ;
    RECT 210.24 42.165 210.45 42.235 ;
    RECT 210.24 42.525 210.45 42.595 ;
    RECT 209.78 41.805 209.99 41.875 ;
    RECT 209.78 42.165 209.99 42.235 ;
    RECT 209.78 42.525 209.99 42.595 ;
    RECT 343.04 41.805 343.25 41.875 ;
    RECT 343.04 42.165 343.25 42.235 ;
    RECT 343.04 42.525 343.25 42.595 ;
    RECT 342.58 41.805 342.79 41.875 ;
    RECT 342.58 42.165 342.79 42.235 ;
    RECT 342.58 42.525 342.79 42.595 ;
    RECT 206.92 41.805 207.13 41.875 ;
    RECT 206.92 42.165 207.13 42.235 ;
    RECT 206.92 42.525 207.13 42.595 ;
    RECT 206.46 41.805 206.67 41.875 ;
    RECT 206.46 42.165 206.67 42.235 ;
    RECT 206.46 42.525 206.67 42.595 ;
    RECT 339.72 41.805 339.93 41.875 ;
    RECT 339.72 42.165 339.93 42.235 ;
    RECT 339.72 42.525 339.93 42.595 ;
    RECT 339.26 41.805 339.47 41.875 ;
    RECT 339.26 42.165 339.47 42.235 ;
    RECT 339.26 42.525 339.47 42.595 ;
    RECT 203.6 41.805 203.81 41.875 ;
    RECT 203.6 42.165 203.81 42.235 ;
    RECT 203.6 42.525 203.81 42.595 ;
    RECT 203.14 41.805 203.35 41.875 ;
    RECT 203.14 42.165 203.35 42.235 ;
    RECT 203.14 42.525 203.35 42.595 ;
    RECT 336.4 41.805 336.61 41.875 ;
    RECT 336.4 42.165 336.61 42.235 ;
    RECT 336.4 42.525 336.61 42.595 ;
    RECT 335.94 41.805 336.15 41.875 ;
    RECT 335.94 42.165 336.15 42.235 ;
    RECT 335.94 42.525 336.15 42.595 ;
    RECT 266.68 41.805 266.89 41.875 ;
    RECT 266.68 42.165 266.89 42.235 ;
    RECT 266.68 42.525 266.89 42.595 ;
    RECT 266.22 41.805 266.43 41.875 ;
    RECT 266.22 42.165 266.43 42.235 ;
    RECT 266.22 42.525 266.43 42.595 ;
    RECT 263.36 41.805 263.57 41.875 ;
    RECT 263.36 42.165 263.57 42.235 ;
    RECT 263.36 42.525 263.57 42.595 ;
    RECT 262.9 41.805 263.11 41.875 ;
    RECT 262.9 42.165 263.11 42.235 ;
    RECT 262.9 42.525 263.11 42.595 ;
    RECT 260.04 41.805 260.25 41.875 ;
    RECT 260.04 42.165 260.25 42.235 ;
    RECT 260.04 42.525 260.25 42.595 ;
    RECT 259.58 41.805 259.79 41.875 ;
    RECT 259.58 42.165 259.79 42.235 ;
    RECT 259.58 42.525 259.79 42.595 ;
    RECT 256.72 41.805 256.93 41.875 ;
    RECT 256.72 42.165 256.93 42.235 ;
    RECT 256.72 42.525 256.93 42.595 ;
    RECT 256.26 41.805 256.47 41.875 ;
    RECT 256.26 42.165 256.47 42.235 ;
    RECT 256.26 42.525 256.47 42.595 ;
    RECT 253.4 41.805 253.61 41.875 ;
    RECT 253.4 42.165 253.61 42.235 ;
    RECT 253.4 42.525 253.61 42.595 ;
    RECT 252.94 41.805 253.15 41.875 ;
    RECT 252.94 42.165 253.15 42.235 ;
    RECT 252.94 42.525 253.15 42.595 ;
    RECT 250.08 41.805 250.29 41.875 ;
    RECT 250.08 42.165 250.29 42.235 ;
    RECT 250.08 42.525 250.29 42.595 ;
    RECT 249.62 41.805 249.83 41.875 ;
    RECT 249.62 42.165 249.83 42.235 ;
    RECT 249.62 42.525 249.83 42.595 ;
    RECT 246.76 41.805 246.97 41.875 ;
    RECT 246.76 42.165 246.97 42.235 ;
    RECT 246.76 42.525 246.97 42.595 ;
    RECT 246.3 41.805 246.51 41.875 ;
    RECT 246.3 42.165 246.51 42.235 ;
    RECT 246.3 42.525 246.51 42.595 ;
    RECT 243.44 41.805 243.65 41.875 ;
    RECT 243.44 42.165 243.65 42.235 ;
    RECT 243.44 42.525 243.65 42.595 ;
    RECT 242.98 41.805 243.19 41.875 ;
    RECT 242.98 42.165 243.19 42.235 ;
    RECT 242.98 42.525 243.19 42.595 ;
    RECT 240.12 41.805 240.33 41.875 ;
    RECT 240.12 42.165 240.33 42.235 ;
    RECT 240.12 42.525 240.33 42.595 ;
    RECT 239.66 41.805 239.87 41.875 ;
    RECT 239.66 42.165 239.87 42.235 ;
    RECT 239.66 42.525 239.87 42.595 ;
    RECT 236.8 41.805 237.01 41.875 ;
    RECT 236.8 42.165 237.01 42.235 ;
    RECT 236.8 42.525 237.01 42.595 ;
    RECT 236.34 41.805 236.55 41.875 ;
    RECT 236.34 42.165 236.55 42.235 ;
    RECT 236.34 42.525 236.55 42.595 ;
    RECT 374.15 42.165 374.22 42.235 ;
    RECT 333.08 41.805 333.29 41.875 ;
    RECT 333.08 42.165 333.29 42.235 ;
    RECT 333.08 42.525 333.29 42.595 ;
    RECT 332.62 41.805 332.83 41.875 ;
    RECT 332.62 42.165 332.83 42.235 ;
    RECT 332.62 42.525 332.83 42.595 ;
    RECT 329.76 41.805 329.97 41.875 ;
    RECT 329.76 42.165 329.97 42.235 ;
    RECT 329.76 42.525 329.97 42.595 ;
    RECT 329.3 41.805 329.51 41.875 ;
    RECT 329.3 42.165 329.51 42.235 ;
    RECT 329.3 42.525 329.51 42.595 ;
    RECT 326.44 41.805 326.65 41.875 ;
    RECT 326.44 42.165 326.65 42.235 ;
    RECT 326.44 42.525 326.65 42.595 ;
    RECT 325.98 41.805 326.19 41.875 ;
    RECT 325.98 42.165 326.19 42.235 ;
    RECT 325.98 42.525 326.19 42.595 ;
    RECT 323.12 41.805 323.33 41.875 ;
    RECT 323.12 42.165 323.33 42.235 ;
    RECT 323.12 42.525 323.33 42.595 ;
    RECT 322.66 41.805 322.87 41.875 ;
    RECT 322.66 42.165 322.87 42.235 ;
    RECT 322.66 42.525 322.87 42.595 ;
    RECT 319.8 41.805 320.01 41.875 ;
    RECT 319.8 42.165 320.01 42.235 ;
    RECT 319.8 42.525 320.01 42.595 ;
    RECT 319.34 41.805 319.55 41.875 ;
    RECT 319.34 42.165 319.55 42.235 ;
    RECT 319.34 42.525 319.55 42.595 ;
    RECT 316.48 41.805 316.69 41.875 ;
    RECT 316.48 42.165 316.69 42.235 ;
    RECT 316.48 42.525 316.69 42.595 ;
    RECT 316.02 41.805 316.23 41.875 ;
    RECT 316.02 42.165 316.23 42.235 ;
    RECT 316.02 42.525 316.23 42.595 ;
    RECT 313.16 41.805 313.37 41.875 ;
    RECT 313.16 42.165 313.37 42.235 ;
    RECT 313.16 42.525 313.37 42.595 ;
    RECT 312.7 41.805 312.91 41.875 ;
    RECT 312.7 42.165 312.91 42.235 ;
    RECT 312.7 42.525 312.91 42.595 ;
    RECT 309.84 41.805 310.05 41.875 ;
    RECT 309.84 42.165 310.05 42.235 ;
    RECT 309.84 42.525 310.05 42.595 ;
    RECT 309.38 41.805 309.59 41.875 ;
    RECT 309.38 42.165 309.59 42.235 ;
    RECT 309.38 42.525 309.59 42.595 ;
    RECT 306.52 41.805 306.73 41.875 ;
    RECT 306.52 42.165 306.73 42.235 ;
    RECT 306.52 42.525 306.73 42.595 ;
    RECT 306.06 41.805 306.27 41.875 ;
    RECT 306.06 42.165 306.27 42.235 ;
    RECT 306.06 42.525 306.27 42.595 ;
    RECT 303.2 41.085 303.41 41.155 ;
    RECT 303.2 41.445 303.41 41.515 ;
    RECT 303.2 41.805 303.41 41.875 ;
    RECT 302.74 41.085 302.95 41.155 ;
    RECT 302.74 41.445 302.95 41.515 ;
    RECT 302.74 41.805 302.95 41.875 ;
    RECT 372.92 41.085 373.13 41.155 ;
    RECT 372.92 41.445 373.13 41.515 ;
    RECT 372.92 41.805 373.13 41.875 ;
    RECT 372.46 41.085 372.67 41.155 ;
    RECT 372.46 41.445 372.67 41.515 ;
    RECT 372.46 41.805 372.67 41.875 ;
    RECT 369.6 41.085 369.81 41.155 ;
    RECT 369.6 41.445 369.81 41.515 ;
    RECT 369.6 41.805 369.81 41.875 ;
    RECT 369.14 41.085 369.35 41.155 ;
    RECT 369.14 41.445 369.35 41.515 ;
    RECT 369.14 41.805 369.35 41.875 ;
    RECT 200.605 41.445 200.675 41.515 ;
    RECT 299.88 41.085 300.09 41.155 ;
    RECT 299.88 41.445 300.09 41.515 ;
    RECT 299.88 41.805 300.09 41.875 ;
    RECT 299.42 41.085 299.63 41.155 ;
    RECT 299.42 41.445 299.63 41.515 ;
    RECT 299.42 41.805 299.63 41.875 ;
    RECT 296.56 41.085 296.77 41.155 ;
    RECT 296.56 41.445 296.77 41.515 ;
    RECT 296.56 41.805 296.77 41.875 ;
    RECT 296.1 41.085 296.31 41.155 ;
    RECT 296.1 41.445 296.31 41.515 ;
    RECT 296.1 41.805 296.31 41.875 ;
    RECT 293.24 41.085 293.45 41.155 ;
    RECT 293.24 41.445 293.45 41.515 ;
    RECT 293.24 41.805 293.45 41.875 ;
    RECT 292.78 41.085 292.99 41.155 ;
    RECT 292.78 41.445 292.99 41.515 ;
    RECT 292.78 41.805 292.99 41.875 ;
    RECT 289.92 41.085 290.13 41.155 ;
    RECT 289.92 41.445 290.13 41.515 ;
    RECT 289.92 41.805 290.13 41.875 ;
    RECT 289.46 41.085 289.67 41.155 ;
    RECT 289.46 41.445 289.67 41.515 ;
    RECT 289.46 41.805 289.67 41.875 ;
    RECT 286.6 41.085 286.81 41.155 ;
    RECT 286.6 41.445 286.81 41.515 ;
    RECT 286.6 41.805 286.81 41.875 ;
    RECT 286.14 41.085 286.35 41.155 ;
    RECT 286.14 41.445 286.35 41.515 ;
    RECT 286.14 41.805 286.35 41.875 ;
    RECT 283.28 41.085 283.49 41.155 ;
    RECT 283.28 41.445 283.49 41.515 ;
    RECT 283.28 41.805 283.49 41.875 ;
    RECT 282.82 41.085 283.03 41.155 ;
    RECT 282.82 41.445 283.03 41.515 ;
    RECT 282.82 41.805 283.03 41.875 ;
    RECT 279.96 41.085 280.17 41.155 ;
    RECT 279.96 41.445 280.17 41.515 ;
    RECT 279.96 41.805 280.17 41.875 ;
    RECT 279.5 41.085 279.71 41.155 ;
    RECT 279.5 41.445 279.71 41.515 ;
    RECT 279.5 41.805 279.71 41.875 ;
    RECT 276.64 41.085 276.85 41.155 ;
    RECT 276.64 41.445 276.85 41.515 ;
    RECT 276.64 41.805 276.85 41.875 ;
    RECT 276.18 41.085 276.39 41.155 ;
    RECT 276.18 41.445 276.39 41.515 ;
    RECT 276.18 41.805 276.39 41.875 ;
    RECT 273.32 41.085 273.53 41.155 ;
    RECT 273.32 41.445 273.53 41.515 ;
    RECT 273.32 41.805 273.53 41.875 ;
    RECT 272.86 41.085 273.07 41.155 ;
    RECT 272.86 41.445 273.07 41.515 ;
    RECT 272.86 41.805 273.07 41.875 ;
    RECT 270.0 41.085 270.21 41.155 ;
    RECT 270.0 41.445 270.21 41.515 ;
    RECT 270.0 41.805 270.21 41.875 ;
    RECT 269.54 41.085 269.75 41.155 ;
    RECT 269.54 41.445 269.75 41.515 ;
    RECT 269.54 41.805 269.75 41.875 ;
    RECT 233.48 41.085 233.69 41.155 ;
    RECT 233.48 41.445 233.69 41.515 ;
    RECT 233.48 41.805 233.69 41.875 ;
    RECT 233.02 41.085 233.23 41.155 ;
    RECT 233.02 41.445 233.23 41.515 ;
    RECT 233.02 41.805 233.23 41.875 ;
    RECT 230.16 41.085 230.37 41.155 ;
    RECT 230.16 41.445 230.37 41.515 ;
    RECT 230.16 41.805 230.37 41.875 ;
    RECT 229.7 41.085 229.91 41.155 ;
    RECT 229.7 41.445 229.91 41.515 ;
    RECT 229.7 41.805 229.91 41.875 ;
    RECT 366.28 41.085 366.49 41.155 ;
    RECT 366.28 41.445 366.49 41.515 ;
    RECT 366.28 41.805 366.49 41.875 ;
    RECT 365.82 41.085 366.03 41.155 ;
    RECT 365.82 41.445 366.03 41.515 ;
    RECT 365.82 41.805 366.03 41.875 ;
    RECT 226.84 41.085 227.05 41.155 ;
    RECT 226.84 41.445 227.05 41.515 ;
    RECT 226.84 41.805 227.05 41.875 ;
    RECT 226.38 41.085 226.59 41.155 ;
    RECT 226.38 41.445 226.59 41.515 ;
    RECT 226.38 41.805 226.59 41.875 ;
    RECT 362.96 41.085 363.17 41.155 ;
    RECT 362.96 41.445 363.17 41.515 ;
    RECT 362.96 41.805 363.17 41.875 ;
    RECT 362.5 41.085 362.71 41.155 ;
    RECT 362.5 41.445 362.71 41.515 ;
    RECT 362.5 41.805 362.71 41.875 ;
    RECT 223.52 41.085 223.73 41.155 ;
    RECT 223.52 41.445 223.73 41.515 ;
    RECT 223.52 41.805 223.73 41.875 ;
    RECT 223.06 41.085 223.27 41.155 ;
    RECT 223.06 41.445 223.27 41.515 ;
    RECT 223.06 41.805 223.27 41.875 ;
    RECT 359.64 41.085 359.85 41.155 ;
    RECT 359.64 41.445 359.85 41.515 ;
    RECT 359.64 41.805 359.85 41.875 ;
    RECT 359.18 41.085 359.39 41.155 ;
    RECT 359.18 41.445 359.39 41.515 ;
    RECT 359.18 41.805 359.39 41.875 ;
    RECT 220.2 41.085 220.41 41.155 ;
    RECT 220.2 41.445 220.41 41.515 ;
    RECT 220.2 41.805 220.41 41.875 ;
    RECT 219.74 41.085 219.95 41.155 ;
    RECT 219.74 41.445 219.95 41.515 ;
    RECT 219.74 41.805 219.95 41.875 ;
    RECT 356.32 41.085 356.53 41.155 ;
    RECT 356.32 41.445 356.53 41.515 ;
    RECT 356.32 41.805 356.53 41.875 ;
    RECT 355.86 41.085 356.07 41.155 ;
    RECT 355.86 41.445 356.07 41.515 ;
    RECT 355.86 41.805 356.07 41.875 ;
    RECT 353.0 41.085 353.21 41.155 ;
    RECT 353.0 41.445 353.21 41.515 ;
    RECT 353.0 41.805 353.21 41.875 ;
    RECT 352.54 41.085 352.75 41.155 ;
    RECT 352.54 41.445 352.75 41.515 ;
    RECT 352.54 41.805 352.75 41.875 ;
    RECT 216.88 41.085 217.09 41.155 ;
    RECT 216.88 41.445 217.09 41.515 ;
    RECT 216.88 41.805 217.09 41.875 ;
    RECT 216.42 41.085 216.63 41.155 ;
    RECT 216.42 41.445 216.63 41.515 ;
    RECT 216.42 41.805 216.63 41.875 ;
    RECT 349.68 41.085 349.89 41.155 ;
    RECT 349.68 41.445 349.89 41.515 ;
    RECT 349.68 41.805 349.89 41.875 ;
    RECT 349.22 41.085 349.43 41.155 ;
    RECT 349.22 41.445 349.43 41.515 ;
    RECT 349.22 41.805 349.43 41.875 ;
    RECT 213.56 41.085 213.77 41.155 ;
    RECT 213.56 41.445 213.77 41.515 ;
    RECT 213.56 41.805 213.77 41.875 ;
    RECT 213.1 41.085 213.31 41.155 ;
    RECT 213.1 41.445 213.31 41.515 ;
    RECT 213.1 41.805 213.31 41.875 ;
    RECT 346.36 41.085 346.57 41.155 ;
    RECT 346.36 41.445 346.57 41.515 ;
    RECT 346.36 41.805 346.57 41.875 ;
    RECT 345.9 41.085 346.11 41.155 ;
    RECT 345.9 41.445 346.11 41.515 ;
    RECT 345.9 41.805 346.11 41.875 ;
    RECT 210.24 41.085 210.45 41.155 ;
    RECT 210.24 41.445 210.45 41.515 ;
    RECT 210.24 41.805 210.45 41.875 ;
    RECT 209.78 41.085 209.99 41.155 ;
    RECT 209.78 41.445 209.99 41.515 ;
    RECT 209.78 41.805 209.99 41.875 ;
    RECT 343.04 41.085 343.25 41.155 ;
    RECT 343.04 41.445 343.25 41.515 ;
    RECT 343.04 41.805 343.25 41.875 ;
    RECT 342.58 41.085 342.79 41.155 ;
    RECT 342.58 41.445 342.79 41.515 ;
    RECT 342.58 41.805 342.79 41.875 ;
    RECT 206.92 41.085 207.13 41.155 ;
    RECT 206.92 41.445 207.13 41.515 ;
    RECT 206.92 41.805 207.13 41.875 ;
    RECT 206.46 41.085 206.67 41.155 ;
    RECT 206.46 41.445 206.67 41.515 ;
    RECT 206.46 41.805 206.67 41.875 ;
    RECT 339.72 41.085 339.93 41.155 ;
    RECT 339.72 41.445 339.93 41.515 ;
    RECT 339.72 41.805 339.93 41.875 ;
    RECT 339.26 41.085 339.47 41.155 ;
    RECT 339.26 41.445 339.47 41.515 ;
    RECT 339.26 41.805 339.47 41.875 ;
    RECT 203.6 41.085 203.81 41.155 ;
    RECT 203.6 41.445 203.81 41.515 ;
    RECT 203.6 41.805 203.81 41.875 ;
    RECT 203.14 41.085 203.35 41.155 ;
    RECT 203.14 41.445 203.35 41.515 ;
    RECT 203.14 41.805 203.35 41.875 ;
    RECT 336.4 41.085 336.61 41.155 ;
    RECT 336.4 41.445 336.61 41.515 ;
    RECT 336.4 41.805 336.61 41.875 ;
    RECT 335.94 41.085 336.15 41.155 ;
    RECT 335.94 41.445 336.15 41.515 ;
    RECT 335.94 41.805 336.15 41.875 ;
    RECT 266.68 41.085 266.89 41.155 ;
    RECT 266.68 41.445 266.89 41.515 ;
    RECT 266.68 41.805 266.89 41.875 ;
    RECT 266.22 41.085 266.43 41.155 ;
    RECT 266.22 41.445 266.43 41.515 ;
    RECT 266.22 41.805 266.43 41.875 ;
    RECT 263.36 41.085 263.57 41.155 ;
    RECT 263.36 41.445 263.57 41.515 ;
    RECT 263.36 41.805 263.57 41.875 ;
    RECT 262.9 41.085 263.11 41.155 ;
    RECT 262.9 41.445 263.11 41.515 ;
    RECT 262.9 41.805 263.11 41.875 ;
    RECT 260.04 41.085 260.25 41.155 ;
    RECT 260.04 41.445 260.25 41.515 ;
    RECT 260.04 41.805 260.25 41.875 ;
    RECT 259.58 41.085 259.79 41.155 ;
    RECT 259.58 41.445 259.79 41.515 ;
    RECT 259.58 41.805 259.79 41.875 ;
    RECT 256.72 41.085 256.93 41.155 ;
    RECT 256.72 41.445 256.93 41.515 ;
    RECT 256.72 41.805 256.93 41.875 ;
    RECT 256.26 41.085 256.47 41.155 ;
    RECT 256.26 41.445 256.47 41.515 ;
    RECT 256.26 41.805 256.47 41.875 ;
    RECT 253.4 41.085 253.61 41.155 ;
    RECT 253.4 41.445 253.61 41.515 ;
    RECT 253.4 41.805 253.61 41.875 ;
    RECT 252.94 41.085 253.15 41.155 ;
    RECT 252.94 41.445 253.15 41.515 ;
    RECT 252.94 41.805 253.15 41.875 ;
    RECT 250.08 41.085 250.29 41.155 ;
    RECT 250.08 41.445 250.29 41.515 ;
    RECT 250.08 41.805 250.29 41.875 ;
    RECT 249.62 41.085 249.83 41.155 ;
    RECT 249.62 41.445 249.83 41.515 ;
    RECT 249.62 41.805 249.83 41.875 ;
    RECT 246.76 41.085 246.97 41.155 ;
    RECT 246.76 41.445 246.97 41.515 ;
    RECT 246.76 41.805 246.97 41.875 ;
    RECT 246.3 41.085 246.51 41.155 ;
    RECT 246.3 41.445 246.51 41.515 ;
    RECT 246.3 41.805 246.51 41.875 ;
    RECT 243.44 41.085 243.65 41.155 ;
    RECT 243.44 41.445 243.65 41.515 ;
    RECT 243.44 41.805 243.65 41.875 ;
    RECT 242.98 41.085 243.19 41.155 ;
    RECT 242.98 41.445 243.19 41.515 ;
    RECT 242.98 41.805 243.19 41.875 ;
    RECT 240.12 41.085 240.33 41.155 ;
    RECT 240.12 41.445 240.33 41.515 ;
    RECT 240.12 41.805 240.33 41.875 ;
    RECT 239.66 41.085 239.87 41.155 ;
    RECT 239.66 41.445 239.87 41.515 ;
    RECT 239.66 41.805 239.87 41.875 ;
    RECT 236.8 41.085 237.01 41.155 ;
    RECT 236.8 41.445 237.01 41.515 ;
    RECT 236.8 41.805 237.01 41.875 ;
    RECT 236.34 41.085 236.55 41.155 ;
    RECT 236.34 41.445 236.55 41.515 ;
    RECT 236.34 41.805 236.55 41.875 ;
    RECT 374.15 41.445 374.22 41.515 ;
    RECT 333.08 41.085 333.29 41.155 ;
    RECT 333.08 41.445 333.29 41.515 ;
    RECT 333.08 41.805 333.29 41.875 ;
    RECT 332.62 41.085 332.83 41.155 ;
    RECT 332.62 41.445 332.83 41.515 ;
    RECT 332.62 41.805 332.83 41.875 ;
    RECT 329.76 41.085 329.97 41.155 ;
    RECT 329.76 41.445 329.97 41.515 ;
    RECT 329.76 41.805 329.97 41.875 ;
    RECT 329.3 41.085 329.51 41.155 ;
    RECT 329.3 41.445 329.51 41.515 ;
    RECT 329.3 41.805 329.51 41.875 ;
    RECT 326.44 41.085 326.65 41.155 ;
    RECT 326.44 41.445 326.65 41.515 ;
    RECT 326.44 41.805 326.65 41.875 ;
    RECT 325.98 41.085 326.19 41.155 ;
    RECT 325.98 41.445 326.19 41.515 ;
    RECT 325.98 41.805 326.19 41.875 ;
    RECT 323.12 41.085 323.33 41.155 ;
    RECT 323.12 41.445 323.33 41.515 ;
    RECT 323.12 41.805 323.33 41.875 ;
    RECT 322.66 41.085 322.87 41.155 ;
    RECT 322.66 41.445 322.87 41.515 ;
    RECT 322.66 41.805 322.87 41.875 ;
    RECT 319.8 41.085 320.01 41.155 ;
    RECT 319.8 41.445 320.01 41.515 ;
    RECT 319.8 41.805 320.01 41.875 ;
    RECT 319.34 41.085 319.55 41.155 ;
    RECT 319.34 41.445 319.55 41.515 ;
    RECT 319.34 41.805 319.55 41.875 ;
    RECT 316.48 41.085 316.69 41.155 ;
    RECT 316.48 41.445 316.69 41.515 ;
    RECT 316.48 41.805 316.69 41.875 ;
    RECT 316.02 41.085 316.23 41.155 ;
    RECT 316.02 41.445 316.23 41.515 ;
    RECT 316.02 41.805 316.23 41.875 ;
    RECT 313.16 41.085 313.37 41.155 ;
    RECT 313.16 41.445 313.37 41.515 ;
    RECT 313.16 41.805 313.37 41.875 ;
    RECT 312.7 41.085 312.91 41.155 ;
    RECT 312.7 41.445 312.91 41.515 ;
    RECT 312.7 41.805 312.91 41.875 ;
    RECT 309.84 41.085 310.05 41.155 ;
    RECT 309.84 41.445 310.05 41.515 ;
    RECT 309.84 41.805 310.05 41.875 ;
    RECT 309.38 41.085 309.59 41.155 ;
    RECT 309.38 41.445 309.59 41.515 ;
    RECT 309.38 41.805 309.59 41.875 ;
    RECT 306.52 41.085 306.73 41.155 ;
    RECT 306.52 41.445 306.73 41.515 ;
    RECT 306.52 41.805 306.73 41.875 ;
    RECT 306.06 41.085 306.27 41.155 ;
    RECT 306.06 41.445 306.27 41.515 ;
    RECT 306.06 41.805 306.27 41.875 ;
    RECT 303.2 40.365 303.41 40.435 ;
    RECT 303.2 40.725 303.41 40.795 ;
    RECT 303.2 41.085 303.41 41.155 ;
    RECT 302.74 40.365 302.95 40.435 ;
    RECT 302.74 40.725 302.95 40.795 ;
    RECT 302.74 41.085 302.95 41.155 ;
    RECT 372.92 40.365 373.13 40.435 ;
    RECT 372.92 40.725 373.13 40.795 ;
    RECT 372.92 41.085 373.13 41.155 ;
    RECT 372.46 40.365 372.67 40.435 ;
    RECT 372.46 40.725 372.67 40.795 ;
    RECT 372.46 41.085 372.67 41.155 ;
    RECT 369.6 40.365 369.81 40.435 ;
    RECT 369.6 40.725 369.81 40.795 ;
    RECT 369.6 41.085 369.81 41.155 ;
    RECT 369.14 40.365 369.35 40.435 ;
    RECT 369.14 40.725 369.35 40.795 ;
    RECT 369.14 41.085 369.35 41.155 ;
    RECT 200.605 40.725 200.675 40.795 ;
    RECT 299.88 40.365 300.09 40.435 ;
    RECT 299.88 40.725 300.09 40.795 ;
    RECT 299.88 41.085 300.09 41.155 ;
    RECT 299.42 40.365 299.63 40.435 ;
    RECT 299.42 40.725 299.63 40.795 ;
    RECT 299.42 41.085 299.63 41.155 ;
    RECT 296.56 40.365 296.77 40.435 ;
    RECT 296.56 40.725 296.77 40.795 ;
    RECT 296.56 41.085 296.77 41.155 ;
    RECT 296.1 40.365 296.31 40.435 ;
    RECT 296.1 40.725 296.31 40.795 ;
    RECT 296.1 41.085 296.31 41.155 ;
    RECT 293.24 40.365 293.45 40.435 ;
    RECT 293.24 40.725 293.45 40.795 ;
    RECT 293.24 41.085 293.45 41.155 ;
    RECT 292.78 40.365 292.99 40.435 ;
    RECT 292.78 40.725 292.99 40.795 ;
    RECT 292.78 41.085 292.99 41.155 ;
    RECT 289.92 40.365 290.13 40.435 ;
    RECT 289.92 40.725 290.13 40.795 ;
    RECT 289.92 41.085 290.13 41.155 ;
    RECT 289.46 40.365 289.67 40.435 ;
    RECT 289.46 40.725 289.67 40.795 ;
    RECT 289.46 41.085 289.67 41.155 ;
    RECT 286.6 40.365 286.81 40.435 ;
    RECT 286.6 40.725 286.81 40.795 ;
    RECT 286.6 41.085 286.81 41.155 ;
    RECT 286.14 40.365 286.35 40.435 ;
    RECT 286.14 40.725 286.35 40.795 ;
    RECT 286.14 41.085 286.35 41.155 ;
    RECT 283.28 40.365 283.49 40.435 ;
    RECT 283.28 40.725 283.49 40.795 ;
    RECT 283.28 41.085 283.49 41.155 ;
    RECT 282.82 40.365 283.03 40.435 ;
    RECT 282.82 40.725 283.03 40.795 ;
    RECT 282.82 41.085 283.03 41.155 ;
    RECT 279.96 40.365 280.17 40.435 ;
    RECT 279.96 40.725 280.17 40.795 ;
    RECT 279.96 41.085 280.17 41.155 ;
    RECT 279.5 40.365 279.71 40.435 ;
    RECT 279.5 40.725 279.71 40.795 ;
    RECT 279.5 41.085 279.71 41.155 ;
    RECT 276.64 40.365 276.85 40.435 ;
    RECT 276.64 40.725 276.85 40.795 ;
    RECT 276.64 41.085 276.85 41.155 ;
    RECT 276.18 40.365 276.39 40.435 ;
    RECT 276.18 40.725 276.39 40.795 ;
    RECT 276.18 41.085 276.39 41.155 ;
    RECT 273.32 40.365 273.53 40.435 ;
    RECT 273.32 40.725 273.53 40.795 ;
    RECT 273.32 41.085 273.53 41.155 ;
    RECT 272.86 40.365 273.07 40.435 ;
    RECT 272.86 40.725 273.07 40.795 ;
    RECT 272.86 41.085 273.07 41.155 ;
    RECT 270.0 40.365 270.21 40.435 ;
    RECT 270.0 40.725 270.21 40.795 ;
    RECT 270.0 41.085 270.21 41.155 ;
    RECT 269.54 40.365 269.75 40.435 ;
    RECT 269.54 40.725 269.75 40.795 ;
    RECT 269.54 41.085 269.75 41.155 ;
    RECT 233.48 40.365 233.69 40.435 ;
    RECT 233.48 40.725 233.69 40.795 ;
    RECT 233.48 41.085 233.69 41.155 ;
    RECT 233.02 40.365 233.23 40.435 ;
    RECT 233.02 40.725 233.23 40.795 ;
    RECT 233.02 41.085 233.23 41.155 ;
    RECT 230.16 40.365 230.37 40.435 ;
    RECT 230.16 40.725 230.37 40.795 ;
    RECT 230.16 41.085 230.37 41.155 ;
    RECT 229.7 40.365 229.91 40.435 ;
    RECT 229.7 40.725 229.91 40.795 ;
    RECT 229.7 41.085 229.91 41.155 ;
    RECT 366.28 40.365 366.49 40.435 ;
    RECT 366.28 40.725 366.49 40.795 ;
    RECT 366.28 41.085 366.49 41.155 ;
    RECT 365.82 40.365 366.03 40.435 ;
    RECT 365.82 40.725 366.03 40.795 ;
    RECT 365.82 41.085 366.03 41.155 ;
    RECT 226.84 40.365 227.05 40.435 ;
    RECT 226.84 40.725 227.05 40.795 ;
    RECT 226.84 41.085 227.05 41.155 ;
    RECT 226.38 40.365 226.59 40.435 ;
    RECT 226.38 40.725 226.59 40.795 ;
    RECT 226.38 41.085 226.59 41.155 ;
    RECT 362.96 40.365 363.17 40.435 ;
    RECT 362.96 40.725 363.17 40.795 ;
    RECT 362.96 41.085 363.17 41.155 ;
    RECT 362.5 40.365 362.71 40.435 ;
    RECT 362.5 40.725 362.71 40.795 ;
    RECT 362.5 41.085 362.71 41.155 ;
    RECT 223.52 40.365 223.73 40.435 ;
    RECT 223.52 40.725 223.73 40.795 ;
    RECT 223.52 41.085 223.73 41.155 ;
    RECT 223.06 40.365 223.27 40.435 ;
    RECT 223.06 40.725 223.27 40.795 ;
    RECT 223.06 41.085 223.27 41.155 ;
    RECT 359.64 40.365 359.85 40.435 ;
    RECT 359.64 40.725 359.85 40.795 ;
    RECT 359.64 41.085 359.85 41.155 ;
    RECT 359.18 40.365 359.39 40.435 ;
    RECT 359.18 40.725 359.39 40.795 ;
    RECT 359.18 41.085 359.39 41.155 ;
    RECT 220.2 40.365 220.41 40.435 ;
    RECT 220.2 40.725 220.41 40.795 ;
    RECT 220.2 41.085 220.41 41.155 ;
    RECT 219.74 40.365 219.95 40.435 ;
    RECT 219.74 40.725 219.95 40.795 ;
    RECT 219.74 41.085 219.95 41.155 ;
    RECT 356.32 40.365 356.53 40.435 ;
    RECT 356.32 40.725 356.53 40.795 ;
    RECT 356.32 41.085 356.53 41.155 ;
    RECT 355.86 40.365 356.07 40.435 ;
    RECT 355.86 40.725 356.07 40.795 ;
    RECT 355.86 41.085 356.07 41.155 ;
    RECT 353.0 40.365 353.21 40.435 ;
    RECT 353.0 40.725 353.21 40.795 ;
    RECT 353.0 41.085 353.21 41.155 ;
    RECT 352.54 40.365 352.75 40.435 ;
    RECT 352.54 40.725 352.75 40.795 ;
    RECT 352.54 41.085 352.75 41.155 ;
    RECT 216.88 40.365 217.09 40.435 ;
    RECT 216.88 40.725 217.09 40.795 ;
    RECT 216.88 41.085 217.09 41.155 ;
    RECT 216.42 40.365 216.63 40.435 ;
    RECT 216.42 40.725 216.63 40.795 ;
    RECT 216.42 41.085 216.63 41.155 ;
    RECT 349.68 40.365 349.89 40.435 ;
    RECT 349.68 40.725 349.89 40.795 ;
    RECT 349.68 41.085 349.89 41.155 ;
    RECT 349.22 40.365 349.43 40.435 ;
    RECT 349.22 40.725 349.43 40.795 ;
    RECT 349.22 41.085 349.43 41.155 ;
    RECT 213.56 40.365 213.77 40.435 ;
    RECT 213.56 40.725 213.77 40.795 ;
    RECT 213.56 41.085 213.77 41.155 ;
    RECT 213.1 40.365 213.31 40.435 ;
    RECT 213.1 40.725 213.31 40.795 ;
    RECT 213.1 41.085 213.31 41.155 ;
    RECT 346.36 40.365 346.57 40.435 ;
    RECT 346.36 40.725 346.57 40.795 ;
    RECT 346.36 41.085 346.57 41.155 ;
    RECT 345.9 40.365 346.11 40.435 ;
    RECT 345.9 40.725 346.11 40.795 ;
    RECT 345.9 41.085 346.11 41.155 ;
    RECT 210.24 40.365 210.45 40.435 ;
    RECT 210.24 40.725 210.45 40.795 ;
    RECT 210.24 41.085 210.45 41.155 ;
    RECT 209.78 40.365 209.99 40.435 ;
    RECT 209.78 40.725 209.99 40.795 ;
    RECT 209.78 41.085 209.99 41.155 ;
    RECT 343.04 40.365 343.25 40.435 ;
    RECT 343.04 40.725 343.25 40.795 ;
    RECT 343.04 41.085 343.25 41.155 ;
    RECT 342.58 40.365 342.79 40.435 ;
    RECT 342.58 40.725 342.79 40.795 ;
    RECT 342.58 41.085 342.79 41.155 ;
    RECT 206.92 40.365 207.13 40.435 ;
    RECT 206.92 40.725 207.13 40.795 ;
    RECT 206.92 41.085 207.13 41.155 ;
    RECT 206.46 40.365 206.67 40.435 ;
    RECT 206.46 40.725 206.67 40.795 ;
    RECT 206.46 41.085 206.67 41.155 ;
    RECT 339.72 40.365 339.93 40.435 ;
    RECT 339.72 40.725 339.93 40.795 ;
    RECT 339.72 41.085 339.93 41.155 ;
    RECT 339.26 40.365 339.47 40.435 ;
    RECT 339.26 40.725 339.47 40.795 ;
    RECT 339.26 41.085 339.47 41.155 ;
    RECT 203.6 40.365 203.81 40.435 ;
    RECT 203.6 40.725 203.81 40.795 ;
    RECT 203.6 41.085 203.81 41.155 ;
    RECT 203.14 40.365 203.35 40.435 ;
    RECT 203.14 40.725 203.35 40.795 ;
    RECT 203.14 41.085 203.35 41.155 ;
    RECT 336.4 40.365 336.61 40.435 ;
    RECT 336.4 40.725 336.61 40.795 ;
    RECT 336.4 41.085 336.61 41.155 ;
    RECT 335.94 40.365 336.15 40.435 ;
    RECT 335.94 40.725 336.15 40.795 ;
    RECT 335.94 41.085 336.15 41.155 ;
    RECT 266.68 40.365 266.89 40.435 ;
    RECT 266.68 40.725 266.89 40.795 ;
    RECT 266.68 41.085 266.89 41.155 ;
    RECT 266.22 40.365 266.43 40.435 ;
    RECT 266.22 40.725 266.43 40.795 ;
    RECT 266.22 41.085 266.43 41.155 ;
    RECT 263.36 40.365 263.57 40.435 ;
    RECT 263.36 40.725 263.57 40.795 ;
    RECT 263.36 41.085 263.57 41.155 ;
    RECT 262.9 40.365 263.11 40.435 ;
    RECT 262.9 40.725 263.11 40.795 ;
    RECT 262.9 41.085 263.11 41.155 ;
    RECT 260.04 40.365 260.25 40.435 ;
    RECT 260.04 40.725 260.25 40.795 ;
    RECT 260.04 41.085 260.25 41.155 ;
    RECT 259.58 40.365 259.79 40.435 ;
    RECT 259.58 40.725 259.79 40.795 ;
    RECT 259.58 41.085 259.79 41.155 ;
    RECT 256.72 40.365 256.93 40.435 ;
    RECT 256.72 40.725 256.93 40.795 ;
    RECT 256.72 41.085 256.93 41.155 ;
    RECT 256.26 40.365 256.47 40.435 ;
    RECT 256.26 40.725 256.47 40.795 ;
    RECT 256.26 41.085 256.47 41.155 ;
    RECT 253.4 40.365 253.61 40.435 ;
    RECT 253.4 40.725 253.61 40.795 ;
    RECT 253.4 41.085 253.61 41.155 ;
    RECT 252.94 40.365 253.15 40.435 ;
    RECT 252.94 40.725 253.15 40.795 ;
    RECT 252.94 41.085 253.15 41.155 ;
    RECT 250.08 40.365 250.29 40.435 ;
    RECT 250.08 40.725 250.29 40.795 ;
    RECT 250.08 41.085 250.29 41.155 ;
    RECT 249.62 40.365 249.83 40.435 ;
    RECT 249.62 40.725 249.83 40.795 ;
    RECT 249.62 41.085 249.83 41.155 ;
    RECT 246.76 40.365 246.97 40.435 ;
    RECT 246.76 40.725 246.97 40.795 ;
    RECT 246.76 41.085 246.97 41.155 ;
    RECT 246.3 40.365 246.51 40.435 ;
    RECT 246.3 40.725 246.51 40.795 ;
    RECT 246.3 41.085 246.51 41.155 ;
    RECT 243.44 40.365 243.65 40.435 ;
    RECT 243.44 40.725 243.65 40.795 ;
    RECT 243.44 41.085 243.65 41.155 ;
    RECT 242.98 40.365 243.19 40.435 ;
    RECT 242.98 40.725 243.19 40.795 ;
    RECT 242.98 41.085 243.19 41.155 ;
    RECT 240.12 40.365 240.33 40.435 ;
    RECT 240.12 40.725 240.33 40.795 ;
    RECT 240.12 41.085 240.33 41.155 ;
    RECT 239.66 40.365 239.87 40.435 ;
    RECT 239.66 40.725 239.87 40.795 ;
    RECT 239.66 41.085 239.87 41.155 ;
    RECT 236.8 40.365 237.01 40.435 ;
    RECT 236.8 40.725 237.01 40.795 ;
    RECT 236.8 41.085 237.01 41.155 ;
    RECT 236.34 40.365 236.55 40.435 ;
    RECT 236.34 40.725 236.55 40.795 ;
    RECT 236.34 41.085 236.55 41.155 ;
    RECT 374.15 40.725 374.22 40.795 ;
    RECT 333.08 40.365 333.29 40.435 ;
    RECT 333.08 40.725 333.29 40.795 ;
    RECT 333.08 41.085 333.29 41.155 ;
    RECT 332.62 40.365 332.83 40.435 ;
    RECT 332.62 40.725 332.83 40.795 ;
    RECT 332.62 41.085 332.83 41.155 ;
    RECT 329.76 40.365 329.97 40.435 ;
    RECT 329.76 40.725 329.97 40.795 ;
    RECT 329.76 41.085 329.97 41.155 ;
    RECT 329.3 40.365 329.51 40.435 ;
    RECT 329.3 40.725 329.51 40.795 ;
    RECT 329.3 41.085 329.51 41.155 ;
    RECT 326.44 40.365 326.65 40.435 ;
    RECT 326.44 40.725 326.65 40.795 ;
    RECT 326.44 41.085 326.65 41.155 ;
    RECT 325.98 40.365 326.19 40.435 ;
    RECT 325.98 40.725 326.19 40.795 ;
    RECT 325.98 41.085 326.19 41.155 ;
    RECT 323.12 40.365 323.33 40.435 ;
    RECT 323.12 40.725 323.33 40.795 ;
    RECT 323.12 41.085 323.33 41.155 ;
    RECT 322.66 40.365 322.87 40.435 ;
    RECT 322.66 40.725 322.87 40.795 ;
    RECT 322.66 41.085 322.87 41.155 ;
    RECT 319.8 40.365 320.01 40.435 ;
    RECT 319.8 40.725 320.01 40.795 ;
    RECT 319.8 41.085 320.01 41.155 ;
    RECT 319.34 40.365 319.55 40.435 ;
    RECT 319.34 40.725 319.55 40.795 ;
    RECT 319.34 41.085 319.55 41.155 ;
    RECT 316.48 40.365 316.69 40.435 ;
    RECT 316.48 40.725 316.69 40.795 ;
    RECT 316.48 41.085 316.69 41.155 ;
    RECT 316.02 40.365 316.23 40.435 ;
    RECT 316.02 40.725 316.23 40.795 ;
    RECT 316.02 41.085 316.23 41.155 ;
    RECT 313.16 40.365 313.37 40.435 ;
    RECT 313.16 40.725 313.37 40.795 ;
    RECT 313.16 41.085 313.37 41.155 ;
    RECT 312.7 40.365 312.91 40.435 ;
    RECT 312.7 40.725 312.91 40.795 ;
    RECT 312.7 41.085 312.91 41.155 ;
    RECT 309.84 40.365 310.05 40.435 ;
    RECT 309.84 40.725 310.05 40.795 ;
    RECT 309.84 41.085 310.05 41.155 ;
    RECT 309.38 40.365 309.59 40.435 ;
    RECT 309.38 40.725 309.59 40.795 ;
    RECT 309.38 41.085 309.59 41.155 ;
    RECT 306.52 40.365 306.73 40.435 ;
    RECT 306.52 40.725 306.73 40.795 ;
    RECT 306.52 41.085 306.73 41.155 ;
    RECT 306.06 40.365 306.27 40.435 ;
    RECT 306.06 40.725 306.27 40.795 ;
    RECT 306.06 41.085 306.27 41.155 ;
    RECT 303.2 58.385 303.41 58.455 ;
    RECT 303.2 58.745 303.41 58.815 ;
    RECT 303.2 59.105 303.41 59.175 ;
    RECT 302.74 58.385 302.95 58.455 ;
    RECT 302.74 58.745 302.95 58.815 ;
    RECT 302.74 59.105 302.95 59.175 ;
    RECT 369.6 58.385 369.81 58.455 ;
    RECT 369.6 58.745 369.81 58.815 ;
    RECT 369.6 59.105 369.81 59.175 ;
    RECT 369.14 58.385 369.35 58.455 ;
    RECT 369.14 58.745 369.35 58.815 ;
    RECT 369.14 59.105 369.35 59.175 ;
    RECT 299.88 58.385 300.09 58.455 ;
    RECT 299.88 58.745 300.09 58.815 ;
    RECT 299.88 59.105 300.09 59.175 ;
    RECT 299.42 58.385 299.63 58.455 ;
    RECT 299.42 58.745 299.63 58.815 ;
    RECT 299.42 59.105 299.63 59.175 ;
    RECT 296.56 58.385 296.77 58.455 ;
    RECT 296.56 58.745 296.77 58.815 ;
    RECT 296.56 59.105 296.77 59.175 ;
    RECT 296.1 58.385 296.31 58.455 ;
    RECT 296.1 58.745 296.31 58.815 ;
    RECT 296.1 59.105 296.31 59.175 ;
    RECT 293.24 58.385 293.45 58.455 ;
    RECT 293.24 58.745 293.45 58.815 ;
    RECT 293.24 59.105 293.45 59.175 ;
    RECT 292.78 58.385 292.99 58.455 ;
    RECT 292.78 58.745 292.99 58.815 ;
    RECT 292.78 59.105 292.99 59.175 ;
    RECT 200.605 58.745 200.675 58.815 ;
    RECT 289.92 58.385 290.13 58.455 ;
    RECT 289.92 58.745 290.13 58.815 ;
    RECT 289.92 59.105 290.13 59.175 ;
    RECT 289.46 58.385 289.67 58.455 ;
    RECT 289.46 58.745 289.67 58.815 ;
    RECT 289.46 59.105 289.67 59.175 ;
    RECT 286.6 58.385 286.81 58.455 ;
    RECT 286.6 58.745 286.81 58.815 ;
    RECT 286.6 59.105 286.81 59.175 ;
    RECT 286.14 58.385 286.35 58.455 ;
    RECT 286.14 58.745 286.35 58.815 ;
    RECT 286.14 59.105 286.35 59.175 ;
    RECT 283.28 58.385 283.49 58.455 ;
    RECT 283.28 58.745 283.49 58.815 ;
    RECT 283.28 59.105 283.49 59.175 ;
    RECT 282.82 58.385 283.03 58.455 ;
    RECT 282.82 58.745 283.03 58.815 ;
    RECT 282.82 59.105 283.03 59.175 ;
    RECT 279.96 58.385 280.17 58.455 ;
    RECT 279.96 58.745 280.17 58.815 ;
    RECT 279.96 59.105 280.17 59.175 ;
    RECT 279.5 58.385 279.71 58.455 ;
    RECT 279.5 58.745 279.71 58.815 ;
    RECT 279.5 59.105 279.71 59.175 ;
    RECT 276.64 58.385 276.85 58.455 ;
    RECT 276.64 58.745 276.85 58.815 ;
    RECT 276.64 59.105 276.85 59.175 ;
    RECT 276.18 58.385 276.39 58.455 ;
    RECT 276.18 58.745 276.39 58.815 ;
    RECT 276.18 59.105 276.39 59.175 ;
    RECT 273.32 58.385 273.53 58.455 ;
    RECT 273.32 58.745 273.53 58.815 ;
    RECT 273.32 59.105 273.53 59.175 ;
    RECT 272.86 58.385 273.07 58.455 ;
    RECT 272.86 58.745 273.07 58.815 ;
    RECT 272.86 59.105 273.07 59.175 ;
    RECT 270.0 58.385 270.21 58.455 ;
    RECT 270.0 58.745 270.21 58.815 ;
    RECT 270.0 59.105 270.21 59.175 ;
    RECT 269.54 58.385 269.75 58.455 ;
    RECT 269.54 58.745 269.75 58.815 ;
    RECT 269.54 59.105 269.75 59.175 ;
    RECT 233.48 58.385 233.69 58.455 ;
    RECT 233.48 58.745 233.69 58.815 ;
    RECT 233.48 59.105 233.69 59.175 ;
    RECT 233.02 58.385 233.23 58.455 ;
    RECT 233.02 58.745 233.23 58.815 ;
    RECT 233.02 59.105 233.23 59.175 ;
    RECT 230.16 58.385 230.37 58.455 ;
    RECT 230.16 58.745 230.37 58.815 ;
    RECT 230.16 59.105 230.37 59.175 ;
    RECT 229.7 58.385 229.91 58.455 ;
    RECT 229.7 58.745 229.91 58.815 ;
    RECT 229.7 59.105 229.91 59.175 ;
    RECT 366.28 58.385 366.49 58.455 ;
    RECT 366.28 58.745 366.49 58.815 ;
    RECT 366.28 59.105 366.49 59.175 ;
    RECT 365.82 58.385 366.03 58.455 ;
    RECT 365.82 58.745 366.03 58.815 ;
    RECT 365.82 59.105 366.03 59.175 ;
    RECT 226.84 58.385 227.05 58.455 ;
    RECT 226.84 58.745 227.05 58.815 ;
    RECT 226.84 59.105 227.05 59.175 ;
    RECT 226.38 58.385 226.59 58.455 ;
    RECT 226.38 58.745 226.59 58.815 ;
    RECT 226.38 59.105 226.59 59.175 ;
    RECT 362.96 58.385 363.17 58.455 ;
    RECT 362.96 58.745 363.17 58.815 ;
    RECT 362.96 59.105 363.17 59.175 ;
    RECT 362.5 58.385 362.71 58.455 ;
    RECT 362.5 58.745 362.71 58.815 ;
    RECT 362.5 59.105 362.71 59.175 ;
    RECT 223.52 58.385 223.73 58.455 ;
    RECT 223.52 58.745 223.73 58.815 ;
    RECT 223.52 59.105 223.73 59.175 ;
    RECT 223.06 58.385 223.27 58.455 ;
    RECT 223.06 58.745 223.27 58.815 ;
    RECT 223.06 59.105 223.27 59.175 ;
    RECT 359.64 58.385 359.85 58.455 ;
    RECT 359.64 58.745 359.85 58.815 ;
    RECT 359.64 59.105 359.85 59.175 ;
    RECT 359.18 58.385 359.39 58.455 ;
    RECT 359.18 58.745 359.39 58.815 ;
    RECT 359.18 59.105 359.39 59.175 ;
    RECT 220.2 58.385 220.41 58.455 ;
    RECT 220.2 58.745 220.41 58.815 ;
    RECT 220.2 59.105 220.41 59.175 ;
    RECT 219.74 58.385 219.95 58.455 ;
    RECT 219.74 58.745 219.95 58.815 ;
    RECT 219.74 59.105 219.95 59.175 ;
    RECT 356.32 58.385 356.53 58.455 ;
    RECT 356.32 58.745 356.53 58.815 ;
    RECT 356.32 59.105 356.53 59.175 ;
    RECT 355.86 58.385 356.07 58.455 ;
    RECT 355.86 58.745 356.07 58.815 ;
    RECT 355.86 59.105 356.07 59.175 ;
    RECT 353.0 58.385 353.21 58.455 ;
    RECT 353.0 58.745 353.21 58.815 ;
    RECT 353.0 59.105 353.21 59.175 ;
    RECT 352.54 58.385 352.75 58.455 ;
    RECT 352.54 58.745 352.75 58.815 ;
    RECT 352.54 59.105 352.75 59.175 ;
    RECT 216.88 58.385 217.09 58.455 ;
    RECT 216.88 58.745 217.09 58.815 ;
    RECT 216.88 59.105 217.09 59.175 ;
    RECT 216.42 58.385 216.63 58.455 ;
    RECT 216.42 58.745 216.63 58.815 ;
    RECT 216.42 59.105 216.63 59.175 ;
    RECT 349.68 58.385 349.89 58.455 ;
    RECT 349.68 58.745 349.89 58.815 ;
    RECT 349.68 59.105 349.89 59.175 ;
    RECT 349.22 58.385 349.43 58.455 ;
    RECT 349.22 58.745 349.43 58.815 ;
    RECT 349.22 59.105 349.43 59.175 ;
    RECT 213.56 58.385 213.77 58.455 ;
    RECT 213.56 58.745 213.77 58.815 ;
    RECT 213.56 59.105 213.77 59.175 ;
    RECT 213.1 58.385 213.31 58.455 ;
    RECT 213.1 58.745 213.31 58.815 ;
    RECT 213.1 59.105 213.31 59.175 ;
    RECT 346.36 58.385 346.57 58.455 ;
    RECT 346.36 58.745 346.57 58.815 ;
    RECT 346.36 59.105 346.57 59.175 ;
    RECT 345.9 58.385 346.11 58.455 ;
    RECT 345.9 58.745 346.11 58.815 ;
    RECT 345.9 59.105 346.11 59.175 ;
    RECT 210.24 58.385 210.45 58.455 ;
    RECT 210.24 58.745 210.45 58.815 ;
    RECT 210.24 59.105 210.45 59.175 ;
    RECT 209.78 58.385 209.99 58.455 ;
    RECT 209.78 58.745 209.99 58.815 ;
    RECT 209.78 59.105 209.99 59.175 ;
    RECT 343.04 58.385 343.25 58.455 ;
    RECT 343.04 58.745 343.25 58.815 ;
    RECT 343.04 59.105 343.25 59.175 ;
    RECT 342.58 58.385 342.79 58.455 ;
    RECT 342.58 58.745 342.79 58.815 ;
    RECT 342.58 59.105 342.79 59.175 ;
    RECT 206.92 58.385 207.13 58.455 ;
    RECT 206.92 58.745 207.13 58.815 ;
    RECT 206.92 59.105 207.13 59.175 ;
    RECT 206.46 58.385 206.67 58.455 ;
    RECT 206.46 58.745 206.67 58.815 ;
    RECT 206.46 59.105 206.67 59.175 ;
    RECT 339.72 58.385 339.93 58.455 ;
    RECT 339.72 58.745 339.93 58.815 ;
    RECT 339.72 59.105 339.93 59.175 ;
    RECT 339.26 58.385 339.47 58.455 ;
    RECT 339.26 58.745 339.47 58.815 ;
    RECT 339.26 59.105 339.47 59.175 ;
    RECT 336.4 58.385 336.61 58.455 ;
    RECT 336.4 58.745 336.61 58.815 ;
    RECT 336.4 59.105 336.61 59.175 ;
    RECT 335.94 58.385 336.15 58.455 ;
    RECT 335.94 58.745 336.15 58.815 ;
    RECT 335.94 59.105 336.15 59.175 ;
    RECT 266.68 58.385 266.89 58.455 ;
    RECT 266.68 58.745 266.89 58.815 ;
    RECT 266.68 59.105 266.89 59.175 ;
    RECT 266.22 58.385 266.43 58.455 ;
    RECT 266.22 58.745 266.43 58.815 ;
    RECT 266.22 59.105 266.43 59.175 ;
    RECT 263.36 58.385 263.57 58.455 ;
    RECT 263.36 58.745 263.57 58.815 ;
    RECT 263.36 59.105 263.57 59.175 ;
    RECT 262.9 58.385 263.11 58.455 ;
    RECT 262.9 58.745 263.11 58.815 ;
    RECT 262.9 59.105 263.11 59.175 ;
    RECT 260.04 58.385 260.25 58.455 ;
    RECT 260.04 58.745 260.25 58.815 ;
    RECT 260.04 59.105 260.25 59.175 ;
    RECT 259.58 58.385 259.79 58.455 ;
    RECT 259.58 58.745 259.79 58.815 ;
    RECT 259.58 59.105 259.79 59.175 ;
    RECT 256.72 58.385 256.93 58.455 ;
    RECT 256.72 58.745 256.93 58.815 ;
    RECT 256.72 59.105 256.93 59.175 ;
    RECT 256.26 58.385 256.47 58.455 ;
    RECT 256.26 58.745 256.47 58.815 ;
    RECT 256.26 59.105 256.47 59.175 ;
    RECT 253.4 58.385 253.61 58.455 ;
    RECT 253.4 58.745 253.61 58.815 ;
    RECT 253.4 59.105 253.61 59.175 ;
    RECT 252.94 58.385 253.15 58.455 ;
    RECT 252.94 58.745 253.15 58.815 ;
    RECT 252.94 59.105 253.15 59.175 ;
    RECT 250.08 58.385 250.29 58.455 ;
    RECT 250.08 58.745 250.29 58.815 ;
    RECT 250.08 59.105 250.29 59.175 ;
    RECT 249.62 58.385 249.83 58.455 ;
    RECT 249.62 58.745 249.83 58.815 ;
    RECT 249.62 59.105 249.83 59.175 ;
    RECT 246.76 58.385 246.97 58.455 ;
    RECT 246.76 58.745 246.97 58.815 ;
    RECT 246.76 59.105 246.97 59.175 ;
    RECT 246.3 58.385 246.51 58.455 ;
    RECT 246.3 58.745 246.51 58.815 ;
    RECT 246.3 59.105 246.51 59.175 ;
    RECT 243.44 58.385 243.65 58.455 ;
    RECT 243.44 58.745 243.65 58.815 ;
    RECT 243.44 59.105 243.65 59.175 ;
    RECT 242.98 58.385 243.19 58.455 ;
    RECT 242.98 58.745 243.19 58.815 ;
    RECT 242.98 59.105 243.19 59.175 ;
    RECT 240.12 58.385 240.33 58.455 ;
    RECT 240.12 58.745 240.33 58.815 ;
    RECT 240.12 59.105 240.33 59.175 ;
    RECT 239.66 58.385 239.87 58.455 ;
    RECT 239.66 58.745 239.87 58.815 ;
    RECT 239.66 59.105 239.87 59.175 ;
    RECT 236.8 58.385 237.01 58.455 ;
    RECT 236.8 58.745 237.01 58.815 ;
    RECT 236.8 59.105 237.01 59.175 ;
    RECT 236.34 58.385 236.55 58.455 ;
    RECT 236.34 58.745 236.55 58.815 ;
    RECT 236.34 59.105 236.55 59.175 ;
    RECT 372.92 58.385 373.13 58.455 ;
    RECT 372.92 58.745 373.13 58.815 ;
    RECT 372.92 59.105 373.13 59.175 ;
    RECT 372.46 58.385 372.67 58.455 ;
    RECT 372.46 58.745 372.67 58.815 ;
    RECT 372.46 59.105 372.67 59.175 ;
    RECT 333.08 58.385 333.29 58.455 ;
    RECT 333.08 58.745 333.29 58.815 ;
    RECT 333.08 59.105 333.29 59.175 ;
    RECT 332.62 58.385 332.83 58.455 ;
    RECT 332.62 58.745 332.83 58.815 ;
    RECT 332.62 59.105 332.83 59.175 ;
    RECT 329.76 58.385 329.97 58.455 ;
    RECT 329.76 58.745 329.97 58.815 ;
    RECT 329.76 59.105 329.97 59.175 ;
    RECT 329.3 58.385 329.51 58.455 ;
    RECT 329.3 58.745 329.51 58.815 ;
    RECT 329.3 59.105 329.51 59.175 ;
    RECT 326.44 58.385 326.65 58.455 ;
    RECT 326.44 58.745 326.65 58.815 ;
    RECT 326.44 59.105 326.65 59.175 ;
    RECT 325.98 58.385 326.19 58.455 ;
    RECT 325.98 58.745 326.19 58.815 ;
    RECT 325.98 59.105 326.19 59.175 ;
    RECT 203.6 58.385 203.81 58.455 ;
    RECT 203.6 58.745 203.81 58.815 ;
    RECT 203.6 59.105 203.81 59.175 ;
    RECT 203.14 58.385 203.35 58.455 ;
    RECT 203.14 58.745 203.35 58.815 ;
    RECT 203.14 59.105 203.35 59.175 ;
    RECT 323.12 58.385 323.33 58.455 ;
    RECT 323.12 58.745 323.33 58.815 ;
    RECT 323.12 59.105 323.33 59.175 ;
    RECT 322.66 58.385 322.87 58.455 ;
    RECT 322.66 58.745 322.87 58.815 ;
    RECT 322.66 59.105 322.87 59.175 ;
    RECT 319.8 58.385 320.01 58.455 ;
    RECT 319.8 58.745 320.01 58.815 ;
    RECT 319.8 59.105 320.01 59.175 ;
    RECT 319.34 58.385 319.55 58.455 ;
    RECT 319.34 58.745 319.55 58.815 ;
    RECT 319.34 59.105 319.55 59.175 ;
    RECT 316.48 58.385 316.69 58.455 ;
    RECT 316.48 58.745 316.69 58.815 ;
    RECT 316.48 59.105 316.69 59.175 ;
    RECT 316.02 58.385 316.23 58.455 ;
    RECT 316.02 58.745 316.23 58.815 ;
    RECT 316.02 59.105 316.23 59.175 ;
    RECT 313.16 58.385 313.37 58.455 ;
    RECT 313.16 58.745 313.37 58.815 ;
    RECT 313.16 59.105 313.37 59.175 ;
    RECT 312.7 58.385 312.91 58.455 ;
    RECT 312.7 58.745 312.91 58.815 ;
    RECT 312.7 59.105 312.91 59.175 ;
    RECT 374.15 58.745 374.22 58.815 ;
    RECT 309.84 58.385 310.05 58.455 ;
    RECT 309.84 58.745 310.05 58.815 ;
    RECT 309.84 59.105 310.05 59.175 ;
    RECT 309.38 58.385 309.59 58.455 ;
    RECT 309.38 58.745 309.59 58.815 ;
    RECT 309.38 59.105 309.59 59.175 ;
    RECT 306.52 58.385 306.73 58.455 ;
    RECT 306.52 58.745 306.73 58.815 ;
    RECT 306.52 59.105 306.73 59.175 ;
    RECT 306.06 58.385 306.27 58.455 ;
    RECT 306.06 58.745 306.27 58.815 ;
    RECT 306.06 59.105 306.27 59.175 ;
    RECT 303.2 39.645 303.41 39.715 ;
    RECT 303.2 40.005 303.41 40.075 ;
    RECT 303.2 40.365 303.41 40.435 ;
    RECT 302.74 39.645 302.95 39.715 ;
    RECT 302.74 40.005 302.95 40.075 ;
    RECT 302.74 40.365 302.95 40.435 ;
    RECT 372.92 39.645 373.13 39.715 ;
    RECT 372.92 40.005 373.13 40.075 ;
    RECT 372.92 40.365 373.13 40.435 ;
    RECT 372.46 39.645 372.67 39.715 ;
    RECT 372.46 40.005 372.67 40.075 ;
    RECT 372.46 40.365 372.67 40.435 ;
    RECT 369.6 39.645 369.81 39.715 ;
    RECT 369.6 40.005 369.81 40.075 ;
    RECT 369.6 40.365 369.81 40.435 ;
    RECT 369.14 39.645 369.35 39.715 ;
    RECT 369.14 40.005 369.35 40.075 ;
    RECT 369.14 40.365 369.35 40.435 ;
    RECT 200.605 40.005 200.675 40.075 ;
    RECT 299.88 39.645 300.09 39.715 ;
    RECT 299.88 40.005 300.09 40.075 ;
    RECT 299.88 40.365 300.09 40.435 ;
    RECT 299.42 39.645 299.63 39.715 ;
    RECT 299.42 40.005 299.63 40.075 ;
    RECT 299.42 40.365 299.63 40.435 ;
    RECT 296.56 39.645 296.77 39.715 ;
    RECT 296.56 40.005 296.77 40.075 ;
    RECT 296.56 40.365 296.77 40.435 ;
    RECT 296.1 39.645 296.31 39.715 ;
    RECT 296.1 40.005 296.31 40.075 ;
    RECT 296.1 40.365 296.31 40.435 ;
    RECT 293.24 39.645 293.45 39.715 ;
    RECT 293.24 40.005 293.45 40.075 ;
    RECT 293.24 40.365 293.45 40.435 ;
    RECT 292.78 39.645 292.99 39.715 ;
    RECT 292.78 40.005 292.99 40.075 ;
    RECT 292.78 40.365 292.99 40.435 ;
    RECT 289.92 39.645 290.13 39.715 ;
    RECT 289.92 40.005 290.13 40.075 ;
    RECT 289.92 40.365 290.13 40.435 ;
    RECT 289.46 39.645 289.67 39.715 ;
    RECT 289.46 40.005 289.67 40.075 ;
    RECT 289.46 40.365 289.67 40.435 ;
    RECT 286.6 39.645 286.81 39.715 ;
    RECT 286.6 40.005 286.81 40.075 ;
    RECT 286.6 40.365 286.81 40.435 ;
    RECT 286.14 39.645 286.35 39.715 ;
    RECT 286.14 40.005 286.35 40.075 ;
    RECT 286.14 40.365 286.35 40.435 ;
    RECT 283.28 39.645 283.49 39.715 ;
    RECT 283.28 40.005 283.49 40.075 ;
    RECT 283.28 40.365 283.49 40.435 ;
    RECT 282.82 39.645 283.03 39.715 ;
    RECT 282.82 40.005 283.03 40.075 ;
    RECT 282.82 40.365 283.03 40.435 ;
    RECT 279.96 39.645 280.17 39.715 ;
    RECT 279.96 40.005 280.17 40.075 ;
    RECT 279.96 40.365 280.17 40.435 ;
    RECT 279.5 39.645 279.71 39.715 ;
    RECT 279.5 40.005 279.71 40.075 ;
    RECT 279.5 40.365 279.71 40.435 ;
    RECT 276.64 39.645 276.85 39.715 ;
    RECT 276.64 40.005 276.85 40.075 ;
    RECT 276.64 40.365 276.85 40.435 ;
    RECT 276.18 39.645 276.39 39.715 ;
    RECT 276.18 40.005 276.39 40.075 ;
    RECT 276.18 40.365 276.39 40.435 ;
    RECT 273.32 39.645 273.53 39.715 ;
    RECT 273.32 40.005 273.53 40.075 ;
    RECT 273.32 40.365 273.53 40.435 ;
    RECT 272.86 39.645 273.07 39.715 ;
    RECT 272.86 40.005 273.07 40.075 ;
    RECT 272.86 40.365 273.07 40.435 ;
    RECT 270.0 39.645 270.21 39.715 ;
    RECT 270.0 40.005 270.21 40.075 ;
    RECT 270.0 40.365 270.21 40.435 ;
    RECT 269.54 39.645 269.75 39.715 ;
    RECT 269.54 40.005 269.75 40.075 ;
    RECT 269.54 40.365 269.75 40.435 ;
    RECT 233.48 39.645 233.69 39.715 ;
    RECT 233.48 40.005 233.69 40.075 ;
    RECT 233.48 40.365 233.69 40.435 ;
    RECT 233.02 39.645 233.23 39.715 ;
    RECT 233.02 40.005 233.23 40.075 ;
    RECT 233.02 40.365 233.23 40.435 ;
    RECT 230.16 39.645 230.37 39.715 ;
    RECT 230.16 40.005 230.37 40.075 ;
    RECT 230.16 40.365 230.37 40.435 ;
    RECT 229.7 39.645 229.91 39.715 ;
    RECT 229.7 40.005 229.91 40.075 ;
    RECT 229.7 40.365 229.91 40.435 ;
    RECT 366.28 39.645 366.49 39.715 ;
    RECT 366.28 40.005 366.49 40.075 ;
    RECT 366.28 40.365 366.49 40.435 ;
    RECT 365.82 39.645 366.03 39.715 ;
    RECT 365.82 40.005 366.03 40.075 ;
    RECT 365.82 40.365 366.03 40.435 ;
    RECT 226.84 39.645 227.05 39.715 ;
    RECT 226.84 40.005 227.05 40.075 ;
    RECT 226.84 40.365 227.05 40.435 ;
    RECT 226.38 39.645 226.59 39.715 ;
    RECT 226.38 40.005 226.59 40.075 ;
    RECT 226.38 40.365 226.59 40.435 ;
    RECT 362.96 39.645 363.17 39.715 ;
    RECT 362.96 40.005 363.17 40.075 ;
    RECT 362.96 40.365 363.17 40.435 ;
    RECT 362.5 39.645 362.71 39.715 ;
    RECT 362.5 40.005 362.71 40.075 ;
    RECT 362.5 40.365 362.71 40.435 ;
    RECT 223.52 39.645 223.73 39.715 ;
    RECT 223.52 40.005 223.73 40.075 ;
    RECT 223.52 40.365 223.73 40.435 ;
    RECT 223.06 39.645 223.27 39.715 ;
    RECT 223.06 40.005 223.27 40.075 ;
    RECT 223.06 40.365 223.27 40.435 ;
    RECT 359.64 39.645 359.85 39.715 ;
    RECT 359.64 40.005 359.85 40.075 ;
    RECT 359.64 40.365 359.85 40.435 ;
    RECT 359.18 39.645 359.39 39.715 ;
    RECT 359.18 40.005 359.39 40.075 ;
    RECT 359.18 40.365 359.39 40.435 ;
    RECT 220.2 39.645 220.41 39.715 ;
    RECT 220.2 40.005 220.41 40.075 ;
    RECT 220.2 40.365 220.41 40.435 ;
    RECT 219.74 39.645 219.95 39.715 ;
    RECT 219.74 40.005 219.95 40.075 ;
    RECT 219.74 40.365 219.95 40.435 ;
    RECT 356.32 39.645 356.53 39.715 ;
    RECT 356.32 40.005 356.53 40.075 ;
    RECT 356.32 40.365 356.53 40.435 ;
    RECT 355.86 39.645 356.07 39.715 ;
    RECT 355.86 40.005 356.07 40.075 ;
    RECT 355.86 40.365 356.07 40.435 ;
    RECT 353.0 39.645 353.21 39.715 ;
    RECT 353.0 40.005 353.21 40.075 ;
    RECT 353.0 40.365 353.21 40.435 ;
    RECT 352.54 39.645 352.75 39.715 ;
    RECT 352.54 40.005 352.75 40.075 ;
    RECT 352.54 40.365 352.75 40.435 ;
    RECT 216.88 39.645 217.09 39.715 ;
    RECT 216.88 40.005 217.09 40.075 ;
    RECT 216.88 40.365 217.09 40.435 ;
    RECT 216.42 39.645 216.63 39.715 ;
    RECT 216.42 40.005 216.63 40.075 ;
    RECT 216.42 40.365 216.63 40.435 ;
    RECT 349.68 39.645 349.89 39.715 ;
    RECT 349.68 40.005 349.89 40.075 ;
    RECT 349.68 40.365 349.89 40.435 ;
    RECT 349.22 39.645 349.43 39.715 ;
    RECT 349.22 40.005 349.43 40.075 ;
    RECT 349.22 40.365 349.43 40.435 ;
    RECT 213.56 39.645 213.77 39.715 ;
    RECT 213.56 40.005 213.77 40.075 ;
    RECT 213.56 40.365 213.77 40.435 ;
    RECT 213.1 39.645 213.31 39.715 ;
    RECT 213.1 40.005 213.31 40.075 ;
    RECT 213.1 40.365 213.31 40.435 ;
    RECT 346.36 39.645 346.57 39.715 ;
    RECT 346.36 40.005 346.57 40.075 ;
    RECT 346.36 40.365 346.57 40.435 ;
    RECT 345.9 39.645 346.11 39.715 ;
    RECT 345.9 40.005 346.11 40.075 ;
    RECT 345.9 40.365 346.11 40.435 ;
    RECT 210.24 39.645 210.45 39.715 ;
    RECT 210.24 40.005 210.45 40.075 ;
    RECT 210.24 40.365 210.45 40.435 ;
    RECT 209.78 39.645 209.99 39.715 ;
    RECT 209.78 40.005 209.99 40.075 ;
    RECT 209.78 40.365 209.99 40.435 ;
    RECT 343.04 39.645 343.25 39.715 ;
    RECT 343.04 40.005 343.25 40.075 ;
    RECT 343.04 40.365 343.25 40.435 ;
    RECT 342.58 39.645 342.79 39.715 ;
    RECT 342.58 40.005 342.79 40.075 ;
    RECT 342.58 40.365 342.79 40.435 ;
    RECT 206.92 39.645 207.13 39.715 ;
    RECT 206.92 40.005 207.13 40.075 ;
    RECT 206.92 40.365 207.13 40.435 ;
    RECT 206.46 39.645 206.67 39.715 ;
    RECT 206.46 40.005 206.67 40.075 ;
    RECT 206.46 40.365 206.67 40.435 ;
    RECT 339.72 39.645 339.93 39.715 ;
    RECT 339.72 40.005 339.93 40.075 ;
    RECT 339.72 40.365 339.93 40.435 ;
    RECT 339.26 39.645 339.47 39.715 ;
    RECT 339.26 40.005 339.47 40.075 ;
    RECT 339.26 40.365 339.47 40.435 ;
    RECT 203.6 39.645 203.81 39.715 ;
    RECT 203.6 40.005 203.81 40.075 ;
    RECT 203.6 40.365 203.81 40.435 ;
    RECT 203.14 39.645 203.35 39.715 ;
    RECT 203.14 40.005 203.35 40.075 ;
    RECT 203.14 40.365 203.35 40.435 ;
    RECT 336.4 39.645 336.61 39.715 ;
    RECT 336.4 40.005 336.61 40.075 ;
    RECT 336.4 40.365 336.61 40.435 ;
    RECT 335.94 39.645 336.15 39.715 ;
    RECT 335.94 40.005 336.15 40.075 ;
    RECT 335.94 40.365 336.15 40.435 ;
    RECT 266.68 39.645 266.89 39.715 ;
    RECT 266.68 40.005 266.89 40.075 ;
    RECT 266.68 40.365 266.89 40.435 ;
    RECT 266.22 39.645 266.43 39.715 ;
    RECT 266.22 40.005 266.43 40.075 ;
    RECT 266.22 40.365 266.43 40.435 ;
    RECT 263.36 39.645 263.57 39.715 ;
    RECT 263.36 40.005 263.57 40.075 ;
    RECT 263.36 40.365 263.57 40.435 ;
    RECT 262.9 39.645 263.11 39.715 ;
    RECT 262.9 40.005 263.11 40.075 ;
    RECT 262.9 40.365 263.11 40.435 ;
    RECT 260.04 39.645 260.25 39.715 ;
    RECT 260.04 40.005 260.25 40.075 ;
    RECT 260.04 40.365 260.25 40.435 ;
    RECT 259.58 39.645 259.79 39.715 ;
    RECT 259.58 40.005 259.79 40.075 ;
    RECT 259.58 40.365 259.79 40.435 ;
    RECT 256.72 39.645 256.93 39.715 ;
    RECT 256.72 40.005 256.93 40.075 ;
    RECT 256.72 40.365 256.93 40.435 ;
    RECT 256.26 39.645 256.47 39.715 ;
    RECT 256.26 40.005 256.47 40.075 ;
    RECT 256.26 40.365 256.47 40.435 ;
    RECT 253.4 39.645 253.61 39.715 ;
    RECT 253.4 40.005 253.61 40.075 ;
    RECT 253.4 40.365 253.61 40.435 ;
    RECT 252.94 39.645 253.15 39.715 ;
    RECT 252.94 40.005 253.15 40.075 ;
    RECT 252.94 40.365 253.15 40.435 ;
    RECT 250.08 39.645 250.29 39.715 ;
    RECT 250.08 40.005 250.29 40.075 ;
    RECT 250.08 40.365 250.29 40.435 ;
    RECT 249.62 39.645 249.83 39.715 ;
    RECT 249.62 40.005 249.83 40.075 ;
    RECT 249.62 40.365 249.83 40.435 ;
    RECT 246.76 39.645 246.97 39.715 ;
    RECT 246.76 40.005 246.97 40.075 ;
    RECT 246.76 40.365 246.97 40.435 ;
    RECT 246.3 39.645 246.51 39.715 ;
    RECT 246.3 40.005 246.51 40.075 ;
    RECT 246.3 40.365 246.51 40.435 ;
    RECT 243.44 39.645 243.65 39.715 ;
    RECT 243.44 40.005 243.65 40.075 ;
    RECT 243.44 40.365 243.65 40.435 ;
    RECT 242.98 39.645 243.19 39.715 ;
    RECT 242.98 40.005 243.19 40.075 ;
    RECT 242.98 40.365 243.19 40.435 ;
    RECT 240.12 39.645 240.33 39.715 ;
    RECT 240.12 40.005 240.33 40.075 ;
    RECT 240.12 40.365 240.33 40.435 ;
    RECT 239.66 39.645 239.87 39.715 ;
    RECT 239.66 40.005 239.87 40.075 ;
    RECT 239.66 40.365 239.87 40.435 ;
    RECT 236.8 39.645 237.01 39.715 ;
    RECT 236.8 40.005 237.01 40.075 ;
    RECT 236.8 40.365 237.01 40.435 ;
    RECT 236.34 39.645 236.55 39.715 ;
    RECT 236.34 40.005 236.55 40.075 ;
    RECT 236.34 40.365 236.55 40.435 ;
    RECT 374.15 40.005 374.22 40.075 ;
    RECT 333.08 39.645 333.29 39.715 ;
    RECT 333.08 40.005 333.29 40.075 ;
    RECT 333.08 40.365 333.29 40.435 ;
    RECT 332.62 39.645 332.83 39.715 ;
    RECT 332.62 40.005 332.83 40.075 ;
    RECT 332.62 40.365 332.83 40.435 ;
    RECT 329.76 39.645 329.97 39.715 ;
    RECT 329.76 40.005 329.97 40.075 ;
    RECT 329.76 40.365 329.97 40.435 ;
    RECT 329.3 39.645 329.51 39.715 ;
    RECT 329.3 40.005 329.51 40.075 ;
    RECT 329.3 40.365 329.51 40.435 ;
    RECT 326.44 39.645 326.65 39.715 ;
    RECT 326.44 40.005 326.65 40.075 ;
    RECT 326.44 40.365 326.65 40.435 ;
    RECT 325.98 39.645 326.19 39.715 ;
    RECT 325.98 40.005 326.19 40.075 ;
    RECT 325.98 40.365 326.19 40.435 ;
    RECT 323.12 39.645 323.33 39.715 ;
    RECT 323.12 40.005 323.33 40.075 ;
    RECT 323.12 40.365 323.33 40.435 ;
    RECT 322.66 39.645 322.87 39.715 ;
    RECT 322.66 40.005 322.87 40.075 ;
    RECT 322.66 40.365 322.87 40.435 ;
    RECT 319.8 39.645 320.01 39.715 ;
    RECT 319.8 40.005 320.01 40.075 ;
    RECT 319.8 40.365 320.01 40.435 ;
    RECT 319.34 39.645 319.55 39.715 ;
    RECT 319.34 40.005 319.55 40.075 ;
    RECT 319.34 40.365 319.55 40.435 ;
    RECT 316.48 39.645 316.69 39.715 ;
    RECT 316.48 40.005 316.69 40.075 ;
    RECT 316.48 40.365 316.69 40.435 ;
    RECT 316.02 39.645 316.23 39.715 ;
    RECT 316.02 40.005 316.23 40.075 ;
    RECT 316.02 40.365 316.23 40.435 ;
    RECT 313.16 39.645 313.37 39.715 ;
    RECT 313.16 40.005 313.37 40.075 ;
    RECT 313.16 40.365 313.37 40.435 ;
    RECT 312.7 39.645 312.91 39.715 ;
    RECT 312.7 40.005 312.91 40.075 ;
    RECT 312.7 40.365 312.91 40.435 ;
    RECT 309.84 39.645 310.05 39.715 ;
    RECT 309.84 40.005 310.05 40.075 ;
    RECT 309.84 40.365 310.05 40.435 ;
    RECT 309.38 39.645 309.59 39.715 ;
    RECT 309.38 40.005 309.59 40.075 ;
    RECT 309.38 40.365 309.59 40.435 ;
    RECT 306.52 39.645 306.73 39.715 ;
    RECT 306.52 40.005 306.73 40.075 ;
    RECT 306.52 40.365 306.73 40.435 ;
    RECT 306.06 39.645 306.27 39.715 ;
    RECT 306.06 40.005 306.27 40.075 ;
    RECT 306.06 40.365 306.27 40.435 ;
    RECT 303.2 38.925 303.41 38.995 ;
    RECT 303.2 39.285 303.41 39.355 ;
    RECT 303.2 39.645 303.41 39.715 ;
    RECT 302.74 38.925 302.95 38.995 ;
    RECT 302.74 39.285 302.95 39.355 ;
    RECT 302.74 39.645 302.95 39.715 ;
    RECT 372.92 38.925 373.13 38.995 ;
    RECT 372.92 39.285 373.13 39.355 ;
    RECT 372.92 39.645 373.13 39.715 ;
    RECT 372.46 38.925 372.67 38.995 ;
    RECT 372.46 39.285 372.67 39.355 ;
    RECT 372.46 39.645 372.67 39.715 ;
    RECT 369.6 38.925 369.81 38.995 ;
    RECT 369.6 39.285 369.81 39.355 ;
    RECT 369.6 39.645 369.81 39.715 ;
    RECT 369.14 38.925 369.35 38.995 ;
    RECT 369.14 39.285 369.35 39.355 ;
    RECT 369.14 39.645 369.35 39.715 ;
    RECT 200.605 39.285 200.675 39.355 ;
    RECT 299.88 38.925 300.09 38.995 ;
    RECT 299.88 39.285 300.09 39.355 ;
    RECT 299.88 39.645 300.09 39.715 ;
    RECT 299.42 38.925 299.63 38.995 ;
    RECT 299.42 39.285 299.63 39.355 ;
    RECT 299.42 39.645 299.63 39.715 ;
    RECT 296.56 38.925 296.77 38.995 ;
    RECT 296.56 39.285 296.77 39.355 ;
    RECT 296.56 39.645 296.77 39.715 ;
    RECT 296.1 38.925 296.31 38.995 ;
    RECT 296.1 39.285 296.31 39.355 ;
    RECT 296.1 39.645 296.31 39.715 ;
    RECT 293.24 38.925 293.45 38.995 ;
    RECT 293.24 39.285 293.45 39.355 ;
    RECT 293.24 39.645 293.45 39.715 ;
    RECT 292.78 38.925 292.99 38.995 ;
    RECT 292.78 39.285 292.99 39.355 ;
    RECT 292.78 39.645 292.99 39.715 ;
    RECT 289.92 38.925 290.13 38.995 ;
    RECT 289.92 39.285 290.13 39.355 ;
    RECT 289.92 39.645 290.13 39.715 ;
    RECT 289.46 38.925 289.67 38.995 ;
    RECT 289.46 39.285 289.67 39.355 ;
    RECT 289.46 39.645 289.67 39.715 ;
    RECT 286.6 38.925 286.81 38.995 ;
    RECT 286.6 39.285 286.81 39.355 ;
    RECT 286.6 39.645 286.81 39.715 ;
    RECT 286.14 38.925 286.35 38.995 ;
    RECT 286.14 39.285 286.35 39.355 ;
    RECT 286.14 39.645 286.35 39.715 ;
    RECT 283.28 38.925 283.49 38.995 ;
    RECT 283.28 39.285 283.49 39.355 ;
    RECT 283.28 39.645 283.49 39.715 ;
    RECT 282.82 38.925 283.03 38.995 ;
    RECT 282.82 39.285 283.03 39.355 ;
    RECT 282.82 39.645 283.03 39.715 ;
    RECT 279.96 38.925 280.17 38.995 ;
    RECT 279.96 39.285 280.17 39.355 ;
    RECT 279.96 39.645 280.17 39.715 ;
    RECT 279.5 38.925 279.71 38.995 ;
    RECT 279.5 39.285 279.71 39.355 ;
    RECT 279.5 39.645 279.71 39.715 ;
    RECT 276.64 38.925 276.85 38.995 ;
    RECT 276.64 39.285 276.85 39.355 ;
    RECT 276.64 39.645 276.85 39.715 ;
    RECT 276.18 38.925 276.39 38.995 ;
    RECT 276.18 39.285 276.39 39.355 ;
    RECT 276.18 39.645 276.39 39.715 ;
    RECT 273.32 38.925 273.53 38.995 ;
    RECT 273.32 39.285 273.53 39.355 ;
    RECT 273.32 39.645 273.53 39.715 ;
    RECT 272.86 38.925 273.07 38.995 ;
    RECT 272.86 39.285 273.07 39.355 ;
    RECT 272.86 39.645 273.07 39.715 ;
    RECT 270.0 38.925 270.21 38.995 ;
    RECT 270.0 39.285 270.21 39.355 ;
    RECT 270.0 39.645 270.21 39.715 ;
    RECT 269.54 38.925 269.75 38.995 ;
    RECT 269.54 39.285 269.75 39.355 ;
    RECT 269.54 39.645 269.75 39.715 ;
    RECT 233.48 38.925 233.69 38.995 ;
    RECT 233.48 39.285 233.69 39.355 ;
    RECT 233.48 39.645 233.69 39.715 ;
    RECT 233.02 38.925 233.23 38.995 ;
    RECT 233.02 39.285 233.23 39.355 ;
    RECT 233.02 39.645 233.23 39.715 ;
    RECT 230.16 38.925 230.37 38.995 ;
    RECT 230.16 39.285 230.37 39.355 ;
    RECT 230.16 39.645 230.37 39.715 ;
    RECT 229.7 38.925 229.91 38.995 ;
    RECT 229.7 39.285 229.91 39.355 ;
    RECT 229.7 39.645 229.91 39.715 ;
    RECT 366.28 38.925 366.49 38.995 ;
    RECT 366.28 39.285 366.49 39.355 ;
    RECT 366.28 39.645 366.49 39.715 ;
    RECT 365.82 38.925 366.03 38.995 ;
    RECT 365.82 39.285 366.03 39.355 ;
    RECT 365.82 39.645 366.03 39.715 ;
    RECT 226.84 38.925 227.05 38.995 ;
    RECT 226.84 39.285 227.05 39.355 ;
    RECT 226.84 39.645 227.05 39.715 ;
    RECT 226.38 38.925 226.59 38.995 ;
    RECT 226.38 39.285 226.59 39.355 ;
    RECT 226.38 39.645 226.59 39.715 ;
    RECT 362.96 38.925 363.17 38.995 ;
    RECT 362.96 39.285 363.17 39.355 ;
    RECT 362.96 39.645 363.17 39.715 ;
    RECT 362.5 38.925 362.71 38.995 ;
    RECT 362.5 39.285 362.71 39.355 ;
    RECT 362.5 39.645 362.71 39.715 ;
    RECT 223.52 38.925 223.73 38.995 ;
    RECT 223.52 39.285 223.73 39.355 ;
    RECT 223.52 39.645 223.73 39.715 ;
    RECT 223.06 38.925 223.27 38.995 ;
    RECT 223.06 39.285 223.27 39.355 ;
    RECT 223.06 39.645 223.27 39.715 ;
    RECT 359.64 38.925 359.85 38.995 ;
    RECT 359.64 39.285 359.85 39.355 ;
    RECT 359.64 39.645 359.85 39.715 ;
    RECT 359.18 38.925 359.39 38.995 ;
    RECT 359.18 39.285 359.39 39.355 ;
    RECT 359.18 39.645 359.39 39.715 ;
    RECT 220.2 38.925 220.41 38.995 ;
    RECT 220.2 39.285 220.41 39.355 ;
    RECT 220.2 39.645 220.41 39.715 ;
    RECT 219.74 38.925 219.95 38.995 ;
    RECT 219.74 39.285 219.95 39.355 ;
    RECT 219.74 39.645 219.95 39.715 ;
    RECT 356.32 38.925 356.53 38.995 ;
    RECT 356.32 39.285 356.53 39.355 ;
    RECT 356.32 39.645 356.53 39.715 ;
    RECT 355.86 38.925 356.07 38.995 ;
    RECT 355.86 39.285 356.07 39.355 ;
    RECT 355.86 39.645 356.07 39.715 ;
    RECT 353.0 38.925 353.21 38.995 ;
    RECT 353.0 39.285 353.21 39.355 ;
    RECT 353.0 39.645 353.21 39.715 ;
    RECT 352.54 38.925 352.75 38.995 ;
    RECT 352.54 39.285 352.75 39.355 ;
    RECT 352.54 39.645 352.75 39.715 ;
    RECT 216.88 38.925 217.09 38.995 ;
    RECT 216.88 39.285 217.09 39.355 ;
    RECT 216.88 39.645 217.09 39.715 ;
    RECT 216.42 38.925 216.63 38.995 ;
    RECT 216.42 39.285 216.63 39.355 ;
    RECT 216.42 39.645 216.63 39.715 ;
    RECT 349.68 38.925 349.89 38.995 ;
    RECT 349.68 39.285 349.89 39.355 ;
    RECT 349.68 39.645 349.89 39.715 ;
    RECT 349.22 38.925 349.43 38.995 ;
    RECT 349.22 39.285 349.43 39.355 ;
    RECT 349.22 39.645 349.43 39.715 ;
    RECT 213.56 38.925 213.77 38.995 ;
    RECT 213.56 39.285 213.77 39.355 ;
    RECT 213.56 39.645 213.77 39.715 ;
    RECT 213.1 38.925 213.31 38.995 ;
    RECT 213.1 39.285 213.31 39.355 ;
    RECT 213.1 39.645 213.31 39.715 ;
    RECT 346.36 38.925 346.57 38.995 ;
    RECT 346.36 39.285 346.57 39.355 ;
    RECT 346.36 39.645 346.57 39.715 ;
    RECT 345.9 38.925 346.11 38.995 ;
    RECT 345.9 39.285 346.11 39.355 ;
    RECT 345.9 39.645 346.11 39.715 ;
    RECT 210.24 38.925 210.45 38.995 ;
    RECT 210.24 39.285 210.45 39.355 ;
    RECT 210.24 39.645 210.45 39.715 ;
    RECT 209.78 38.925 209.99 38.995 ;
    RECT 209.78 39.285 209.99 39.355 ;
    RECT 209.78 39.645 209.99 39.715 ;
    RECT 343.04 38.925 343.25 38.995 ;
    RECT 343.04 39.285 343.25 39.355 ;
    RECT 343.04 39.645 343.25 39.715 ;
    RECT 342.58 38.925 342.79 38.995 ;
    RECT 342.58 39.285 342.79 39.355 ;
    RECT 342.58 39.645 342.79 39.715 ;
    RECT 206.92 38.925 207.13 38.995 ;
    RECT 206.92 39.285 207.13 39.355 ;
    RECT 206.92 39.645 207.13 39.715 ;
    RECT 206.46 38.925 206.67 38.995 ;
    RECT 206.46 39.285 206.67 39.355 ;
    RECT 206.46 39.645 206.67 39.715 ;
    RECT 339.72 38.925 339.93 38.995 ;
    RECT 339.72 39.285 339.93 39.355 ;
    RECT 339.72 39.645 339.93 39.715 ;
    RECT 339.26 38.925 339.47 38.995 ;
    RECT 339.26 39.285 339.47 39.355 ;
    RECT 339.26 39.645 339.47 39.715 ;
    RECT 203.6 38.925 203.81 38.995 ;
    RECT 203.6 39.285 203.81 39.355 ;
    RECT 203.6 39.645 203.81 39.715 ;
    RECT 203.14 38.925 203.35 38.995 ;
    RECT 203.14 39.285 203.35 39.355 ;
    RECT 203.14 39.645 203.35 39.715 ;
    RECT 336.4 38.925 336.61 38.995 ;
    RECT 336.4 39.285 336.61 39.355 ;
    RECT 336.4 39.645 336.61 39.715 ;
    RECT 335.94 38.925 336.15 38.995 ;
    RECT 335.94 39.285 336.15 39.355 ;
    RECT 335.94 39.645 336.15 39.715 ;
    RECT 266.68 38.925 266.89 38.995 ;
    RECT 266.68 39.285 266.89 39.355 ;
    RECT 266.68 39.645 266.89 39.715 ;
    RECT 266.22 38.925 266.43 38.995 ;
    RECT 266.22 39.285 266.43 39.355 ;
    RECT 266.22 39.645 266.43 39.715 ;
    RECT 263.36 38.925 263.57 38.995 ;
    RECT 263.36 39.285 263.57 39.355 ;
    RECT 263.36 39.645 263.57 39.715 ;
    RECT 262.9 38.925 263.11 38.995 ;
    RECT 262.9 39.285 263.11 39.355 ;
    RECT 262.9 39.645 263.11 39.715 ;
    RECT 260.04 38.925 260.25 38.995 ;
    RECT 260.04 39.285 260.25 39.355 ;
    RECT 260.04 39.645 260.25 39.715 ;
    RECT 259.58 38.925 259.79 38.995 ;
    RECT 259.58 39.285 259.79 39.355 ;
    RECT 259.58 39.645 259.79 39.715 ;
    RECT 256.72 38.925 256.93 38.995 ;
    RECT 256.72 39.285 256.93 39.355 ;
    RECT 256.72 39.645 256.93 39.715 ;
    RECT 256.26 38.925 256.47 38.995 ;
    RECT 256.26 39.285 256.47 39.355 ;
    RECT 256.26 39.645 256.47 39.715 ;
    RECT 253.4 38.925 253.61 38.995 ;
    RECT 253.4 39.285 253.61 39.355 ;
    RECT 253.4 39.645 253.61 39.715 ;
    RECT 252.94 38.925 253.15 38.995 ;
    RECT 252.94 39.285 253.15 39.355 ;
    RECT 252.94 39.645 253.15 39.715 ;
    RECT 250.08 38.925 250.29 38.995 ;
    RECT 250.08 39.285 250.29 39.355 ;
    RECT 250.08 39.645 250.29 39.715 ;
    RECT 249.62 38.925 249.83 38.995 ;
    RECT 249.62 39.285 249.83 39.355 ;
    RECT 249.62 39.645 249.83 39.715 ;
    RECT 246.76 38.925 246.97 38.995 ;
    RECT 246.76 39.285 246.97 39.355 ;
    RECT 246.76 39.645 246.97 39.715 ;
    RECT 246.3 38.925 246.51 38.995 ;
    RECT 246.3 39.285 246.51 39.355 ;
    RECT 246.3 39.645 246.51 39.715 ;
    RECT 243.44 38.925 243.65 38.995 ;
    RECT 243.44 39.285 243.65 39.355 ;
    RECT 243.44 39.645 243.65 39.715 ;
    RECT 242.98 38.925 243.19 38.995 ;
    RECT 242.98 39.285 243.19 39.355 ;
    RECT 242.98 39.645 243.19 39.715 ;
    RECT 240.12 38.925 240.33 38.995 ;
    RECT 240.12 39.285 240.33 39.355 ;
    RECT 240.12 39.645 240.33 39.715 ;
    RECT 239.66 38.925 239.87 38.995 ;
    RECT 239.66 39.285 239.87 39.355 ;
    RECT 239.66 39.645 239.87 39.715 ;
    RECT 236.8 38.925 237.01 38.995 ;
    RECT 236.8 39.285 237.01 39.355 ;
    RECT 236.8 39.645 237.01 39.715 ;
    RECT 236.34 38.925 236.55 38.995 ;
    RECT 236.34 39.285 236.55 39.355 ;
    RECT 236.34 39.645 236.55 39.715 ;
    RECT 374.15 39.285 374.22 39.355 ;
    RECT 333.08 38.925 333.29 38.995 ;
    RECT 333.08 39.285 333.29 39.355 ;
    RECT 333.08 39.645 333.29 39.715 ;
    RECT 332.62 38.925 332.83 38.995 ;
    RECT 332.62 39.285 332.83 39.355 ;
    RECT 332.62 39.645 332.83 39.715 ;
    RECT 329.76 38.925 329.97 38.995 ;
    RECT 329.76 39.285 329.97 39.355 ;
    RECT 329.76 39.645 329.97 39.715 ;
    RECT 329.3 38.925 329.51 38.995 ;
    RECT 329.3 39.285 329.51 39.355 ;
    RECT 329.3 39.645 329.51 39.715 ;
    RECT 326.44 38.925 326.65 38.995 ;
    RECT 326.44 39.285 326.65 39.355 ;
    RECT 326.44 39.645 326.65 39.715 ;
    RECT 325.98 38.925 326.19 38.995 ;
    RECT 325.98 39.285 326.19 39.355 ;
    RECT 325.98 39.645 326.19 39.715 ;
    RECT 323.12 38.925 323.33 38.995 ;
    RECT 323.12 39.285 323.33 39.355 ;
    RECT 323.12 39.645 323.33 39.715 ;
    RECT 322.66 38.925 322.87 38.995 ;
    RECT 322.66 39.285 322.87 39.355 ;
    RECT 322.66 39.645 322.87 39.715 ;
    RECT 319.8 38.925 320.01 38.995 ;
    RECT 319.8 39.285 320.01 39.355 ;
    RECT 319.8 39.645 320.01 39.715 ;
    RECT 319.34 38.925 319.55 38.995 ;
    RECT 319.34 39.285 319.55 39.355 ;
    RECT 319.34 39.645 319.55 39.715 ;
    RECT 316.48 38.925 316.69 38.995 ;
    RECT 316.48 39.285 316.69 39.355 ;
    RECT 316.48 39.645 316.69 39.715 ;
    RECT 316.02 38.925 316.23 38.995 ;
    RECT 316.02 39.285 316.23 39.355 ;
    RECT 316.02 39.645 316.23 39.715 ;
    RECT 313.16 38.925 313.37 38.995 ;
    RECT 313.16 39.285 313.37 39.355 ;
    RECT 313.16 39.645 313.37 39.715 ;
    RECT 312.7 38.925 312.91 38.995 ;
    RECT 312.7 39.285 312.91 39.355 ;
    RECT 312.7 39.645 312.91 39.715 ;
    RECT 309.84 38.925 310.05 38.995 ;
    RECT 309.84 39.285 310.05 39.355 ;
    RECT 309.84 39.645 310.05 39.715 ;
    RECT 309.38 38.925 309.59 38.995 ;
    RECT 309.38 39.285 309.59 39.355 ;
    RECT 309.38 39.645 309.59 39.715 ;
    RECT 306.52 38.925 306.73 38.995 ;
    RECT 306.52 39.285 306.73 39.355 ;
    RECT 306.52 39.645 306.73 39.715 ;
    RECT 306.06 38.925 306.27 38.995 ;
    RECT 306.06 39.285 306.27 39.355 ;
    RECT 306.06 39.645 306.27 39.715 ;
    RECT 303.2 38.205 303.41 38.275 ;
    RECT 303.2 38.565 303.41 38.635 ;
    RECT 303.2 38.925 303.41 38.995 ;
    RECT 302.74 38.205 302.95 38.275 ;
    RECT 302.74 38.565 302.95 38.635 ;
    RECT 302.74 38.925 302.95 38.995 ;
    RECT 372.92 38.205 373.13 38.275 ;
    RECT 372.92 38.565 373.13 38.635 ;
    RECT 372.92 38.925 373.13 38.995 ;
    RECT 372.46 38.205 372.67 38.275 ;
    RECT 372.46 38.565 372.67 38.635 ;
    RECT 372.46 38.925 372.67 38.995 ;
    RECT 369.6 38.205 369.81 38.275 ;
    RECT 369.6 38.565 369.81 38.635 ;
    RECT 369.6 38.925 369.81 38.995 ;
    RECT 369.14 38.205 369.35 38.275 ;
    RECT 369.14 38.565 369.35 38.635 ;
    RECT 369.14 38.925 369.35 38.995 ;
    RECT 200.605 38.565 200.675 38.635 ;
    RECT 299.88 38.205 300.09 38.275 ;
    RECT 299.88 38.565 300.09 38.635 ;
    RECT 299.88 38.925 300.09 38.995 ;
    RECT 299.42 38.205 299.63 38.275 ;
    RECT 299.42 38.565 299.63 38.635 ;
    RECT 299.42 38.925 299.63 38.995 ;
    RECT 296.56 38.205 296.77 38.275 ;
    RECT 296.56 38.565 296.77 38.635 ;
    RECT 296.56 38.925 296.77 38.995 ;
    RECT 296.1 38.205 296.31 38.275 ;
    RECT 296.1 38.565 296.31 38.635 ;
    RECT 296.1 38.925 296.31 38.995 ;
    RECT 293.24 38.205 293.45 38.275 ;
    RECT 293.24 38.565 293.45 38.635 ;
    RECT 293.24 38.925 293.45 38.995 ;
    RECT 292.78 38.205 292.99 38.275 ;
    RECT 292.78 38.565 292.99 38.635 ;
    RECT 292.78 38.925 292.99 38.995 ;
    RECT 289.92 38.205 290.13 38.275 ;
    RECT 289.92 38.565 290.13 38.635 ;
    RECT 289.92 38.925 290.13 38.995 ;
    RECT 289.46 38.205 289.67 38.275 ;
    RECT 289.46 38.565 289.67 38.635 ;
    RECT 289.46 38.925 289.67 38.995 ;
    RECT 286.6 38.205 286.81 38.275 ;
    RECT 286.6 38.565 286.81 38.635 ;
    RECT 286.6 38.925 286.81 38.995 ;
    RECT 286.14 38.205 286.35 38.275 ;
    RECT 286.14 38.565 286.35 38.635 ;
    RECT 286.14 38.925 286.35 38.995 ;
    RECT 283.28 38.205 283.49 38.275 ;
    RECT 283.28 38.565 283.49 38.635 ;
    RECT 283.28 38.925 283.49 38.995 ;
    RECT 282.82 38.205 283.03 38.275 ;
    RECT 282.82 38.565 283.03 38.635 ;
    RECT 282.82 38.925 283.03 38.995 ;
    RECT 279.96 38.205 280.17 38.275 ;
    RECT 279.96 38.565 280.17 38.635 ;
    RECT 279.96 38.925 280.17 38.995 ;
    RECT 279.5 38.205 279.71 38.275 ;
    RECT 279.5 38.565 279.71 38.635 ;
    RECT 279.5 38.925 279.71 38.995 ;
    RECT 276.64 38.205 276.85 38.275 ;
    RECT 276.64 38.565 276.85 38.635 ;
    RECT 276.64 38.925 276.85 38.995 ;
    RECT 276.18 38.205 276.39 38.275 ;
    RECT 276.18 38.565 276.39 38.635 ;
    RECT 276.18 38.925 276.39 38.995 ;
    RECT 273.32 38.205 273.53 38.275 ;
    RECT 273.32 38.565 273.53 38.635 ;
    RECT 273.32 38.925 273.53 38.995 ;
    RECT 272.86 38.205 273.07 38.275 ;
    RECT 272.86 38.565 273.07 38.635 ;
    RECT 272.86 38.925 273.07 38.995 ;
    RECT 270.0 38.205 270.21 38.275 ;
    RECT 270.0 38.565 270.21 38.635 ;
    RECT 270.0 38.925 270.21 38.995 ;
    RECT 269.54 38.205 269.75 38.275 ;
    RECT 269.54 38.565 269.75 38.635 ;
    RECT 269.54 38.925 269.75 38.995 ;
    RECT 233.48 38.205 233.69 38.275 ;
    RECT 233.48 38.565 233.69 38.635 ;
    RECT 233.48 38.925 233.69 38.995 ;
    RECT 233.02 38.205 233.23 38.275 ;
    RECT 233.02 38.565 233.23 38.635 ;
    RECT 233.02 38.925 233.23 38.995 ;
    RECT 230.16 38.205 230.37 38.275 ;
    RECT 230.16 38.565 230.37 38.635 ;
    RECT 230.16 38.925 230.37 38.995 ;
    RECT 229.7 38.205 229.91 38.275 ;
    RECT 229.7 38.565 229.91 38.635 ;
    RECT 229.7 38.925 229.91 38.995 ;
    RECT 366.28 38.205 366.49 38.275 ;
    RECT 366.28 38.565 366.49 38.635 ;
    RECT 366.28 38.925 366.49 38.995 ;
    RECT 365.82 38.205 366.03 38.275 ;
    RECT 365.82 38.565 366.03 38.635 ;
    RECT 365.82 38.925 366.03 38.995 ;
    RECT 226.84 38.205 227.05 38.275 ;
    RECT 226.84 38.565 227.05 38.635 ;
    RECT 226.84 38.925 227.05 38.995 ;
    RECT 226.38 38.205 226.59 38.275 ;
    RECT 226.38 38.565 226.59 38.635 ;
    RECT 226.38 38.925 226.59 38.995 ;
    RECT 362.96 38.205 363.17 38.275 ;
    RECT 362.96 38.565 363.17 38.635 ;
    RECT 362.96 38.925 363.17 38.995 ;
    RECT 362.5 38.205 362.71 38.275 ;
    RECT 362.5 38.565 362.71 38.635 ;
    RECT 362.5 38.925 362.71 38.995 ;
    RECT 223.52 38.205 223.73 38.275 ;
    RECT 223.52 38.565 223.73 38.635 ;
    RECT 223.52 38.925 223.73 38.995 ;
    RECT 223.06 38.205 223.27 38.275 ;
    RECT 223.06 38.565 223.27 38.635 ;
    RECT 223.06 38.925 223.27 38.995 ;
    RECT 359.64 38.205 359.85 38.275 ;
    RECT 359.64 38.565 359.85 38.635 ;
    RECT 359.64 38.925 359.85 38.995 ;
    RECT 359.18 38.205 359.39 38.275 ;
    RECT 359.18 38.565 359.39 38.635 ;
    RECT 359.18 38.925 359.39 38.995 ;
    RECT 220.2 38.205 220.41 38.275 ;
    RECT 220.2 38.565 220.41 38.635 ;
    RECT 220.2 38.925 220.41 38.995 ;
    RECT 219.74 38.205 219.95 38.275 ;
    RECT 219.74 38.565 219.95 38.635 ;
    RECT 219.74 38.925 219.95 38.995 ;
    RECT 356.32 38.205 356.53 38.275 ;
    RECT 356.32 38.565 356.53 38.635 ;
    RECT 356.32 38.925 356.53 38.995 ;
    RECT 355.86 38.205 356.07 38.275 ;
    RECT 355.86 38.565 356.07 38.635 ;
    RECT 355.86 38.925 356.07 38.995 ;
    RECT 353.0 38.205 353.21 38.275 ;
    RECT 353.0 38.565 353.21 38.635 ;
    RECT 353.0 38.925 353.21 38.995 ;
    RECT 352.54 38.205 352.75 38.275 ;
    RECT 352.54 38.565 352.75 38.635 ;
    RECT 352.54 38.925 352.75 38.995 ;
    RECT 216.88 38.205 217.09 38.275 ;
    RECT 216.88 38.565 217.09 38.635 ;
    RECT 216.88 38.925 217.09 38.995 ;
    RECT 216.42 38.205 216.63 38.275 ;
    RECT 216.42 38.565 216.63 38.635 ;
    RECT 216.42 38.925 216.63 38.995 ;
    RECT 349.68 38.205 349.89 38.275 ;
    RECT 349.68 38.565 349.89 38.635 ;
    RECT 349.68 38.925 349.89 38.995 ;
    RECT 349.22 38.205 349.43 38.275 ;
    RECT 349.22 38.565 349.43 38.635 ;
    RECT 349.22 38.925 349.43 38.995 ;
    RECT 213.56 38.205 213.77 38.275 ;
    RECT 213.56 38.565 213.77 38.635 ;
    RECT 213.56 38.925 213.77 38.995 ;
    RECT 213.1 38.205 213.31 38.275 ;
    RECT 213.1 38.565 213.31 38.635 ;
    RECT 213.1 38.925 213.31 38.995 ;
    RECT 346.36 38.205 346.57 38.275 ;
    RECT 346.36 38.565 346.57 38.635 ;
    RECT 346.36 38.925 346.57 38.995 ;
    RECT 345.9 38.205 346.11 38.275 ;
    RECT 345.9 38.565 346.11 38.635 ;
    RECT 345.9 38.925 346.11 38.995 ;
    RECT 210.24 38.205 210.45 38.275 ;
    RECT 210.24 38.565 210.45 38.635 ;
    RECT 210.24 38.925 210.45 38.995 ;
    RECT 209.78 38.205 209.99 38.275 ;
    RECT 209.78 38.565 209.99 38.635 ;
    RECT 209.78 38.925 209.99 38.995 ;
    RECT 343.04 38.205 343.25 38.275 ;
    RECT 343.04 38.565 343.25 38.635 ;
    RECT 343.04 38.925 343.25 38.995 ;
    RECT 342.58 38.205 342.79 38.275 ;
    RECT 342.58 38.565 342.79 38.635 ;
    RECT 342.58 38.925 342.79 38.995 ;
    RECT 206.92 38.205 207.13 38.275 ;
    RECT 206.92 38.565 207.13 38.635 ;
    RECT 206.92 38.925 207.13 38.995 ;
    RECT 206.46 38.205 206.67 38.275 ;
    RECT 206.46 38.565 206.67 38.635 ;
    RECT 206.46 38.925 206.67 38.995 ;
    RECT 339.72 38.205 339.93 38.275 ;
    RECT 339.72 38.565 339.93 38.635 ;
    RECT 339.72 38.925 339.93 38.995 ;
    RECT 339.26 38.205 339.47 38.275 ;
    RECT 339.26 38.565 339.47 38.635 ;
    RECT 339.26 38.925 339.47 38.995 ;
    RECT 203.6 38.205 203.81 38.275 ;
    RECT 203.6 38.565 203.81 38.635 ;
    RECT 203.6 38.925 203.81 38.995 ;
    RECT 203.14 38.205 203.35 38.275 ;
    RECT 203.14 38.565 203.35 38.635 ;
    RECT 203.14 38.925 203.35 38.995 ;
    RECT 336.4 38.205 336.61 38.275 ;
    RECT 336.4 38.565 336.61 38.635 ;
    RECT 336.4 38.925 336.61 38.995 ;
    RECT 335.94 38.205 336.15 38.275 ;
    RECT 335.94 38.565 336.15 38.635 ;
    RECT 335.94 38.925 336.15 38.995 ;
    RECT 266.68 38.205 266.89 38.275 ;
    RECT 266.68 38.565 266.89 38.635 ;
    RECT 266.68 38.925 266.89 38.995 ;
    RECT 266.22 38.205 266.43 38.275 ;
    RECT 266.22 38.565 266.43 38.635 ;
    RECT 266.22 38.925 266.43 38.995 ;
    RECT 263.36 38.205 263.57 38.275 ;
    RECT 263.36 38.565 263.57 38.635 ;
    RECT 263.36 38.925 263.57 38.995 ;
    RECT 262.9 38.205 263.11 38.275 ;
    RECT 262.9 38.565 263.11 38.635 ;
    RECT 262.9 38.925 263.11 38.995 ;
    RECT 260.04 38.205 260.25 38.275 ;
    RECT 260.04 38.565 260.25 38.635 ;
    RECT 260.04 38.925 260.25 38.995 ;
    RECT 259.58 38.205 259.79 38.275 ;
    RECT 259.58 38.565 259.79 38.635 ;
    RECT 259.58 38.925 259.79 38.995 ;
    RECT 256.72 38.205 256.93 38.275 ;
    RECT 256.72 38.565 256.93 38.635 ;
    RECT 256.72 38.925 256.93 38.995 ;
    RECT 256.26 38.205 256.47 38.275 ;
    RECT 256.26 38.565 256.47 38.635 ;
    RECT 256.26 38.925 256.47 38.995 ;
    RECT 253.4 38.205 253.61 38.275 ;
    RECT 253.4 38.565 253.61 38.635 ;
    RECT 253.4 38.925 253.61 38.995 ;
    RECT 252.94 38.205 253.15 38.275 ;
    RECT 252.94 38.565 253.15 38.635 ;
    RECT 252.94 38.925 253.15 38.995 ;
    RECT 250.08 38.205 250.29 38.275 ;
    RECT 250.08 38.565 250.29 38.635 ;
    RECT 250.08 38.925 250.29 38.995 ;
    RECT 249.62 38.205 249.83 38.275 ;
    RECT 249.62 38.565 249.83 38.635 ;
    RECT 249.62 38.925 249.83 38.995 ;
    RECT 246.76 38.205 246.97 38.275 ;
    RECT 246.76 38.565 246.97 38.635 ;
    RECT 246.76 38.925 246.97 38.995 ;
    RECT 246.3 38.205 246.51 38.275 ;
    RECT 246.3 38.565 246.51 38.635 ;
    RECT 246.3 38.925 246.51 38.995 ;
    RECT 243.44 38.205 243.65 38.275 ;
    RECT 243.44 38.565 243.65 38.635 ;
    RECT 243.44 38.925 243.65 38.995 ;
    RECT 242.98 38.205 243.19 38.275 ;
    RECT 242.98 38.565 243.19 38.635 ;
    RECT 242.98 38.925 243.19 38.995 ;
    RECT 240.12 38.205 240.33 38.275 ;
    RECT 240.12 38.565 240.33 38.635 ;
    RECT 240.12 38.925 240.33 38.995 ;
    RECT 239.66 38.205 239.87 38.275 ;
    RECT 239.66 38.565 239.87 38.635 ;
    RECT 239.66 38.925 239.87 38.995 ;
    RECT 236.8 38.205 237.01 38.275 ;
    RECT 236.8 38.565 237.01 38.635 ;
    RECT 236.8 38.925 237.01 38.995 ;
    RECT 236.34 38.205 236.55 38.275 ;
    RECT 236.34 38.565 236.55 38.635 ;
    RECT 236.34 38.925 236.55 38.995 ;
    RECT 374.15 38.565 374.22 38.635 ;
    RECT 333.08 38.205 333.29 38.275 ;
    RECT 333.08 38.565 333.29 38.635 ;
    RECT 333.08 38.925 333.29 38.995 ;
    RECT 332.62 38.205 332.83 38.275 ;
    RECT 332.62 38.565 332.83 38.635 ;
    RECT 332.62 38.925 332.83 38.995 ;
    RECT 329.76 38.205 329.97 38.275 ;
    RECT 329.76 38.565 329.97 38.635 ;
    RECT 329.76 38.925 329.97 38.995 ;
    RECT 329.3 38.205 329.51 38.275 ;
    RECT 329.3 38.565 329.51 38.635 ;
    RECT 329.3 38.925 329.51 38.995 ;
    RECT 326.44 38.205 326.65 38.275 ;
    RECT 326.44 38.565 326.65 38.635 ;
    RECT 326.44 38.925 326.65 38.995 ;
    RECT 325.98 38.205 326.19 38.275 ;
    RECT 325.98 38.565 326.19 38.635 ;
    RECT 325.98 38.925 326.19 38.995 ;
    RECT 323.12 38.205 323.33 38.275 ;
    RECT 323.12 38.565 323.33 38.635 ;
    RECT 323.12 38.925 323.33 38.995 ;
    RECT 322.66 38.205 322.87 38.275 ;
    RECT 322.66 38.565 322.87 38.635 ;
    RECT 322.66 38.925 322.87 38.995 ;
    RECT 319.8 38.205 320.01 38.275 ;
    RECT 319.8 38.565 320.01 38.635 ;
    RECT 319.8 38.925 320.01 38.995 ;
    RECT 319.34 38.205 319.55 38.275 ;
    RECT 319.34 38.565 319.55 38.635 ;
    RECT 319.34 38.925 319.55 38.995 ;
    RECT 316.48 38.205 316.69 38.275 ;
    RECT 316.48 38.565 316.69 38.635 ;
    RECT 316.48 38.925 316.69 38.995 ;
    RECT 316.02 38.205 316.23 38.275 ;
    RECT 316.02 38.565 316.23 38.635 ;
    RECT 316.02 38.925 316.23 38.995 ;
    RECT 313.16 38.205 313.37 38.275 ;
    RECT 313.16 38.565 313.37 38.635 ;
    RECT 313.16 38.925 313.37 38.995 ;
    RECT 312.7 38.205 312.91 38.275 ;
    RECT 312.7 38.565 312.91 38.635 ;
    RECT 312.7 38.925 312.91 38.995 ;
    RECT 309.84 38.205 310.05 38.275 ;
    RECT 309.84 38.565 310.05 38.635 ;
    RECT 309.84 38.925 310.05 38.995 ;
    RECT 309.38 38.205 309.59 38.275 ;
    RECT 309.38 38.565 309.59 38.635 ;
    RECT 309.38 38.925 309.59 38.995 ;
    RECT 306.52 38.205 306.73 38.275 ;
    RECT 306.52 38.565 306.73 38.635 ;
    RECT 306.52 38.925 306.73 38.995 ;
    RECT 306.06 38.205 306.27 38.275 ;
    RECT 306.06 38.565 306.27 38.635 ;
    RECT 306.06 38.925 306.27 38.995 ;
    RECT 303.2 37.485 303.41 37.555 ;
    RECT 303.2 37.845 303.41 37.915 ;
    RECT 303.2 38.205 303.41 38.275 ;
    RECT 302.74 37.485 302.95 37.555 ;
    RECT 302.74 37.845 302.95 37.915 ;
    RECT 302.74 38.205 302.95 38.275 ;
    RECT 372.92 37.485 373.13 37.555 ;
    RECT 372.92 37.845 373.13 37.915 ;
    RECT 372.92 38.205 373.13 38.275 ;
    RECT 372.46 37.485 372.67 37.555 ;
    RECT 372.46 37.845 372.67 37.915 ;
    RECT 372.46 38.205 372.67 38.275 ;
    RECT 369.6 37.485 369.81 37.555 ;
    RECT 369.6 37.845 369.81 37.915 ;
    RECT 369.6 38.205 369.81 38.275 ;
    RECT 369.14 37.485 369.35 37.555 ;
    RECT 369.14 37.845 369.35 37.915 ;
    RECT 369.14 38.205 369.35 38.275 ;
    RECT 200.605 37.845 200.675 37.915 ;
    RECT 299.88 37.485 300.09 37.555 ;
    RECT 299.88 37.845 300.09 37.915 ;
    RECT 299.88 38.205 300.09 38.275 ;
    RECT 299.42 37.485 299.63 37.555 ;
    RECT 299.42 37.845 299.63 37.915 ;
    RECT 299.42 38.205 299.63 38.275 ;
    RECT 296.56 37.485 296.77 37.555 ;
    RECT 296.56 37.845 296.77 37.915 ;
    RECT 296.56 38.205 296.77 38.275 ;
    RECT 296.1 37.485 296.31 37.555 ;
    RECT 296.1 37.845 296.31 37.915 ;
    RECT 296.1 38.205 296.31 38.275 ;
    RECT 293.24 37.485 293.45 37.555 ;
    RECT 293.24 37.845 293.45 37.915 ;
    RECT 293.24 38.205 293.45 38.275 ;
    RECT 292.78 37.485 292.99 37.555 ;
    RECT 292.78 37.845 292.99 37.915 ;
    RECT 292.78 38.205 292.99 38.275 ;
    RECT 289.92 37.485 290.13 37.555 ;
    RECT 289.92 37.845 290.13 37.915 ;
    RECT 289.92 38.205 290.13 38.275 ;
    RECT 289.46 37.485 289.67 37.555 ;
    RECT 289.46 37.845 289.67 37.915 ;
    RECT 289.46 38.205 289.67 38.275 ;
    RECT 286.6 37.485 286.81 37.555 ;
    RECT 286.6 37.845 286.81 37.915 ;
    RECT 286.6 38.205 286.81 38.275 ;
    RECT 286.14 37.485 286.35 37.555 ;
    RECT 286.14 37.845 286.35 37.915 ;
    RECT 286.14 38.205 286.35 38.275 ;
    RECT 283.28 37.485 283.49 37.555 ;
    RECT 283.28 37.845 283.49 37.915 ;
    RECT 283.28 38.205 283.49 38.275 ;
    RECT 282.82 37.485 283.03 37.555 ;
    RECT 282.82 37.845 283.03 37.915 ;
    RECT 282.82 38.205 283.03 38.275 ;
    RECT 279.96 37.485 280.17 37.555 ;
    RECT 279.96 37.845 280.17 37.915 ;
    RECT 279.96 38.205 280.17 38.275 ;
    RECT 279.5 37.485 279.71 37.555 ;
    RECT 279.5 37.845 279.71 37.915 ;
    RECT 279.5 38.205 279.71 38.275 ;
    RECT 276.64 37.485 276.85 37.555 ;
    RECT 276.64 37.845 276.85 37.915 ;
    RECT 276.64 38.205 276.85 38.275 ;
    RECT 276.18 37.485 276.39 37.555 ;
    RECT 276.18 37.845 276.39 37.915 ;
    RECT 276.18 38.205 276.39 38.275 ;
    RECT 273.32 37.485 273.53 37.555 ;
    RECT 273.32 37.845 273.53 37.915 ;
    RECT 273.32 38.205 273.53 38.275 ;
    RECT 272.86 37.485 273.07 37.555 ;
    RECT 272.86 37.845 273.07 37.915 ;
    RECT 272.86 38.205 273.07 38.275 ;
    RECT 270.0 37.485 270.21 37.555 ;
    RECT 270.0 37.845 270.21 37.915 ;
    RECT 270.0 38.205 270.21 38.275 ;
    RECT 269.54 37.485 269.75 37.555 ;
    RECT 269.54 37.845 269.75 37.915 ;
    RECT 269.54 38.205 269.75 38.275 ;
    RECT 233.48 37.485 233.69 37.555 ;
    RECT 233.48 37.845 233.69 37.915 ;
    RECT 233.48 38.205 233.69 38.275 ;
    RECT 233.02 37.485 233.23 37.555 ;
    RECT 233.02 37.845 233.23 37.915 ;
    RECT 233.02 38.205 233.23 38.275 ;
    RECT 230.16 37.485 230.37 37.555 ;
    RECT 230.16 37.845 230.37 37.915 ;
    RECT 230.16 38.205 230.37 38.275 ;
    RECT 229.7 37.485 229.91 37.555 ;
    RECT 229.7 37.845 229.91 37.915 ;
    RECT 229.7 38.205 229.91 38.275 ;
    RECT 366.28 37.485 366.49 37.555 ;
    RECT 366.28 37.845 366.49 37.915 ;
    RECT 366.28 38.205 366.49 38.275 ;
    RECT 365.82 37.485 366.03 37.555 ;
    RECT 365.82 37.845 366.03 37.915 ;
    RECT 365.82 38.205 366.03 38.275 ;
    RECT 226.84 37.485 227.05 37.555 ;
    RECT 226.84 37.845 227.05 37.915 ;
    RECT 226.84 38.205 227.05 38.275 ;
    RECT 226.38 37.485 226.59 37.555 ;
    RECT 226.38 37.845 226.59 37.915 ;
    RECT 226.38 38.205 226.59 38.275 ;
    RECT 362.96 37.485 363.17 37.555 ;
    RECT 362.96 37.845 363.17 37.915 ;
    RECT 362.96 38.205 363.17 38.275 ;
    RECT 362.5 37.485 362.71 37.555 ;
    RECT 362.5 37.845 362.71 37.915 ;
    RECT 362.5 38.205 362.71 38.275 ;
    RECT 223.52 37.485 223.73 37.555 ;
    RECT 223.52 37.845 223.73 37.915 ;
    RECT 223.52 38.205 223.73 38.275 ;
    RECT 223.06 37.485 223.27 37.555 ;
    RECT 223.06 37.845 223.27 37.915 ;
    RECT 223.06 38.205 223.27 38.275 ;
    RECT 359.64 37.485 359.85 37.555 ;
    RECT 359.64 37.845 359.85 37.915 ;
    RECT 359.64 38.205 359.85 38.275 ;
    RECT 359.18 37.485 359.39 37.555 ;
    RECT 359.18 37.845 359.39 37.915 ;
    RECT 359.18 38.205 359.39 38.275 ;
    RECT 220.2 37.485 220.41 37.555 ;
    RECT 220.2 37.845 220.41 37.915 ;
    RECT 220.2 38.205 220.41 38.275 ;
    RECT 219.74 37.485 219.95 37.555 ;
    RECT 219.74 37.845 219.95 37.915 ;
    RECT 219.74 38.205 219.95 38.275 ;
    RECT 356.32 37.485 356.53 37.555 ;
    RECT 356.32 37.845 356.53 37.915 ;
    RECT 356.32 38.205 356.53 38.275 ;
    RECT 355.86 37.485 356.07 37.555 ;
    RECT 355.86 37.845 356.07 37.915 ;
    RECT 355.86 38.205 356.07 38.275 ;
    RECT 353.0 37.485 353.21 37.555 ;
    RECT 353.0 37.845 353.21 37.915 ;
    RECT 353.0 38.205 353.21 38.275 ;
    RECT 352.54 37.485 352.75 37.555 ;
    RECT 352.54 37.845 352.75 37.915 ;
    RECT 352.54 38.205 352.75 38.275 ;
    RECT 216.88 37.485 217.09 37.555 ;
    RECT 216.88 37.845 217.09 37.915 ;
    RECT 216.88 38.205 217.09 38.275 ;
    RECT 216.42 37.485 216.63 37.555 ;
    RECT 216.42 37.845 216.63 37.915 ;
    RECT 216.42 38.205 216.63 38.275 ;
    RECT 349.68 37.485 349.89 37.555 ;
    RECT 349.68 37.845 349.89 37.915 ;
    RECT 349.68 38.205 349.89 38.275 ;
    RECT 349.22 37.485 349.43 37.555 ;
    RECT 349.22 37.845 349.43 37.915 ;
    RECT 349.22 38.205 349.43 38.275 ;
    RECT 213.56 37.485 213.77 37.555 ;
    RECT 213.56 37.845 213.77 37.915 ;
    RECT 213.56 38.205 213.77 38.275 ;
    RECT 213.1 37.485 213.31 37.555 ;
    RECT 213.1 37.845 213.31 37.915 ;
    RECT 213.1 38.205 213.31 38.275 ;
    RECT 346.36 37.485 346.57 37.555 ;
    RECT 346.36 37.845 346.57 37.915 ;
    RECT 346.36 38.205 346.57 38.275 ;
    RECT 345.9 37.485 346.11 37.555 ;
    RECT 345.9 37.845 346.11 37.915 ;
    RECT 345.9 38.205 346.11 38.275 ;
    RECT 210.24 37.485 210.45 37.555 ;
    RECT 210.24 37.845 210.45 37.915 ;
    RECT 210.24 38.205 210.45 38.275 ;
    RECT 209.78 37.485 209.99 37.555 ;
    RECT 209.78 37.845 209.99 37.915 ;
    RECT 209.78 38.205 209.99 38.275 ;
    RECT 343.04 37.485 343.25 37.555 ;
    RECT 343.04 37.845 343.25 37.915 ;
    RECT 343.04 38.205 343.25 38.275 ;
    RECT 342.58 37.485 342.79 37.555 ;
    RECT 342.58 37.845 342.79 37.915 ;
    RECT 342.58 38.205 342.79 38.275 ;
    RECT 206.92 37.485 207.13 37.555 ;
    RECT 206.92 37.845 207.13 37.915 ;
    RECT 206.92 38.205 207.13 38.275 ;
    RECT 206.46 37.485 206.67 37.555 ;
    RECT 206.46 37.845 206.67 37.915 ;
    RECT 206.46 38.205 206.67 38.275 ;
    RECT 339.72 37.485 339.93 37.555 ;
    RECT 339.72 37.845 339.93 37.915 ;
    RECT 339.72 38.205 339.93 38.275 ;
    RECT 339.26 37.485 339.47 37.555 ;
    RECT 339.26 37.845 339.47 37.915 ;
    RECT 339.26 38.205 339.47 38.275 ;
    RECT 203.6 37.485 203.81 37.555 ;
    RECT 203.6 37.845 203.81 37.915 ;
    RECT 203.6 38.205 203.81 38.275 ;
    RECT 203.14 37.485 203.35 37.555 ;
    RECT 203.14 37.845 203.35 37.915 ;
    RECT 203.14 38.205 203.35 38.275 ;
    RECT 336.4 37.485 336.61 37.555 ;
    RECT 336.4 37.845 336.61 37.915 ;
    RECT 336.4 38.205 336.61 38.275 ;
    RECT 335.94 37.485 336.15 37.555 ;
    RECT 335.94 37.845 336.15 37.915 ;
    RECT 335.94 38.205 336.15 38.275 ;
    RECT 266.68 37.485 266.89 37.555 ;
    RECT 266.68 37.845 266.89 37.915 ;
    RECT 266.68 38.205 266.89 38.275 ;
    RECT 266.22 37.485 266.43 37.555 ;
    RECT 266.22 37.845 266.43 37.915 ;
    RECT 266.22 38.205 266.43 38.275 ;
    RECT 263.36 37.485 263.57 37.555 ;
    RECT 263.36 37.845 263.57 37.915 ;
    RECT 263.36 38.205 263.57 38.275 ;
    RECT 262.9 37.485 263.11 37.555 ;
    RECT 262.9 37.845 263.11 37.915 ;
    RECT 262.9 38.205 263.11 38.275 ;
    RECT 260.04 37.485 260.25 37.555 ;
    RECT 260.04 37.845 260.25 37.915 ;
    RECT 260.04 38.205 260.25 38.275 ;
    RECT 259.58 37.485 259.79 37.555 ;
    RECT 259.58 37.845 259.79 37.915 ;
    RECT 259.58 38.205 259.79 38.275 ;
    RECT 256.72 37.485 256.93 37.555 ;
    RECT 256.72 37.845 256.93 37.915 ;
    RECT 256.72 38.205 256.93 38.275 ;
    RECT 256.26 37.485 256.47 37.555 ;
    RECT 256.26 37.845 256.47 37.915 ;
    RECT 256.26 38.205 256.47 38.275 ;
    RECT 253.4 37.485 253.61 37.555 ;
    RECT 253.4 37.845 253.61 37.915 ;
    RECT 253.4 38.205 253.61 38.275 ;
    RECT 252.94 37.485 253.15 37.555 ;
    RECT 252.94 37.845 253.15 37.915 ;
    RECT 252.94 38.205 253.15 38.275 ;
    RECT 250.08 37.485 250.29 37.555 ;
    RECT 250.08 37.845 250.29 37.915 ;
    RECT 250.08 38.205 250.29 38.275 ;
    RECT 249.62 37.485 249.83 37.555 ;
    RECT 249.62 37.845 249.83 37.915 ;
    RECT 249.62 38.205 249.83 38.275 ;
    RECT 246.76 37.485 246.97 37.555 ;
    RECT 246.76 37.845 246.97 37.915 ;
    RECT 246.76 38.205 246.97 38.275 ;
    RECT 246.3 37.485 246.51 37.555 ;
    RECT 246.3 37.845 246.51 37.915 ;
    RECT 246.3 38.205 246.51 38.275 ;
    RECT 243.44 37.485 243.65 37.555 ;
    RECT 243.44 37.845 243.65 37.915 ;
    RECT 243.44 38.205 243.65 38.275 ;
    RECT 242.98 37.485 243.19 37.555 ;
    RECT 242.98 37.845 243.19 37.915 ;
    RECT 242.98 38.205 243.19 38.275 ;
    RECT 240.12 37.485 240.33 37.555 ;
    RECT 240.12 37.845 240.33 37.915 ;
    RECT 240.12 38.205 240.33 38.275 ;
    RECT 239.66 37.485 239.87 37.555 ;
    RECT 239.66 37.845 239.87 37.915 ;
    RECT 239.66 38.205 239.87 38.275 ;
    RECT 236.8 37.485 237.01 37.555 ;
    RECT 236.8 37.845 237.01 37.915 ;
    RECT 236.8 38.205 237.01 38.275 ;
    RECT 236.34 37.485 236.55 37.555 ;
    RECT 236.34 37.845 236.55 37.915 ;
    RECT 236.34 38.205 236.55 38.275 ;
    RECT 374.15 37.845 374.22 37.915 ;
    RECT 333.08 37.485 333.29 37.555 ;
    RECT 333.08 37.845 333.29 37.915 ;
    RECT 333.08 38.205 333.29 38.275 ;
    RECT 332.62 37.485 332.83 37.555 ;
    RECT 332.62 37.845 332.83 37.915 ;
    RECT 332.62 38.205 332.83 38.275 ;
    RECT 329.76 37.485 329.97 37.555 ;
    RECT 329.76 37.845 329.97 37.915 ;
    RECT 329.76 38.205 329.97 38.275 ;
    RECT 329.3 37.485 329.51 37.555 ;
    RECT 329.3 37.845 329.51 37.915 ;
    RECT 329.3 38.205 329.51 38.275 ;
    RECT 326.44 37.485 326.65 37.555 ;
    RECT 326.44 37.845 326.65 37.915 ;
    RECT 326.44 38.205 326.65 38.275 ;
    RECT 325.98 37.485 326.19 37.555 ;
    RECT 325.98 37.845 326.19 37.915 ;
    RECT 325.98 38.205 326.19 38.275 ;
    RECT 323.12 37.485 323.33 37.555 ;
    RECT 323.12 37.845 323.33 37.915 ;
    RECT 323.12 38.205 323.33 38.275 ;
    RECT 322.66 37.485 322.87 37.555 ;
    RECT 322.66 37.845 322.87 37.915 ;
    RECT 322.66 38.205 322.87 38.275 ;
    RECT 319.8 37.485 320.01 37.555 ;
    RECT 319.8 37.845 320.01 37.915 ;
    RECT 319.8 38.205 320.01 38.275 ;
    RECT 319.34 37.485 319.55 37.555 ;
    RECT 319.34 37.845 319.55 37.915 ;
    RECT 319.34 38.205 319.55 38.275 ;
    RECT 316.48 37.485 316.69 37.555 ;
    RECT 316.48 37.845 316.69 37.915 ;
    RECT 316.48 38.205 316.69 38.275 ;
    RECT 316.02 37.485 316.23 37.555 ;
    RECT 316.02 37.845 316.23 37.915 ;
    RECT 316.02 38.205 316.23 38.275 ;
    RECT 313.16 37.485 313.37 37.555 ;
    RECT 313.16 37.845 313.37 37.915 ;
    RECT 313.16 38.205 313.37 38.275 ;
    RECT 312.7 37.485 312.91 37.555 ;
    RECT 312.7 37.845 312.91 37.915 ;
    RECT 312.7 38.205 312.91 38.275 ;
    RECT 309.84 37.485 310.05 37.555 ;
    RECT 309.84 37.845 310.05 37.915 ;
    RECT 309.84 38.205 310.05 38.275 ;
    RECT 309.38 37.485 309.59 37.555 ;
    RECT 309.38 37.845 309.59 37.915 ;
    RECT 309.38 38.205 309.59 38.275 ;
    RECT 306.52 37.485 306.73 37.555 ;
    RECT 306.52 37.845 306.73 37.915 ;
    RECT 306.52 38.205 306.73 38.275 ;
    RECT 306.06 37.485 306.27 37.555 ;
    RECT 306.06 37.845 306.27 37.915 ;
    RECT 306.06 38.205 306.27 38.275 ;
    RECT 303.2 36.765 303.41 36.835 ;
    RECT 303.2 37.125 303.41 37.195 ;
    RECT 303.2 37.485 303.41 37.555 ;
    RECT 302.74 36.765 302.95 36.835 ;
    RECT 302.74 37.125 302.95 37.195 ;
    RECT 302.74 37.485 302.95 37.555 ;
    RECT 372.92 36.765 373.13 36.835 ;
    RECT 372.92 37.125 373.13 37.195 ;
    RECT 372.92 37.485 373.13 37.555 ;
    RECT 372.46 36.765 372.67 36.835 ;
    RECT 372.46 37.125 372.67 37.195 ;
    RECT 372.46 37.485 372.67 37.555 ;
    RECT 369.6 36.765 369.81 36.835 ;
    RECT 369.6 37.125 369.81 37.195 ;
    RECT 369.6 37.485 369.81 37.555 ;
    RECT 369.14 36.765 369.35 36.835 ;
    RECT 369.14 37.125 369.35 37.195 ;
    RECT 369.14 37.485 369.35 37.555 ;
    RECT 200.605 37.125 200.675 37.195 ;
    RECT 299.88 36.765 300.09 36.835 ;
    RECT 299.88 37.125 300.09 37.195 ;
    RECT 299.88 37.485 300.09 37.555 ;
    RECT 299.42 36.765 299.63 36.835 ;
    RECT 299.42 37.125 299.63 37.195 ;
    RECT 299.42 37.485 299.63 37.555 ;
    RECT 296.56 36.765 296.77 36.835 ;
    RECT 296.56 37.125 296.77 37.195 ;
    RECT 296.56 37.485 296.77 37.555 ;
    RECT 296.1 36.765 296.31 36.835 ;
    RECT 296.1 37.125 296.31 37.195 ;
    RECT 296.1 37.485 296.31 37.555 ;
    RECT 293.24 36.765 293.45 36.835 ;
    RECT 293.24 37.125 293.45 37.195 ;
    RECT 293.24 37.485 293.45 37.555 ;
    RECT 292.78 36.765 292.99 36.835 ;
    RECT 292.78 37.125 292.99 37.195 ;
    RECT 292.78 37.485 292.99 37.555 ;
    RECT 289.92 36.765 290.13 36.835 ;
    RECT 289.92 37.125 290.13 37.195 ;
    RECT 289.92 37.485 290.13 37.555 ;
    RECT 289.46 36.765 289.67 36.835 ;
    RECT 289.46 37.125 289.67 37.195 ;
    RECT 289.46 37.485 289.67 37.555 ;
    RECT 286.6 36.765 286.81 36.835 ;
    RECT 286.6 37.125 286.81 37.195 ;
    RECT 286.6 37.485 286.81 37.555 ;
    RECT 286.14 36.765 286.35 36.835 ;
    RECT 286.14 37.125 286.35 37.195 ;
    RECT 286.14 37.485 286.35 37.555 ;
    RECT 283.28 36.765 283.49 36.835 ;
    RECT 283.28 37.125 283.49 37.195 ;
    RECT 283.28 37.485 283.49 37.555 ;
    RECT 282.82 36.765 283.03 36.835 ;
    RECT 282.82 37.125 283.03 37.195 ;
    RECT 282.82 37.485 283.03 37.555 ;
    RECT 279.96 36.765 280.17 36.835 ;
    RECT 279.96 37.125 280.17 37.195 ;
    RECT 279.96 37.485 280.17 37.555 ;
    RECT 279.5 36.765 279.71 36.835 ;
    RECT 279.5 37.125 279.71 37.195 ;
    RECT 279.5 37.485 279.71 37.555 ;
    RECT 276.64 36.765 276.85 36.835 ;
    RECT 276.64 37.125 276.85 37.195 ;
    RECT 276.64 37.485 276.85 37.555 ;
    RECT 276.18 36.765 276.39 36.835 ;
    RECT 276.18 37.125 276.39 37.195 ;
    RECT 276.18 37.485 276.39 37.555 ;
    RECT 273.32 36.765 273.53 36.835 ;
    RECT 273.32 37.125 273.53 37.195 ;
    RECT 273.32 37.485 273.53 37.555 ;
    RECT 272.86 36.765 273.07 36.835 ;
    RECT 272.86 37.125 273.07 37.195 ;
    RECT 272.86 37.485 273.07 37.555 ;
    RECT 270.0 36.765 270.21 36.835 ;
    RECT 270.0 37.125 270.21 37.195 ;
    RECT 270.0 37.485 270.21 37.555 ;
    RECT 269.54 36.765 269.75 36.835 ;
    RECT 269.54 37.125 269.75 37.195 ;
    RECT 269.54 37.485 269.75 37.555 ;
    RECT 233.48 36.765 233.69 36.835 ;
    RECT 233.48 37.125 233.69 37.195 ;
    RECT 233.48 37.485 233.69 37.555 ;
    RECT 233.02 36.765 233.23 36.835 ;
    RECT 233.02 37.125 233.23 37.195 ;
    RECT 233.02 37.485 233.23 37.555 ;
    RECT 230.16 36.765 230.37 36.835 ;
    RECT 230.16 37.125 230.37 37.195 ;
    RECT 230.16 37.485 230.37 37.555 ;
    RECT 229.7 36.765 229.91 36.835 ;
    RECT 229.7 37.125 229.91 37.195 ;
    RECT 229.7 37.485 229.91 37.555 ;
    RECT 366.28 36.765 366.49 36.835 ;
    RECT 366.28 37.125 366.49 37.195 ;
    RECT 366.28 37.485 366.49 37.555 ;
    RECT 365.82 36.765 366.03 36.835 ;
    RECT 365.82 37.125 366.03 37.195 ;
    RECT 365.82 37.485 366.03 37.555 ;
    RECT 226.84 36.765 227.05 36.835 ;
    RECT 226.84 37.125 227.05 37.195 ;
    RECT 226.84 37.485 227.05 37.555 ;
    RECT 226.38 36.765 226.59 36.835 ;
    RECT 226.38 37.125 226.59 37.195 ;
    RECT 226.38 37.485 226.59 37.555 ;
    RECT 362.96 36.765 363.17 36.835 ;
    RECT 362.96 37.125 363.17 37.195 ;
    RECT 362.96 37.485 363.17 37.555 ;
    RECT 362.5 36.765 362.71 36.835 ;
    RECT 362.5 37.125 362.71 37.195 ;
    RECT 362.5 37.485 362.71 37.555 ;
    RECT 223.52 36.765 223.73 36.835 ;
    RECT 223.52 37.125 223.73 37.195 ;
    RECT 223.52 37.485 223.73 37.555 ;
    RECT 223.06 36.765 223.27 36.835 ;
    RECT 223.06 37.125 223.27 37.195 ;
    RECT 223.06 37.485 223.27 37.555 ;
    RECT 359.64 36.765 359.85 36.835 ;
    RECT 359.64 37.125 359.85 37.195 ;
    RECT 359.64 37.485 359.85 37.555 ;
    RECT 359.18 36.765 359.39 36.835 ;
    RECT 359.18 37.125 359.39 37.195 ;
    RECT 359.18 37.485 359.39 37.555 ;
    RECT 220.2 36.765 220.41 36.835 ;
    RECT 220.2 37.125 220.41 37.195 ;
    RECT 220.2 37.485 220.41 37.555 ;
    RECT 219.74 36.765 219.95 36.835 ;
    RECT 219.74 37.125 219.95 37.195 ;
    RECT 219.74 37.485 219.95 37.555 ;
    RECT 356.32 36.765 356.53 36.835 ;
    RECT 356.32 37.125 356.53 37.195 ;
    RECT 356.32 37.485 356.53 37.555 ;
    RECT 355.86 36.765 356.07 36.835 ;
    RECT 355.86 37.125 356.07 37.195 ;
    RECT 355.86 37.485 356.07 37.555 ;
    RECT 353.0 36.765 353.21 36.835 ;
    RECT 353.0 37.125 353.21 37.195 ;
    RECT 353.0 37.485 353.21 37.555 ;
    RECT 352.54 36.765 352.75 36.835 ;
    RECT 352.54 37.125 352.75 37.195 ;
    RECT 352.54 37.485 352.75 37.555 ;
    RECT 216.88 36.765 217.09 36.835 ;
    RECT 216.88 37.125 217.09 37.195 ;
    RECT 216.88 37.485 217.09 37.555 ;
    RECT 216.42 36.765 216.63 36.835 ;
    RECT 216.42 37.125 216.63 37.195 ;
    RECT 216.42 37.485 216.63 37.555 ;
    RECT 349.68 36.765 349.89 36.835 ;
    RECT 349.68 37.125 349.89 37.195 ;
    RECT 349.68 37.485 349.89 37.555 ;
    RECT 349.22 36.765 349.43 36.835 ;
    RECT 349.22 37.125 349.43 37.195 ;
    RECT 349.22 37.485 349.43 37.555 ;
    RECT 213.56 36.765 213.77 36.835 ;
    RECT 213.56 37.125 213.77 37.195 ;
    RECT 213.56 37.485 213.77 37.555 ;
    RECT 213.1 36.765 213.31 36.835 ;
    RECT 213.1 37.125 213.31 37.195 ;
    RECT 213.1 37.485 213.31 37.555 ;
    RECT 346.36 36.765 346.57 36.835 ;
    RECT 346.36 37.125 346.57 37.195 ;
    RECT 346.36 37.485 346.57 37.555 ;
    RECT 345.9 36.765 346.11 36.835 ;
    RECT 345.9 37.125 346.11 37.195 ;
    RECT 345.9 37.485 346.11 37.555 ;
    RECT 210.24 36.765 210.45 36.835 ;
    RECT 210.24 37.125 210.45 37.195 ;
    RECT 210.24 37.485 210.45 37.555 ;
    RECT 209.78 36.765 209.99 36.835 ;
    RECT 209.78 37.125 209.99 37.195 ;
    RECT 209.78 37.485 209.99 37.555 ;
    RECT 343.04 36.765 343.25 36.835 ;
    RECT 343.04 37.125 343.25 37.195 ;
    RECT 343.04 37.485 343.25 37.555 ;
    RECT 342.58 36.765 342.79 36.835 ;
    RECT 342.58 37.125 342.79 37.195 ;
    RECT 342.58 37.485 342.79 37.555 ;
    RECT 206.92 36.765 207.13 36.835 ;
    RECT 206.92 37.125 207.13 37.195 ;
    RECT 206.92 37.485 207.13 37.555 ;
    RECT 206.46 36.765 206.67 36.835 ;
    RECT 206.46 37.125 206.67 37.195 ;
    RECT 206.46 37.485 206.67 37.555 ;
    RECT 339.72 36.765 339.93 36.835 ;
    RECT 339.72 37.125 339.93 37.195 ;
    RECT 339.72 37.485 339.93 37.555 ;
    RECT 339.26 36.765 339.47 36.835 ;
    RECT 339.26 37.125 339.47 37.195 ;
    RECT 339.26 37.485 339.47 37.555 ;
    RECT 203.6 36.765 203.81 36.835 ;
    RECT 203.6 37.125 203.81 37.195 ;
    RECT 203.6 37.485 203.81 37.555 ;
    RECT 203.14 36.765 203.35 36.835 ;
    RECT 203.14 37.125 203.35 37.195 ;
    RECT 203.14 37.485 203.35 37.555 ;
    RECT 336.4 36.765 336.61 36.835 ;
    RECT 336.4 37.125 336.61 37.195 ;
    RECT 336.4 37.485 336.61 37.555 ;
    RECT 335.94 36.765 336.15 36.835 ;
    RECT 335.94 37.125 336.15 37.195 ;
    RECT 335.94 37.485 336.15 37.555 ;
    RECT 266.68 36.765 266.89 36.835 ;
    RECT 266.68 37.125 266.89 37.195 ;
    RECT 266.68 37.485 266.89 37.555 ;
    RECT 266.22 36.765 266.43 36.835 ;
    RECT 266.22 37.125 266.43 37.195 ;
    RECT 266.22 37.485 266.43 37.555 ;
    RECT 263.36 36.765 263.57 36.835 ;
    RECT 263.36 37.125 263.57 37.195 ;
    RECT 263.36 37.485 263.57 37.555 ;
    RECT 262.9 36.765 263.11 36.835 ;
    RECT 262.9 37.125 263.11 37.195 ;
    RECT 262.9 37.485 263.11 37.555 ;
    RECT 260.04 36.765 260.25 36.835 ;
    RECT 260.04 37.125 260.25 37.195 ;
    RECT 260.04 37.485 260.25 37.555 ;
    RECT 259.58 36.765 259.79 36.835 ;
    RECT 259.58 37.125 259.79 37.195 ;
    RECT 259.58 37.485 259.79 37.555 ;
    RECT 256.72 36.765 256.93 36.835 ;
    RECT 256.72 37.125 256.93 37.195 ;
    RECT 256.72 37.485 256.93 37.555 ;
    RECT 256.26 36.765 256.47 36.835 ;
    RECT 256.26 37.125 256.47 37.195 ;
    RECT 256.26 37.485 256.47 37.555 ;
    RECT 253.4 36.765 253.61 36.835 ;
    RECT 253.4 37.125 253.61 37.195 ;
    RECT 253.4 37.485 253.61 37.555 ;
    RECT 252.94 36.765 253.15 36.835 ;
    RECT 252.94 37.125 253.15 37.195 ;
    RECT 252.94 37.485 253.15 37.555 ;
    RECT 250.08 36.765 250.29 36.835 ;
    RECT 250.08 37.125 250.29 37.195 ;
    RECT 250.08 37.485 250.29 37.555 ;
    RECT 249.62 36.765 249.83 36.835 ;
    RECT 249.62 37.125 249.83 37.195 ;
    RECT 249.62 37.485 249.83 37.555 ;
    RECT 246.76 36.765 246.97 36.835 ;
    RECT 246.76 37.125 246.97 37.195 ;
    RECT 246.76 37.485 246.97 37.555 ;
    RECT 246.3 36.765 246.51 36.835 ;
    RECT 246.3 37.125 246.51 37.195 ;
    RECT 246.3 37.485 246.51 37.555 ;
    RECT 243.44 36.765 243.65 36.835 ;
    RECT 243.44 37.125 243.65 37.195 ;
    RECT 243.44 37.485 243.65 37.555 ;
    RECT 242.98 36.765 243.19 36.835 ;
    RECT 242.98 37.125 243.19 37.195 ;
    RECT 242.98 37.485 243.19 37.555 ;
    RECT 240.12 36.765 240.33 36.835 ;
    RECT 240.12 37.125 240.33 37.195 ;
    RECT 240.12 37.485 240.33 37.555 ;
    RECT 239.66 36.765 239.87 36.835 ;
    RECT 239.66 37.125 239.87 37.195 ;
    RECT 239.66 37.485 239.87 37.555 ;
    RECT 236.8 36.765 237.01 36.835 ;
    RECT 236.8 37.125 237.01 37.195 ;
    RECT 236.8 37.485 237.01 37.555 ;
    RECT 236.34 36.765 236.55 36.835 ;
    RECT 236.34 37.125 236.55 37.195 ;
    RECT 236.34 37.485 236.55 37.555 ;
    RECT 374.15 37.125 374.22 37.195 ;
    RECT 333.08 36.765 333.29 36.835 ;
    RECT 333.08 37.125 333.29 37.195 ;
    RECT 333.08 37.485 333.29 37.555 ;
    RECT 332.62 36.765 332.83 36.835 ;
    RECT 332.62 37.125 332.83 37.195 ;
    RECT 332.62 37.485 332.83 37.555 ;
    RECT 329.76 36.765 329.97 36.835 ;
    RECT 329.76 37.125 329.97 37.195 ;
    RECT 329.76 37.485 329.97 37.555 ;
    RECT 329.3 36.765 329.51 36.835 ;
    RECT 329.3 37.125 329.51 37.195 ;
    RECT 329.3 37.485 329.51 37.555 ;
    RECT 326.44 36.765 326.65 36.835 ;
    RECT 326.44 37.125 326.65 37.195 ;
    RECT 326.44 37.485 326.65 37.555 ;
    RECT 325.98 36.765 326.19 36.835 ;
    RECT 325.98 37.125 326.19 37.195 ;
    RECT 325.98 37.485 326.19 37.555 ;
    RECT 323.12 36.765 323.33 36.835 ;
    RECT 323.12 37.125 323.33 37.195 ;
    RECT 323.12 37.485 323.33 37.555 ;
    RECT 322.66 36.765 322.87 36.835 ;
    RECT 322.66 37.125 322.87 37.195 ;
    RECT 322.66 37.485 322.87 37.555 ;
    RECT 319.8 36.765 320.01 36.835 ;
    RECT 319.8 37.125 320.01 37.195 ;
    RECT 319.8 37.485 320.01 37.555 ;
    RECT 319.34 36.765 319.55 36.835 ;
    RECT 319.34 37.125 319.55 37.195 ;
    RECT 319.34 37.485 319.55 37.555 ;
    RECT 316.48 36.765 316.69 36.835 ;
    RECT 316.48 37.125 316.69 37.195 ;
    RECT 316.48 37.485 316.69 37.555 ;
    RECT 316.02 36.765 316.23 36.835 ;
    RECT 316.02 37.125 316.23 37.195 ;
    RECT 316.02 37.485 316.23 37.555 ;
    RECT 313.16 36.765 313.37 36.835 ;
    RECT 313.16 37.125 313.37 37.195 ;
    RECT 313.16 37.485 313.37 37.555 ;
    RECT 312.7 36.765 312.91 36.835 ;
    RECT 312.7 37.125 312.91 37.195 ;
    RECT 312.7 37.485 312.91 37.555 ;
    RECT 309.84 36.765 310.05 36.835 ;
    RECT 309.84 37.125 310.05 37.195 ;
    RECT 309.84 37.485 310.05 37.555 ;
    RECT 309.38 36.765 309.59 36.835 ;
    RECT 309.38 37.125 309.59 37.195 ;
    RECT 309.38 37.485 309.59 37.555 ;
    RECT 306.52 36.765 306.73 36.835 ;
    RECT 306.52 37.125 306.73 37.195 ;
    RECT 306.52 37.485 306.73 37.555 ;
    RECT 306.06 36.765 306.27 36.835 ;
    RECT 306.06 37.125 306.27 37.195 ;
    RECT 306.06 37.485 306.27 37.555 ;
    RECT 303.2 36.045 303.41 36.115 ;
    RECT 303.2 36.405 303.41 36.475 ;
    RECT 303.2 36.765 303.41 36.835 ;
    RECT 302.74 36.045 302.95 36.115 ;
    RECT 302.74 36.405 302.95 36.475 ;
    RECT 302.74 36.765 302.95 36.835 ;
    RECT 372.92 36.045 373.13 36.115 ;
    RECT 372.92 36.405 373.13 36.475 ;
    RECT 372.92 36.765 373.13 36.835 ;
    RECT 372.46 36.045 372.67 36.115 ;
    RECT 372.46 36.405 372.67 36.475 ;
    RECT 372.46 36.765 372.67 36.835 ;
    RECT 369.6 36.045 369.81 36.115 ;
    RECT 369.6 36.405 369.81 36.475 ;
    RECT 369.6 36.765 369.81 36.835 ;
    RECT 369.14 36.045 369.35 36.115 ;
    RECT 369.14 36.405 369.35 36.475 ;
    RECT 369.14 36.765 369.35 36.835 ;
    RECT 200.605 36.405 200.675 36.475 ;
    RECT 299.88 36.045 300.09 36.115 ;
    RECT 299.88 36.405 300.09 36.475 ;
    RECT 299.88 36.765 300.09 36.835 ;
    RECT 299.42 36.045 299.63 36.115 ;
    RECT 299.42 36.405 299.63 36.475 ;
    RECT 299.42 36.765 299.63 36.835 ;
    RECT 296.56 36.045 296.77 36.115 ;
    RECT 296.56 36.405 296.77 36.475 ;
    RECT 296.56 36.765 296.77 36.835 ;
    RECT 296.1 36.045 296.31 36.115 ;
    RECT 296.1 36.405 296.31 36.475 ;
    RECT 296.1 36.765 296.31 36.835 ;
    RECT 293.24 36.045 293.45 36.115 ;
    RECT 293.24 36.405 293.45 36.475 ;
    RECT 293.24 36.765 293.45 36.835 ;
    RECT 292.78 36.045 292.99 36.115 ;
    RECT 292.78 36.405 292.99 36.475 ;
    RECT 292.78 36.765 292.99 36.835 ;
    RECT 289.92 36.045 290.13 36.115 ;
    RECT 289.92 36.405 290.13 36.475 ;
    RECT 289.92 36.765 290.13 36.835 ;
    RECT 289.46 36.045 289.67 36.115 ;
    RECT 289.46 36.405 289.67 36.475 ;
    RECT 289.46 36.765 289.67 36.835 ;
    RECT 286.6 36.045 286.81 36.115 ;
    RECT 286.6 36.405 286.81 36.475 ;
    RECT 286.6 36.765 286.81 36.835 ;
    RECT 286.14 36.045 286.35 36.115 ;
    RECT 286.14 36.405 286.35 36.475 ;
    RECT 286.14 36.765 286.35 36.835 ;
    RECT 283.28 36.045 283.49 36.115 ;
    RECT 283.28 36.405 283.49 36.475 ;
    RECT 283.28 36.765 283.49 36.835 ;
    RECT 282.82 36.045 283.03 36.115 ;
    RECT 282.82 36.405 283.03 36.475 ;
    RECT 282.82 36.765 283.03 36.835 ;
    RECT 279.96 36.045 280.17 36.115 ;
    RECT 279.96 36.405 280.17 36.475 ;
    RECT 279.96 36.765 280.17 36.835 ;
    RECT 279.5 36.045 279.71 36.115 ;
    RECT 279.5 36.405 279.71 36.475 ;
    RECT 279.5 36.765 279.71 36.835 ;
    RECT 276.64 36.045 276.85 36.115 ;
    RECT 276.64 36.405 276.85 36.475 ;
    RECT 276.64 36.765 276.85 36.835 ;
    RECT 276.18 36.045 276.39 36.115 ;
    RECT 276.18 36.405 276.39 36.475 ;
    RECT 276.18 36.765 276.39 36.835 ;
    RECT 273.32 36.045 273.53 36.115 ;
    RECT 273.32 36.405 273.53 36.475 ;
    RECT 273.32 36.765 273.53 36.835 ;
    RECT 272.86 36.045 273.07 36.115 ;
    RECT 272.86 36.405 273.07 36.475 ;
    RECT 272.86 36.765 273.07 36.835 ;
    RECT 270.0 36.045 270.21 36.115 ;
    RECT 270.0 36.405 270.21 36.475 ;
    RECT 270.0 36.765 270.21 36.835 ;
    RECT 269.54 36.045 269.75 36.115 ;
    RECT 269.54 36.405 269.75 36.475 ;
    RECT 269.54 36.765 269.75 36.835 ;
    RECT 233.48 36.045 233.69 36.115 ;
    RECT 233.48 36.405 233.69 36.475 ;
    RECT 233.48 36.765 233.69 36.835 ;
    RECT 233.02 36.045 233.23 36.115 ;
    RECT 233.02 36.405 233.23 36.475 ;
    RECT 233.02 36.765 233.23 36.835 ;
    RECT 230.16 36.045 230.37 36.115 ;
    RECT 230.16 36.405 230.37 36.475 ;
    RECT 230.16 36.765 230.37 36.835 ;
    RECT 229.7 36.045 229.91 36.115 ;
    RECT 229.7 36.405 229.91 36.475 ;
    RECT 229.7 36.765 229.91 36.835 ;
    RECT 366.28 36.045 366.49 36.115 ;
    RECT 366.28 36.405 366.49 36.475 ;
    RECT 366.28 36.765 366.49 36.835 ;
    RECT 365.82 36.045 366.03 36.115 ;
    RECT 365.82 36.405 366.03 36.475 ;
    RECT 365.82 36.765 366.03 36.835 ;
    RECT 226.84 36.045 227.05 36.115 ;
    RECT 226.84 36.405 227.05 36.475 ;
    RECT 226.84 36.765 227.05 36.835 ;
    RECT 226.38 36.045 226.59 36.115 ;
    RECT 226.38 36.405 226.59 36.475 ;
    RECT 226.38 36.765 226.59 36.835 ;
    RECT 362.96 36.045 363.17 36.115 ;
    RECT 362.96 36.405 363.17 36.475 ;
    RECT 362.96 36.765 363.17 36.835 ;
    RECT 362.5 36.045 362.71 36.115 ;
    RECT 362.5 36.405 362.71 36.475 ;
    RECT 362.5 36.765 362.71 36.835 ;
    RECT 223.52 36.045 223.73 36.115 ;
    RECT 223.52 36.405 223.73 36.475 ;
    RECT 223.52 36.765 223.73 36.835 ;
    RECT 223.06 36.045 223.27 36.115 ;
    RECT 223.06 36.405 223.27 36.475 ;
    RECT 223.06 36.765 223.27 36.835 ;
    RECT 359.64 36.045 359.85 36.115 ;
    RECT 359.64 36.405 359.85 36.475 ;
    RECT 359.64 36.765 359.85 36.835 ;
    RECT 359.18 36.045 359.39 36.115 ;
    RECT 359.18 36.405 359.39 36.475 ;
    RECT 359.18 36.765 359.39 36.835 ;
    RECT 220.2 36.045 220.41 36.115 ;
    RECT 220.2 36.405 220.41 36.475 ;
    RECT 220.2 36.765 220.41 36.835 ;
    RECT 219.74 36.045 219.95 36.115 ;
    RECT 219.74 36.405 219.95 36.475 ;
    RECT 219.74 36.765 219.95 36.835 ;
    RECT 356.32 36.045 356.53 36.115 ;
    RECT 356.32 36.405 356.53 36.475 ;
    RECT 356.32 36.765 356.53 36.835 ;
    RECT 355.86 36.045 356.07 36.115 ;
    RECT 355.86 36.405 356.07 36.475 ;
    RECT 355.86 36.765 356.07 36.835 ;
    RECT 353.0 36.045 353.21 36.115 ;
    RECT 353.0 36.405 353.21 36.475 ;
    RECT 353.0 36.765 353.21 36.835 ;
    RECT 352.54 36.045 352.75 36.115 ;
    RECT 352.54 36.405 352.75 36.475 ;
    RECT 352.54 36.765 352.75 36.835 ;
    RECT 216.88 36.045 217.09 36.115 ;
    RECT 216.88 36.405 217.09 36.475 ;
    RECT 216.88 36.765 217.09 36.835 ;
    RECT 216.42 36.045 216.63 36.115 ;
    RECT 216.42 36.405 216.63 36.475 ;
    RECT 216.42 36.765 216.63 36.835 ;
    RECT 349.68 36.045 349.89 36.115 ;
    RECT 349.68 36.405 349.89 36.475 ;
    RECT 349.68 36.765 349.89 36.835 ;
    RECT 349.22 36.045 349.43 36.115 ;
    RECT 349.22 36.405 349.43 36.475 ;
    RECT 349.22 36.765 349.43 36.835 ;
    RECT 213.56 36.045 213.77 36.115 ;
    RECT 213.56 36.405 213.77 36.475 ;
    RECT 213.56 36.765 213.77 36.835 ;
    RECT 213.1 36.045 213.31 36.115 ;
    RECT 213.1 36.405 213.31 36.475 ;
    RECT 213.1 36.765 213.31 36.835 ;
    RECT 346.36 36.045 346.57 36.115 ;
    RECT 346.36 36.405 346.57 36.475 ;
    RECT 346.36 36.765 346.57 36.835 ;
    RECT 345.9 36.045 346.11 36.115 ;
    RECT 345.9 36.405 346.11 36.475 ;
    RECT 345.9 36.765 346.11 36.835 ;
    RECT 210.24 36.045 210.45 36.115 ;
    RECT 210.24 36.405 210.45 36.475 ;
    RECT 210.24 36.765 210.45 36.835 ;
    RECT 209.78 36.045 209.99 36.115 ;
    RECT 209.78 36.405 209.99 36.475 ;
    RECT 209.78 36.765 209.99 36.835 ;
    RECT 343.04 36.045 343.25 36.115 ;
    RECT 343.04 36.405 343.25 36.475 ;
    RECT 343.04 36.765 343.25 36.835 ;
    RECT 342.58 36.045 342.79 36.115 ;
    RECT 342.58 36.405 342.79 36.475 ;
    RECT 342.58 36.765 342.79 36.835 ;
    RECT 206.92 36.045 207.13 36.115 ;
    RECT 206.92 36.405 207.13 36.475 ;
    RECT 206.92 36.765 207.13 36.835 ;
    RECT 206.46 36.045 206.67 36.115 ;
    RECT 206.46 36.405 206.67 36.475 ;
    RECT 206.46 36.765 206.67 36.835 ;
    RECT 339.72 36.045 339.93 36.115 ;
    RECT 339.72 36.405 339.93 36.475 ;
    RECT 339.72 36.765 339.93 36.835 ;
    RECT 339.26 36.045 339.47 36.115 ;
    RECT 339.26 36.405 339.47 36.475 ;
    RECT 339.26 36.765 339.47 36.835 ;
    RECT 203.6 36.045 203.81 36.115 ;
    RECT 203.6 36.405 203.81 36.475 ;
    RECT 203.6 36.765 203.81 36.835 ;
    RECT 203.14 36.045 203.35 36.115 ;
    RECT 203.14 36.405 203.35 36.475 ;
    RECT 203.14 36.765 203.35 36.835 ;
    RECT 336.4 36.045 336.61 36.115 ;
    RECT 336.4 36.405 336.61 36.475 ;
    RECT 336.4 36.765 336.61 36.835 ;
    RECT 335.94 36.045 336.15 36.115 ;
    RECT 335.94 36.405 336.15 36.475 ;
    RECT 335.94 36.765 336.15 36.835 ;
    RECT 266.68 36.045 266.89 36.115 ;
    RECT 266.68 36.405 266.89 36.475 ;
    RECT 266.68 36.765 266.89 36.835 ;
    RECT 266.22 36.045 266.43 36.115 ;
    RECT 266.22 36.405 266.43 36.475 ;
    RECT 266.22 36.765 266.43 36.835 ;
    RECT 263.36 36.045 263.57 36.115 ;
    RECT 263.36 36.405 263.57 36.475 ;
    RECT 263.36 36.765 263.57 36.835 ;
    RECT 262.9 36.045 263.11 36.115 ;
    RECT 262.9 36.405 263.11 36.475 ;
    RECT 262.9 36.765 263.11 36.835 ;
    RECT 260.04 36.045 260.25 36.115 ;
    RECT 260.04 36.405 260.25 36.475 ;
    RECT 260.04 36.765 260.25 36.835 ;
    RECT 259.58 36.045 259.79 36.115 ;
    RECT 259.58 36.405 259.79 36.475 ;
    RECT 259.58 36.765 259.79 36.835 ;
    RECT 256.72 36.045 256.93 36.115 ;
    RECT 256.72 36.405 256.93 36.475 ;
    RECT 256.72 36.765 256.93 36.835 ;
    RECT 256.26 36.045 256.47 36.115 ;
    RECT 256.26 36.405 256.47 36.475 ;
    RECT 256.26 36.765 256.47 36.835 ;
    RECT 253.4 36.045 253.61 36.115 ;
    RECT 253.4 36.405 253.61 36.475 ;
    RECT 253.4 36.765 253.61 36.835 ;
    RECT 252.94 36.045 253.15 36.115 ;
    RECT 252.94 36.405 253.15 36.475 ;
    RECT 252.94 36.765 253.15 36.835 ;
    RECT 250.08 36.045 250.29 36.115 ;
    RECT 250.08 36.405 250.29 36.475 ;
    RECT 250.08 36.765 250.29 36.835 ;
    RECT 249.62 36.045 249.83 36.115 ;
    RECT 249.62 36.405 249.83 36.475 ;
    RECT 249.62 36.765 249.83 36.835 ;
    RECT 246.76 36.045 246.97 36.115 ;
    RECT 246.76 36.405 246.97 36.475 ;
    RECT 246.76 36.765 246.97 36.835 ;
    RECT 246.3 36.045 246.51 36.115 ;
    RECT 246.3 36.405 246.51 36.475 ;
    RECT 246.3 36.765 246.51 36.835 ;
    RECT 243.44 36.045 243.65 36.115 ;
    RECT 243.44 36.405 243.65 36.475 ;
    RECT 243.44 36.765 243.65 36.835 ;
    RECT 242.98 36.045 243.19 36.115 ;
    RECT 242.98 36.405 243.19 36.475 ;
    RECT 242.98 36.765 243.19 36.835 ;
    RECT 240.12 36.045 240.33 36.115 ;
    RECT 240.12 36.405 240.33 36.475 ;
    RECT 240.12 36.765 240.33 36.835 ;
    RECT 239.66 36.045 239.87 36.115 ;
    RECT 239.66 36.405 239.87 36.475 ;
    RECT 239.66 36.765 239.87 36.835 ;
    RECT 236.8 36.045 237.01 36.115 ;
    RECT 236.8 36.405 237.01 36.475 ;
    RECT 236.8 36.765 237.01 36.835 ;
    RECT 236.34 36.045 236.55 36.115 ;
    RECT 236.34 36.405 236.55 36.475 ;
    RECT 236.34 36.765 236.55 36.835 ;
    RECT 374.15 36.405 374.22 36.475 ;
    RECT 333.08 36.045 333.29 36.115 ;
    RECT 333.08 36.405 333.29 36.475 ;
    RECT 333.08 36.765 333.29 36.835 ;
    RECT 332.62 36.045 332.83 36.115 ;
    RECT 332.62 36.405 332.83 36.475 ;
    RECT 332.62 36.765 332.83 36.835 ;
    RECT 329.76 36.045 329.97 36.115 ;
    RECT 329.76 36.405 329.97 36.475 ;
    RECT 329.76 36.765 329.97 36.835 ;
    RECT 329.3 36.045 329.51 36.115 ;
    RECT 329.3 36.405 329.51 36.475 ;
    RECT 329.3 36.765 329.51 36.835 ;
    RECT 326.44 36.045 326.65 36.115 ;
    RECT 326.44 36.405 326.65 36.475 ;
    RECT 326.44 36.765 326.65 36.835 ;
    RECT 325.98 36.045 326.19 36.115 ;
    RECT 325.98 36.405 326.19 36.475 ;
    RECT 325.98 36.765 326.19 36.835 ;
    RECT 323.12 36.045 323.33 36.115 ;
    RECT 323.12 36.405 323.33 36.475 ;
    RECT 323.12 36.765 323.33 36.835 ;
    RECT 322.66 36.045 322.87 36.115 ;
    RECT 322.66 36.405 322.87 36.475 ;
    RECT 322.66 36.765 322.87 36.835 ;
    RECT 319.8 36.045 320.01 36.115 ;
    RECT 319.8 36.405 320.01 36.475 ;
    RECT 319.8 36.765 320.01 36.835 ;
    RECT 319.34 36.045 319.55 36.115 ;
    RECT 319.34 36.405 319.55 36.475 ;
    RECT 319.34 36.765 319.55 36.835 ;
    RECT 316.48 36.045 316.69 36.115 ;
    RECT 316.48 36.405 316.69 36.475 ;
    RECT 316.48 36.765 316.69 36.835 ;
    RECT 316.02 36.045 316.23 36.115 ;
    RECT 316.02 36.405 316.23 36.475 ;
    RECT 316.02 36.765 316.23 36.835 ;
    RECT 313.16 36.045 313.37 36.115 ;
    RECT 313.16 36.405 313.37 36.475 ;
    RECT 313.16 36.765 313.37 36.835 ;
    RECT 312.7 36.045 312.91 36.115 ;
    RECT 312.7 36.405 312.91 36.475 ;
    RECT 312.7 36.765 312.91 36.835 ;
    RECT 309.84 36.045 310.05 36.115 ;
    RECT 309.84 36.405 310.05 36.475 ;
    RECT 309.84 36.765 310.05 36.835 ;
    RECT 309.38 36.045 309.59 36.115 ;
    RECT 309.38 36.405 309.59 36.475 ;
    RECT 309.38 36.765 309.59 36.835 ;
    RECT 306.52 36.045 306.73 36.115 ;
    RECT 306.52 36.405 306.73 36.475 ;
    RECT 306.52 36.765 306.73 36.835 ;
    RECT 306.06 36.045 306.27 36.115 ;
    RECT 306.06 36.405 306.27 36.475 ;
    RECT 306.06 36.765 306.27 36.835 ;
    RECT 61.25 49.725 61.46 49.795 ;
    RECT 61.25 50.085 61.46 50.155 ;
    RECT 61.25 50.445 61.46 50.515 ;
    RECT 61.71 49.725 61.92 49.795 ;
    RECT 61.71 50.085 61.92 50.155 ;
    RECT 61.71 50.445 61.92 50.515 ;
    RECT 57.93 49.725 58.14 49.795 ;
    RECT 57.93 50.085 58.14 50.155 ;
    RECT 57.93 50.445 58.14 50.515 ;
    RECT 58.39 49.725 58.6 49.795 ;
    RECT 58.39 50.085 58.6 50.155 ;
    RECT 58.39 50.445 58.6 50.515 ;
    RECT 54.61 49.725 54.82 49.795 ;
    RECT 54.61 50.085 54.82 50.155 ;
    RECT 54.61 50.445 54.82 50.515 ;
    RECT 55.07 49.725 55.28 49.795 ;
    RECT 55.07 50.085 55.28 50.155 ;
    RECT 55.07 50.445 55.28 50.515 ;
    RECT 51.29 49.725 51.5 49.795 ;
    RECT 51.29 50.085 51.5 50.155 ;
    RECT 51.29 50.445 51.5 50.515 ;
    RECT 51.75 49.725 51.96 49.795 ;
    RECT 51.75 50.085 51.96 50.155 ;
    RECT 51.75 50.445 51.96 50.515 ;
    RECT 47.97 49.725 48.18 49.795 ;
    RECT 47.97 50.085 48.18 50.155 ;
    RECT 47.97 50.445 48.18 50.515 ;
    RECT 48.43 49.725 48.64 49.795 ;
    RECT 48.43 50.085 48.64 50.155 ;
    RECT 48.43 50.445 48.64 50.515 ;
    RECT 44.65 49.725 44.86 49.795 ;
    RECT 44.65 50.085 44.86 50.155 ;
    RECT 44.65 50.445 44.86 50.515 ;
    RECT 45.11 49.725 45.32 49.795 ;
    RECT 45.11 50.085 45.32 50.155 ;
    RECT 45.11 50.445 45.32 50.515 ;
    RECT 41.33 49.725 41.54 49.795 ;
    RECT 41.33 50.085 41.54 50.155 ;
    RECT 41.33 50.445 41.54 50.515 ;
    RECT 41.79 49.725 42.0 49.795 ;
    RECT 41.79 50.085 42.0 50.155 ;
    RECT 41.79 50.445 42.0 50.515 ;
    RECT 38.01 49.725 38.22 49.795 ;
    RECT 38.01 50.085 38.22 50.155 ;
    RECT 38.01 50.445 38.22 50.515 ;
    RECT 38.47 49.725 38.68 49.795 ;
    RECT 38.47 50.085 38.68 50.155 ;
    RECT 38.47 50.445 38.68 50.515 ;
    RECT 34.69 49.725 34.9 49.795 ;
    RECT 34.69 50.085 34.9 50.155 ;
    RECT 34.69 50.445 34.9 50.515 ;
    RECT 35.15 49.725 35.36 49.795 ;
    RECT 35.15 50.085 35.36 50.155 ;
    RECT 35.15 50.445 35.36 50.515 ;
    RECT 173.945 50.085 174.015 50.155 ;
    RECT 130.97 49.725 131.18 49.795 ;
    RECT 130.97 50.085 131.18 50.155 ;
    RECT 130.97 50.445 131.18 50.515 ;
    RECT 131.43 49.725 131.64 49.795 ;
    RECT 131.43 50.085 131.64 50.155 ;
    RECT 131.43 50.445 131.64 50.515 ;
    RECT 127.65 49.725 127.86 49.795 ;
    RECT 127.65 50.085 127.86 50.155 ;
    RECT 127.65 50.445 127.86 50.515 ;
    RECT 128.11 49.725 128.32 49.795 ;
    RECT 128.11 50.085 128.32 50.155 ;
    RECT 128.11 50.445 128.32 50.515 ;
    RECT 124.33 49.725 124.54 49.795 ;
    RECT 124.33 50.085 124.54 50.155 ;
    RECT 124.33 50.445 124.54 50.515 ;
    RECT 124.79 49.725 125.0 49.795 ;
    RECT 124.79 50.085 125.0 50.155 ;
    RECT 124.79 50.445 125.0 50.515 ;
    RECT 121.01 49.725 121.22 49.795 ;
    RECT 121.01 50.085 121.22 50.155 ;
    RECT 121.01 50.445 121.22 50.515 ;
    RECT 121.47 49.725 121.68 49.795 ;
    RECT 121.47 50.085 121.68 50.155 ;
    RECT 121.47 50.445 121.68 50.515 ;
    RECT 117.69 49.725 117.9 49.795 ;
    RECT 117.69 50.085 117.9 50.155 ;
    RECT 117.69 50.445 117.9 50.515 ;
    RECT 118.15 49.725 118.36 49.795 ;
    RECT 118.15 50.085 118.36 50.155 ;
    RECT 118.15 50.445 118.36 50.515 ;
    RECT 114.37 49.725 114.58 49.795 ;
    RECT 114.37 50.085 114.58 50.155 ;
    RECT 114.37 50.445 114.58 50.515 ;
    RECT 114.83 49.725 115.04 49.795 ;
    RECT 114.83 50.085 115.04 50.155 ;
    RECT 114.83 50.445 115.04 50.515 ;
    RECT 111.05 49.725 111.26 49.795 ;
    RECT 111.05 50.085 111.26 50.155 ;
    RECT 111.05 50.445 111.26 50.515 ;
    RECT 111.51 49.725 111.72 49.795 ;
    RECT 111.51 50.085 111.72 50.155 ;
    RECT 111.51 50.445 111.72 50.515 ;
    RECT 107.73 49.725 107.94 49.795 ;
    RECT 107.73 50.085 107.94 50.155 ;
    RECT 107.73 50.445 107.94 50.515 ;
    RECT 108.19 49.725 108.4 49.795 ;
    RECT 108.19 50.085 108.4 50.155 ;
    RECT 108.19 50.445 108.4 50.515 ;
    RECT 104.41 49.725 104.62 49.795 ;
    RECT 104.41 50.085 104.62 50.155 ;
    RECT 104.41 50.445 104.62 50.515 ;
    RECT 104.87 49.725 105.08 49.795 ;
    RECT 104.87 50.085 105.08 50.155 ;
    RECT 104.87 50.445 105.08 50.515 ;
    RECT 101.09 49.725 101.3 49.795 ;
    RECT 101.09 50.085 101.3 50.155 ;
    RECT 101.09 50.445 101.3 50.515 ;
    RECT 101.55 49.725 101.76 49.795 ;
    RECT 101.55 50.085 101.76 50.155 ;
    RECT 101.55 50.445 101.76 50.515 ;
    RECT 0.4 50.085 0.47 50.155 ;
    RECT 170.81 49.725 171.02 49.795 ;
    RECT 170.81 50.085 171.02 50.155 ;
    RECT 170.81 50.445 171.02 50.515 ;
    RECT 171.27 49.725 171.48 49.795 ;
    RECT 171.27 50.085 171.48 50.155 ;
    RECT 171.27 50.445 171.48 50.515 ;
    RECT 167.49 49.725 167.7 49.795 ;
    RECT 167.49 50.085 167.7 50.155 ;
    RECT 167.49 50.445 167.7 50.515 ;
    RECT 167.95 49.725 168.16 49.795 ;
    RECT 167.95 50.085 168.16 50.155 ;
    RECT 167.95 50.445 168.16 50.515 ;
    RECT 97.77 49.725 97.98 49.795 ;
    RECT 97.77 50.085 97.98 50.155 ;
    RECT 97.77 50.445 97.98 50.515 ;
    RECT 98.23 49.725 98.44 49.795 ;
    RECT 98.23 50.085 98.44 50.155 ;
    RECT 98.23 50.445 98.44 50.515 ;
    RECT 94.45 49.725 94.66 49.795 ;
    RECT 94.45 50.085 94.66 50.155 ;
    RECT 94.45 50.445 94.66 50.515 ;
    RECT 94.91 49.725 95.12 49.795 ;
    RECT 94.91 50.085 95.12 50.155 ;
    RECT 94.91 50.445 95.12 50.515 ;
    RECT 91.13 49.725 91.34 49.795 ;
    RECT 91.13 50.085 91.34 50.155 ;
    RECT 91.13 50.445 91.34 50.515 ;
    RECT 91.59 49.725 91.8 49.795 ;
    RECT 91.59 50.085 91.8 50.155 ;
    RECT 91.59 50.445 91.8 50.515 ;
    RECT 87.81 49.725 88.02 49.795 ;
    RECT 87.81 50.085 88.02 50.155 ;
    RECT 87.81 50.445 88.02 50.515 ;
    RECT 88.27 49.725 88.48 49.795 ;
    RECT 88.27 50.085 88.48 50.155 ;
    RECT 88.27 50.445 88.48 50.515 ;
    RECT 84.49 49.725 84.7 49.795 ;
    RECT 84.49 50.085 84.7 50.155 ;
    RECT 84.49 50.445 84.7 50.515 ;
    RECT 84.95 49.725 85.16 49.795 ;
    RECT 84.95 50.085 85.16 50.155 ;
    RECT 84.95 50.445 85.16 50.515 ;
    RECT 81.17 49.725 81.38 49.795 ;
    RECT 81.17 50.085 81.38 50.155 ;
    RECT 81.17 50.445 81.38 50.515 ;
    RECT 81.63 49.725 81.84 49.795 ;
    RECT 81.63 50.085 81.84 50.155 ;
    RECT 81.63 50.445 81.84 50.515 ;
    RECT 77.85 49.725 78.06 49.795 ;
    RECT 77.85 50.085 78.06 50.155 ;
    RECT 77.85 50.445 78.06 50.515 ;
    RECT 78.31 49.725 78.52 49.795 ;
    RECT 78.31 50.085 78.52 50.155 ;
    RECT 78.31 50.445 78.52 50.515 ;
    RECT 74.53 49.725 74.74 49.795 ;
    RECT 74.53 50.085 74.74 50.155 ;
    RECT 74.53 50.445 74.74 50.515 ;
    RECT 74.99 49.725 75.2 49.795 ;
    RECT 74.99 50.085 75.2 50.155 ;
    RECT 74.99 50.445 75.2 50.515 ;
    RECT 71.21 49.725 71.42 49.795 ;
    RECT 71.21 50.085 71.42 50.155 ;
    RECT 71.21 50.445 71.42 50.515 ;
    RECT 71.67 49.725 71.88 49.795 ;
    RECT 71.67 50.085 71.88 50.155 ;
    RECT 71.67 50.445 71.88 50.515 ;
    RECT 31.37 49.725 31.58 49.795 ;
    RECT 31.37 50.085 31.58 50.155 ;
    RECT 31.37 50.445 31.58 50.515 ;
    RECT 31.83 49.725 32.04 49.795 ;
    RECT 31.83 50.085 32.04 50.155 ;
    RECT 31.83 50.445 32.04 50.515 ;
    RECT 67.89 49.725 68.1 49.795 ;
    RECT 67.89 50.085 68.1 50.155 ;
    RECT 67.89 50.445 68.1 50.515 ;
    RECT 68.35 49.725 68.56 49.795 ;
    RECT 68.35 50.085 68.56 50.155 ;
    RECT 68.35 50.445 68.56 50.515 ;
    RECT 28.05 49.725 28.26 49.795 ;
    RECT 28.05 50.085 28.26 50.155 ;
    RECT 28.05 50.445 28.26 50.515 ;
    RECT 28.51 49.725 28.72 49.795 ;
    RECT 28.51 50.085 28.72 50.155 ;
    RECT 28.51 50.445 28.72 50.515 ;
    RECT 24.73 49.725 24.94 49.795 ;
    RECT 24.73 50.085 24.94 50.155 ;
    RECT 24.73 50.445 24.94 50.515 ;
    RECT 25.19 49.725 25.4 49.795 ;
    RECT 25.19 50.085 25.4 50.155 ;
    RECT 25.19 50.445 25.4 50.515 ;
    RECT 21.41 49.725 21.62 49.795 ;
    RECT 21.41 50.085 21.62 50.155 ;
    RECT 21.41 50.445 21.62 50.515 ;
    RECT 21.87 49.725 22.08 49.795 ;
    RECT 21.87 50.085 22.08 50.155 ;
    RECT 21.87 50.445 22.08 50.515 ;
    RECT 18.09 49.725 18.3 49.795 ;
    RECT 18.09 50.085 18.3 50.155 ;
    RECT 18.09 50.445 18.3 50.515 ;
    RECT 18.55 49.725 18.76 49.795 ;
    RECT 18.55 50.085 18.76 50.155 ;
    RECT 18.55 50.445 18.76 50.515 ;
    RECT 14.77 49.725 14.98 49.795 ;
    RECT 14.77 50.085 14.98 50.155 ;
    RECT 14.77 50.445 14.98 50.515 ;
    RECT 15.23 49.725 15.44 49.795 ;
    RECT 15.23 50.085 15.44 50.155 ;
    RECT 15.23 50.445 15.44 50.515 ;
    RECT 11.45 49.725 11.66 49.795 ;
    RECT 11.45 50.085 11.66 50.155 ;
    RECT 11.45 50.445 11.66 50.515 ;
    RECT 11.91 49.725 12.12 49.795 ;
    RECT 11.91 50.085 12.12 50.155 ;
    RECT 11.91 50.445 12.12 50.515 ;
    RECT 8.13 49.725 8.34 49.795 ;
    RECT 8.13 50.085 8.34 50.155 ;
    RECT 8.13 50.445 8.34 50.515 ;
    RECT 8.59 49.725 8.8 49.795 ;
    RECT 8.59 50.085 8.8 50.155 ;
    RECT 8.59 50.445 8.8 50.515 ;
    RECT 4.81 49.725 5.02 49.795 ;
    RECT 4.81 50.085 5.02 50.155 ;
    RECT 4.81 50.445 5.02 50.515 ;
    RECT 5.27 49.725 5.48 49.795 ;
    RECT 5.27 50.085 5.48 50.155 ;
    RECT 5.27 50.445 5.48 50.515 ;
    RECT 164.17 49.725 164.38 49.795 ;
    RECT 164.17 50.085 164.38 50.155 ;
    RECT 164.17 50.445 164.38 50.515 ;
    RECT 164.63 49.725 164.84 49.795 ;
    RECT 164.63 50.085 164.84 50.155 ;
    RECT 164.63 50.445 164.84 50.515 ;
    RECT 1.49 49.725 1.7 49.795 ;
    RECT 1.49 50.085 1.7 50.155 ;
    RECT 1.49 50.445 1.7 50.515 ;
    RECT 1.95 49.725 2.16 49.795 ;
    RECT 1.95 50.085 2.16 50.155 ;
    RECT 1.95 50.445 2.16 50.515 ;
    RECT 160.85 49.725 161.06 49.795 ;
    RECT 160.85 50.085 161.06 50.155 ;
    RECT 160.85 50.445 161.06 50.515 ;
    RECT 161.31 49.725 161.52 49.795 ;
    RECT 161.31 50.085 161.52 50.155 ;
    RECT 161.31 50.445 161.52 50.515 ;
    RECT 157.53 49.725 157.74 49.795 ;
    RECT 157.53 50.085 157.74 50.155 ;
    RECT 157.53 50.445 157.74 50.515 ;
    RECT 157.99 49.725 158.2 49.795 ;
    RECT 157.99 50.085 158.2 50.155 ;
    RECT 157.99 50.445 158.2 50.515 ;
    RECT 154.21 49.725 154.42 49.795 ;
    RECT 154.21 50.085 154.42 50.155 ;
    RECT 154.21 50.445 154.42 50.515 ;
    RECT 154.67 49.725 154.88 49.795 ;
    RECT 154.67 50.085 154.88 50.155 ;
    RECT 154.67 50.445 154.88 50.515 ;
    RECT 150.89 49.725 151.1 49.795 ;
    RECT 150.89 50.085 151.1 50.155 ;
    RECT 150.89 50.445 151.1 50.515 ;
    RECT 151.35 49.725 151.56 49.795 ;
    RECT 151.35 50.085 151.56 50.155 ;
    RECT 151.35 50.445 151.56 50.515 ;
    RECT 147.57 49.725 147.78 49.795 ;
    RECT 147.57 50.085 147.78 50.155 ;
    RECT 147.57 50.445 147.78 50.515 ;
    RECT 148.03 49.725 148.24 49.795 ;
    RECT 148.03 50.085 148.24 50.155 ;
    RECT 148.03 50.445 148.24 50.515 ;
    RECT 144.25 49.725 144.46 49.795 ;
    RECT 144.25 50.085 144.46 50.155 ;
    RECT 144.25 50.445 144.46 50.515 ;
    RECT 144.71 49.725 144.92 49.795 ;
    RECT 144.71 50.085 144.92 50.155 ;
    RECT 144.71 50.445 144.92 50.515 ;
    RECT 140.93 49.725 141.14 49.795 ;
    RECT 140.93 50.085 141.14 50.155 ;
    RECT 140.93 50.445 141.14 50.515 ;
    RECT 141.39 49.725 141.6 49.795 ;
    RECT 141.39 50.085 141.6 50.155 ;
    RECT 141.39 50.445 141.6 50.515 ;
    RECT 137.61 49.725 137.82 49.795 ;
    RECT 137.61 50.085 137.82 50.155 ;
    RECT 137.61 50.445 137.82 50.515 ;
    RECT 138.07 49.725 138.28 49.795 ;
    RECT 138.07 50.085 138.28 50.155 ;
    RECT 138.07 50.445 138.28 50.515 ;
    RECT 134.29 49.725 134.5 49.795 ;
    RECT 134.29 50.085 134.5 50.155 ;
    RECT 134.29 50.445 134.5 50.515 ;
    RECT 134.75 49.725 134.96 49.795 ;
    RECT 134.75 50.085 134.96 50.155 ;
    RECT 134.75 50.445 134.96 50.515 ;
    RECT 64.57 49.725 64.78 49.795 ;
    RECT 64.57 50.085 64.78 50.155 ;
    RECT 64.57 50.445 64.78 50.515 ;
    RECT 65.03 49.725 65.24 49.795 ;
    RECT 65.03 50.085 65.24 50.155 ;
    RECT 65.03 50.445 65.24 50.515 ;
    RECT 61.25 49.005 61.46 49.075 ;
    RECT 61.25 49.365 61.46 49.435 ;
    RECT 61.25 49.725 61.46 49.795 ;
    RECT 61.71 49.005 61.92 49.075 ;
    RECT 61.71 49.365 61.92 49.435 ;
    RECT 61.71 49.725 61.92 49.795 ;
    RECT 57.93 49.005 58.14 49.075 ;
    RECT 57.93 49.365 58.14 49.435 ;
    RECT 57.93 49.725 58.14 49.795 ;
    RECT 58.39 49.005 58.6 49.075 ;
    RECT 58.39 49.365 58.6 49.435 ;
    RECT 58.39 49.725 58.6 49.795 ;
    RECT 54.61 49.005 54.82 49.075 ;
    RECT 54.61 49.365 54.82 49.435 ;
    RECT 54.61 49.725 54.82 49.795 ;
    RECT 55.07 49.005 55.28 49.075 ;
    RECT 55.07 49.365 55.28 49.435 ;
    RECT 55.07 49.725 55.28 49.795 ;
    RECT 51.29 49.005 51.5 49.075 ;
    RECT 51.29 49.365 51.5 49.435 ;
    RECT 51.29 49.725 51.5 49.795 ;
    RECT 51.75 49.005 51.96 49.075 ;
    RECT 51.75 49.365 51.96 49.435 ;
    RECT 51.75 49.725 51.96 49.795 ;
    RECT 47.97 49.005 48.18 49.075 ;
    RECT 47.97 49.365 48.18 49.435 ;
    RECT 47.97 49.725 48.18 49.795 ;
    RECT 48.43 49.005 48.64 49.075 ;
    RECT 48.43 49.365 48.64 49.435 ;
    RECT 48.43 49.725 48.64 49.795 ;
    RECT 44.65 49.005 44.86 49.075 ;
    RECT 44.65 49.365 44.86 49.435 ;
    RECT 44.65 49.725 44.86 49.795 ;
    RECT 45.11 49.005 45.32 49.075 ;
    RECT 45.11 49.365 45.32 49.435 ;
    RECT 45.11 49.725 45.32 49.795 ;
    RECT 41.33 49.005 41.54 49.075 ;
    RECT 41.33 49.365 41.54 49.435 ;
    RECT 41.33 49.725 41.54 49.795 ;
    RECT 41.79 49.005 42.0 49.075 ;
    RECT 41.79 49.365 42.0 49.435 ;
    RECT 41.79 49.725 42.0 49.795 ;
    RECT 38.01 49.005 38.22 49.075 ;
    RECT 38.01 49.365 38.22 49.435 ;
    RECT 38.01 49.725 38.22 49.795 ;
    RECT 38.47 49.005 38.68 49.075 ;
    RECT 38.47 49.365 38.68 49.435 ;
    RECT 38.47 49.725 38.68 49.795 ;
    RECT 34.69 49.005 34.9 49.075 ;
    RECT 34.69 49.365 34.9 49.435 ;
    RECT 34.69 49.725 34.9 49.795 ;
    RECT 35.15 49.005 35.36 49.075 ;
    RECT 35.15 49.365 35.36 49.435 ;
    RECT 35.15 49.725 35.36 49.795 ;
    RECT 173.945 49.365 174.015 49.435 ;
    RECT 130.97 49.005 131.18 49.075 ;
    RECT 130.97 49.365 131.18 49.435 ;
    RECT 130.97 49.725 131.18 49.795 ;
    RECT 131.43 49.005 131.64 49.075 ;
    RECT 131.43 49.365 131.64 49.435 ;
    RECT 131.43 49.725 131.64 49.795 ;
    RECT 127.65 49.005 127.86 49.075 ;
    RECT 127.65 49.365 127.86 49.435 ;
    RECT 127.65 49.725 127.86 49.795 ;
    RECT 128.11 49.005 128.32 49.075 ;
    RECT 128.11 49.365 128.32 49.435 ;
    RECT 128.11 49.725 128.32 49.795 ;
    RECT 124.33 49.005 124.54 49.075 ;
    RECT 124.33 49.365 124.54 49.435 ;
    RECT 124.33 49.725 124.54 49.795 ;
    RECT 124.79 49.005 125.0 49.075 ;
    RECT 124.79 49.365 125.0 49.435 ;
    RECT 124.79 49.725 125.0 49.795 ;
    RECT 121.01 49.005 121.22 49.075 ;
    RECT 121.01 49.365 121.22 49.435 ;
    RECT 121.01 49.725 121.22 49.795 ;
    RECT 121.47 49.005 121.68 49.075 ;
    RECT 121.47 49.365 121.68 49.435 ;
    RECT 121.47 49.725 121.68 49.795 ;
    RECT 117.69 49.005 117.9 49.075 ;
    RECT 117.69 49.365 117.9 49.435 ;
    RECT 117.69 49.725 117.9 49.795 ;
    RECT 118.15 49.005 118.36 49.075 ;
    RECT 118.15 49.365 118.36 49.435 ;
    RECT 118.15 49.725 118.36 49.795 ;
    RECT 114.37 49.005 114.58 49.075 ;
    RECT 114.37 49.365 114.58 49.435 ;
    RECT 114.37 49.725 114.58 49.795 ;
    RECT 114.83 49.005 115.04 49.075 ;
    RECT 114.83 49.365 115.04 49.435 ;
    RECT 114.83 49.725 115.04 49.795 ;
    RECT 111.05 49.005 111.26 49.075 ;
    RECT 111.05 49.365 111.26 49.435 ;
    RECT 111.05 49.725 111.26 49.795 ;
    RECT 111.51 49.005 111.72 49.075 ;
    RECT 111.51 49.365 111.72 49.435 ;
    RECT 111.51 49.725 111.72 49.795 ;
    RECT 107.73 49.005 107.94 49.075 ;
    RECT 107.73 49.365 107.94 49.435 ;
    RECT 107.73 49.725 107.94 49.795 ;
    RECT 108.19 49.005 108.4 49.075 ;
    RECT 108.19 49.365 108.4 49.435 ;
    RECT 108.19 49.725 108.4 49.795 ;
    RECT 104.41 49.005 104.62 49.075 ;
    RECT 104.41 49.365 104.62 49.435 ;
    RECT 104.41 49.725 104.62 49.795 ;
    RECT 104.87 49.005 105.08 49.075 ;
    RECT 104.87 49.365 105.08 49.435 ;
    RECT 104.87 49.725 105.08 49.795 ;
    RECT 101.09 49.005 101.3 49.075 ;
    RECT 101.09 49.365 101.3 49.435 ;
    RECT 101.09 49.725 101.3 49.795 ;
    RECT 101.55 49.005 101.76 49.075 ;
    RECT 101.55 49.365 101.76 49.435 ;
    RECT 101.55 49.725 101.76 49.795 ;
    RECT 0.4 49.365 0.47 49.435 ;
    RECT 170.81 49.005 171.02 49.075 ;
    RECT 170.81 49.365 171.02 49.435 ;
    RECT 170.81 49.725 171.02 49.795 ;
    RECT 171.27 49.005 171.48 49.075 ;
    RECT 171.27 49.365 171.48 49.435 ;
    RECT 171.27 49.725 171.48 49.795 ;
    RECT 167.49 49.005 167.7 49.075 ;
    RECT 167.49 49.365 167.7 49.435 ;
    RECT 167.49 49.725 167.7 49.795 ;
    RECT 167.95 49.005 168.16 49.075 ;
    RECT 167.95 49.365 168.16 49.435 ;
    RECT 167.95 49.725 168.16 49.795 ;
    RECT 97.77 49.005 97.98 49.075 ;
    RECT 97.77 49.365 97.98 49.435 ;
    RECT 97.77 49.725 97.98 49.795 ;
    RECT 98.23 49.005 98.44 49.075 ;
    RECT 98.23 49.365 98.44 49.435 ;
    RECT 98.23 49.725 98.44 49.795 ;
    RECT 94.45 49.005 94.66 49.075 ;
    RECT 94.45 49.365 94.66 49.435 ;
    RECT 94.45 49.725 94.66 49.795 ;
    RECT 94.91 49.005 95.12 49.075 ;
    RECT 94.91 49.365 95.12 49.435 ;
    RECT 94.91 49.725 95.12 49.795 ;
    RECT 91.13 49.005 91.34 49.075 ;
    RECT 91.13 49.365 91.34 49.435 ;
    RECT 91.13 49.725 91.34 49.795 ;
    RECT 91.59 49.005 91.8 49.075 ;
    RECT 91.59 49.365 91.8 49.435 ;
    RECT 91.59 49.725 91.8 49.795 ;
    RECT 87.81 49.005 88.02 49.075 ;
    RECT 87.81 49.365 88.02 49.435 ;
    RECT 87.81 49.725 88.02 49.795 ;
    RECT 88.27 49.005 88.48 49.075 ;
    RECT 88.27 49.365 88.48 49.435 ;
    RECT 88.27 49.725 88.48 49.795 ;
    RECT 84.49 49.005 84.7 49.075 ;
    RECT 84.49 49.365 84.7 49.435 ;
    RECT 84.49 49.725 84.7 49.795 ;
    RECT 84.95 49.005 85.16 49.075 ;
    RECT 84.95 49.365 85.16 49.435 ;
    RECT 84.95 49.725 85.16 49.795 ;
    RECT 81.17 49.005 81.38 49.075 ;
    RECT 81.17 49.365 81.38 49.435 ;
    RECT 81.17 49.725 81.38 49.795 ;
    RECT 81.63 49.005 81.84 49.075 ;
    RECT 81.63 49.365 81.84 49.435 ;
    RECT 81.63 49.725 81.84 49.795 ;
    RECT 77.85 49.005 78.06 49.075 ;
    RECT 77.85 49.365 78.06 49.435 ;
    RECT 77.85 49.725 78.06 49.795 ;
    RECT 78.31 49.005 78.52 49.075 ;
    RECT 78.31 49.365 78.52 49.435 ;
    RECT 78.31 49.725 78.52 49.795 ;
    RECT 74.53 49.005 74.74 49.075 ;
    RECT 74.53 49.365 74.74 49.435 ;
    RECT 74.53 49.725 74.74 49.795 ;
    RECT 74.99 49.005 75.2 49.075 ;
    RECT 74.99 49.365 75.2 49.435 ;
    RECT 74.99 49.725 75.2 49.795 ;
    RECT 71.21 49.005 71.42 49.075 ;
    RECT 71.21 49.365 71.42 49.435 ;
    RECT 71.21 49.725 71.42 49.795 ;
    RECT 71.67 49.005 71.88 49.075 ;
    RECT 71.67 49.365 71.88 49.435 ;
    RECT 71.67 49.725 71.88 49.795 ;
    RECT 31.37 49.005 31.58 49.075 ;
    RECT 31.37 49.365 31.58 49.435 ;
    RECT 31.37 49.725 31.58 49.795 ;
    RECT 31.83 49.005 32.04 49.075 ;
    RECT 31.83 49.365 32.04 49.435 ;
    RECT 31.83 49.725 32.04 49.795 ;
    RECT 67.89 49.005 68.1 49.075 ;
    RECT 67.89 49.365 68.1 49.435 ;
    RECT 67.89 49.725 68.1 49.795 ;
    RECT 68.35 49.005 68.56 49.075 ;
    RECT 68.35 49.365 68.56 49.435 ;
    RECT 68.35 49.725 68.56 49.795 ;
    RECT 28.05 49.005 28.26 49.075 ;
    RECT 28.05 49.365 28.26 49.435 ;
    RECT 28.05 49.725 28.26 49.795 ;
    RECT 28.51 49.005 28.72 49.075 ;
    RECT 28.51 49.365 28.72 49.435 ;
    RECT 28.51 49.725 28.72 49.795 ;
    RECT 24.73 49.005 24.94 49.075 ;
    RECT 24.73 49.365 24.94 49.435 ;
    RECT 24.73 49.725 24.94 49.795 ;
    RECT 25.19 49.005 25.4 49.075 ;
    RECT 25.19 49.365 25.4 49.435 ;
    RECT 25.19 49.725 25.4 49.795 ;
    RECT 21.41 49.005 21.62 49.075 ;
    RECT 21.41 49.365 21.62 49.435 ;
    RECT 21.41 49.725 21.62 49.795 ;
    RECT 21.87 49.005 22.08 49.075 ;
    RECT 21.87 49.365 22.08 49.435 ;
    RECT 21.87 49.725 22.08 49.795 ;
    RECT 18.09 49.005 18.3 49.075 ;
    RECT 18.09 49.365 18.3 49.435 ;
    RECT 18.09 49.725 18.3 49.795 ;
    RECT 18.55 49.005 18.76 49.075 ;
    RECT 18.55 49.365 18.76 49.435 ;
    RECT 18.55 49.725 18.76 49.795 ;
    RECT 14.77 49.005 14.98 49.075 ;
    RECT 14.77 49.365 14.98 49.435 ;
    RECT 14.77 49.725 14.98 49.795 ;
    RECT 15.23 49.005 15.44 49.075 ;
    RECT 15.23 49.365 15.44 49.435 ;
    RECT 15.23 49.725 15.44 49.795 ;
    RECT 11.45 49.005 11.66 49.075 ;
    RECT 11.45 49.365 11.66 49.435 ;
    RECT 11.45 49.725 11.66 49.795 ;
    RECT 11.91 49.005 12.12 49.075 ;
    RECT 11.91 49.365 12.12 49.435 ;
    RECT 11.91 49.725 12.12 49.795 ;
    RECT 8.13 49.005 8.34 49.075 ;
    RECT 8.13 49.365 8.34 49.435 ;
    RECT 8.13 49.725 8.34 49.795 ;
    RECT 8.59 49.005 8.8 49.075 ;
    RECT 8.59 49.365 8.8 49.435 ;
    RECT 8.59 49.725 8.8 49.795 ;
    RECT 4.81 49.005 5.02 49.075 ;
    RECT 4.81 49.365 5.02 49.435 ;
    RECT 4.81 49.725 5.02 49.795 ;
    RECT 5.27 49.005 5.48 49.075 ;
    RECT 5.27 49.365 5.48 49.435 ;
    RECT 5.27 49.725 5.48 49.795 ;
    RECT 164.17 49.005 164.38 49.075 ;
    RECT 164.17 49.365 164.38 49.435 ;
    RECT 164.17 49.725 164.38 49.795 ;
    RECT 164.63 49.005 164.84 49.075 ;
    RECT 164.63 49.365 164.84 49.435 ;
    RECT 164.63 49.725 164.84 49.795 ;
    RECT 1.49 49.005 1.7 49.075 ;
    RECT 1.49 49.365 1.7 49.435 ;
    RECT 1.49 49.725 1.7 49.795 ;
    RECT 1.95 49.005 2.16 49.075 ;
    RECT 1.95 49.365 2.16 49.435 ;
    RECT 1.95 49.725 2.16 49.795 ;
    RECT 160.85 49.005 161.06 49.075 ;
    RECT 160.85 49.365 161.06 49.435 ;
    RECT 160.85 49.725 161.06 49.795 ;
    RECT 161.31 49.005 161.52 49.075 ;
    RECT 161.31 49.365 161.52 49.435 ;
    RECT 161.31 49.725 161.52 49.795 ;
    RECT 157.53 49.005 157.74 49.075 ;
    RECT 157.53 49.365 157.74 49.435 ;
    RECT 157.53 49.725 157.74 49.795 ;
    RECT 157.99 49.005 158.2 49.075 ;
    RECT 157.99 49.365 158.2 49.435 ;
    RECT 157.99 49.725 158.2 49.795 ;
    RECT 154.21 49.005 154.42 49.075 ;
    RECT 154.21 49.365 154.42 49.435 ;
    RECT 154.21 49.725 154.42 49.795 ;
    RECT 154.67 49.005 154.88 49.075 ;
    RECT 154.67 49.365 154.88 49.435 ;
    RECT 154.67 49.725 154.88 49.795 ;
    RECT 150.89 49.005 151.1 49.075 ;
    RECT 150.89 49.365 151.1 49.435 ;
    RECT 150.89 49.725 151.1 49.795 ;
    RECT 151.35 49.005 151.56 49.075 ;
    RECT 151.35 49.365 151.56 49.435 ;
    RECT 151.35 49.725 151.56 49.795 ;
    RECT 147.57 49.005 147.78 49.075 ;
    RECT 147.57 49.365 147.78 49.435 ;
    RECT 147.57 49.725 147.78 49.795 ;
    RECT 148.03 49.005 148.24 49.075 ;
    RECT 148.03 49.365 148.24 49.435 ;
    RECT 148.03 49.725 148.24 49.795 ;
    RECT 144.25 49.005 144.46 49.075 ;
    RECT 144.25 49.365 144.46 49.435 ;
    RECT 144.25 49.725 144.46 49.795 ;
    RECT 144.71 49.005 144.92 49.075 ;
    RECT 144.71 49.365 144.92 49.435 ;
    RECT 144.71 49.725 144.92 49.795 ;
    RECT 140.93 49.005 141.14 49.075 ;
    RECT 140.93 49.365 141.14 49.435 ;
    RECT 140.93 49.725 141.14 49.795 ;
    RECT 141.39 49.005 141.6 49.075 ;
    RECT 141.39 49.365 141.6 49.435 ;
    RECT 141.39 49.725 141.6 49.795 ;
    RECT 137.61 49.005 137.82 49.075 ;
    RECT 137.61 49.365 137.82 49.435 ;
    RECT 137.61 49.725 137.82 49.795 ;
    RECT 138.07 49.005 138.28 49.075 ;
    RECT 138.07 49.365 138.28 49.435 ;
    RECT 138.07 49.725 138.28 49.795 ;
    RECT 134.29 49.005 134.5 49.075 ;
    RECT 134.29 49.365 134.5 49.435 ;
    RECT 134.29 49.725 134.5 49.795 ;
    RECT 134.75 49.005 134.96 49.075 ;
    RECT 134.75 49.365 134.96 49.435 ;
    RECT 134.75 49.725 134.96 49.795 ;
    RECT 64.57 49.005 64.78 49.075 ;
    RECT 64.57 49.365 64.78 49.435 ;
    RECT 64.57 49.725 64.78 49.795 ;
    RECT 65.03 49.005 65.24 49.075 ;
    RECT 65.03 49.365 65.24 49.435 ;
    RECT 65.03 49.725 65.24 49.795 ;
    RECT 61.25 48.285 61.46 48.355 ;
    RECT 61.25 48.645 61.46 48.715 ;
    RECT 61.25 49.005 61.46 49.075 ;
    RECT 61.71 48.285 61.92 48.355 ;
    RECT 61.71 48.645 61.92 48.715 ;
    RECT 61.71 49.005 61.92 49.075 ;
    RECT 57.93 48.285 58.14 48.355 ;
    RECT 57.93 48.645 58.14 48.715 ;
    RECT 57.93 49.005 58.14 49.075 ;
    RECT 58.39 48.285 58.6 48.355 ;
    RECT 58.39 48.645 58.6 48.715 ;
    RECT 58.39 49.005 58.6 49.075 ;
    RECT 54.61 48.285 54.82 48.355 ;
    RECT 54.61 48.645 54.82 48.715 ;
    RECT 54.61 49.005 54.82 49.075 ;
    RECT 55.07 48.285 55.28 48.355 ;
    RECT 55.07 48.645 55.28 48.715 ;
    RECT 55.07 49.005 55.28 49.075 ;
    RECT 51.29 48.285 51.5 48.355 ;
    RECT 51.29 48.645 51.5 48.715 ;
    RECT 51.29 49.005 51.5 49.075 ;
    RECT 51.75 48.285 51.96 48.355 ;
    RECT 51.75 48.645 51.96 48.715 ;
    RECT 51.75 49.005 51.96 49.075 ;
    RECT 47.97 48.285 48.18 48.355 ;
    RECT 47.97 48.645 48.18 48.715 ;
    RECT 47.97 49.005 48.18 49.075 ;
    RECT 48.43 48.285 48.64 48.355 ;
    RECT 48.43 48.645 48.64 48.715 ;
    RECT 48.43 49.005 48.64 49.075 ;
    RECT 44.65 48.285 44.86 48.355 ;
    RECT 44.65 48.645 44.86 48.715 ;
    RECT 44.65 49.005 44.86 49.075 ;
    RECT 45.11 48.285 45.32 48.355 ;
    RECT 45.11 48.645 45.32 48.715 ;
    RECT 45.11 49.005 45.32 49.075 ;
    RECT 41.33 48.285 41.54 48.355 ;
    RECT 41.33 48.645 41.54 48.715 ;
    RECT 41.33 49.005 41.54 49.075 ;
    RECT 41.79 48.285 42.0 48.355 ;
    RECT 41.79 48.645 42.0 48.715 ;
    RECT 41.79 49.005 42.0 49.075 ;
    RECT 38.01 48.285 38.22 48.355 ;
    RECT 38.01 48.645 38.22 48.715 ;
    RECT 38.01 49.005 38.22 49.075 ;
    RECT 38.47 48.285 38.68 48.355 ;
    RECT 38.47 48.645 38.68 48.715 ;
    RECT 38.47 49.005 38.68 49.075 ;
    RECT 34.69 48.285 34.9 48.355 ;
    RECT 34.69 48.645 34.9 48.715 ;
    RECT 34.69 49.005 34.9 49.075 ;
    RECT 35.15 48.285 35.36 48.355 ;
    RECT 35.15 48.645 35.36 48.715 ;
    RECT 35.15 49.005 35.36 49.075 ;
    RECT 173.945 48.645 174.015 48.715 ;
    RECT 130.97 48.285 131.18 48.355 ;
    RECT 130.97 48.645 131.18 48.715 ;
    RECT 130.97 49.005 131.18 49.075 ;
    RECT 131.43 48.285 131.64 48.355 ;
    RECT 131.43 48.645 131.64 48.715 ;
    RECT 131.43 49.005 131.64 49.075 ;
    RECT 127.65 48.285 127.86 48.355 ;
    RECT 127.65 48.645 127.86 48.715 ;
    RECT 127.65 49.005 127.86 49.075 ;
    RECT 128.11 48.285 128.32 48.355 ;
    RECT 128.11 48.645 128.32 48.715 ;
    RECT 128.11 49.005 128.32 49.075 ;
    RECT 124.33 48.285 124.54 48.355 ;
    RECT 124.33 48.645 124.54 48.715 ;
    RECT 124.33 49.005 124.54 49.075 ;
    RECT 124.79 48.285 125.0 48.355 ;
    RECT 124.79 48.645 125.0 48.715 ;
    RECT 124.79 49.005 125.0 49.075 ;
    RECT 121.01 48.285 121.22 48.355 ;
    RECT 121.01 48.645 121.22 48.715 ;
    RECT 121.01 49.005 121.22 49.075 ;
    RECT 121.47 48.285 121.68 48.355 ;
    RECT 121.47 48.645 121.68 48.715 ;
    RECT 121.47 49.005 121.68 49.075 ;
    RECT 117.69 48.285 117.9 48.355 ;
    RECT 117.69 48.645 117.9 48.715 ;
    RECT 117.69 49.005 117.9 49.075 ;
    RECT 118.15 48.285 118.36 48.355 ;
    RECT 118.15 48.645 118.36 48.715 ;
    RECT 118.15 49.005 118.36 49.075 ;
    RECT 114.37 48.285 114.58 48.355 ;
    RECT 114.37 48.645 114.58 48.715 ;
    RECT 114.37 49.005 114.58 49.075 ;
    RECT 114.83 48.285 115.04 48.355 ;
    RECT 114.83 48.645 115.04 48.715 ;
    RECT 114.83 49.005 115.04 49.075 ;
    RECT 111.05 48.285 111.26 48.355 ;
    RECT 111.05 48.645 111.26 48.715 ;
    RECT 111.05 49.005 111.26 49.075 ;
    RECT 111.51 48.285 111.72 48.355 ;
    RECT 111.51 48.645 111.72 48.715 ;
    RECT 111.51 49.005 111.72 49.075 ;
    RECT 107.73 48.285 107.94 48.355 ;
    RECT 107.73 48.645 107.94 48.715 ;
    RECT 107.73 49.005 107.94 49.075 ;
    RECT 108.19 48.285 108.4 48.355 ;
    RECT 108.19 48.645 108.4 48.715 ;
    RECT 108.19 49.005 108.4 49.075 ;
    RECT 104.41 48.285 104.62 48.355 ;
    RECT 104.41 48.645 104.62 48.715 ;
    RECT 104.41 49.005 104.62 49.075 ;
    RECT 104.87 48.285 105.08 48.355 ;
    RECT 104.87 48.645 105.08 48.715 ;
    RECT 104.87 49.005 105.08 49.075 ;
    RECT 101.09 48.285 101.3 48.355 ;
    RECT 101.09 48.645 101.3 48.715 ;
    RECT 101.09 49.005 101.3 49.075 ;
    RECT 101.55 48.285 101.76 48.355 ;
    RECT 101.55 48.645 101.76 48.715 ;
    RECT 101.55 49.005 101.76 49.075 ;
    RECT 0.4 48.645 0.47 48.715 ;
    RECT 170.81 48.285 171.02 48.355 ;
    RECT 170.81 48.645 171.02 48.715 ;
    RECT 170.81 49.005 171.02 49.075 ;
    RECT 171.27 48.285 171.48 48.355 ;
    RECT 171.27 48.645 171.48 48.715 ;
    RECT 171.27 49.005 171.48 49.075 ;
    RECT 167.49 48.285 167.7 48.355 ;
    RECT 167.49 48.645 167.7 48.715 ;
    RECT 167.49 49.005 167.7 49.075 ;
    RECT 167.95 48.285 168.16 48.355 ;
    RECT 167.95 48.645 168.16 48.715 ;
    RECT 167.95 49.005 168.16 49.075 ;
    RECT 97.77 48.285 97.98 48.355 ;
    RECT 97.77 48.645 97.98 48.715 ;
    RECT 97.77 49.005 97.98 49.075 ;
    RECT 98.23 48.285 98.44 48.355 ;
    RECT 98.23 48.645 98.44 48.715 ;
    RECT 98.23 49.005 98.44 49.075 ;
    RECT 94.45 48.285 94.66 48.355 ;
    RECT 94.45 48.645 94.66 48.715 ;
    RECT 94.45 49.005 94.66 49.075 ;
    RECT 94.91 48.285 95.12 48.355 ;
    RECT 94.91 48.645 95.12 48.715 ;
    RECT 94.91 49.005 95.12 49.075 ;
    RECT 91.13 48.285 91.34 48.355 ;
    RECT 91.13 48.645 91.34 48.715 ;
    RECT 91.13 49.005 91.34 49.075 ;
    RECT 91.59 48.285 91.8 48.355 ;
    RECT 91.59 48.645 91.8 48.715 ;
    RECT 91.59 49.005 91.8 49.075 ;
    RECT 87.81 48.285 88.02 48.355 ;
    RECT 87.81 48.645 88.02 48.715 ;
    RECT 87.81 49.005 88.02 49.075 ;
    RECT 88.27 48.285 88.48 48.355 ;
    RECT 88.27 48.645 88.48 48.715 ;
    RECT 88.27 49.005 88.48 49.075 ;
    RECT 84.49 48.285 84.7 48.355 ;
    RECT 84.49 48.645 84.7 48.715 ;
    RECT 84.49 49.005 84.7 49.075 ;
    RECT 84.95 48.285 85.16 48.355 ;
    RECT 84.95 48.645 85.16 48.715 ;
    RECT 84.95 49.005 85.16 49.075 ;
    RECT 81.17 48.285 81.38 48.355 ;
    RECT 81.17 48.645 81.38 48.715 ;
    RECT 81.17 49.005 81.38 49.075 ;
    RECT 81.63 48.285 81.84 48.355 ;
    RECT 81.63 48.645 81.84 48.715 ;
    RECT 81.63 49.005 81.84 49.075 ;
    RECT 77.85 48.285 78.06 48.355 ;
    RECT 77.85 48.645 78.06 48.715 ;
    RECT 77.85 49.005 78.06 49.075 ;
    RECT 78.31 48.285 78.52 48.355 ;
    RECT 78.31 48.645 78.52 48.715 ;
    RECT 78.31 49.005 78.52 49.075 ;
    RECT 74.53 48.285 74.74 48.355 ;
    RECT 74.53 48.645 74.74 48.715 ;
    RECT 74.53 49.005 74.74 49.075 ;
    RECT 74.99 48.285 75.2 48.355 ;
    RECT 74.99 48.645 75.2 48.715 ;
    RECT 74.99 49.005 75.2 49.075 ;
    RECT 71.21 48.285 71.42 48.355 ;
    RECT 71.21 48.645 71.42 48.715 ;
    RECT 71.21 49.005 71.42 49.075 ;
    RECT 71.67 48.285 71.88 48.355 ;
    RECT 71.67 48.645 71.88 48.715 ;
    RECT 71.67 49.005 71.88 49.075 ;
    RECT 31.37 48.285 31.58 48.355 ;
    RECT 31.37 48.645 31.58 48.715 ;
    RECT 31.37 49.005 31.58 49.075 ;
    RECT 31.83 48.285 32.04 48.355 ;
    RECT 31.83 48.645 32.04 48.715 ;
    RECT 31.83 49.005 32.04 49.075 ;
    RECT 67.89 48.285 68.1 48.355 ;
    RECT 67.89 48.645 68.1 48.715 ;
    RECT 67.89 49.005 68.1 49.075 ;
    RECT 68.35 48.285 68.56 48.355 ;
    RECT 68.35 48.645 68.56 48.715 ;
    RECT 68.35 49.005 68.56 49.075 ;
    RECT 28.05 48.285 28.26 48.355 ;
    RECT 28.05 48.645 28.26 48.715 ;
    RECT 28.05 49.005 28.26 49.075 ;
    RECT 28.51 48.285 28.72 48.355 ;
    RECT 28.51 48.645 28.72 48.715 ;
    RECT 28.51 49.005 28.72 49.075 ;
    RECT 24.73 48.285 24.94 48.355 ;
    RECT 24.73 48.645 24.94 48.715 ;
    RECT 24.73 49.005 24.94 49.075 ;
    RECT 25.19 48.285 25.4 48.355 ;
    RECT 25.19 48.645 25.4 48.715 ;
    RECT 25.19 49.005 25.4 49.075 ;
    RECT 21.41 48.285 21.62 48.355 ;
    RECT 21.41 48.645 21.62 48.715 ;
    RECT 21.41 49.005 21.62 49.075 ;
    RECT 21.87 48.285 22.08 48.355 ;
    RECT 21.87 48.645 22.08 48.715 ;
    RECT 21.87 49.005 22.08 49.075 ;
    RECT 18.09 48.285 18.3 48.355 ;
    RECT 18.09 48.645 18.3 48.715 ;
    RECT 18.09 49.005 18.3 49.075 ;
    RECT 18.55 48.285 18.76 48.355 ;
    RECT 18.55 48.645 18.76 48.715 ;
    RECT 18.55 49.005 18.76 49.075 ;
    RECT 14.77 48.285 14.98 48.355 ;
    RECT 14.77 48.645 14.98 48.715 ;
    RECT 14.77 49.005 14.98 49.075 ;
    RECT 15.23 48.285 15.44 48.355 ;
    RECT 15.23 48.645 15.44 48.715 ;
    RECT 15.23 49.005 15.44 49.075 ;
    RECT 11.45 48.285 11.66 48.355 ;
    RECT 11.45 48.645 11.66 48.715 ;
    RECT 11.45 49.005 11.66 49.075 ;
    RECT 11.91 48.285 12.12 48.355 ;
    RECT 11.91 48.645 12.12 48.715 ;
    RECT 11.91 49.005 12.12 49.075 ;
    RECT 8.13 48.285 8.34 48.355 ;
    RECT 8.13 48.645 8.34 48.715 ;
    RECT 8.13 49.005 8.34 49.075 ;
    RECT 8.59 48.285 8.8 48.355 ;
    RECT 8.59 48.645 8.8 48.715 ;
    RECT 8.59 49.005 8.8 49.075 ;
    RECT 4.81 48.285 5.02 48.355 ;
    RECT 4.81 48.645 5.02 48.715 ;
    RECT 4.81 49.005 5.02 49.075 ;
    RECT 5.27 48.285 5.48 48.355 ;
    RECT 5.27 48.645 5.48 48.715 ;
    RECT 5.27 49.005 5.48 49.075 ;
    RECT 164.17 48.285 164.38 48.355 ;
    RECT 164.17 48.645 164.38 48.715 ;
    RECT 164.17 49.005 164.38 49.075 ;
    RECT 164.63 48.285 164.84 48.355 ;
    RECT 164.63 48.645 164.84 48.715 ;
    RECT 164.63 49.005 164.84 49.075 ;
    RECT 1.49 48.285 1.7 48.355 ;
    RECT 1.49 48.645 1.7 48.715 ;
    RECT 1.49 49.005 1.7 49.075 ;
    RECT 1.95 48.285 2.16 48.355 ;
    RECT 1.95 48.645 2.16 48.715 ;
    RECT 1.95 49.005 2.16 49.075 ;
    RECT 160.85 48.285 161.06 48.355 ;
    RECT 160.85 48.645 161.06 48.715 ;
    RECT 160.85 49.005 161.06 49.075 ;
    RECT 161.31 48.285 161.52 48.355 ;
    RECT 161.31 48.645 161.52 48.715 ;
    RECT 161.31 49.005 161.52 49.075 ;
    RECT 157.53 48.285 157.74 48.355 ;
    RECT 157.53 48.645 157.74 48.715 ;
    RECT 157.53 49.005 157.74 49.075 ;
    RECT 157.99 48.285 158.2 48.355 ;
    RECT 157.99 48.645 158.2 48.715 ;
    RECT 157.99 49.005 158.2 49.075 ;
    RECT 154.21 48.285 154.42 48.355 ;
    RECT 154.21 48.645 154.42 48.715 ;
    RECT 154.21 49.005 154.42 49.075 ;
    RECT 154.67 48.285 154.88 48.355 ;
    RECT 154.67 48.645 154.88 48.715 ;
    RECT 154.67 49.005 154.88 49.075 ;
    RECT 150.89 48.285 151.1 48.355 ;
    RECT 150.89 48.645 151.1 48.715 ;
    RECT 150.89 49.005 151.1 49.075 ;
    RECT 151.35 48.285 151.56 48.355 ;
    RECT 151.35 48.645 151.56 48.715 ;
    RECT 151.35 49.005 151.56 49.075 ;
    RECT 147.57 48.285 147.78 48.355 ;
    RECT 147.57 48.645 147.78 48.715 ;
    RECT 147.57 49.005 147.78 49.075 ;
    RECT 148.03 48.285 148.24 48.355 ;
    RECT 148.03 48.645 148.24 48.715 ;
    RECT 148.03 49.005 148.24 49.075 ;
    RECT 144.25 48.285 144.46 48.355 ;
    RECT 144.25 48.645 144.46 48.715 ;
    RECT 144.25 49.005 144.46 49.075 ;
    RECT 144.71 48.285 144.92 48.355 ;
    RECT 144.71 48.645 144.92 48.715 ;
    RECT 144.71 49.005 144.92 49.075 ;
    RECT 140.93 48.285 141.14 48.355 ;
    RECT 140.93 48.645 141.14 48.715 ;
    RECT 140.93 49.005 141.14 49.075 ;
    RECT 141.39 48.285 141.6 48.355 ;
    RECT 141.39 48.645 141.6 48.715 ;
    RECT 141.39 49.005 141.6 49.075 ;
    RECT 137.61 48.285 137.82 48.355 ;
    RECT 137.61 48.645 137.82 48.715 ;
    RECT 137.61 49.005 137.82 49.075 ;
    RECT 138.07 48.285 138.28 48.355 ;
    RECT 138.07 48.645 138.28 48.715 ;
    RECT 138.07 49.005 138.28 49.075 ;
    RECT 134.29 48.285 134.5 48.355 ;
    RECT 134.29 48.645 134.5 48.715 ;
    RECT 134.29 49.005 134.5 49.075 ;
    RECT 134.75 48.285 134.96 48.355 ;
    RECT 134.75 48.645 134.96 48.715 ;
    RECT 134.75 49.005 134.96 49.075 ;
    RECT 64.57 48.285 64.78 48.355 ;
    RECT 64.57 48.645 64.78 48.715 ;
    RECT 64.57 49.005 64.78 49.075 ;
    RECT 65.03 48.285 65.24 48.355 ;
    RECT 65.03 48.645 65.24 48.715 ;
    RECT 65.03 49.005 65.24 49.075 ;
    RECT 61.25 47.565 61.46 47.635 ;
    RECT 61.25 47.925 61.46 47.995 ;
    RECT 61.25 48.285 61.46 48.355 ;
    RECT 61.71 47.565 61.92 47.635 ;
    RECT 61.71 47.925 61.92 47.995 ;
    RECT 61.71 48.285 61.92 48.355 ;
    RECT 57.93 47.565 58.14 47.635 ;
    RECT 57.93 47.925 58.14 47.995 ;
    RECT 57.93 48.285 58.14 48.355 ;
    RECT 58.39 47.565 58.6 47.635 ;
    RECT 58.39 47.925 58.6 47.995 ;
    RECT 58.39 48.285 58.6 48.355 ;
    RECT 54.61 47.565 54.82 47.635 ;
    RECT 54.61 47.925 54.82 47.995 ;
    RECT 54.61 48.285 54.82 48.355 ;
    RECT 55.07 47.565 55.28 47.635 ;
    RECT 55.07 47.925 55.28 47.995 ;
    RECT 55.07 48.285 55.28 48.355 ;
    RECT 51.29 47.565 51.5 47.635 ;
    RECT 51.29 47.925 51.5 47.995 ;
    RECT 51.29 48.285 51.5 48.355 ;
    RECT 51.75 47.565 51.96 47.635 ;
    RECT 51.75 47.925 51.96 47.995 ;
    RECT 51.75 48.285 51.96 48.355 ;
    RECT 47.97 47.565 48.18 47.635 ;
    RECT 47.97 47.925 48.18 47.995 ;
    RECT 47.97 48.285 48.18 48.355 ;
    RECT 48.43 47.565 48.64 47.635 ;
    RECT 48.43 47.925 48.64 47.995 ;
    RECT 48.43 48.285 48.64 48.355 ;
    RECT 44.65 47.565 44.86 47.635 ;
    RECT 44.65 47.925 44.86 47.995 ;
    RECT 44.65 48.285 44.86 48.355 ;
    RECT 45.11 47.565 45.32 47.635 ;
    RECT 45.11 47.925 45.32 47.995 ;
    RECT 45.11 48.285 45.32 48.355 ;
    RECT 41.33 47.565 41.54 47.635 ;
    RECT 41.33 47.925 41.54 47.995 ;
    RECT 41.33 48.285 41.54 48.355 ;
    RECT 41.79 47.565 42.0 47.635 ;
    RECT 41.79 47.925 42.0 47.995 ;
    RECT 41.79 48.285 42.0 48.355 ;
    RECT 38.01 47.565 38.22 47.635 ;
    RECT 38.01 47.925 38.22 47.995 ;
    RECT 38.01 48.285 38.22 48.355 ;
    RECT 38.47 47.565 38.68 47.635 ;
    RECT 38.47 47.925 38.68 47.995 ;
    RECT 38.47 48.285 38.68 48.355 ;
    RECT 34.69 47.565 34.9 47.635 ;
    RECT 34.69 47.925 34.9 47.995 ;
    RECT 34.69 48.285 34.9 48.355 ;
    RECT 35.15 47.565 35.36 47.635 ;
    RECT 35.15 47.925 35.36 47.995 ;
    RECT 35.15 48.285 35.36 48.355 ;
    RECT 173.945 47.925 174.015 47.995 ;
    RECT 130.97 47.565 131.18 47.635 ;
    RECT 130.97 47.925 131.18 47.995 ;
    RECT 130.97 48.285 131.18 48.355 ;
    RECT 131.43 47.565 131.64 47.635 ;
    RECT 131.43 47.925 131.64 47.995 ;
    RECT 131.43 48.285 131.64 48.355 ;
    RECT 127.65 47.565 127.86 47.635 ;
    RECT 127.65 47.925 127.86 47.995 ;
    RECT 127.65 48.285 127.86 48.355 ;
    RECT 128.11 47.565 128.32 47.635 ;
    RECT 128.11 47.925 128.32 47.995 ;
    RECT 128.11 48.285 128.32 48.355 ;
    RECT 124.33 47.565 124.54 47.635 ;
    RECT 124.33 47.925 124.54 47.995 ;
    RECT 124.33 48.285 124.54 48.355 ;
    RECT 124.79 47.565 125.0 47.635 ;
    RECT 124.79 47.925 125.0 47.995 ;
    RECT 124.79 48.285 125.0 48.355 ;
    RECT 121.01 47.565 121.22 47.635 ;
    RECT 121.01 47.925 121.22 47.995 ;
    RECT 121.01 48.285 121.22 48.355 ;
    RECT 121.47 47.565 121.68 47.635 ;
    RECT 121.47 47.925 121.68 47.995 ;
    RECT 121.47 48.285 121.68 48.355 ;
    RECT 117.69 47.565 117.9 47.635 ;
    RECT 117.69 47.925 117.9 47.995 ;
    RECT 117.69 48.285 117.9 48.355 ;
    RECT 118.15 47.565 118.36 47.635 ;
    RECT 118.15 47.925 118.36 47.995 ;
    RECT 118.15 48.285 118.36 48.355 ;
    RECT 114.37 47.565 114.58 47.635 ;
    RECT 114.37 47.925 114.58 47.995 ;
    RECT 114.37 48.285 114.58 48.355 ;
    RECT 114.83 47.565 115.04 47.635 ;
    RECT 114.83 47.925 115.04 47.995 ;
    RECT 114.83 48.285 115.04 48.355 ;
    RECT 111.05 47.565 111.26 47.635 ;
    RECT 111.05 47.925 111.26 47.995 ;
    RECT 111.05 48.285 111.26 48.355 ;
    RECT 111.51 47.565 111.72 47.635 ;
    RECT 111.51 47.925 111.72 47.995 ;
    RECT 111.51 48.285 111.72 48.355 ;
    RECT 107.73 47.565 107.94 47.635 ;
    RECT 107.73 47.925 107.94 47.995 ;
    RECT 107.73 48.285 107.94 48.355 ;
    RECT 108.19 47.565 108.4 47.635 ;
    RECT 108.19 47.925 108.4 47.995 ;
    RECT 108.19 48.285 108.4 48.355 ;
    RECT 104.41 47.565 104.62 47.635 ;
    RECT 104.41 47.925 104.62 47.995 ;
    RECT 104.41 48.285 104.62 48.355 ;
    RECT 104.87 47.565 105.08 47.635 ;
    RECT 104.87 47.925 105.08 47.995 ;
    RECT 104.87 48.285 105.08 48.355 ;
    RECT 101.09 47.565 101.3 47.635 ;
    RECT 101.09 47.925 101.3 47.995 ;
    RECT 101.09 48.285 101.3 48.355 ;
    RECT 101.55 47.565 101.76 47.635 ;
    RECT 101.55 47.925 101.76 47.995 ;
    RECT 101.55 48.285 101.76 48.355 ;
    RECT 0.4 47.925 0.47 47.995 ;
    RECT 170.81 47.565 171.02 47.635 ;
    RECT 170.81 47.925 171.02 47.995 ;
    RECT 170.81 48.285 171.02 48.355 ;
    RECT 171.27 47.565 171.48 47.635 ;
    RECT 171.27 47.925 171.48 47.995 ;
    RECT 171.27 48.285 171.48 48.355 ;
    RECT 167.49 47.565 167.7 47.635 ;
    RECT 167.49 47.925 167.7 47.995 ;
    RECT 167.49 48.285 167.7 48.355 ;
    RECT 167.95 47.565 168.16 47.635 ;
    RECT 167.95 47.925 168.16 47.995 ;
    RECT 167.95 48.285 168.16 48.355 ;
    RECT 97.77 47.565 97.98 47.635 ;
    RECT 97.77 47.925 97.98 47.995 ;
    RECT 97.77 48.285 97.98 48.355 ;
    RECT 98.23 47.565 98.44 47.635 ;
    RECT 98.23 47.925 98.44 47.995 ;
    RECT 98.23 48.285 98.44 48.355 ;
    RECT 94.45 47.565 94.66 47.635 ;
    RECT 94.45 47.925 94.66 47.995 ;
    RECT 94.45 48.285 94.66 48.355 ;
    RECT 94.91 47.565 95.12 47.635 ;
    RECT 94.91 47.925 95.12 47.995 ;
    RECT 94.91 48.285 95.12 48.355 ;
    RECT 91.13 47.565 91.34 47.635 ;
    RECT 91.13 47.925 91.34 47.995 ;
    RECT 91.13 48.285 91.34 48.355 ;
    RECT 91.59 47.565 91.8 47.635 ;
    RECT 91.59 47.925 91.8 47.995 ;
    RECT 91.59 48.285 91.8 48.355 ;
    RECT 87.81 47.565 88.02 47.635 ;
    RECT 87.81 47.925 88.02 47.995 ;
    RECT 87.81 48.285 88.02 48.355 ;
    RECT 88.27 47.565 88.48 47.635 ;
    RECT 88.27 47.925 88.48 47.995 ;
    RECT 88.27 48.285 88.48 48.355 ;
    RECT 84.49 47.565 84.7 47.635 ;
    RECT 84.49 47.925 84.7 47.995 ;
    RECT 84.49 48.285 84.7 48.355 ;
    RECT 84.95 47.565 85.16 47.635 ;
    RECT 84.95 47.925 85.16 47.995 ;
    RECT 84.95 48.285 85.16 48.355 ;
    RECT 81.17 47.565 81.38 47.635 ;
    RECT 81.17 47.925 81.38 47.995 ;
    RECT 81.17 48.285 81.38 48.355 ;
    RECT 81.63 47.565 81.84 47.635 ;
    RECT 81.63 47.925 81.84 47.995 ;
    RECT 81.63 48.285 81.84 48.355 ;
    RECT 77.85 47.565 78.06 47.635 ;
    RECT 77.85 47.925 78.06 47.995 ;
    RECT 77.85 48.285 78.06 48.355 ;
    RECT 78.31 47.565 78.52 47.635 ;
    RECT 78.31 47.925 78.52 47.995 ;
    RECT 78.31 48.285 78.52 48.355 ;
    RECT 74.53 47.565 74.74 47.635 ;
    RECT 74.53 47.925 74.74 47.995 ;
    RECT 74.53 48.285 74.74 48.355 ;
    RECT 74.99 47.565 75.2 47.635 ;
    RECT 74.99 47.925 75.2 47.995 ;
    RECT 74.99 48.285 75.2 48.355 ;
    RECT 71.21 47.565 71.42 47.635 ;
    RECT 71.21 47.925 71.42 47.995 ;
    RECT 71.21 48.285 71.42 48.355 ;
    RECT 71.67 47.565 71.88 47.635 ;
    RECT 71.67 47.925 71.88 47.995 ;
    RECT 71.67 48.285 71.88 48.355 ;
    RECT 31.37 47.565 31.58 47.635 ;
    RECT 31.37 47.925 31.58 47.995 ;
    RECT 31.37 48.285 31.58 48.355 ;
    RECT 31.83 47.565 32.04 47.635 ;
    RECT 31.83 47.925 32.04 47.995 ;
    RECT 31.83 48.285 32.04 48.355 ;
    RECT 67.89 47.565 68.1 47.635 ;
    RECT 67.89 47.925 68.1 47.995 ;
    RECT 67.89 48.285 68.1 48.355 ;
    RECT 68.35 47.565 68.56 47.635 ;
    RECT 68.35 47.925 68.56 47.995 ;
    RECT 68.35 48.285 68.56 48.355 ;
    RECT 28.05 47.565 28.26 47.635 ;
    RECT 28.05 47.925 28.26 47.995 ;
    RECT 28.05 48.285 28.26 48.355 ;
    RECT 28.51 47.565 28.72 47.635 ;
    RECT 28.51 47.925 28.72 47.995 ;
    RECT 28.51 48.285 28.72 48.355 ;
    RECT 24.73 47.565 24.94 47.635 ;
    RECT 24.73 47.925 24.94 47.995 ;
    RECT 24.73 48.285 24.94 48.355 ;
    RECT 25.19 47.565 25.4 47.635 ;
    RECT 25.19 47.925 25.4 47.995 ;
    RECT 25.19 48.285 25.4 48.355 ;
    RECT 21.41 47.565 21.62 47.635 ;
    RECT 21.41 47.925 21.62 47.995 ;
    RECT 21.41 48.285 21.62 48.355 ;
    RECT 21.87 47.565 22.08 47.635 ;
    RECT 21.87 47.925 22.08 47.995 ;
    RECT 21.87 48.285 22.08 48.355 ;
    RECT 18.09 47.565 18.3 47.635 ;
    RECT 18.09 47.925 18.3 47.995 ;
    RECT 18.09 48.285 18.3 48.355 ;
    RECT 18.55 47.565 18.76 47.635 ;
    RECT 18.55 47.925 18.76 47.995 ;
    RECT 18.55 48.285 18.76 48.355 ;
    RECT 14.77 47.565 14.98 47.635 ;
    RECT 14.77 47.925 14.98 47.995 ;
    RECT 14.77 48.285 14.98 48.355 ;
    RECT 15.23 47.565 15.44 47.635 ;
    RECT 15.23 47.925 15.44 47.995 ;
    RECT 15.23 48.285 15.44 48.355 ;
    RECT 11.45 47.565 11.66 47.635 ;
    RECT 11.45 47.925 11.66 47.995 ;
    RECT 11.45 48.285 11.66 48.355 ;
    RECT 11.91 47.565 12.12 47.635 ;
    RECT 11.91 47.925 12.12 47.995 ;
    RECT 11.91 48.285 12.12 48.355 ;
    RECT 8.13 47.565 8.34 47.635 ;
    RECT 8.13 47.925 8.34 47.995 ;
    RECT 8.13 48.285 8.34 48.355 ;
    RECT 8.59 47.565 8.8 47.635 ;
    RECT 8.59 47.925 8.8 47.995 ;
    RECT 8.59 48.285 8.8 48.355 ;
    RECT 4.81 47.565 5.02 47.635 ;
    RECT 4.81 47.925 5.02 47.995 ;
    RECT 4.81 48.285 5.02 48.355 ;
    RECT 5.27 47.565 5.48 47.635 ;
    RECT 5.27 47.925 5.48 47.995 ;
    RECT 5.27 48.285 5.48 48.355 ;
    RECT 164.17 47.565 164.38 47.635 ;
    RECT 164.17 47.925 164.38 47.995 ;
    RECT 164.17 48.285 164.38 48.355 ;
    RECT 164.63 47.565 164.84 47.635 ;
    RECT 164.63 47.925 164.84 47.995 ;
    RECT 164.63 48.285 164.84 48.355 ;
    RECT 1.49 47.565 1.7 47.635 ;
    RECT 1.49 47.925 1.7 47.995 ;
    RECT 1.49 48.285 1.7 48.355 ;
    RECT 1.95 47.565 2.16 47.635 ;
    RECT 1.95 47.925 2.16 47.995 ;
    RECT 1.95 48.285 2.16 48.355 ;
    RECT 160.85 47.565 161.06 47.635 ;
    RECT 160.85 47.925 161.06 47.995 ;
    RECT 160.85 48.285 161.06 48.355 ;
    RECT 161.31 47.565 161.52 47.635 ;
    RECT 161.31 47.925 161.52 47.995 ;
    RECT 161.31 48.285 161.52 48.355 ;
    RECT 157.53 47.565 157.74 47.635 ;
    RECT 157.53 47.925 157.74 47.995 ;
    RECT 157.53 48.285 157.74 48.355 ;
    RECT 157.99 47.565 158.2 47.635 ;
    RECT 157.99 47.925 158.2 47.995 ;
    RECT 157.99 48.285 158.2 48.355 ;
    RECT 154.21 47.565 154.42 47.635 ;
    RECT 154.21 47.925 154.42 47.995 ;
    RECT 154.21 48.285 154.42 48.355 ;
    RECT 154.67 47.565 154.88 47.635 ;
    RECT 154.67 47.925 154.88 47.995 ;
    RECT 154.67 48.285 154.88 48.355 ;
    RECT 150.89 47.565 151.1 47.635 ;
    RECT 150.89 47.925 151.1 47.995 ;
    RECT 150.89 48.285 151.1 48.355 ;
    RECT 151.35 47.565 151.56 47.635 ;
    RECT 151.35 47.925 151.56 47.995 ;
    RECT 151.35 48.285 151.56 48.355 ;
    RECT 147.57 47.565 147.78 47.635 ;
    RECT 147.57 47.925 147.78 47.995 ;
    RECT 147.57 48.285 147.78 48.355 ;
    RECT 148.03 47.565 148.24 47.635 ;
    RECT 148.03 47.925 148.24 47.995 ;
    RECT 148.03 48.285 148.24 48.355 ;
    RECT 144.25 47.565 144.46 47.635 ;
    RECT 144.25 47.925 144.46 47.995 ;
    RECT 144.25 48.285 144.46 48.355 ;
    RECT 144.71 47.565 144.92 47.635 ;
    RECT 144.71 47.925 144.92 47.995 ;
    RECT 144.71 48.285 144.92 48.355 ;
    RECT 140.93 47.565 141.14 47.635 ;
    RECT 140.93 47.925 141.14 47.995 ;
    RECT 140.93 48.285 141.14 48.355 ;
    RECT 141.39 47.565 141.6 47.635 ;
    RECT 141.39 47.925 141.6 47.995 ;
    RECT 141.39 48.285 141.6 48.355 ;
    RECT 137.61 47.565 137.82 47.635 ;
    RECT 137.61 47.925 137.82 47.995 ;
    RECT 137.61 48.285 137.82 48.355 ;
    RECT 138.07 47.565 138.28 47.635 ;
    RECT 138.07 47.925 138.28 47.995 ;
    RECT 138.07 48.285 138.28 48.355 ;
    RECT 134.29 47.565 134.5 47.635 ;
    RECT 134.29 47.925 134.5 47.995 ;
    RECT 134.29 48.285 134.5 48.355 ;
    RECT 134.75 47.565 134.96 47.635 ;
    RECT 134.75 47.925 134.96 47.995 ;
    RECT 134.75 48.285 134.96 48.355 ;
    RECT 64.57 47.565 64.78 47.635 ;
    RECT 64.57 47.925 64.78 47.995 ;
    RECT 64.57 48.285 64.78 48.355 ;
    RECT 65.03 47.565 65.24 47.635 ;
    RECT 65.03 47.925 65.24 47.995 ;
    RECT 65.03 48.285 65.24 48.355 ;
    RECT 61.25 11.565 61.46 11.635 ;
    RECT 61.25 11.925 61.46 11.995 ;
    RECT 61.25 12.285 61.46 12.355 ;
    RECT 61.71 11.565 61.92 11.635 ;
    RECT 61.71 11.925 61.92 11.995 ;
    RECT 61.71 12.285 61.92 12.355 ;
    RECT 57.93 11.565 58.14 11.635 ;
    RECT 57.93 11.925 58.14 11.995 ;
    RECT 57.93 12.285 58.14 12.355 ;
    RECT 58.39 11.565 58.6 11.635 ;
    RECT 58.39 11.925 58.6 11.995 ;
    RECT 58.39 12.285 58.6 12.355 ;
    RECT 54.61 11.565 54.82 11.635 ;
    RECT 54.61 11.925 54.82 11.995 ;
    RECT 54.61 12.285 54.82 12.355 ;
    RECT 55.07 11.565 55.28 11.635 ;
    RECT 55.07 11.925 55.28 11.995 ;
    RECT 55.07 12.285 55.28 12.355 ;
    RECT 51.29 11.565 51.5 11.635 ;
    RECT 51.29 11.925 51.5 11.995 ;
    RECT 51.29 12.285 51.5 12.355 ;
    RECT 51.75 11.565 51.96 11.635 ;
    RECT 51.75 11.925 51.96 11.995 ;
    RECT 51.75 12.285 51.96 12.355 ;
    RECT 47.97 11.565 48.18 11.635 ;
    RECT 47.97 11.925 48.18 11.995 ;
    RECT 47.97 12.285 48.18 12.355 ;
    RECT 48.43 11.565 48.64 11.635 ;
    RECT 48.43 11.925 48.64 11.995 ;
    RECT 48.43 12.285 48.64 12.355 ;
    RECT 44.65 11.565 44.86 11.635 ;
    RECT 44.65 11.925 44.86 11.995 ;
    RECT 44.65 12.285 44.86 12.355 ;
    RECT 45.11 11.565 45.32 11.635 ;
    RECT 45.11 11.925 45.32 11.995 ;
    RECT 45.11 12.285 45.32 12.355 ;
    RECT 41.33 11.565 41.54 11.635 ;
    RECT 41.33 11.925 41.54 11.995 ;
    RECT 41.33 12.285 41.54 12.355 ;
    RECT 41.79 11.565 42.0 11.635 ;
    RECT 41.79 11.925 42.0 11.995 ;
    RECT 41.79 12.285 42.0 12.355 ;
    RECT 38.01 11.565 38.22 11.635 ;
    RECT 38.01 11.925 38.22 11.995 ;
    RECT 38.01 12.285 38.22 12.355 ;
    RECT 38.47 11.565 38.68 11.635 ;
    RECT 38.47 11.925 38.68 11.995 ;
    RECT 38.47 12.285 38.68 12.355 ;
    RECT 34.69 11.565 34.9 11.635 ;
    RECT 34.69 11.925 34.9 11.995 ;
    RECT 34.69 12.285 34.9 12.355 ;
    RECT 35.15 11.565 35.36 11.635 ;
    RECT 35.15 11.925 35.36 11.995 ;
    RECT 35.15 12.285 35.36 12.355 ;
    RECT 130.97 11.565 131.18 11.635 ;
    RECT 130.97 11.925 131.18 11.995 ;
    RECT 130.97 12.285 131.18 12.355 ;
    RECT 131.43 11.565 131.64 11.635 ;
    RECT 131.43 11.925 131.64 11.995 ;
    RECT 131.43 12.285 131.64 12.355 ;
    RECT 127.65 11.565 127.86 11.635 ;
    RECT 127.65 11.925 127.86 11.995 ;
    RECT 127.65 12.285 127.86 12.355 ;
    RECT 128.11 11.565 128.32 11.635 ;
    RECT 128.11 11.925 128.32 11.995 ;
    RECT 128.11 12.285 128.32 12.355 ;
    RECT 124.33 11.565 124.54 11.635 ;
    RECT 124.33 11.925 124.54 11.995 ;
    RECT 124.33 12.285 124.54 12.355 ;
    RECT 124.79 11.565 125.0 11.635 ;
    RECT 124.79 11.925 125.0 11.995 ;
    RECT 124.79 12.285 125.0 12.355 ;
    RECT 121.01 11.565 121.22 11.635 ;
    RECT 121.01 11.925 121.22 11.995 ;
    RECT 121.01 12.285 121.22 12.355 ;
    RECT 121.47 11.565 121.68 11.635 ;
    RECT 121.47 11.925 121.68 11.995 ;
    RECT 121.47 12.285 121.68 12.355 ;
    RECT 117.69 11.565 117.9 11.635 ;
    RECT 117.69 11.925 117.9 11.995 ;
    RECT 117.69 12.285 117.9 12.355 ;
    RECT 118.15 11.565 118.36 11.635 ;
    RECT 118.15 11.925 118.36 11.995 ;
    RECT 118.15 12.285 118.36 12.355 ;
    RECT 114.37 11.565 114.58 11.635 ;
    RECT 114.37 11.925 114.58 11.995 ;
    RECT 114.37 12.285 114.58 12.355 ;
    RECT 114.83 11.565 115.04 11.635 ;
    RECT 114.83 11.925 115.04 11.995 ;
    RECT 114.83 12.285 115.04 12.355 ;
    RECT 111.05 11.565 111.26 11.635 ;
    RECT 111.05 11.925 111.26 11.995 ;
    RECT 111.05 12.285 111.26 12.355 ;
    RECT 111.51 11.565 111.72 11.635 ;
    RECT 111.51 11.925 111.72 11.995 ;
    RECT 111.51 12.285 111.72 12.355 ;
    RECT 107.73 11.565 107.94 11.635 ;
    RECT 107.73 11.925 107.94 11.995 ;
    RECT 107.73 12.285 107.94 12.355 ;
    RECT 108.19 11.565 108.4 11.635 ;
    RECT 108.19 11.925 108.4 11.995 ;
    RECT 108.19 12.285 108.4 12.355 ;
    RECT 104.41 11.565 104.62 11.635 ;
    RECT 104.41 11.925 104.62 11.995 ;
    RECT 104.41 12.285 104.62 12.355 ;
    RECT 104.87 11.565 105.08 11.635 ;
    RECT 104.87 11.925 105.08 11.995 ;
    RECT 104.87 12.285 105.08 12.355 ;
    RECT 101.09 11.565 101.3 11.635 ;
    RECT 101.09 11.925 101.3 11.995 ;
    RECT 101.09 12.285 101.3 12.355 ;
    RECT 101.55 11.565 101.76 11.635 ;
    RECT 101.55 11.925 101.76 11.995 ;
    RECT 101.55 12.285 101.76 12.355 ;
    RECT 173.945 11.925 174.015 11.995 ;
    RECT 167.49 11.565 167.7 11.635 ;
    RECT 167.49 11.925 167.7 11.995 ;
    RECT 167.49 12.285 167.7 12.355 ;
    RECT 167.95 11.565 168.16 11.635 ;
    RECT 167.95 11.925 168.16 11.995 ;
    RECT 167.95 12.285 168.16 12.355 ;
    RECT 97.77 11.565 97.98 11.635 ;
    RECT 97.77 11.925 97.98 11.995 ;
    RECT 97.77 12.285 97.98 12.355 ;
    RECT 98.23 11.565 98.44 11.635 ;
    RECT 98.23 11.925 98.44 11.995 ;
    RECT 98.23 12.285 98.44 12.355 ;
    RECT 94.45 11.565 94.66 11.635 ;
    RECT 94.45 11.925 94.66 11.995 ;
    RECT 94.45 12.285 94.66 12.355 ;
    RECT 94.91 11.565 95.12 11.635 ;
    RECT 94.91 11.925 95.12 11.995 ;
    RECT 94.91 12.285 95.12 12.355 ;
    RECT 91.13 11.565 91.34 11.635 ;
    RECT 91.13 11.925 91.34 11.995 ;
    RECT 91.13 12.285 91.34 12.355 ;
    RECT 91.59 11.565 91.8 11.635 ;
    RECT 91.59 11.925 91.8 11.995 ;
    RECT 91.59 12.285 91.8 12.355 ;
    RECT 87.81 11.565 88.02 11.635 ;
    RECT 87.81 11.925 88.02 11.995 ;
    RECT 87.81 12.285 88.02 12.355 ;
    RECT 88.27 11.565 88.48 11.635 ;
    RECT 88.27 11.925 88.48 11.995 ;
    RECT 88.27 12.285 88.48 12.355 ;
    RECT 84.49 11.565 84.7 11.635 ;
    RECT 84.49 11.925 84.7 11.995 ;
    RECT 84.49 12.285 84.7 12.355 ;
    RECT 84.95 11.565 85.16 11.635 ;
    RECT 84.95 11.925 85.16 11.995 ;
    RECT 84.95 12.285 85.16 12.355 ;
    RECT 81.17 11.565 81.38 11.635 ;
    RECT 81.17 11.925 81.38 11.995 ;
    RECT 81.17 12.285 81.38 12.355 ;
    RECT 81.63 11.565 81.84 11.635 ;
    RECT 81.63 11.925 81.84 11.995 ;
    RECT 81.63 12.285 81.84 12.355 ;
    RECT 77.85 11.565 78.06 11.635 ;
    RECT 77.85 11.925 78.06 11.995 ;
    RECT 77.85 12.285 78.06 12.355 ;
    RECT 78.31 11.565 78.52 11.635 ;
    RECT 78.31 11.925 78.52 11.995 ;
    RECT 78.31 12.285 78.52 12.355 ;
    RECT 74.53 11.565 74.74 11.635 ;
    RECT 74.53 11.925 74.74 11.995 ;
    RECT 74.53 12.285 74.74 12.355 ;
    RECT 74.99 11.565 75.2 11.635 ;
    RECT 74.99 11.925 75.2 11.995 ;
    RECT 74.99 12.285 75.2 12.355 ;
    RECT 71.21 11.565 71.42 11.635 ;
    RECT 71.21 11.925 71.42 11.995 ;
    RECT 71.21 12.285 71.42 12.355 ;
    RECT 71.67 11.565 71.88 11.635 ;
    RECT 71.67 11.925 71.88 11.995 ;
    RECT 71.67 12.285 71.88 12.355 ;
    RECT 31.37 11.565 31.58 11.635 ;
    RECT 31.37 11.925 31.58 11.995 ;
    RECT 31.37 12.285 31.58 12.355 ;
    RECT 31.83 11.565 32.04 11.635 ;
    RECT 31.83 11.925 32.04 11.995 ;
    RECT 31.83 12.285 32.04 12.355 ;
    RECT 67.89 11.565 68.1 11.635 ;
    RECT 67.89 11.925 68.1 11.995 ;
    RECT 67.89 12.285 68.1 12.355 ;
    RECT 68.35 11.565 68.56 11.635 ;
    RECT 68.35 11.925 68.56 11.995 ;
    RECT 68.35 12.285 68.56 12.355 ;
    RECT 28.05 11.565 28.26 11.635 ;
    RECT 28.05 11.925 28.26 11.995 ;
    RECT 28.05 12.285 28.26 12.355 ;
    RECT 28.51 11.565 28.72 11.635 ;
    RECT 28.51 11.925 28.72 11.995 ;
    RECT 28.51 12.285 28.72 12.355 ;
    RECT 24.73 11.565 24.94 11.635 ;
    RECT 24.73 11.925 24.94 11.995 ;
    RECT 24.73 12.285 24.94 12.355 ;
    RECT 25.19 11.565 25.4 11.635 ;
    RECT 25.19 11.925 25.4 11.995 ;
    RECT 25.19 12.285 25.4 12.355 ;
    RECT 21.41 11.565 21.62 11.635 ;
    RECT 21.41 11.925 21.62 11.995 ;
    RECT 21.41 12.285 21.62 12.355 ;
    RECT 21.87 11.565 22.08 11.635 ;
    RECT 21.87 11.925 22.08 11.995 ;
    RECT 21.87 12.285 22.08 12.355 ;
    RECT 18.09 11.565 18.3 11.635 ;
    RECT 18.09 11.925 18.3 11.995 ;
    RECT 18.09 12.285 18.3 12.355 ;
    RECT 18.55 11.565 18.76 11.635 ;
    RECT 18.55 11.925 18.76 11.995 ;
    RECT 18.55 12.285 18.76 12.355 ;
    RECT 14.77 11.565 14.98 11.635 ;
    RECT 14.77 11.925 14.98 11.995 ;
    RECT 14.77 12.285 14.98 12.355 ;
    RECT 15.23 11.565 15.44 11.635 ;
    RECT 15.23 11.925 15.44 11.995 ;
    RECT 15.23 12.285 15.44 12.355 ;
    RECT 11.45 11.565 11.66 11.635 ;
    RECT 11.45 11.925 11.66 11.995 ;
    RECT 11.45 12.285 11.66 12.355 ;
    RECT 11.91 11.565 12.12 11.635 ;
    RECT 11.91 11.925 12.12 11.995 ;
    RECT 11.91 12.285 12.12 12.355 ;
    RECT 8.13 11.565 8.34 11.635 ;
    RECT 8.13 11.925 8.34 11.995 ;
    RECT 8.13 12.285 8.34 12.355 ;
    RECT 8.59 11.565 8.8 11.635 ;
    RECT 8.59 11.925 8.8 11.995 ;
    RECT 8.59 12.285 8.8 12.355 ;
    RECT 0.4 11.925 0.47 11.995 ;
    RECT 4.81 11.565 5.02 11.635 ;
    RECT 4.81 11.925 5.02 11.995 ;
    RECT 4.81 12.285 5.02 12.355 ;
    RECT 5.27 11.565 5.48 11.635 ;
    RECT 5.27 11.925 5.48 11.995 ;
    RECT 5.27 12.285 5.48 12.355 ;
    RECT 164.17 11.565 164.38 11.635 ;
    RECT 164.17 11.925 164.38 11.995 ;
    RECT 164.17 12.285 164.38 12.355 ;
    RECT 164.63 11.565 164.84 11.635 ;
    RECT 164.63 11.925 164.84 11.995 ;
    RECT 164.63 12.285 164.84 12.355 ;
    RECT 160.85 11.565 161.06 11.635 ;
    RECT 160.85 11.925 161.06 11.995 ;
    RECT 160.85 12.285 161.06 12.355 ;
    RECT 161.31 11.565 161.52 11.635 ;
    RECT 161.31 11.925 161.52 11.995 ;
    RECT 161.31 12.285 161.52 12.355 ;
    RECT 157.53 11.565 157.74 11.635 ;
    RECT 157.53 11.925 157.74 11.995 ;
    RECT 157.53 12.285 157.74 12.355 ;
    RECT 157.99 11.565 158.2 11.635 ;
    RECT 157.99 11.925 158.2 11.995 ;
    RECT 157.99 12.285 158.2 12.355 ;
    RECT 154.21 11.565 154.42 11.635 ;
    RECT 154.21 11.925 154.42 11.995 ;
    RECT 154.21 12.285 154.42 12.355 ;
    RECT 154.67 11.565 154.88 11.635 ;
    RECT 154.67 11.925 154.88 11.995 ;
    RECT 154.67 12.285 154.88 12.355 ;
    RECT 150.89 11.565 151.1 11.635 ;
    RECT 150.89 11.925 151.1 11.995 ;
    RECT 150.89 12.285 151.1 12.355 ;
    RECT 151.35 11.565 151.56 11.635 ;
    RECT 151.35 11.925 151.56 11.995 ;
    RECT 151.35 12.285 151.56 12.355 ;
    RECT 170.81 11.565 171.02 11.635 ;
    RECT 170.81 11.925 171.02 11.995 ;
    RECT 170.81 12.285 171.02 12.355 ;
    RECT 171.27 11.565 171.48 11.635 ;
    RECT 171.27 11.925 171.48 11.995 ;
    RECT 171.27 12.285 171.48 12.355 ;
    RECT 147.57 11.565 147.78 11.635 ;
    RECT 147.57 11.925 147.78 11.995 ;
    RECT 147.57 12.285 147.78 12.355 ;
    RECT 148.03 11.565 148.24 11.635 ;
    RECT 148.03 11.925 148.24 11.995 ;
    RECT 148.03 12.285 148.24 12.355 ;
    RECT 144.25 11.565 144.46 11.635 ;
    RECT 144.25 11.925 144.46 11.995 ;
    RECT 144.25 12.285 144.46 12.355 ;
    RECT 144.71 11.565 144.92 11.635 ;
    RECT 144.71 11.925 144.92 11.995 ;
    RECT 144.71 12.285 144.92 12.355 ;
    RECT 140.93 11.565 141.14 11.635 ;
    RECT 140.93 11.925 141.14 11.995 ;
    RECT 140.93 12.285 141.14 12.355 ;
    RECT 141.39 11.565 141.6 11.635 ;
    RECT 141.39 11.925 141.6 11.995 ;
    RECT 141.39 12.285 141.6 12.355 ;
    RECT 137.61 11.565 137.82 11.635 ;
    RECT 137.61 11.925 137.82 11.995 ;
    RECT 137.61 12.285 137.82 12.355 ;
    RECT 138.07 11.565 138.28 11.635 ;
    RECT 138.07 11.925 138.28 11.995 ;
    RECT 138.07 12.285 138.28 12.355 ;
    RECT 134.29 11.565 134.5 11.635 ;
    RECT 134.29 11.925 134.5 11.995 ;
    RECT 134.29 12.285 134.5 12.355 ;
    RECT 134.75 11.565 134.96 11.635 ;
    RECT 134.75 11.925 134.96 11.995 ;
    RECT 134.75 12.285 134.96 12.355 ;
    RECT 1.49 11.565 1.7 11.635 ;
    RECT 1.49 11.925 1.7 11.995 ;
    RECT 1.49 12.285 1.7 12.355 ;
    RECT 1.95 11.565 2.16 11.635 ;
    RECT 1.95 11.925 2.16 11.995 ;
    RECT 1.95 12.285 2.16 12.355 ;
    RECT 64.57 11.565 64.78 11.635 ;
    RECT 64.57 11.925 64.78 11.995 ;
    RECT 64.57 12.285 64.78 12.355 ;
    RECT 65.03 11.565 65.24 11.635 ;
    RECT 65.03 11.925 65.24 11.995 ;
    RECT 65.03 12.285 65.24 12.355 ;
    RECT 61.25 18.045 61.46 18.115 ;
    RECT 61.25 18.405 61.46 18.475 ;
    RECT 61.25 18.765 61.46 18.835 ;
    RECT 61.71 18.045 61.92 18.115 ;
    RECT 61.71 18.405 61.92 18.475 ;
    RECT 61.71 18.765 61.92 18.835 ;
    RECT 57.93 18.045 58.14 18.115 ;
    RECT 57.93 18.405 58.14 18.475 ;
    RECT 57.93 18.765 58.14 18.835 ;
    RECT 58.39 18.045 58.6 18.115 ;
    RECT 58.39 18.405 58.6 18.475 ;
    RECT 58.39 18.765 58.6 18.835 ;
    RECT 54.61 18.045 54.82 18.115 ;
    RECT 54.61 18.405 54.82 18.475 ;
    RECT 54.61 18.765 54.82 18.835 ;
    RECT 55.07 18.045 55.28 18.115 ;
    RECT 55.07 18.405 55.28 18.475 ;
    RECT 55.07 18.765 55.28 18.835 ;
    RECT 51.29 18.045 51.5 18.115 ;
    RECT 51.29 18.405 51.5 18.475 ;
    RECT 51.29 18.765 51.5 18.835 ;
    RECT 51.75 18.045 51.96 18.115 ;
    RECT 51.75 18.405 51.96 18.475 ;
    RECT 51.75 18.765 51.96 18.835 ;
    RECT 47.97 18.045 48.18 18.115 ;
    RECT 47.97 18.405 48.18 18.475 ;
    RECT 47.97 18.765 48.18 18.835 ;
    RECT 48.43 18.045 48.64 18.115 ;
    RECT 48.43 18.405 48.64 18.475 ;
    RECT 48.43 18.765 48.64 18.835 ;
    RECT 44.65 18.045 44.86 18.115 ;
    RECT 44.65 18.405 44.86 18.475 ;
    RECT 44.65 18.765 44.86 18.835 ;
    RECT 45.11 18.045 45.32 18.115 ;
    RECT 45.11 18.405 45.32 18.475 ;
    RECT 45.11 18.765 45.32 18.835 ;
    RECT 41.33 18.045 41.54 18.115 ;
    RECT 41.33 18.405 41.54 18.475 ;
    RECT 41.33 18.765 41.54 18.835 ;
    RECT 41.79 18.045 42.0 18.115 ;
    RECT 41.79 18.405 42.0 18.475 ;
    RECT 41.79 18.765 42.0 18.835 ;
    RECT 38.01 18.045 38.22 18.115 ;
    RECT 38.01 18.405 38.22 18.475 ;
    RECT 38.01 18.765 38.22 18.835 ;
    RECT 38.47 18.045 38.68 18.115 ;
    RECT 38.47 18.405 38.68 18.475 ;
    RECT 38.47 18.765 38.68 18.835 ;
    RECT 34.69 18.045 34.9 18.115 ;
    RECT 34.69 18.405 34.9 18.475 ;
    RECT 34.69 18.765 34.9 18.835 ;
    RECT 35.15 18.045 35.36 18.115 ;
    RECT 35.15 18.405 35.36 18.475 ;
    RECT 35.15 18.765 35.36 18.835 ;
    RECT 173.945 18.405 174.015 18.475 ;
    RECT 130.97 18.045 131.18 18.115 ;
    RECT 130.97 18.405 131.18 18.475 ;
    RECT 130.97 18.765 131.18 18.835 ;
    RECT 131.43 18.045 131.64 18.115 ;
    RECT 131.43 18.405 131.64 18.475 ;
    RECT 131.43 18.765 131.64 18.835 ;
    RECT 127.65 18.045 127.86 18.115 ;
    RECT 127.65 18.405 127.86 18.475 ;
    RECT 127.65 18.765 127.86 18.835 ;
    RECT 128.11 18.045 128.32 18.115 ;
    RECT 128.11 18.405 128.32 18.475 ;
    RECT 128.11 18.765 128.32 18.835 ;
    RECT 124.33 18.045 124.54 18.115 ;
    RECT 124.33 18.405 124.54 18.475 ;
    RECT 124.33 18.765 124.54 18.835 ;
    RECT 124.79 18.045 125.0 18.115 ;
    RECT 124.79 18.405 125.0 18.475 ;
    RECT 124.79 18.765 125.0 18.835 ;
    RECT 121.01 18.045 121.22 18.115 ;
    RECT 121.01 18.405 121.22 18.475 ;
    RECT 121.01 18.765 121.22 18.835 ;
    RECT 121.47 18.045 121.68 18.115 ;
    RECT 121.47 18.405 121.68 18.475 ;
    RECT 121.47 18.765 121.68 18.835 ;
    RECT 117.69 18.045 117.9 18.115 ;
    RECT 117.69 18.405 117.9 18.475 ;
    RECT 117.69 18.765 117.9 18.835 ;
    RECT 118.15 18.045 118.36 18.115 ;
    RECT 118.15 18.405 118.36 18.475 ;
    RECT 118.15 18.765 118.36 18.835 ;
    RECT 114.37 18.045 114.58 18.115 ;
    RECT 114.37 18.405 114.58 18.475 ;
    RECT 114.37 18.765 114.58 18.835 ;
    RECT 114.83 18.045 115.04 18.115 ;
    RECT 114.83 18.405 115.04 18.475 ;
    RECT 114.83 18.765 115.04 18.835 ;
    RECT 111.05 18.045 111.26 18.115 ;
    RECT 111.05 18.405 111.26 18.475 ;
    RECT 111.05 18.765 111.26 18.835 ;
    RECT 111.51 18.045 111.72 18.115 ;
    RECT 111.51 18.405 111.72 18.475 ;
    RECT 111.51 18.765 111.72 18.835 ;
    RECT 107.73 18.045 107.94 18.115 ;
    RECT 107.73 18.405 107.94 18.475 ;
    RECT 107.73 18.765 107.94 18.835 ;
    RECT 108.19 18.045 108.4 18.115 ;
    RECT 108.19 18.405 108.4 18.475 ;
    RECT 108.19 18.765 108.4 18.835 ;
    RECT 104.41 18.045 104.62 18.115 ;
    RECT 104.41 18.405 104.62 18.475 ;
    RECT 104.41 18.765 104.62 18.835 ;
    RECT 104.87 18.045 105.08 18.115 ;
    RECT 104.87 18.405 105.08 18.475 ;
    RECT 104.87 18.765 105.08 18.835 ;
    RECT 101.09 18.045 101.3 18.115 ;
    RECT 101.09 18.405 101.3 18.475 ;
    RECT 101.09 18.765 101.3 18.835 ;
    RECT 101.55 18.045 101.76 18.115 ;
    RECT 101.55 18.405 101.76 18.475 ;
    RECT 101.55 18.765 101.76 18.835 ;
    RECT 0.4 18.405 0.47 18.475 ;
    RECT 170.81 18.045 171.02 18.115 ;
    RECT 170.81 18.405 171.02 18.475 ;
    RECT 170.81 18.765 171.02 18.835 ;
    RECT 171.27 18.045 171.48 18.115 ;
    RECT 171.27 18.405 171.48 18.475 ;
    RECT 171.27 18.765 171.48 18.835 ;
    RECT 167.49 18.045 167.7 18.115 ;
    RECT 167.49 18.405 167.7 18.475 ;
    RECT 167.49 18.765 167.7 18.835 ;
    RECT 167.95 18.045 168.16 18.115 ;
    RECT 167.95 18.405 168.16 18.475 ;
    RECT 167.95 18.765 168.16 18.835 ;
    RECT 97.77 18.045 97.98 18.115 ;
    RECT 97.77 18.405 97.98 18.475 ;
    RECT 97.77 18.765 97.98 18.835 ;
    RECT 98.23 18.045 98.44 18.115 ;
    RECT 98.23 18.405 98.44 18.475 ;
    RECT 98.23 18.765 98.44 18.835 ;
    RECT 94.45 18.045 94.66 18.115 ;
    RECT 94.45 18.405 94.66 18.475 ;
    RECT 94.45 18.765 94.66 18.835 ;
    RECT 94.91 18.045 95.12 18.115 ;
    RECT 94.91 18.405 95.12 18.475 ;
    RECT 94.91 18.765 95.12 18.835 ;
    RECT 91.13 18.045 91.34 18.115 ;
    RECT 91.13 18.405 91.34 18.475 ;
    RECT 91.13 18.765 91.34 18.835 ;
    RECT 91.59 18.045 91.8 18.115 ;
    RECT 91.59 18.405 91.8 18.475 ;
    RECT 91.59 18.765 91.8 18.835 ;
    RECT 87.81 18.045 88.02 18.115 ;
    RECT 87.81 18.405 88.02 18.475 ;
    RECT 87.81 18.765 88.02 18.835 ;
    RECT 88.27 18.045 88.48 18.115 ;
    RECT 88.27 18.405 88.48 18.475 ;
    RECT 88.27 18.765 88.48 18.835 ;
    RECT 84.49 18.045 84.7 18.115 ;
    RECT 84.49 18.405 84.7 18.475 ;
    RECT 84.49 18.765 84.7 18.835 ;
    RECT 84.95 18.045 85.16 18.115 ;
    RECT 84.95 18.405 85.16 18.475 ;
    RECT 84.95 18.765 85.16 18.835 ;
    RECT 81.17 18.045 81.38 18.115 ;
    RECT 81.17 18.405 81.38 18.475 ;
    RECT 81.17 18.765 81.38 18.835 ;
    RECT 81.63 18.045 81.84 18.115 ;
    RECT 81.63 18.405 81.84 18.475 ;
    RECT 81.63 18.765 81.84 18.835 ;
    RECT 77.85 18.045 78.06 18.115 ;
    RECT 77.85 18.405 78.06 18.475 ;
    RECT 77.85 18.765 78.06 18.835 ;
    RECT 78.31 18.045 78.52 18.115 ;
    RECT 78.31 18.405 78.52 18.475 ;
    RECT 78.31 18.765 78.52 18.835 ;
    RECT 74.53 18.045 74.74 18.115 ;
    RECT 74.53 18.405 74.74 18.475 ;
    RECT 74.53 18.765 74.74 18.835 ;
    RECT 74.99 18.045 75.2 18.115 ;
    RECT 74.99 18.405 75.2 18.475 ;
    RECT 74.99 18.765 75.2 18.835 ;
    RECT 71.21 18.045 71.42 18.115 ;
    RECT 71.21 18.405 71.42 18.475 ;
    RECT 71.21 18.765 71.42 18.835 ;
    RECT 71.67 18.045 71.88 18.115 ;
    RECT 71.67 18.405 71.88 18.475 ;
    RECT 71.67 18.765 71.88 18.835 ;
    RECT 31.37 18.045 31.58 18.115 ;
    RECT 31.37 18.405 31.58 18.475 ;
    RECT 31.37 18.765 31.58 18.835 ;
    RECT 31.83 18.045 32.04 18.115 ;
    RECT 31.83 18.405 32.04 18.475 ;
    RECT 31.83 18.765 32.04 18.835 ;
    RECT 67.89 18.045 68.1 18.115 ;
    RECT 67.89 18.405 68.1 18.475 ;
    RECT 67.89 18.765 68.1 18.835 ;
    RECT 68.35 18.045 68.56 18.115 ;
    RECT 68.35 18.405 68.56 18.475 ;
    RECT 68.35 18.765 68.56 18.835 ;
    RECT 28.05 18.045 28.26 18.115 ;
    RECT 28.05 18.405 28.26 18.475 ;
    RECT 28.05 18.765 28.26 18.835 ;
    RECT 28.51 18.045 28.72 18.115 ;
    RECT 28.51 18.405 28.72 18.475 ;
    RECT 28.51 18.765 28.72 18.835 ;
    RECT 24.73 18.045 24.94 18.115 ;
    RECT 24.73 18.405 24.94 18.475 ;
    RECT 24.73 18.765 24.94 18.835 ;
    RECT 25.19 18.045 25.4 18.115 ;
    RECT 25.19 18.405 25.4 18.475 ;
    RECT 25.19 18.765 25.4 18.835 ;
    RECT 21.41 18.045 21.62 18.115 ;
    RECT 21.41 18.405 21.62 18.475 ;
    RECT 21.41 18.765 21.62 18.835 ;
    RECT 21.87 18.045 22.08 18.115 ;
    RECT 21.87 18.405 22.08 18.475 ;
    RECT 21.87 18.765 22.08 18.835 ;
    RECT 18.09 18.045 18.3 18.115 ;
    RECT 18.09 18.405 18.3 18.475 ;
    RECT 18.09 18.765 18.3 18.835 ;
    RECT 18.55 18.045 18.76 18.115 ;
    RECT 18.55 18.405 18.76 18.475 ;
    RECT 18.55 18.765 18.76 18.835 ;
    RECT 14.77 18.045 14.98 18.115 ;
    RECT 14.77 18.405 14.98 18.475 ;
    RECT 14.77 18.765 14.98 18.835 ;
    RECT 15.23 18.045 15.44 18.115 ;
    RECT 15.23 18.405 15.44 18.475 ;
    RECT 15.23 18.765 15.44 18.835 ;
    RECT 11.45 18.045 11.66 18.115 ;
    RECT 11.45 18.405 11.66 18.475 ;
    RECT 11.45 18.765 11.66 18.835 ;
    RECT 11.91 18.045 12.12 18.115 ;
    RECT 11.91 18.405 12.12 18.475 ;
    RECT 11.91 18.765 12.12 18.835 ;
    RECT 8.13 18.045 8.34 18.115 ;
    RECT 8.13 18.405 8.34 18.475 ;
    RECT 8.13 18.765 8.34 18.835 ;
    RECT 8.59 18.045 8.8 18.115 ;
    RECT 8.59 18.405 8.8 18.475 ;
    RECT 8.59 18.765 8.8 18.835 ;
    RECT 4.81 18.045 5.02 18.115 ;
    RECT 4.81 18.405 5.02 18.475 ;
    RECT 4.81 18.765 5.02 18.835 ;
    RECT 5.27 18.045 5.48 18.115 ;
    RECT 5.27 18.405 5.48 18.475 ;
    RECT 5.27 18.765 5.48 18.835 ;
    RECT 164.17 18.045 164.38 18.115 ;
    RECT 164.17 18.405 164.38 18.475 ;
    RECT 164.17 18.765 164.38 18.835 ;
    RECT 164.63 18.045 164.84 18.115 ;
    RECT 164.63 18.405 164.84 18.475 ;
    RECT 164.63 18.765 164.84 18.835 ;
    RECT 1.49 18.045 1.7 18.115 ;
    RECT 1.49 18.405 1.7 18.475 ;
    RECT 1.49 18.765 1.7 18.835 ;
    RECT 1.95 18.045 2.16 18.115 ;
    RECT 1.95 18.405 2.16 18.475 ;
    RECT 1.95 18.765 2.16 18.835 ;
    RECT 160.85 18.045 161.06 18.115 ;
    RECT 160.85 18.405 161.06 18.475 ;
    RECT 160.85 18.765 161.06 18.835 ;
    RECT 161.31 18.045 161.52 18.115 ;
    RECT 161.31 18.405 161.52 18.475 ;
    RECT 161.31 18.765 161.52 18.835 ;
    RECT 157.53 18.045 157.74 18.115 ;
    RECT 157.53 18.405 157.74 18.475 ;
    RECT 157.53 18.765 157.74 18.835 ;
    RECT 157.99 18.045 158.2 18.115 ;
    RECT 157.99 18.405 158.2 18.475 ;
    RECT 157.99 18.765 158.2 18.835 ;
    RECT 154.21 18.045 154.42 18.115 ;
    RECT 154.21 18.405 154.42 18.475 ;
    RECT 154.21 18.765 154.42 18.835 ;
    RECT 154.67 18.045 154.88 18.115 ;
    RECT 154.67 18.405 154.88 18.475 ;
    RECT 154.67 18.765 154.88 18.835 ;
    RECT 150.89 18.045 151.1 18.115 ;
    RECT 150.89 18.405 151.1 18.475 ;
    RECT 150.89 18.765 151.1 18.835 ;
    RECT 151.35 18.045 151.56 18.115 ;
    RECT 151.35 18.405 151.56 18.475 ;
    RECT 151.35 18.765 151.56 18.835 ;
    RECT 147.57 18.045 147.78 18.115 ;
    RECT 147.57 18.405 147.78 18.475 ;
    RECT 147.57 18.765 147.78 18.835 ;
    RECT 148.03 18.045 148.24 18.115 ;
    RECT 148.03 18.405 148.24 18.475 ;
    RECT 148.03 18.765 148.24 18.835 ;
    RECT 144.25 18.045 144.46 18.115 ;
    RECT 144.25 18.405 144.46 18.475 ;
    RECT 144.25 18.765 144.46 18.835 ;
    RECT 144.71 18.045 144.92 18.115 ;
    RECT 144.71 18.405 144.92 18.475 ;
    RECT 144.71 18.765 144.92 18.835 ;
    RECT 140.93 18.045 141.14 18.115 ;
    RECT 140.93 18.405 141.14 18.475 ;
    RECT 140.93 18.765 141.14 18.835 ;
    RECT 141.39 18.045 141.6 18.115 ;
    RECT 141.39 18.405 141.6 18.475 ;
    RECT 141.39 18.765 141.6 18.835 ;
    RECT 137.61 18.045 137.82 18.115 ;
    RECT 137.61 18.405 137.82 18.475 ;
    RECT 137.61 18.765 137.82 18.835 ;
    RECT 138.07 18.045 138.28 18.115 ;
    RECT 138.07 18.405 138.28 18.475 ;
    RECT 138.07 18.765 138.28 18.835 ;
    RECT 134.29 18.045 134.5 18.115 ;
    RECT 134.29 18.405 134.5 18.475 ;
    RECT 134.29 18.765 134.5 18.835 ;
    RECT 134.75 18.045 134.96 18.115 ;
    RECT 134.75 18.405 134.96 18.475 ;
    RECT 134.75 18.765 134.96 18.835 ;
    RECT 64.57 18.045 64.78 18.115 ;
    RECT 64.57 18.405 64.78 18.475 ;
    RECT 64.57 18.765 64.78 18.835 ;
    RECT 65.03 18.045 65.24 18.115 ;
    RECT 65.03 18.405 65.24 18.475 ;
    RECT 65.03 18.765 65.24 18.835 ;
    RECT 61.25 17.325 61.46 17.395 ;
    RECT 61.25 17.685 61.46 17.755 ;
    RECT 61.25 18.045 61.46 18.115 ;
    RECT 61.71 17.325 61.92 17.395 ;
    RECT 61.71 17.685 61.92 17.755 ;
    RECT 61.71 18.045 61.92 18.115 ;
    RECT 57.93 17.325 58.14 17.395 ;
    RECT 57.93 17.685 58.14 17.755 ;
    RECT 57.93 18.045 58.14 18.115 ;
    RECT 58.39 17.325 58.6 17.395 ;
    RECT 58.39 17.685 58.6 17.755 ;
    RECT 58.39 18.045 58.6 18.115 ;
    RECT 54.61 17.325 54.82 17.395 ;
    RECT 54.61 17.685 54.82 17.755 ;
    RECT 54.61 18.045 54.82 18.115 ;
    RECT 55.07 17.325 55.28 17.395 ;
    RECT 55.07 17.685 55.28 17.755 ;
    RECT 55.07 18.045 55.28 18.115 ;
    RECT 51.29 17.325 51.5 17.395 ;
    RECT 51.29 17.685 51.5 17.755 ;
    RECT 51.29 18.045 51.5 18.115 ;
    RECT 51.75 17.325 51.96 17.395 ;
    RECT 51.75 17.685 51.96 17.755 ;
    RECT 51.75 18.045 51.96 18.115 ;
    RECT 47.97 17.325 48.18 17.395 ;
    RECT 47.97 17.685 48.18 17.755 ;
    RECT 47.97 18.045 48.18 18.115 ;
    RECT 48.43 17.325 48.64 17.395 ;
    RECT 48.43 17.685 48.64 17.755 ;
    RECT 48.43 18.045 48.64 18.115 ;
    RECT 44.65 17.325 44.86 17.395 ;
    RECT 44.65 17.685 44.86 17.755 ;
    RECT 44.65 18.045 44.86 18.115 ;
    RECT 45.11 17.325 45.32 17.395 ;
    RECT 45.11 17.685 45.32 17.755 ;
    RECT 45.11 18.045 45.32 18.115 ;
    RECT 41.33 17.325 41.54 17.395 ;
    RECT 41.33 17.685 41.54 17.755 ;
    RECT 41.33 18.045 41.54 18.115 ;
    RECT 41.79 17.325 42.0 17.395 ;
    RECT 41.79 17.685 42.0 17.755 ;
    RECT 41.79 18.045 42.0 18.115 ;
    RECT 38.01 17.325 38.22 17.395 ;
    RECT 38.01 17.685 38.22 17.755 ;
    RECT 38.01 18.045 38.22 18.115 ;
    RECT 38.47 17.325 38.68 17.395 ;
    RECT 38.47 17.685 38.68 17.755 ;
    RECT 38.47 18.045 38.68 18.115 ;
    RECT 34.69 17.325 34.9 17.395 ;
    RECT 34.69 17.685 34.9 17.755 ;
    RECT 34.69 18.045 34.9 18.115 ;
    RECT 35.15 17.325 35.36 17.395 ;
    RECT 35.15 17.685 35.36 17.755 ;
    RECT 35.15 18.045 35.36 18.115 ;
    RECT 173.945 17.685 174.015 17.755 ;
    RECT 130.97 17.325 131.18 17.395 ;
    RECT 130.97 17.685 131.18 17.755 ;
    RECT 130.97 18.045 131.18 18.115 ;
    RECT 131.43 17.325 131.64 17.395 ;
    RECT 131.43 17.685 131.64 17.755 ;
    RECT 131.43 18.045 131.64 18.115 ;
    RECT 127.65 17.325 127.86 17.395 ;
    RECT 127.65 17.685 127.86 17.755 ;
    RECT 127.65 18.045 127.86 18.115 ;
    RECT 128.11 17.325 128.32 17.395 ;
    RECT 128.11 17.685 128.32 17.755 ;
    RECT 128.11 18.045 128.32 18.115 ;
    RECT 124.33 17.325 124.54 17.395 ;
    RECT 124.33 17.685 124.54 17.755 ;
    RECT 124.33 18.045 124.54 18.115 ;
    RECT 124.79 17.325 125.0 17.395 ;
    RECT 124.79 17.685 125.0 17.755 ;
    RECT 124.79 18.045 125.0 18.115 ;
    RECT 121.01 17.325 121.22 17.395 ;
    RECT 121.01 17.685 121.22 17.755 ;
    RECT 121.01 18.045 121.22 18.115 ;
    RECT 121.47 17.325 121.68 17.395 ;
    RECT 121.47 17.685 121.68 17.755 ;
    RECT 121.47 18.045 121.68 18.115 ;
    RECT 117.69 17.325 117.9 17.395 ;
    RECT 117.69 17.685 117.9 17.755 ;
    RECT 117.69 18.045 117.9 18.115 ;
    RECT 118.15 17.325 118.36 17.395 ;
    RECT 118.15 17.685 118.36 17.755 ;
    RECT 118.15 18.045 118.36 18.115 ;
    RECT 114.37 17.325 114.58 17.395 ;
    RECT 114.37 17.685 114.58 17.755 ;
    RECT 114.37 18.045 114.58 18.115 ;
    RECT 114.83 17.325 115.04 17.395 ;
    RECT 114.83 17.685 115.04 17.755 ;
    RECT 114.83 18.045 115.04 18.115 ;
    RECT 111.05 17.325 111.26 17.395 ;
    RECT 111.05 17.685 111.26 17.755 ;
    RECT 111.05 18.045 111.26 18.115 ;
    RECT 111.51 17.325 111.72 17.395 ;
    RECT 111.51 17.685 111.72 17.755 ;
    RECT 111.51 18.045 111.72 18.115 ;
    RECT 107.73 17.325 107.94 17.395 ;
    RECT 107.73 17.685 107.94 17.755 ;
    RECT 107.73 18.045 107.94 18.115 ;
    RECT 108.19 17.325 108.4 17.395 ;
    RECT 108.19 17.685 108.4 17.755 ;
    RECT 108.19 18.045 108.4 18.115 ;
    RECT 104.41 17.325 104.62 17.395 ;
    RECT 104.41 17.685 104.62 17.755 ;
    RECT 104.41 18.045 104.62 18.115 ;
    RECT 104.87 17.325 105.08 17.395 ;
    RECT 104.87 17.685 105.08 17.755 ;
    RECT 104.87 18.045 105.08 18.115 ;
    RECT 101.09 17.325 101.3 17.395 ;
    RECT 101.09 17.685 101.3 17.755 ;
    RECT 101.09 18.045 101.3 18.115 ;
    RECT 101.55 17.325 101.76 17.395 ;
    RECT 101.55 17.685 101.76 17.755 ;
    RECT 101.55 18.045 101.76 18.115 ;
    RECT 0.4 17.685 0.47 17.755 ;
    RECT 170.81 17.325 171.02 17.395 ;
    RECT 170.81 17.685 171.02 17.755 ;
    RECT 170.81 18.045 171.02 18.115 ;
    RECT 171.27 17.325 171.48 17.395 ;
    RECT 171.27 17.685 171.48 17.755 ;
    RECT 171.27 18.045 171.48 18.115 ;
    RECT 167.49 17.325 167.7 17.395 ;
    RECT 167.49 17.685 167.7 17.755 ;
    RECT 167.49 18.045 167.7 18.115 ;
    RECT 167.95 17.325 168.16 17.395 ;
    RECT 167.95 17.685 168.16 17.755 ;
    RECT 167.95 18.045 168.16 18.115 ;
    RECT 97.77 17.325 97.98 17.395 ;
    RECT 97.77 17.685 97.98 17.755 ;
    RECT 97.77 18.045 97.98 18.115 ;
    RECT 98.23 17.325 98.44 17.395 ;
    RECT 98.23 17.685 98.44 17.755 ;
    RECT 98.23 18.045 98.44 18.115 ;
    RECT 94.45 17.325 94.66 17.395 ;
    RECT 94.45 17.685 94.66 17.755 ;
    RECT 94.45 18.045 94.66 18.115 ;
    RECT 94.91 17.325 95.12 17.395 ;
    RECT 94.91 17.685 95.12 17.755 ;
    RECT 94.91 18.045 95.12 18.115 ;
    RECT 91.13 17.325 91.34 17.395 ;
    RECT 91.13 17.685 91.34 17.755 ;
    RECT 91.13 18.045 91.34 18.115 ;
    RECT 91.59 17.325 91.8 17.395 ;
    RECT 91.59 17.685 91.8 17.755 ;
    RECT 91.59 18.045 91.8 18.115 ;
    RECT 87.81 17.325 88.02 17.395 ;
    RECT 87.81 17.685 88.02 17.755 ;
    RECT 87.81 18.045 88.02 18.115 ;
    RECT 88.27 17.325 88.48 17.395 ;
    RECT 88.27 17.685 88.48 17.755 ;
    RECT 88.27 18.045 88.48 18.115 ;
    RECT 84.49 17.325 84.7 17.395 ;
    RECT 84.49 17.685 84.7 17.755 ;
    RECT 84.49 18.045 84.7 18.115 ;
    RECT 84.95 17.325 85.16 17.395 ;
    RECT 84.95 17.685 85.16 17.755 ;
    RECT 84.95 18.045 85.16 18.115 ;
    RECT 81.17 17.325 81.38 17.395 ;
    RECT 81.17 17.685 81.38 17.755 ;
    RECT 81.17 18.045 81.38 18.115 ;
    RECT 81.63 17.325 81.84 17.395 ;
    RECT 81.63 17.685 81.84 17.755 ;
    RECT 81.63 18.045 81.84 18.115 ;
    RECT 77.85 17.325 78.06 17.395 ;
    RECT 77.85 17.685 78.06 17.755 ;
    RECT 77.85 18.045 78.06 18.115 ;
    RECT 78.31 17.325 78.52 17.395 ;
    RECT 78.31 17.685 78.52 17.755 ;
    RECT 78.31 18.045 78.52 18.115 ;
    RECT 74.53 17.325 74.74 17.395 ;
    RECT 74.53 17.685 74.74 17.755 ;
    RECT 74.53 18.045 74.74 18.115 ;
    RECT 74.99 17.325 75.2 17.395 ;
    RECT 74.99 17.685 75.2 17.755 ;
    RECT 74.99 18.045 75.2 18.115 ;
    RECT 71.21 17.325 71.42 17.395 ;
    RECT 71.21 17.685 71.42 17.755 ;
    RECT 71.21 18.045 71.42 18.115 ;
    RECT 71.67 17.325 71.88 17.395 ;
    RECT 71.67 17.685 71.88 17.755 ;
    RECT 71.67 18.045 71.88 18.115 ;
    RECT 31.37 17.325 31.58 17.395 ;
    RECT 31.37 17.685 31.58 17.755 ;
    RECT 31.37 18.045 31.58 18.115 ;
    RECT 31.83 17.325 32.04 17.395 ;
    RECT 31.83 17.685 32.04 17.755 ;
    RECT 31.83 18.045 32.04 18.115 ;
    RECT 67.89 17.325 68.1 17.395 ;
    RECT 67.89 17.685 68.1 17.755 ;
    RECT 67.89 18.045 68.1 18.115 ;
    RECT 68.35 17.325 68.56 17.395 ;
    RECT 68.35 17.685 68.56 17.755 ;
    RECT 68.35 18.045 68.56 18.115 ;
    RECT 28.05 17.325 28.26 17.395 ;
    RECT 28.05 17.685 28.26 17.755 ;
    RECT 28.05 18.045 28.26 18.115 ;
    RECT 28.51 17.325 28.72 17.395 ;
    RECT 28.51 17.685 28.72 17.755 ;
    RECT 28.51 18.045 28.72 18.115 ;
    RECT 24.73 17.325 24.94 17.395 ;
    RECT 24.73 17.685 24.94 17.755 ;
    RECT 24.73 18.045 24.94 18.115 ;
    RECT 25.19 17.325 25.4 17.395 ;
    RECT 25.19 17.685 25.4 17.755 ;
    RECT 25.19 18.045 25.4 18.115 ;
    RECT 21.41 17.325 21.62 17.395 ;
    RECT 21.41 17.685 21.62 17.755 ;
    RECT 21.41 18.045 21.62 18.115 ;
    RECT 21.87 17.325 22.08 17.395 ;
    RECT 21.87 17.685 22.08 17.755 ;
    RECT 21.87 18.045 22.08 18.115 ;
    RECT 18.09 17.325 18.3 17.395 ;
    RECT 18.09 17.685 18.3 17.755 ;
    RECT 18.09 18.045 18.3 18.115 ;
    RECT 18.55 17.325 18.76 17.395 ;
    RECT 18.55 17.685 18.76 17.755 ;
    RECT 18.55 18.045 18.76 18.115 ;
    RECT 14.77 17.325 14.98 17.395 ;
    RECT 14.77 17.685 14.98 17.755 ;
    RECT 14.77 18.045 14.98 18.115 ;
    RECT 15.23 17.325 15.44 17.395 ;
    RECT 15.23 17.685 15.44 17.755 ;
    RECT 15.23 18.045 15.44 18.115 ;
    RECT 11.45 17.325 11.66 17.395 ;
    RECT 11.45 17.685 11.66 17.755 ;
    RECT 11.45 18.045 11.66 18.115 ;
    RECT 11.91 17.325 12.12 17.395 ;
    RECT 11.91 17.685 12.12 17.755 ;
    RECT 11.91 18.045 12.12 18.115 ;
    RECT 8.13 17.325 8.34 17.395 ;
    RECT 8.13 17.685 8.34 17.755 ;
    RECT 8.13 18.045 8.34 18.115 ;
    RECT 8.59 17.325 8.8 17.395 ;
    RECT 8.59 17.685 8.8 17.755 ;
    RECT 8.59 18.045 8.8 18.115 ;
    RECT 4.81 17.325 5.02 17.395 ;
    RECT 4.81 17.685 5.02 17.755 ;
    RECT 4.81 18.045 5.02 18.115 ;
    RECT 5.27 17.325 5.48 17.395 ;
    RECT 5.27 17.685 5.48 17.755 ;
    RECT 5.27 18.045 5.48 18.115 ;
    RECT 164.17 17.325 164.38 17.395 ;
    RECT 164.17 17.685 164.38 17.755 ;
    RECT 164.17 18.045 164.38 18.115 ;
    RECT 164.63 17.325 164.84 17.395 ;
    RECT 164.63 17.685 164.84 17.755 ;
    RECT 164.63 18.045 164.84 18.115 ;
    RECT 1.49 17.325 1.7 17.395 ;
    RECT 1.49 17.685 1.7 17.755 ;
    RECT 1.49 18.045 1.7 18.115 ;
    RECT 1.95 17.325 2.16 17.395 ;
    RECT 1.95 17.685 2.16 17.755 ;
    RECT 1.95 18.045 2.16 18.115 ;
    RECT 160.85 17.325 161.06 17.395 ;
    RECT 160.85 17.685 161.06 17.755 ;
    RECT 160.85 18.045 161.06 18.115 ;
    RECT 161.31 17.325 161.52 17.395 ;
    RECT 161.31 17.685 161.52 17.755 ;
    RECT 161.31 18.045 161.52 18.115 ;
    RECT 157.53 17.325 157.74 17.395 ;
    RECT 157.53 17.685 157.74 17.755 ;
    RECT 157.53 18.045 157.74 18.115 ;
    RECT 157.99 17.325 158.2 17.395 ;
    RECT 157.99 17.685 158.2 17.755 ;
    RECT 157.99 18.045 158.2 18.115 ;
    RECT 154.21 17.325 154.42 17.395 ;
    RECT 154.21 17.685 154.42 17.755 ;
    RECT 154.21 18.045 154.42 18.115 ;
    RECT 154.67 17.325 154.88 17.395 ;
    RECT 154.67 17.685 154.88 17.755 ;
    RECT 154.67 18.045 154.88 18.115 ;
    RECT 150.89 17.325 151.1 17.395 ;
    RECT 150.89 17.685 151.1 17.755 ;
    RECT 150.89 18.045 151.1 18.115 ;
    RECT 151.35 17.325 151.56 17.395 ;
    RECT 151.35 17.685 151.56 17.755 ;
    RECT 151.35 18.045 151.56 18.115 ;
    RECT 147.57 17.325 147.78 17.395 ;
    RECT 147.57 17.685 147.78 17.755 ;
    RECT 147.57 18.045 147.78 18.115 ;
    RECT 148.03 17.325 148.24 17.395 ;
    RECT 148.03 17.685 148.24 17.755 ;
    RECT 148.03 18.045 148.24 18.115 ;
    RECT 144.25 17.325 144.46 17.395 ;
    RECT 144.25 17.685 144.46 17.755 ;
    RECT 144.25 18.045 144.46 18.115 ;
    RECT 144.71 17.325 144.92 17.395 ;
    RECT 144.71 17.685 144.92 17.755 ;
    RECT 144.71 18.045 144.92 18.115 ;
    RECT 140.93 17.325 141.14 17.395 ;
    RECT 140.93 17.685 141.14 17.755 ;
    RECT 140.93 18.045 141.14 18.115 ;
    RECT 141.39 17.325 141.6 17.395 ;
    RECT 141.39 17.685 141.6 17.755 ;
    RECT 141.39 18.045 141.6 18.115 ;
    RECT 137.61 17.325 137.82 17.395 ;
    RECT 137.61 17.685 137.82 17.755 ;
    RECT 137.61 18.045 137.82 18.115 ;
    RECT 138.07 17.325 138.28 17.395 ;
    RECT 138.07 17.685 138.28 17.755 ;
    RECT 138.07 18.045 138.28 18.115 ;
    RECT 134.29 17.325 134.5 17.395 ;
    RECT 134.29 17.685 134.5 17.755 ;
    RECT 134.29 18.045 134.5 18.115 ;
    RECT 134.75 17.325 134.96 17.395 ;
    RECT 134.75 17.685 134.96 17.755 ;
    RECT 134.75 18.045 134.96 18.115 ;
    RECT 64.57 17.325 64.78 17.395 ;
    RECT 64.57 17.685 64.78 17.755 ;
    RECT 64.57 18.045 64.78 18.115 ;
    RECT 65.03 17.325 65.24 17.395 ;
    RECT 65.03 17.685 65.24 17.755 ;
    RECT 65.03 18.045 65.24 18.115 ;
    RECT 61.25 16.605 61.46 16.675 ;
    RECT 61.25 16.965 61.46 17.035 ;
    RECT 61.25 17.325 61.46 17.395 ;
    RECT 61.71 16.605 61.92 16.675 ;
    RECT 61.71 16.965 61.92 17.035 ;
    RECT 61.71 17.325 61.92 17.395 ;
    RECT 57.93 16.605 58.14 16.675 ;
    RECT 57.93 16.965 58.14 17.035 ;
    RECT 57.93 17.325 58.14 17.395 ;
    RECT 58.39 16.605 58.6 16.675 ;
    RECT 58.39 16.965 58.6 17.035 ;
    RECT 58.39 17.325 58.6 17.395 ;
    RECT 54.61 16.605 54.82 16.675 ;
    RECT 54.61 16.965 54.82 17.035 ;
    RECT 54.61 17.325 54.82 17.395 ;
    RECT 55.07 16.605 55.28 16.675 ;
    RECT 55.07 16.965 55.28 17.035 ;
    RECT 55.07 17.325 55.28 17.395 ;
    RECT 51.29 16.605 51.5 16.675 ;
    RECT 51.29 16.965 51.5 17.035 ;
    RECT 51.29 17.325 51.5 17.395 ;
    RECT 51.75 16.605 51.96 16.675 ;
    RECT 51.75 16.965 51.96 17.035 ;
    RECT 51.75 17.325 51.96 17.395 ;
    RECT 47.97 16.605 48.18 16.675 ;
    RECT 47.97 16.965 48.18 17.035 ;
    RECT 47.97 17.325 48.18 17.395 ;
    RECT 48.43 16.605 48.64 16.675 ;
    RECT 48.43 16.965 48.64 17.035 ;
    RECT 48.43 17.325 48.64 17.395 ;
    RECT 44.65 16.605 44.86 16.675 ;
    RECT 44.65 16.965 44.86 17.035 ;
    RECT 44.65 17.325 44.86 17.395 ;
    RECT 45.11 16.605 45.32 16.675 ;
    RECT 45.11 16.965 45.32 17.035 ;
    RECT 45.11 17.325 45.32 17.395 ;
    RECT 41.33 16.605 41.54 16.675 ;
    RECT 41.33 16.965 41.54 17.035 ;
    RECT 41.33 17.325 41.54 17.395 ;
    RECT 41.79 16.605 42.0 16.675 ;
    RECT 41.79 16.965 42.0 17.035 ;
    RECT 41.79 17.325 42.0 17.395 ;
    RECT 38.01 16.605 38.22 16.675 ;
    RECT 38.01 16.965 38.22 17.035 ;
    RECT 38.01 17.325 38.22 17.395 ;
    RECT 38.47 16.605 38.68 16.675 ;
    RECT 38.47 16.965 38.68 17.035 ;
    RECT 38.47 17.325 38.68 17.395 ;
    RECT 34.69 16.605 34.9 16.675 ;
    RECT 34.69 16.965 34.9 17.035 ;
    RECT 34.69 17.325 34.9 17.395 ;
    RECT 35.15 16.605 35.36 16.675 ;
    RECT 35.15 16.965 35.36 17.035 ;
    RECT 35.15 17.325 35.36 17.395 ;
    RECT 173.945 16.965 174.015 17.035 ;
    RECT 130.97 16.605 131.18 16.675 ;
    RECT 130.97 16.965 131.18 17.035 ;
    RECT 130.97 17.325 131.18 17.395 ;
    RECT 131.43 16.605 131.64 16.675 ;
    RECT 131.43 16.965 131.64 17.035 ;
    RECT 131.43 17.325 131.64 17.395 ;
    RECT 127.65 16.605 127.86 16.675 ;
    RECT 127.65 16.965 127.86 17.035 ;
    RECT 127.65 17.325 127.86 17.395 ;
    RECT 128.11 16.605 128.32 16.675 ;
    RECT 128.11 16.965 128.32 17.035 ;
    RECT 128.11 17.325 128.32 17.395 ;
    RECT 124.33 16.605 124.54 16.675 ;
    RECT 124.33 16.965 124.54 17.035 ;
    RECT 124.33 17.325 124.54 17.395 ;
    RECT 124.79 16.605 125.0 16.675 ;
    RECT 124.79 16.965 125.0 17.035 ;
    RECT 124.79 17.325 125.0 17.395 ;
    RECT 121.01 16.605 121.22 16.675 ;
    RECT 121.01 16.965 121.22 17.035 ;
    RECT 121.01 17.325 121.22 17.395 ;
    RECT 121.47 16.605 121.68 16.675 ;
    RECT 121.47 16.965 121.68 17.035 ;
    RECT 121.47 17.325 121.68 17.395 ;
    RECT 117.69 16.605 117.9 16.675 ;
    RECT 117.69 16.965 117.9 17.035 ;
    RECT 117.69 17.325 117.9 17.395 ;
    RECT 118.15 16.605 118.36 16.675 ;
    RECT 118.15 16.965 118.36 17.035 ;
    RECT 118.15 17.325 118.36 17.395 ;
    RECT 114.37 16.605 114.58 16.675 ;
    RECT 114.37 16.965 114.58 17.035 ;
    RECT 114.37 17.325 114.58 17.395 ;
    RECT 114.83 16.605 115.04 16.675 ;
    RECT 114.83 16.965 115.04 17.035 ;
    RECT 114.83 17.325 115.04 17.395 ;
    RECT 111.05 16.605 111.26 16.675 ;
    RECT 111.05 16.965 111.26 17.035 ;
    RECT 111.05 17.325 111.26 17.395 ;
    RECT 111.51 16.605 111.72 16.675 ;
    RECT 111.51 16.965 111.72 17.035 ;
    RECT 111.51 17.325 111.72 17.395 ;
    RECT 107.73 16.605 107.94 16.675 ;
    RECT 107.73 16.965 107.94 17.035 ;
    RECT 107.73 17.325 107.94 17.395 ;
    RECT 108.19 16.605 108.4 16.675 ;
    RECT 108.19 16.965 108.4 17.035 ;
    RECT 108.19 17.325 108.4 17.395 ;
    RECT 104.41 16.605 104.62 16.675 ;
    RECT 104.41 16.965 104.62 17.035 ;
    RECT 104.41 17.325 104.62 17.395 ;
    RECT 104.87 16.605 105.08 16.675 ;
    RECT 104.87 16.965 105.08 17.035 ;
    RECT 104.87 17.325 105.08 17.395 ;
    RECT 101.09 16.605 101.3 16.675 ;
    RECT 101.09 16.965 101.3 17.035 ;
    RECT 101.09 17.325 101.3 17.395 ;
    RECT 101.55 16.605 101.76 16.675 ;
    RECT 101.55 16.965 101.76 17.035 ;
    RECT 101.55 17.325 101.76 17.395 ;
    RECT 0.4 16.965 0.47 17.035 ;
    RECT 170.81 16.605 171.02 16.675 ;
    RECT 170.81 16.965 171.02 17.035 ;
    RECT 170.81 17.325 171.02 17.395 ;
    RECT 171.27 16.605 171.48 16.675 ;
    RECT 171.27 16.965 171.48 17.035 ;
    RECT 171.27 17.325 171.48 17.395 ;
    RECT 167.49 16.605 167.7 16.675 ;
    RECT 167.49 16.965 167.7 17.035 ;
    RECT 167.49 17.325 167.7 17.395 ;
    RECT 167.95 16.605 168.16 16.675 ;
    RECT 167.95 16.965 168.16 17.035 ;
    RECT 167.95 17.325 168.16 17.395 ;
    RECT 97.77 16.605 97.98 16.675 ;
    RECT 97.77 16.965 97.98 17.035 ;
    RECT 97.77 17.325 97.98 17.395 ;
    RECT 98.23 16.605 98.44 16.675 ;
    RECT 98.23 16.965 98.44 17.035 ;
    RECT 98.23 17.325 98.44 17.395 ;
    RECT 94.45 16.605 94.66 16.675 ;
    RECT 94.45 16.965 94.66 17.035 ;
    RECT 94.45 17.325 94.66 17.395 ;
    RECT 94.91 16.605 95.12 16.675 ;
    RECT 94.91 16.965 95.12 17.035 ;
    RECT 94.91 17.325 95.12 17.395 ;
    RECT 91.13 16.605 91.34 16.675 ;
    RECT 91.13 16.965 91.34 17.035 ;
    RECT 91.13 17.325 91.34 17.395 ;
    RECT 91.59 16.605 91.8 16.675 ;
    RECT 91.59 16.965 91.8 17.035 ;
    RECT 91.59 17.325 91.8 17.395 ;
    RECT 87.81 16.605 88.02 16.675 ;
    RECT 87.81 16.965 88.02 17.035 ;
    RECT 87.81 17.325 88.02 17.395 ;
    RECT 88.27 16.605 88.48 16.675 ;
    RECT 88.27 16.965 88.48 17.035 ;
    RECT 88.27 17.325 88.48 17.395 ;
    RECT 84.49 16.605 84.7 16.675 ;
    RECT 84.49 16.965 84.7 17.035 ;
    RECT 84.49 17.325 84.7 17.395 ;
    RECT 84.95 16.605 85.16 16.675 ;
    RECT 84.95 16.965 85.16 17.035 ;
    RECT 84.95 17.325 85.16 17.395 ;
    RECT 81.17 16.605 81.38 16.675 ;
    RECT 81.17 16.965 81.38 17.035 ;
    RECT 81.17 17.325 81.38 17.395 ;
    RECT 81.63 16.605 81.84 16.675 ;
    RECT 81.63 16.965 81.84 17.035 ;
    RECT 81.63 17.325 81.84 17.395 ;
    RECT 77.85 16.605 78.06 16.675 ;
    RECT 77.85 16.965 78.06 17.035 ;
    RECT 77.85 17.325 78.06 17.395 ;
    RECT 78.31 16.605 78.52 16.675 ;
    RECT 78.31 16.965 78.52 17.035 ;
    RECT 78.31 17.325 78.52 17.395 ;
    RECT 74.53 16.605 74.74 16.675 ;
    RECT 74.53 16.965 74.74 17.035 ;
    RECT 74.53 17.325 74.74 17.395 ;
    RECT 74.99 16.605 75.2 16.675 ;
    RECT 74.99 16.965 75.2 17.035 ;
    RECT 74.99 17.325 75.2 17.395 ;
    RECT 71.21 16.605 71.42 16.675 ;
    RECT 71.21 16.965 71.42 17.035 ;
    RECT 71.21 17.325 71.42 17.395 ;
    RECT 71.67 16.605 71.88 16.675 ;
    RECT 71.67 16.965 71.88 17.035 ;
    RECT 71.67 17.325 71.88 17.395 ;
    RECT 31.37 16.605 31.58 16.675 ;
    RECT 31.37 16.965 31.58 17.035 ;
    RECT 31.37 17.325 31.58 17.395 ;
    RECT 31.83 16.605 32.04 16.675 ;
    RECT 31.83 16.965 32.04 17.035 ;
    RECT 31.83 17.325 32.04 17.395 ;
    RECT 67.89 16.605 68.1 16.675 ;
    RECT 67.89 16.965 68.1 17.035 ;
    RECT 67.89 17.325 68.1 17.395 ;
    RECT 68.35 16.605 68.56 16.675 ;
    RECT 68.35 16.965 68.56 17.035 ;
    RECT 68.35 17.325 68.56 17.395 ;
    RECT 28.05 16.605 28.26 16.675 ;
    RECT 28.05 16.965 28.26 17.035 ;
    RECT 28.05 17.325 28.26 17.395 ;
    RECT 28.51 16.605 28.72 16.675 ;
    RECT 28.51 16.965 28.72 17.035 ;
    RECT 28.51 17.325 28.72 17.395 ;
    RECT 24.73 16.605 24.94 16.675 ;
    RECT 24.73 16.965 24.94 17.035 ;
    RECT 24.73 17.325 24.94 17.395 ;
    RECT 25.19 16.605 25.4 16.675 ;
    RECT 25.19 16.965 25.4 17.035 ;
    RECT 25.19 17.325 25.4 17.395 ;
    RECT 21.41 16.605 21.62 16.675 ;
    RECT 21.41 16.965 21.62 17.035 ;
    RECT 21.41 17.325 21.62 17.395 ;
    RECT 21.87 16.605 22.08 16.675 ;
    RECT 21.87 16.965 22.08 17.035 ;
    RECT 21.87 17.325 22.08 17.395 ;
    RECT 18.09 16.605 18.3 16.675 ;
    RECT 18.09 16.965 18.3 17.035 ;
    RECT 18.09 17.325 18.3 17.395 ;
    RECT 18.55 16.605 18.76 16.675 ;
    RECT 18.55 16.965 18.76 17.035 ;
    RECT 18.55 17.325 18.76 17.395 ;
    RECT 14.77 16.605 14.98 16.675 ;
    RECT 14.77 16.965 14.98 17.035 ;
    RECT 14.77 17.325 14.98 17.395 ;
    RECT 15.23 16.605 15.44 16.675 ;
    RECT 15.23 16.965 15.44 17.035 ;
    RECT 15.23 17.325 15.44 17.395 ;
    RECT 11.45 16.605 11.66 16.675 ;
    RECT 11.45 16.965 11.66 17.035 ;
    RECT 11.45 17.325 11.66 17.395 ;
    RECT 11.91 16.605 12.12 16.675 ;
    RECT 11.91 16.965 12.12 17.035 ;
    RECT 11.91 17.325 12.12 17.395 ;
    RECT 8.13 16.605 8.34 16.675 ;
    RECT 8.13 16.965 8.34 17.035 ;
    RECT 8.13 17.325 8.34 17.395 ;
    RECT 8.59 16.605 8.8 16.675 ;
    RECT 8.59 16.965 8.8 17.035 ;
    RECT 8.59 17.325 8.8 17.395 ;
    RECT 4.81 16.605 5.02 16.675 ;
    RECT 4.81 16.965 5.02 17.035 ;
    RECT 4.81 17.325 5.02 17.395 ;
    RECT 5.27 16.605 5.48 16.675 ;
    RECT 5.27 16.965 5.48 17.035 ;
    RECT 5.27 17.325 5.48 17.395 ;
    RECT 164.17 16.605 164.38 16.675 ;
    RECT 164.17 16.965 164.38 17.035 ;
    RECT 164.17 17.325 164.38 17.395 ;
    RECT 164.63 16.605 164.84 16.675 ;
    RECT 164.63 16.965 164.84 17.035 ;
    RECT 164.63 17.325 164.84 17.395 ;
    RECT 1.49 16.605 1.7 16.675 ;
    RECT 1.49 16.965 1.7 17.035 ;
    RECT 1.49 17.325 1.7 17.395 ;
    RECT 1.95 16.605 2.16 16.675 ;
    RECT 1.95 16.965 2.16 17.035 ;
    RECT 1.95 17.325 2.16 17.395 ;
    RECT 160.85 16.605 161.06 16.675 ;
    RECT 160.85 16.965 161.06 17.035 ;
    RECT 160.85 17.325 161.06 17.395 ;
    RECT 161.31 16.605 161.52 16.675 ;
    RECT 161.31 16.965 161.52 17.035 ;
    RECT 161.31 17.325 161.52 17.395 ;
    RECT 157.53 16.605 157.74 16.675 ;
    RECT 157.53 16.965 157.74 17.035 ;
    RECT 157.53 17.325 157.74 17.395 ;
    RECT 157.99 16.605 158.2 16.675 ;
    RECT 157.99 16.965 158.2 17.035 ;
    RECT 157.99 17.325 158.2 17.395 ;
    RECT 154.21 16.605 154.42 16.675 ;
    RECT 154.21 16.965 154.42 17.035 ;
    RECT 154.21 17.325 154.42 17.395 ;
    RECT 154.67 16.605 154.88 16.675 ;
    RECT 154.67 16.965 154.88 17.035 ;
    RECT 154.67 17.325 154.88 17.395 ;
    RECT 150.89 16.605 151.1 16.675 ;
    RECT 150.89 16.965 151.1 17.035 ;
    RECT 150.89 17.325 151.1 17.395 ;
    RECT 151.35 16.605 151.56 16.675 ;
    RECT 151.35 16.965 151.56 17.035 ;
    RECT 151.35 17.325 151.56 17.395 ;
    RECT 147.57 16.605 147.78 16.675 ;
    RECT 147.57 16.965 147.78 17.035 ;
    RECT 147.57 17.325 147.78 17.395 ;
    RECT 148.03 16.605 148.24 16.675 ;
    RECT 148.03 16.965 148.24 17.035 ;
    RECT 148.03 17.325 148.24 17.395 ;
    RECT 144.25 16.605 144.46 16.675 ;
    RECT 144.25 16.965 144.46 17.035 ;
    RECT 144.25 17.325 144.46 17.395 ;
    RECT 144.71 16.605 144.92 16.675 ;
    RECT 144.71 16.965 144.92 17.035 ;
    RECT 144.71 17.325 144.92 17.395 ;
    RECT 140.93 16.605 141.14 16.675 ;
    RECT 140.93 16.965 141.14 17.035 ;
    RECT 140.93 17.325 141.14 17.395 ;
    RECT 141.39 16.605 141.6 16.675 ;
    RECT 141.39 16.965 141.6 17.035 ;
    RECT 141.39 17.325 141.6 17.395 ;
    RECT 137.61 16.605 137.82 16.675 ;
    RECT 137.61 16.965 137.82 17.035 ;
    RECT 137.61 17.325 137.82 17.395 ;
    RECT 138.07 16.605 138.28 16.675 ;
    RECT 138.07 16.965 138.28 17.035 ;
    RECT 138.07 17.325 138.28 17.395 ;
    RECT 134.29 16.605 134.5 16.675 ;
    RECT 134.29 16.965 134.5 17.035 ;
    RECT 134.29 17.325 134.5 17.395 ;
    RECT 134.75 16.605 134.96 16.675 ;
    RECT 134.75 16.965 134.96 17.035 ;
    RECT 134.75 17.325 134.96 17.395 ;
    RECT 64.57 16.605 64.78 16.675 ;
    RECT 64.57 16.965 64.78 17.035 ;
    RECT 64.57 17.325 64.78 17.395 ;
    RECT 65.03 16.605 65.24 16.675 ;
    RECT 65.03 16.965 65.24 17.035 ;
    RECT 65.03 17.325 65.24 17.395 ;
    RECT 61.25 15.885 61.46 15.955 ;
    RECT 61.25 16.245 61.46 16.315 ;
    RECT 61.25 16.605 61.46 16.675 ;
    RECT 61.71 15.885 61.92 15.955 ;
    RECT 61.71 16.245 61.92 16.315 ;
    RECT 61.71 16.605 61.92 16.675 ;
    RECT 57.93 15.885 58.14 15.955 ;
    RECT 57.93 16.245 58.14 16.315 ;
    RECT 57.93 16.605 58.14 16.675 ;
    RECT 58.39 15.885 58.6 15.955 ;
    RECT 58.39 16.245 58.6 16.315 ;
    RECT 58.39 16.605 58.6 16.675 ;
    RECT 54.61 15.885 54.82 15.955 ;
    RECT 54.61 16.245 54.82 16.315 ;
    RECT 54.61 16.605 54.82 16.675 ;
    RECT 55.07 15.885 55.28 15.955 ;
    RECT 55.07 16.245 55.28 16.315 ;
    RECT 55.07 16.605 55.28 16.675 ;
    RECT 51.29 15.885 51.5 15.955 ;
    RECT 51.29 16.245 51.5 16.315 ;
    RECT 51.29 16.605 51.5 16.675 ;
    RECT 51.75 15.885 51.96 15.955 ;
    RECT 51.75 16.245 51.96 16.315 ;
    RECT 51.75 16.605 51.96 16.675 ;
    RECT 47.97 15.885 48.18 15.955 ;
    RECT 47.97 16.245 48.18 16.315 ;
    RECT 47.97 16.605 48.18 16.675 ;
    RECT 48.43 15.885 48.64 15.955 ;
    RECT 48.43 16.245 48.64 16.315 ;
    RECT 48.43 16.605 48.64 16.675 ;
    RECT 44.65 15.885 44.86 15.955 ;
    RECT 44.65 16.245 44.86 16.315 ;
    RECT 44.65 16.605 44.86 16.675 ;
    RECT 45.11 15.885 45.32 15.955 ;
    RECT 45.11 16.245 45.32 16.315 ;
    RECT 45.11 16.605 45.32 16.675 ;
    RECT 41.33 15.885 41.54 15.955 ;
    RECT 41.33 16.245 41.54 16.315 ;
    RECT 41.33 16.605 41.54 16.675 ;
    RECT 41.79 15.885 42.0 15.955 ;
    RECT 41.79 16.245 42.0 16.315 ;
    RECT 41.79 16.605 42.0 16.675 ;
    RECT 38.01 15.885 38.22 15.955 ;
    RECT 38.01 16.245 38.22 16.315 ;
    RECT 38.01 16.605 38.22 16.675 ;
    RECT 38.47 15.885 38.68 15.955 ;
    RECT 38.47 16.245 38.68 16.315 ;
    RECT 38.47 16.605 38.68 16.675 ;
    RECT 34.69 15.885 34.9 15.955 ;
    RECT 34.69 16.245 34.9 16.315 ;
    RECT 34.69 16.605 34.9 16.675 ;
    RECT 35.15 15.885 35.36 15.955 ;
    RECT 35.15 16.245 35.36 16.315 ;
    RECT 35.15 16.605 35.36 16.675 ;
    RECT 173.945 16.245 174.015 16.315 ;
    RECT 130.97 15.885 131.18 15.955 ;
    RECT 130.97 16.245 131.18 16.315 ;
    RECT 130.97 16.605 131.18 16.675 ;
    RECT 131.43 15.885 131.64 15.955 ;
    RECT 131.43 16.245 131.64 16.315 ;
    RECT 131.43 16.605 131.64 16.675 ;
    RECT 127.65 15.885 127.86 15.955 ;
    RECT 127.65 16.245 127.86 16.315 ;
    RECT 127.65 16.605 127.86 16.675 ;
    RECT 128.11 15.885 128.32 15.955 ;
    RECT 128.11 16.245 128.32 16.315 ;
    RECT 128.11 16.605 128.32 16.675 ;
    RECT 124.33 15.885 124.54 15.955 ;
    RECT 124.33 16.245 124.54 16.315 ;
    RECT 124.33 16.605 124.54 16.675 ;
    RECT 124.79 15.885 125.0 15.955 ;
    RECT 124.79 16.245 125.0 16.315 ;
    RECT 124.79 16.605 125.0 16.675 ;
    RECT 121.01 15.885 121.22 15.955 ;
    RECT 121.01 16.245 121.22 16.315 ;
    RECT 121.01 16.605 121.22 16.675 ;
    RECT 121.47 15.885 121.68 15.955 ;
    RECT 121.47 16.245 121.68 16.315 ;
    RECT 121.47 16.605 121.68 16.675 ;
    RECT 117.69 15.885 117.9 15.955 ;
    RECT 117.69 16.245 117.9 16.315 ;
    RECT 117.69 16.605 117.9 16.675 ;
    RECT 118.15 15.885 118.36 15.955 ;
    RECT 118.15 16.245 118.36 16.315 ;
    RECT 118.15 16.605 118.36 16.675 ;
    RECT 114.37 15.885 114.58 15.955 ;
    RECT 114.37 16.245 114.58 16.315 ;
    RECT 114.37 16.605 114.58 16.675 ;
    RECT 114.83 15.885 115.04 15.955 ;
    RECT 114.83 16.245 115.04 16.315 ;
    RECT 114.83 16.605 115.04 16.675 ;
    RECT 111.05 15.885 111.26 15.955 ;
    RECT 111.05 16.245 111.26 16.315 ;
    RECT 111.05 16.605 111.26 16.675 ;
    RECT 111.51 15.885 111.72 15.955 ;
    RECT 111.51 16.245 111.72 16.315 ;
    RECT 111.51 16.605 111.72 16.675 ;
    RECT 107.73 15.885 107.94 15.955 ;
    RECT 107.73 16.245 107.94 16.315 ;
    RECT 107.73 16.605 107.94 16.675 ;
    RECT 108.19 15.885 108.4 15.955 ;
    RECT 108.19 16.245 108.4 16.315 ;
    RECT 108.19 16.605 108.4 16.675 ;
    RECT 104.41 15.885 104.62 15.955 ;
    RECT 104.41 16.245 104.62 16.315 ;
    RECT 104.41 16.605 104.62 16.675 ;
    RECT 104.87 15.885 105.08 15.955 ;
    RECT 104.87 16.245 105.08 16.315 ;
    RECT 104.87 16.605 105.08 16.675 ;
    RECT 101.09 15.885 101.3 15.955 ;
    RECT 101.09 16.245 101.3 16.315 ;
    RECT 101.09 16.605 101.3 16.675 ;
    RECT 101.55 15.885 101.76 15.955 ;
    RECT 101.55 16.245 101.76 16.315 ;
    RECT 101.55 16.605 101.76 16.675 ;
    RECT 0.4 16.245 0.47 16.315 ;
    RECT 170.81 15.885 171.02 15.955 ;
    RECT 170.81 16.245 171.02 16.315 ;
    RECT 170.81 16.605 171.02 16.675 ;
    RECT 171.27 15.885 171.48 15.955 ;
    RECT 171.27 16.245 171.48 16.315 ;
    RECT 171.27 16.605 171.48 16.675 ;
    RECT 167.49 15.885 167.7 15.955 ;
    RECT 167.49 16.245 167.7 16.315 ;
    RECT 167.49 16.605 167.7 16.675 ;
    RECT 167.95 15.885 168.16 15.955 ;
    RECT 167.95 16.245 168.16 16.315 ;
    RECT 167.95 16.605 168.16 16.675 ;
    RECT 97.77 15.885 97.98 15.955 ;
    RECT 97.77 16.245 97.98 16.315 ;
    RECT 97.77 16.605 97.98 16.675 ;
    RECT 98.23 15.885 98.44 15.955 ;
    RECT 98.23 16.245 98.44 16.315 ;
    RECT 98.23 16.605 98.44 16.675 ;
    RECT 94.45 15.885 94.66 15.955 ;
    RECT 94.45 16.245 94.66 16.315 ;
    RECT 94.45 16.605 94.66 16.675 ;
    RECT 94.91 15.885 95.12 15.955 ;
    RECT 94.91 16.245 95.12 16.315 ;
    RECT 94.91 16.605 95.12 16.675 ;
    RECT 91.13 15.885 91.34 15.955 ;
    RECT 91.13 16.245 91.34 16.315 ;
    RECT 91.13 16.605 91.34 16.675 ;
    RECT 91.59 15.885 91.8 15.955 ;
    RECT 91.59 16.245 91.8 16.315 ;
    RECT 91.59 16.605 91.8 16.675 ;
    RECT 87.81 15.885 88.02 15.955 ;
    RECT 87.81 16.245 88.02 16.315 ;
    RECT 87.81 16.605 88.02 16.675 ;
    RECT 88.27 15.885 88.48 15.955 ;
    RECT 88.27 16.245 88.48 16.315 ;
    RECT 88.27 16.605 88.48 16.675 ;
    RECT 84.49 15.885 84.7 15.955 ;
    RECT 84.49 16.245 84.7 16.315 ;
    RECT 84.49 16.605 84.7 16.675 ;
    RECT 84.95 15.885 85.16 15.955 ;
    RECT 84.95 16.245 85.16 16.315 ;
    RECT 84.95 16.605 85.16 16.675 ;
    RECT 81.17 15.885 81.38 15.955 ;
    RECT 81.17 16.245 81.38 16.315 ;
    RECT 81.17 16.605 81.38 16.675 ;
    RECT 81.63 15.885 81.84 15.955 ;
    RECT 81.63 16.245 81.84 16.315 ;
    RECT 81.63 16.605 81.84 16.675 ;
    RECT 77.85 15.885 78.06 15.955 ;
    RECT 77.85 16.245 78.06 16.315 ;
    RECT 77.85 16.605 78.06 16.675 ;
    RECT 78.31 15.885 78.52 15.955 ;
    RECT 78.31 16.245 78.52 16.315 ;
    RECT 78.31 16.605 78.52 16.675 ;
    RECT 74.53 15.885 74.74 15.955 ;
    RECT 74.53 16.245 74.74 16.315 ;
    RECT 74.53 16.605 74.74 16.675 ;
    RECT 74.99 15.885 75.2 15.955 ;
    RECT 74.99 16.245 75.2 16.315 ;
    RECT 74.99 16.605 75.2 16.675 ;
    RECT 71.21 15.885 71.42 15.955 ;
    RECT 71.21 16.245 71.42 16.315 ;
    RECT 71.21 16.605 71.42 16.675 ;
    RECT 71.67 15.885 71.88 15.955 ;
    RECT 71.67 16.245 71.88 16.315 ;
    RECT 71.67 16.605 71.88 16.675 ;
    RECT 31.37 15.885 31.58 15.955 ;
    RECT 31.37 16.245 31.58 16.315 ;
    RECT 31.37 16.605 31.58 16.675 ;
    RECT 31.83 15.885 32.04 15.955 ;
    RECT 31.83 16.245 32.04 16.315 ;
    RECT 31.83 16.605 32.04 16.675 ;
    RECT 67.89 15.885 68.1 15.955 ;
    RECT 67.89 16.245 68.1 16.315 ;
    RECT 67.89 16.605 68.1 16.675 ;
    RECT 68.35 15.885 68.56 15.955 ;
    RECT 68.35 16.245 68.56 16.315 ;
    RECT 68.35 16.605 68.56 16.675 ;
    RECT 28.05 15.885 28.26 15.955 ;
    RECT 28.05 16.245 28.26 16.315 ;
    RECT 28.05 16.605 28.26 16.675 ;
    RECT 28.51 15.885 28.72 15.955 ;
    RECT 28.51 16.245 28.72 16.315 ;
    RECT 28.51 16.605 28.72 16.675 ;
    RECT 24.73 15.885 24.94 15.955 ;
    RECT 24.73 16.245 24.94 16.315 ;
    RECT 24.73 16.605 24.94 16.675 ;
    RECT 25.19 15.885 25.4 15.955 ;
    RECT 25.19 16.245 25.4 16.315 ;
    RECT 25.19 16.605 25.4 16.675 ;
    RECT 21.41 15.885 21.62 15.955 ;
    RECT 21.41 16.245 21.62 16.315 ;
    RECT 21.41 16.605 21.62 16.675 ;
    RECT 21.87 15.885 22.08 15.955 ;
    RECT 21.87 16.245 22.08 16.315 ;
    RECT 21.87 16.605 22.08 16.675 ;
    RECT 18.09 15.885 18.3 15.955 ;
    RECT 18.09 16.245 18.3 16.315 ;
    RECT 18.09 16.605 18.3 16.675 ;
    RECT 18.55 15.885 18.76 15.955 ;
    RECT 18.55 16.245 18.76 16.315 ;
    RECT 18.55 16.605 18.76 16.675 ;
    RECT 14.77 15.885 14.98 15.955 ;
    RECT 14.77 16.245 14.98 16.315 ;
    RECT 14.77 16.605 14.98 16.675 ;
    RECT 15.23 15.885 15.44 15.955 ;
    RECT 15.23 16.245 15.44 16.315 ;
    RECT 15.23 16.605 15.44 16.675 ;
    RECT 11.45 15.885 11.66 15.955 ;
    RECT 11.45 16.245 11.66 16.315 ;
    RECT 11.45 16.605 11.66 16.675 ;
    RECT 11.91 15.885 12.12 15.955 ;
    RECT 11.91 16.245 12.12 16.315 ;
    RECT 11.91 16.605 12.12 16.675 ;
    RECT 8.13 15.885 8.34 15.955 ;
    RECT 8.13 16.245 8.34 16.315 ;
    RECT 8.13 16.605 8.34 16.675 ;
    RECT 8.59 15.885 8.8 15.955 ;
    RECT 8.59 16.245 8.8 16.315 ;
    RECT 8.59 16.605 8.8 16.675 ;
    RECT 4.81 15.885 5.02 15.955 ;
    RECT 4.81 16.245 5.02 16.315 ;
    RECT 4.81 16.605 5.02 16.675 ;
    RECT 5.27 15.885 5.48 15.955 ;
    RECT 5.27 16.245 5.48 16.315 ;
    RECT 5.27 16.605 5.48 16.675 ;
    RECT 164.17 15.885 164.38 15.955 ;
    RECT 164.17 16.245 164.38 16.315 ;
    RECT 164.17 16.605 164.38 16.675 ;
    RECT 164.63 15.885 164.84 15.955 ;
    RECT 164.63 16.245 164.84 16.315 ;
    RECT 164.63 16.605 164.84 16.675 ;
    RECT 1.49 15.885 1.7 15.955 ;
    RECT 1.49 16.245 1.7 16.315 ;
    RECT 1.49 16.605 1.7 16.675 ;
    RECT 1.95 15.885 2.16 15.955 ;
    RECT 1.95 16.245 2.16 16.315 ;
    RECT 1.95 16.605 2.16 16.675 ;
    RECT 160.85 15.885 161.06 15.955 ;
    RECT 160.85 16.245 161.06 16.315 ;
    RECT 160.85 16.605 161.06 16.675 ;
    RECT 161.31 15.885 161.52 15.955 ;
    RECT 161.31 16.245 161.52 16.315 ;
    RECT 161.31 16.605 161.52 16.675 ;
    RECT 157.53 15.885 157.74 15.955 ;
    RECT 157.53 16.245 157.74 16.315 ;
    RECT 157.53 16.605 157.74 16.675 ;
    RECT 157.99 15.885 158.2 15.955 ;
    RECT 157.99 16.245 158.2 16.315 ;
    RECT 157.99 16.605 158.2 16.675 ;
    RECT 154.21 15.885 154.42 15.955 ;
    RECT 154.21 16.245 154.42 16.315 ;
    RECT 154.21 16.605 154.42 16.675 ;
    RECT 154.67 15.885 154.88 15.955 ;
    RECT 154.67 16.245 154.88 16.315 ;
    RECT 154.67 16.605 154.88 16.675 ;
    RECT 150.89 15.885 151.1 15.955 ;
    RECT 150.89 16.245 151.1 16.315 ;
    RECT 150.89 16.605 151.1 16.675 ;
    RECT 151.35 15.885 151.56 15.955 ;
    RECT 151.35 16.245 151.56 16.315 ;
    RECT 151.35 16.605 151.56 16.675 ;
    RECT 147.57 15.885 147.78 15.955 ;
    RECT 147.57 16.245 147.78 16.315 ;
    RECT 147.57 16.605 147.78 16.675 ;
    RECT 148.03 15.885 148.24 15.955 ;
    RECT 148.03 16.245 148.24 16.315 ;
    RECT 148.03 16.605 148.24 16.675 ;
    RECT 144.25 15.885 144.46 15.955 ;
    RECT 144.25 16.245 144.46 16.315 ;
    RECT 144.25 16.605 144.46 16.675 ;
    RECT 144.71 15.885 144.92 15.955 ;
    RECT 144.71 16.245 144.92 16.315 ;
    RECT 144.71 16.605 144.92 16.675 ;
    RECT 140.93 15.885 141.14 15.955 ;
    RECT 140.93 16.245 141.14 16.315 ;
    RECT 140.93 16.605 141.14 16.675 ;
    RECT 141.39 15.885 141.6 15.955 ;
    RECT 141.39 16.245 141.6 16.315 ;
    RECT 141.39 16.605 141.6 16.675 ;
    RECT 137.61 15.885 137.82 15.955 ;
    RECT 137.61 16.245 137.82 16.315 ;
    RECT 137.61 16.605 137.82 16.675 ;
    RECT 138.07 15.885 138.28 15.955 ;
    RECT 138.07 16.245 138.28 16.315 ;
    RECT 138.07 16.605 138.28 16.675 ;
    RECT 134.29 15.885 134.5 15.955 ;
    RECT 134.29 16.245 134.5 16.315 ;
    RECT 134.29 16.605 134.5 16.675 ;
    RECT 134.75 15.885 134.96 15.955 ;
    RECT 134.75 16.245 134.96 16.315 ;
    RECT 134.75 16.605 134.96 16.675 ;
    RECT 64.57 15.885 64.78 15.955 ;
    RECT 64.57 16.245 64.78 16.315 ;
    RECT 64.57 16.605 64.78 16.675 ;
    RECT 65.03 15.885 65.24 15.955 ;
    RECT 65.03 16.245 65.24 16.315 ;
    RECT 65.03 16.605 65.24 16.675 ;
    RECT 61.25 46.845 61.46 46.915 ;
    RECT 61.25 47.205 61.46 47.275 ;
    RECT 61.25 47.565 61.46 47.635 ;
    RECT 61.71 46.845 61.92 46.915 ;
    RECT 61.71 47.205 61.92 47.275 ;
    RECT 61.71 47.565 61.92 47.635 ;
    RECT 57.93 46.845 58.14 46.915 ;
    RECT 57.93 47.205 58.14 47.275 ;
    RECT 57.93 47.565 58.14 47.635 ;
    RECT 58.39 46.845 58.6 46.915 ;
    RECT 58.39 47.205 58.6 47.275 ;
    RECT 58.39 47.565 58.6 47.635 ;
    RECT 54.61 46.845 54.82 46.915 ;
    RECT 54.61 47.205 54.82 47.275 ;
    RECT 54.61 47.565 54.82 47.635 ;
    RECT 55.07 46.845 55.28 46.915 ;
    RECT 55.07 47.205 55.28 47.275 ;
    RECT 55.07 47.565 55.28 47.635 ;
    RECT 51.29 46.845 51.5 46.915 ;
    RECT 51.29 47.205 51.5 47.275 ;
    RECT 51.29 47.565 51.5 47.635 ;
    RECT 51.75 46.845 51.96 46.915 ;
    RECT 51.75 47.205 51.96 47.275 ;
    RECT 51.75 47.565 51.96 47.635 ;
    RECT 47.97 46.845 48.18 46.915 ;
    RECT 47.97 47.205 48.18 47.275 ;
    RECT 47.97 47.565 48.18 47.635 ;
    RECT 48.43 46.845 48.64 46.915 ;
    RECT 48.43 47.205 48.64 47.275 ;
    RECT 48.43 47.565 48.64 47.635 ;
    RECT 44.65 46.845 44.86 46.915 ;
    RECT 44.65 47.205 44.86 47.275 ;
    RECT 44.65 47.565 44.86 47.635 ;
    RECT 45.11 46.845 45.32 46.915 ;
    RECT 45.11 47.205 45.32 47.275 ;
    RECT 45.11 47.565 45.32 47.635 ;
    RECT 41.33 46.845 41.54 46.915 ;
    RECT 41.33 47.205 41.54 47.275 ;
    RECT 41.33 47.565 41.54 47.635 ;
    RECT 41.79 46.845 42.0 46.915 ;
    RECT 41.79 47.205 42.0 47.275 ;
    RECT 41.79 47.565 42.0 47.635 ;
    RECT 38.01 46.845 38.22 46.915 ;
    RECT 38.01 47.205 38.22 47.275 ;
    RECT 38.01 47.565 38.22 47.635 ;
    RECT 38.47 46.845 38.68 46.915 ;
    RECT 38.47 47.205 38.68 47.275 ;
    RECT 38.47 47.565 38.68 47.635 ;
    RECT 34.69 46.845 34.9 46.915 ;
    RECT 34.69 47.205 34.9 47.275 ;
    RECT 34.69 47.565 34.9 47.635 ;
    RECT 35.15 46.845 35.36 46.915 ;
    RECT 35.15 47.205 35.36 47.275 ;
    RECT 35.15 47.565 35.36 47.635 ;
    RECT 173.945 47.205 174.015 47.275 ;
    RECT 130.97 46.845 131.18 46.915 ;
    RECT 130.97 47.205 131.18 47.275 ;
    RECT 130.97 47.565 131.18 47.635 ;
    RECT 131.43 46.845 131.64 46.915 ;
    RECT 131.43 47.205 131.64 47.275 ;
    RECT 131.43 47.565 131.64 47.635 ;
    RECT 127.65 46.845 127.86 46.915 ;
    RECT 127.65 47.205 127.86 47.275 ;
    RECT 127.65 47.565 127.86 47.635 ;
    RECT 128.11 46.845 128.32 46.915 ;
    RECT 128.11 47.205 128.32 47.275 ;
    RECT 128.11 47.565 128.32 47.635 ;
    RECT 124.33 46.845 124.54 46.915 ;
    RECT 124.33 47.205 124.54 47.275 ;
    RECT 124.33 47.565 124.54 47.635 ;
    RECT 124.79 46.845 125.0 46.915 ;
    RECT 124.79 47.205 125.0 47.275 ;
    RECT 124.79 47.565 125.0 47.635 ;
    RECT 121.01 46.845 121.22 46.915 ;
    RECT 121.01 47.205 121.22 47.275 ;
    RECT 121.01 47.565 121.22 47.635 ;
    RECT 121.47 46.845 121.68 46.915 ;
    RECT 121.47 47.205 121.68 47.275 ;
    RECT 121.47 47.565 121.68 47.635 ;
    RECT 117.69 46.845 117.9 46.915 ;
    RECT 117.69 47.205 117.9 47.275 ;
    RECT 117.69 47.565 117.9 47.635 ;
    RECT 118.15 46.845 118.36 46.915 ;
    RECT 118.15 47.205 118.36 47.275 ;
    RECT 118.15 47.565 118.36 47.635 ;
    RECT 114.37 46.845 114.58 46.915 ;
    RECT 114.37 47.205 114.58 47.275 ;
    RECT 114.37 47.565 114.58 47.635 ;
    RECT 114.83 46.845 115.04 46.915 ;
    RECT 114.83 47.205 115.04 47.275 ;
    RECT 114.83 47.565 115.04 47.635 ;
    RECT 111.05 46.845 111.26 46.915 ;
    RECT 111.05 47.205 111.26 47.275 ;
    RECT 111.05 47.565 111.26 47.635 ;
    RECT 111.51 46.845 111.72 46.915 ;
    RECT 111.51 47.205 111.72 47.275 ;
    RECT 111.51 47.565 111.72 47.635 ;
    RECT 107.73 46.845 107.94 46.915 ;
    RECT 107.73 47.205 107.94 47.275 ;
    RECT 107.73 47.565 107.94 47.635 ;
    RECT 108.19 46.845 108.4 46.915 ;
    RECT 108.19 47.205 108.4 47.275 ;
    RECT 108.19 47.565 108.4 47.635 ;
    RECT 104.41 46.845 104.62 46.915 ;
    RECT 104.41 47.205 104.62 47.275 ;
    RECT 104.41 47.565 104.62 47.635 ;
    RECT 104.87 46.845 105.08 46.915 ;
    RECT 104.87 47.205 105.08 47.275 ;
    RECT 104.87 47.565 105.08 47.635 ;
    RECT 101.09 46.845 101.3 46.915 ;
    RECT 101.09 47.205 101.3 47.275 ;
    RECT 101.09 47.565 101.3 47.635 ;
    RECT 101.55 46.845 101.76 46.915 ;
    RECT 101.55 47.205 101.76 47.275 ;
    RECT 101.55 47.565 101.76 47.635 ;
    RECT 0.4 47.205 0.47 47.275 ;
    RECT 170.81 46.845 171.02 46.915 ;
    RECT 170.81 47.205 171.02 47.275 ;
    RECT 170.81 47.565 171.02 47.635 ;
    RECT 171.27 46.845 171.48 46.915 ;
    RECT 171.27 47.205 171.48 47.275 ;
    RECT 171.27 47.565 171.48 47.635 ;
    RECT 167.49 46.845 167.7 46.915 ;
    RECT 167.49 47.205 167.7 47.275 ;
    RECT 167.49 47.565 167.7 47.635 ;
    RECT 167.95 46.845 168.16 46.915 ;
    RECT 167.95 47.205 168.16 47.275 ;
    RECT 167.95 47.565 168.16 47.635 ;
    RECT 97.77 46.845 97.98 46.915 ;
    RECT 97.77 47.205 97.98 47.275 ;
    RECT 97.77 47.565 97.98 47.635 ;
    RECT 98.23 46.845 98.44 46.915 ;
    RECT 98.23 47.205 98.44 47.275 ;
    RECT 98.23 47.565 98.44 47.635 ;
    RECT 94.45 46.845 94.66 46.915 ;
    RECT 94.45 47.205 94.66 47.275 ;
    RECT 94.45 47.565 94.66 47.635 ;
    RECT 94.91 46.845 95.12 46.915 ;
    RECT 94.91 47.205 95.12 47.275 ;
    RECT 94.91 47.565 95.12 47.635 ;
    RECT 91.13 46.845 91.34 46.915 ;
    RECT 91.13 47.205 91.34 47.275 ;
    RECT 91.13 47.565 91.34 47.635 ;
    RECT 91.59 46.845 91.8 46.915 ;
    RECT 91.59 47.205 91.8 47.275 ;
    RECT 91.59 47.565 91.8 47.635 ;
    RECT 87.81 46.845 88.02 46.915 ;
    RECT 87.81 47.205 88.02 47.275 ;
    RECT 87.81 47.565 88.02 47.635 ;
    RECT 88.27 46.845 88.48 46.915 ;
    RECT 88.27 47.205 88.48 47.275 ;
    RECT 88.27 47.565 88.48 47.635 ;
    RECT 84.49 46.845 84.7 46.915 ;
    RECT 84.49 47.205 84.7 47.275 ;
    RECT 84.49 47.565 84.7 47.635 ;
    RECT 84.95 46.845 85.16 46.915 ;
    RECT 84.95 47.205 85.16 47.275 ;
    RECT 84.95 47.565 85.16 47.635 ;
    RECT 81.17 46.845 81.38 46.915 ;
    RECT 81.17 47.205 81.38 47.275 ;
    RECT 81.17 47.565 81.38 47.635 ;
    RECT 81.63 46.845 81.84 46.915 ;
    RECT 81.63 47.205 81.84 47.275 ;
    RECT 81.63 47.565 81.84 47.635 ;
    RECT 77.85 46.845 78.06 46.915 ;
    RECT 77.85 47.205 78.06 47.275 ;
    RECT 77.85 47.565 78.06 47.635 ;
    RECT 78.31 46.845 78.52 46.915 ;
    RECT 78.31 47.205 78.52 47.275 ;
    RECT 78.31 47.565 78.52 47.635 ;
    RECT 74.53 46.845 74.74 46.915 ;
    RECT 74.53 47.205 74.74 47.275 ;
    RECT 74.53 47.565 74.74 47.635 ;
    RECT 74.99 46.845 75.2 46.915 ;
    RECT 74.99 47.205 75.2 47.275 ;
    RECT 74.99 47.565 75.2 47.635 ;
    RECT 71.21 46.845 71.42 46.915 ;
    RECT 71.21 47.205 71.42 47.275 ;
    RECT 71.21 47.565 71.42 47.635 ;
    RECT 71.67 46.845 71.88 46.915 ;
    RECT 71.67 47.205 71.88 47.275 ;
    RECT 71.67 47.565 71.88 47.635 ;
    RECT 31.37 46.845 31.58 46.915 ;
    RECT 31.37 47.205 31.58 47.275 ;
    RECT 31.37 47.565 31.58 47.635 ;
    RECT 31.83 46.845 32.04 46.915 ;
    RECT 31.83 47.205 32.04 47.275 ;
    RECT 31.83 47.565 32.04 47.635 ;
    RECT 67.89 46.845 68.1 46.915 ;
    RECT 67.89 47.205 68.1 47.275 ;
    RECT 67.89 47.565 68.1 47.635 ;
    RECT 68.35 46.845 68.56 46.915 ;
    RECT 68.35 47.205 68.56 47.275 ;
    RECT 68.35 47.565 68.56 47.635 ;
    RECT 28.05 46.845 28.26 46.915 ;
    RECT 28.05 47.205 28.26 47.275 ;
    RECT 28.05 47.565 28.26 47.635 ;
    RECT 28.51 46.845 28.72 46.915 ;
    RECT 28.51 47.205 28.72 47.275 ;
    RECT 28.51 47.565 28.72 47.635 ;
    RECT 24.73 46.845 24.94 46.915 ;
    RECT 24.73 47.205 24.94 47.275 ;
    RECT 24.73 47.565 24.94 47.635 ;
    RECT 25.19 46.845 25.4 46.915 ;
    RECT 25.19 47.205 25.4 47.275 ;
    RECT 25.19 47.565 25.4 47.635 ;
    RECT 21.41 46.845 21.62 46.915 ;
    RECT 21.41 47.205 21.62 47.275 ;
    RECT 21.41 47.565 21.62 47.635 ;
    RECT 21.87 46.845 22.08 46.915 ;
    RECT 21.87 47.205 22.08 47.275 ;
    RECT 21.87 47.565 22.08 47.635 ;
    RECT 18.09 46.845 18.3 46.915 ;
    RECT 18.09 47.205 18.3 47.275 ;
    RECT 18.09 47.565 18.3 47.635 ;
    RECT 18.55 46.845 18.76 46.915 ;
    RECT 18.55 47.205 18.76 47.275 ;
    RECT 18.55 47.565 18.76 47.635 ;
    RECT 14.77 46.845 14.98 46.915 ;
    RECT 14.77 47.205 14.98 47.275 ;
    RECT 14.77 47.565 14.98 47.635 ;
    RECT 15.23 46.845 15.44 46.915 ;
    RECT 15.23 47.205 15.44 47.275 ;
    RECT 15.23 47.565 15.44 47.635 ;
    RECT 11.45 46.845 11.66 46.915 ;
    RECT 11.45 47.205 11.66 47.275 ;
    RECT 11.45 47.565 11.66 47.635 ;
    RECT 11.91 46.845 12.12 46.915 ;
    RECT 11.91 47.205 12.12 47.275 ;
    RECT 11.91 47.565 12.12 47.635 ;
    RECT 8.13 46.845 8.34 46.915 ;
    RECT 8.13 47.205 8.34 47.275 ;
    RECT 8.13 47.565 8.34 47.635 ;
    RECT 8.59 46.845 8.8 46.915 ;
    RECT 8.59 47.205 8.8 47.275 ;
    RECT 8.59 47.565 8.8 47.635 ;
    RECT 4.81 46.845 5.02 46.915 ;
    RECT 4.81 47.205 5.02 47.275 ;
    RECT 4.81 47.565 5.02 47.635 ;
    RECT 5.27 46.845 5.48 46.915 ;
    RECT 5.27 47.205 5.48 47.275 ;
    RECT 5.27 47.565 5.48 47.635 ;
    RECT 164.17 46.845 164.38 46.915 ;
    RECT 164.17 47.205 164.38 47.275 ;
    RECT 164.17 47.565 164.38 47.635 ;
    RECT 164.63 46.845 164.84 46.915 ;
    RECT 164.63 47.205 164.84 47.275 ;
    RECT 164.63 47.565 164.84 47.635 ;
    RECT 1.49 46.845 1.7 46.915 ;
    RECT 1.49 47.205 1.7 47.275 ;
    RECT 1.49 47.565 1.7 47.635 ;
    RECT 1.95 46.845 2.16 46.915 ;
    RECT 1.95 47.205 2.16 47.275 ;
    RECT 1.95 47.565 2.16 47.635 ;
    RECT 160.85 46.845 161.06 46.915 ;
    RECT 160.85 47.205 161.06 47.275 ;
    RECT 160.85 47.565 161.06 47.635 ;
    RECT 161.31 46.845 161.52 46.915 ;
    RECT 161.31 47.205 161.52 47.275 ;
    RECT 161.31 47.565 161.52 47.635 ;
    RECT 157.53 46.845 157.74 46.915 ;
    RECT 157.53 47.205 157.74 47.275 ;
    RECT 157.53 47.565 157.74 47.635 ;
    RECT 157.99 46.845 158.2 46.915 ;
    RECT 157.99 47.205 158.2 47.275 ;
    RECT 157.99 47.565 158.2 47.635 ;
    RECT 154.21 46.845 154.42 46.915 ;
    RECT 154.21 47.205 154.42 47.275 ;
    RECT 154.21 47.565 154.42 47.635 ;
    RECT 154.67 46.845 154.88 46.915 ;
    RECT 154.67 47.205 154.88 47.275 ;
    RECT 154.67 47.565 154.88 47.635 ;
    RECT 150.89 46.845 151.1 46.915 ;
    RECT 150.89 47.205 151.1 47.275 ;
    RECT 150.89 47.565 151.1 47.635 ;
    RECT 151.35 46.845 151.56 46.915 ;
    RECT 151.35 47.205 151.56 47.275 ;
    RECT 151.35 47.565 151.56 47.635 ;
    RECT 147.57 46.845 147.78 46.915 ;
    RECT 147.57 47.205 147.78 47.275 ;
    RECT 147.57 47.565 147.78 47.635 ;
    RECT 148.03 46.845 148.24 46.915 ;
    RECT 148.03 47.205 148.24 47.275 ;
    RECT 148.03 47.565 148.24 47.635 ;
    RECT 144.25 46.845 144.46 46.915 ;
    RECT 144.25 47.205 144.46 47.275 ;
    RECT 144.25 47.565 144.46 47.635 ;
    RECT 144.71 46.845 144.92 46.915 ;
    RECT 144.71 47.205 144.92 47.275 ;
    RECT 144.71 47.565 144.92 47.635 ;
    RECT 140.93 46.845 141.14 46.915 ;
    RECT 140.93 47.205 141.14 47.275 ;
    RECT 140.93 47.565 141.14 47.635 ;
    RECT 141.39 46.845 141.6 46.915 ;
    RECT 141.39 47.205 141.6 47.275 ;
    RECT 141.39 47.565 141.6 47.635 ;
    RECT 137.61 46.845 137.82 46.915 ;
    RECT 137.61 47.205 137.82 47.275 ;
    RECT 137.61 47.565 137.82 47.635 ;
    RECT 138.07 46.845 138.28 46.915 ;
    RECT 138.07 47.205 138.28 47.275 ;
    RECT 138.07 47.565 138.28 47.635 ;
    RECT 134.29 46.845 134.5 46.915 ;
    RECT 134.29 47.205 134.5 47.275 ;
    RECT 134.29 47.565 134.5 47.635 ;
    RECT 134.75 46.845 134.96 46.915 ;
    RECT 134.75 47.205 134.96 47.275 ;
    RECT 134.75 47.565 134.96 47.635 ;
    RECT 64.57 46.845 64.78 46.915 ;
    RECT 64.57 47.205 64.78 47.275 ;
    RECT 64.57 47.565 64.78 47.635 ;
    RECT 65.03 46.845 65.24 46.915 ;
    RECT 65.03 47.205 65.24 47.275 ;
    RECT 65.03 47.565 65.24 47.635 ;
    RECT 61.25 15.165 61.46 15.235 ;
    RECT 61.25 15.525 61.46 15.595 ;
    RECT 61.25 15.885 61.46 15.955 ;
    RECT 61.71 15.165 61.92 15.235 ;
    RECT 61.71 15.525 61.92 15.595 ;
    RECT 61.71 15.885 61.92 15.955 ;
    RECT 57.93 15.165 58.14 15.235 ;
    RECT 57.93 15.525 58.14 15.595 ;
    RECT 57.93 15.885 58.14 15.955 ;
    RECT 58.39 15.165 58.6 15.235 ;
    RECT 58.39 15.525 58.6 15.595 ;
    RECT 58.39 15.885 58.6 15.955 ;
    RECT 54.61 15.165 54.82 15.235 ;
    RECT 54.61 15.525 54.82 15.595 ;
    RECT 54.61 15.885 54.82 15.955 ;
    RECT 55.07 15.165 55.28 15.235 ;
    RECT 55.07 15.525 55.28 15.595 ;
    RECT 55.07 15.885 55.28 15.955 ;
    RECT 51.29 15.165 51.5 15.235 ;
    RECT 51.29 15.525 51.5 15.595 ;
    RECT 51.29 15.885 51.5 15.955 ;
    RECT 51.75 15.165 51.96 15.235 ;
    RECT 51.75 15.525 51.96 15.595 ;
    RECT 51.75 15.885 51.96 15.955 ;
    RECT 47.97 15.165 48.18 15.235 ;
    RECT 47.97 15.525 48.18 15.595 ;
    RECT 47.97 15.885 48.18 15.955 ;
    RECT 48.43 15.165 48.64 15.235 ;
    RECT 48.43 15.525 48.64 15.595 ;
    RECT 48.43 15.885 48.64 15.955 ;
    RECT 44.65 15.165 44.86 15.235 ;
    RECT 44.65 15.525 44.86 15.595 ;
    RECT 44.65 15.885 44.86 15.955 ;
    RECT 45.11 15.165 45.32 15.235 ;
    RECT 45.11 15.525 45.32 15.595 ;
    RECT 45.11 15.885 45.32 15.955 ;
    RECT 41.33 15.165 41.54 15.235 ;
    RECT 41.33 15.525 41.54 15.595 ;
    RECT 41.33 15.885 41.54 15.955 ;
    RECT 41.79 15.165 42.0 15.235 ;
    RECT 41.79 15.525 42.0 15.595 ;
    RECT 41.79 15.885 42.0 15.955 ;
    RECT 38.01 15.165 38.22 15.235 ;
    RECT 38.01 15.525 38.22 15.595 ;
    RECT 38.01 15.885 38.22 15.955 ;
    RECT 38.47 15.165 38.68 15.235 ;
    RECT 38.47 15.525 38.68 15.595 ;
    RECT 38.47 15.885 38.68 15.955 ;
    RECT 34.69 15.165 34.9 15.235 ;
    RECT 34.69 15.525 34.9 15.595 ;
    RECT 34.69 15.885 34.9 15.955 ;
    RECT 35.15 15.165 35.36 15.235 ;
    RECT 35.15 15.525 35.36 15.595 ;
    RECT 35.15 15.885 35.36 15.955 ;
    RECT 173.945 15.525 174.015 15.595 ;
    RECT 130.97 15.165 131.18 15.235 ;
    RECT 130.97 15.525 131.18 15.595 ;
    RECT 130.97 15.885 131.18 15.955 ;
    RECT 131.43 15.165 131.64 15.235 ;
    RECT 131.43 15.525 131.64 15.595 ;
    RECT 131.43 15.885 131.64 15.955 ;
    RECT 127.65 15.165 127.86 15.235 ;
    RECT 127.65 15.525 127.86 15.595 ;
    RECT 127.65 15.885 127.86 15.955 ;
    RECT 128.11 15.165 128.32 15.235 ;
    RECT 128.11 15.525 128.32 15.595 ;
    RECT 128.11 15.885 128.32 15.955 ;
    RECT 124.33 15.165 124.54 15.235 ;
    RECT 124.33 15.525 124.54 15.595 ;
    RECT 124.33 15.885 124.54 15.955 ;
    RECT 124.79 15.165 125.0 15.235 ;
    RECT 124.79 15.525 125.0 15.595 ;
    RECT 124.79 15.885 125.0 15.955 ;
    RECT 121.01 15.165 121.22 15.235 ;
    RECT 121.01 15.525 121.22 15.595 ;
    RECT 121.01 15.885 121.22 15.955 ;
    RECT 121.47 15.165 121.68 15.235 ;
    RECT 121.47 15.525 121.68 15.595 ;
    RECT 121.47 15.885 121.68 15.955 ;
    RECT 117.69 15.165 117.9 15.235 ;
    RECT 117.69 15.525 117.9 15.595 ;
    RECT 117.69 15.885 117.9 15.955 ;
    RECT 118.15 15.165 118.36 15.235 ;
    RECT 118.15 15.525 118.36 15.595 ;
    RECT 118.15 15.885 118.36 15.955 ;
    RECT 114.37 15.165 114.58 15.235 ;
    RECT 114.37 15.525 114.58 15.595 ;
    RECT 114.37 15.885 114.58 15.955 ;
    RECT 114.83 15.165 115.04 15.235 ;
    RECT 114.83 15.525 115.04 15.595 ;
    RECT 114.83 15.885 115.04 15.955 ;
    RECT 111.05 15.165 111.26 15.235 ;
    RECT 111.05 15.525 111.26 15.595 ;
    RECT 111.05 15.885 111.26 15.955 ;
    RECT 111.51 15.165 111.72 15.235 ;
    RECT 111.51 15.525 111.72 15.595 ;
    RECT 111.51 15.885 111.72 15.955 ;
    RECT 107.73 15.165 107.94 15.235 ;
    RECT 107.73 15.525 107.94 15.595 ;
    RECT 107.73 15.885 107.94 15.955 ;
    RECT 108.19 15.165 108.4 15.235 ;
    RECT 108.19 15.525 108.4 15.595 ;
    RECT 108.19 15.885 108.4 15.955 ;
    RECT 104.41 15.165 104.62 15.235 ;
    RECT 104.41 15.525 104.62 15.595 ;
    RECT 104.41 15.885 104.62 15.955 ;
    RECT 104.87 15.165 105.08 15.235 ;
    RECT 104.87 15.525 105.08 15.595 ;
    RECT 104.87 15.885 105.08 15.955 ;
    RECT 101.09 15.165 101.3 15.235 ;
    RECT 101.09 15.525 101.3 15.595 ;
    RECT 101.09 15.885 101.3 15.955 ;
    RECT 101.55 15.165 101.76 15.235 ;
    RECT 101.55 15.525 101.76 15.595 ;
    RECT 101.55 15.885 101.76 15.955 ;
    RECT 0.4 15.525 0.47 15.595 ;
    RECT 170.81 15.165 171.02 15.235 ;
    RECT 170.81 15.525 171.02 15.595 ;
    RECT 170.81 15.885 171.02 15.955 ;
    RECT 171.27 15.165 171.48 15.235 ;
    RECT 171.27 15.525 171.48 15.595 ;
    RECT 171.27 15.885 171.48 15.955 ;
    RECT 167.49 15.165 167.7 15.235 ;
    RECT 167.49 15.525 167.7 15.595 ;
    RECT 167.49 15.885 167.7 15.955 ;
    RECT 167.95 15.165 168.16 15.235 ;
    RECT 167.95 15.525 168.16 15.595 ;
    RECT 167.95 15.885 168.16 15.955 ;
    RECT 97.77 15.165 97.98 15.235 ;
    RECT 97.77 15.525 97.98 15.595 ;
    RECT 97.77 15.885 97.98 15.955 ;
    RECT 98.23 15.165 98.44 15.235 ;
    RECT 98.23 15.525 98.44 15.595 ;
    RECT 98.23 15.885 98.44 15.955 ;
    RECT 94.45 15.165 94.66 15.235 ;
    RECT 94.45 15.525 94.66 15.595 ;
    RECT 94.45 15.885 94.66 15.955 ;
    RECT 94.91 15.165 95.12 15.235 ;
    RECT 94.91 15.525 95.12 15.595 ;
    RECT 94.91 15.885 95.12 15.955 ;
    RECT 91.13 15.165 91.34 15.235 ;
    RECT 91.13 15.525 91.34 15.595 ;
    RECT 91.13 15.885 91.34 15.955 ;
    RECT 91.59 15.165 91.8 15.235 ;
    RECT 91.59 15.525 91.8 15.595 ;
    RECT 91.59 15.885 91.8 15.955 ;
    RECT 87.81 15.165 88.02 15.235 ;
    RECT 87.81 15.525 88.02 15.595 ;
    RECT 87.81 15.885 88.02 15.955 ;
    RECT 88.27 15.165 88.48 15.235 ;
    RECT 88.27 15.525 88.48 15.595 ;
    RECT 88.27 15.885 88.48 15.955 ;
    RECT 84.49 15.165 84.7 15.235 ;
    RECT 84.49 15.525 84.7 15.595 ;
    RECT 84.49 15.885 84.7 15.955 ;
    RECT 84.95 15.165 85.16 15.235 ;
    RECT 84.95 15.525 85.16 15.595 ;
    RECT 84.95 15.885 85.16 15.955 ;
    RECT 81.17 15.165 81.38 15.235 ;
    RECT 81.17 15.525 81.38 15.595 ;
    RECT 81.17 15.885 81.38 15.955 ;
    RECT 81.63 15.165 81.84 15.235 ;
    RECT 81.63 15.525 81.84 15.595 ;
    RECT 81.63 15.885 81.84 15.955 ;
    RECT 77.85 15.165 78.06 15.235 ;
    RECT 77.85 15.525 78.06 15.595 ;
    RECT 77.85 15.885 78.06 15.955 ;
    RECT 78.31 15.165 78.52 15.235 ;
    RECT 78.31 15.525 78.52 15.595 ;
    RECT 78.31 15.885 78.52 15.955 ;
    RECT 74.53 15.165 74.74 15.235 ;
    RECT 74.53 15.525 74.74 15.595 ;
    RECT 74.53 15.885 74.74 15.955 ;
    RECT 74.99 15.165 75.2 15.235 ;
    RECT 74.99 15.525 75.2 15.595 ;
    RECT 74.99 15.885 75.2 15.955 ;
    RECT 71.21 15.165 71.42 15.235 ;
    RECT 71.21 15.525 71.42 15.595 ;
    RECT 71.21 15.885 71.42 15.955 ;
    RECT 71.67 15.165 71.88 15.235 ;
    RECT 71.67 15.525 71.88 15.595 ;
    RECT 71.67 15.885 71.88 15.955 ;
    RECT 31.37 15.165 31.58 15.235 ;
    RECT 31.37 15.525 31.58 15.595 ;
    RECT 31.37 15.885 31.58 15.955 ;
    RECT 31.83 15.165 32.04 15.235 ;
    RECT 31.83 15.525 32.04 15.595 ;
    RECT 31.83 15.885 32.04 15.955 ;
    RECT 67.89 15.165 68.1 15.235 ;
    RECT 67.89 15.525 68.1 15.595 ;
    RECT 67.89 15.885 68.1 15.955 ;
    RECT 68.35 15.165 68.56 15.235 ;
    RECT 68.35 15.525 68.56 15.595 ;
    RECT 68.35 15.885 68.56 15.955 ;
    RECT 28.05 15.165 28.26 15.235 ;
    RECT 28.05 15.525 28.26 15.595 ;
    RECT 28.05 15.885 28.26 15.955 ;
    RECT 28.51 15.165 28.72 15.235 ;
    RECT 28.51 15.525 28.72 15.595 ;
    RECT 28.51 15.885 28.72 15.955 ;
    RECT 24.73 15.165 24.94 15.235 ;
    RECT 24.73 15.525 24.94 15.595 ;
    RECT 24.73 15.885 24.94 15.955 ;
    RECT 25.19 15.165 25.4 15.235 ;
    RECT 25.19 15.525 25.4 15.595 ;
    RECT 25.19 15.885 25.4 15.955 ;
    RECT 21.41 15.165 21.62 15.235 ;
    RECT 21.41 15.525 21.62 15.595 ;
    RECT 21.41 15.885 21.62 15.955 ;
    RECT 21.87 15.165 22.08 15.235 ;
    RECT 21.87 15.525 22.08 15.595 ;
    RECT 21.87 15.885 22.08 15.955 ;
    RECT 18.09 15.165 18.3 15.235 ;
    RECT 18.09 15.525 18.3 15.595 ;
    RECT 18.09 15.885 18.3 15.955 ;
    RECT 18.55 15.165 18.76 15.235 ;
    RECT 18.55 15.525 18.76 15.595 ;
    RECT 18.55 15.885 18.76 15.955 ;
    RECT 14.77 15.165 14.98 15.235 ;
    RECT 14.77 15.525 14.98 15.595 ;
    RECT 14.77 15.885 14.98 15.955 ;
    RECT 15.23 15.165 15.44 15.235 ;
    RECT 15.23 15.525 15.44 15.595 ;
    RECT 15.23 15.885 15.44 15.955 ;
    RECT 11.45 15.165 11.66 15.235 ;
    RECT 11.45 15.525 11.66 15.595 ;
    RECT 11.45 15.885 11.66 15.955 ;
    RECT 11.91 15.165 12.12 15.235 ;
    RECT 11.91 15.525 12.12 15.595 ;
    RECT 11.91 15.885 12.12 15.955 ;
    RECT 8.13 15.165 8.34 15.235 ;
    RECT 8.13 15.525 8.34 15.595 ;
    RECT 8.13 15.885 8.34 15.955 ;
    RECT 8.59 15.165 8.8 15.235 ;
    RECT 8.59 15.525 8.8 15.595 ;
    RECT 8.59 15.885 8.8 15.955 ;
    RECT 4.81 15.165 5.02 15.235 ;
    RECT 4.81 15.525 5.02 15.595 ;
    RECT 4.81 15.885 5.02 15.955 ;
    RECT 5.27 15.165 5.48 15.235 ;
    RECT 5.27 15.525 5.48 15.595 ;
    RECT 5.27 15.885 5.48 15.955 ;
    RECT 164.17 15.165 164.38 15.235 ;
    RECT 164.17 15.525 164.38 15.595 ;
    RECT 164.17 15.885 164.38 15.955 ;
    RECT 164.63 15.165 164.84 15.235 ;
    RECT 164.63 15.525 164.84 15.595 ;
    RECT 164.63 15.885 164.84 15.955 ;
    RECT 1.49 15.165 1.7 15.235 ;
    RECT 1.49 15.525 1.7 15.595 ;
    RECT 1.49 15.885 1.7 15.955 ;
    RECT 1.95 15.165 2.16 15.235 ;
    RECT 1.95 15.525 2.16 15.595 ;
    RECT 1.95 15.885 2.16 15.955 ;
    RECT 160.85 15.165 161.06 15.235 ;
    RECT 160.85 15.525 161.06 15.595 ;
    RECT 160.85 15.885 161.06 15.955 ;
    RECT 161.31 15.165 161.52 15.235 ;
    RECT 161.31 15.525 161.52 15.595 ;
    RECT 161.31 15.885 161.52 15.955 ;
    RECT 157.53 15.165 157.74 15.235 ;
    RECT 157.53 15.525 157.74 15.595 ;
    RECT 157.53 15.885 157.74 15.955 ;
    RECT 157.99 15.165 158.2 15.235 ;
    RECT 157.99 15.525 158.2 15.595 ;
    RECT 157.99 15.885 158.2 15.955 ;
    RECT 154.21 15.165 154.42 15.235 ;
    RECT 154.21 15.525 154.42 15.595 ;
    RECT 154.21 15.885 154.42 15.955 ;
    RECT 154.67 15.165 154.88 15.235 ;
    RECT 154.67 15.525 154.88 15.595 ;
    RECT 154.67 15.885 154.88 15.955 ;
    RECT 150.89 15.165 151.1 15.235 ;
    RECT 150.89 15.525 151.1 15.595 ;
    RECT 150.89 15.885 151.1 15.955 ;
    RECT 151.35 15.165 151.56 15.235 ;
    RECT 151.35 15.525 151.56 15.595 ;
    RECT 151.35 15.885 151.56 15.955 ;
    RECT 147.57 15.165 147.78 15.235 ;
    RECT 147.57 15.525 147.78 15.595 ;
    RECT 147.57 15.885 147.78 15.955 ;
    RECT 148.03 15.165 148.24 15.235 ;
    RECT 148.03 15.525 148.24 15.595 ;
    RECT 148.03 15.885 148.24 15.955 ;
    RECT 144.25 15.165 144.46 15.235 ;
    RECT 144.25 15.525 144.46 15.595 ;
    RECT 144.25 15.885 144.46 15.955 ;
    RECT 144.71 15.165 144.92 15.235 ;
    RECT 144.71 15.525 144.92 15.595 ;
    RECT 144.71 15.885 144.92 15.955 ;
    RECT 140.93 15.165 141.14 15.235 ;
    RECT 140.93 15.525 141.14 15.595 ;
    RECT 140.93 15.885 141.14 15.955 ;
    RECT 141.39 15.165 141.6 15.235 ;
    RECT 141.39 15.525 141.6 15.595 ;
    RECT 141.39 15.885 141.6 15.955 ;
    RECT 137.61 15.165 137.82 15.235 ;
    RECT 137.61 15.525 137.82 15.595 ;
    RECT 137.61 15.885 137.82 15.955 ;
    RECT 138.07 15.165 138.28 15.235 ;
    RECT 138.07 15.525 138.28 15.595 ;
    RECT 138.07 15.885 138.28 15.955 ;
    RECT 134.29 15.165 134.5 15.235 ;
    RECT 134.29 15.525 134.5 15.595 ;
    RECT 134.29 15.885 134.5 15.955 ;
    RECT 134.75 15.165 134.96 15.235 ;
    RECT 134.75 15.525 134.96 15.595 ;
    RECT 134.75 15.885 134.96 15.955 ;
    RECT 64.57 15.165 64.78 15.235 ;
    RECT 64.57 15.525 64.78 15.595 ;
    RECT 64.57 15.885 64.78 15.955 ;
    RECT 65.03 15.165 65.24 15.235 ;
    RECT 65.03 15.525 65.24 15.595 ;
    RECT 65.03 15.885 65.24 15.955 ;
    RECT 61.25 46.125 61.46 46.195 ;
    RECT 61.25 46.485 61.46 46.555 ;
    RECT 61.25 46.845 61.46 46.915 ;
    RECT 61.71 46.125 61.92 46.195 ;
    RECT 61.71 46.485 61.92 46.555 ;
    RECT 61.71 46.845 61.92 46.915 ;
    RECT 57.93 46.125 58.14 46.195 ;
    RECT 57.93 46.485 58.14 46.555 ;
    RECT 57.93 46.845 58.14 46.915 ;
    RECT 58.39 46.125 58.6 46.195 ;
    RECT 58.39 46.485 58.6 46.555 ;
    RECT 58.39 46.845 58.6 46.915 ;
    RECT 54.61 46.125 54.82 46.195 ;
    RECT 54.61 46.485 54.82 46.555 ;
    RECT 54.61 46.845 54.82 46.915 ;
    RECT 55.07 46.125 55.28 46.195 ;
    RECT 55.07 46.485 55.28 46.555 ;
    RECT 55.07 46.845 55.28 46.915 ;
    RECT 51.29 46.125 51.5 46.195 ;
    RECT 51.29 46.485 51.5 46.555 ;
    RECT 51.29 46.845 51.5 46.915 ;
    RECT 51.75 46.125 51.96 46.195 ;
    RECT 51.75 46.485 51.96 46.555 ;
    RECT 51.75 46.845 51.96 46.915 ;
    RECT 47.97 46.125 48.18 46.195 ;
    RECT 47.97 46.485 48.18 46.555 ;
    RECT 47.97 46.845 48.18 46.915 ;
    RECT 48.43 46.125 48.64 46.195 ;
    RECT 48.43 46.485 48.64 46.555 ;
    RECT 48.43 46.845 48.64 46.915 ;
    RECT 44.65 46.125 44.86 46.195 ;
    RECT 44.65 46.485 44.86 46.555 ;
    RECT 44.65 46.845 44.86 46.915 ;
    RECT 45.11 46.125 45.32 46.195 ;
    RECT 45.11 46.485 45.32 46.555 ;
    RECT 45.11 46.845 45.32 46.915 ;
    RECT 41.33 46.125 41.54 46.195 ;
    RECT 41.33 46.485 41.54 46.555 ;
    RECT 41.33 46.845 41.54 46.915 ;
    RECT 41.79 46.125 42.0 46.195 ;
    RECT 41.79 46.485 42.0 46.555 ;
    RECT 41.79 46.845 42.0 46.915 ;
    RECT 38.01 46.125 38.22 46.195 ;
    RECT 38.01 46.485 38.22 46.555 ;
    RECT 38.01 46.845 38.22 46.915 ;
    RECT 38.47 46.125 38.68 46.195 ;
    RECT 38.47 46.485 38.68 46.555 ;
    RECT 38.47 46.845 38.68 46.915 ;
    RECT 34.69 46.125 34.9 46.195 ;
    RECT 34.69 46.485 34.9 46.555 ;
    RECT 34.69 46.845 34.9 46.915 ;
    RECT 35.15 46.125 35.36 46.195 ;
    RECT 35.15 46.485 35.36 46.555 ;
    RECT 35.15 46.845 35.36 46.915 ;
    RECT 173.945 46.485 174.015 46.555 ;
    RECT 130.97 46.125 131.18 46.195 ;
    RECT 130.97 46.485 131.18 46.555 ;
    RECT 130.97 46.845 131.18 46.915 ;
    RECT 131.43 46.125 131.64 46.195 ;
    RECT 131.43 46.485 131.64 46.555 ;
    RECT 131.43 46.845 131.64 46.915 ;
    RECT 127.65 46.125 127.86 46.195 ;
    RECT 127.65 46.485 127.86 46.555 ;
    RECT 127.65 46.845 127.86 46.915 ;
    RECT 128.11 46.125 128.32 46.195 ;
    RECT 128.11 46.485 128.32 46.555 ;
    RECT 128.11 46.845 128.32 46.915 ;
    RECT 124.33 46.125 124.54 46.195 ;
    RECT 124.33 46.485 124.54 46.555 ;
    RECT 124.33 46.845 124.54 46.915 ;
    RECT 124.79 46.125 125.0 46.195 ;
    RECT 124.79 46.485 125.0 46.555 ;
    RECT 124.79 46.845 125.0 46.915 ;
    RECT 121.01 46.125 121.22 46.195 ;
    RECT 121.01 46.485 121.22 46.555 ;
    RECT 121.01 46.845 121.22 46.915 ;
    RECT 121.47 46.125 121.68 46.195 ;
    RECT 121.47 46.485 121.68 46.555 ;
    RECT 121.47 46.845 121.68 46.915 ;
    RECT 117.69 46.125 117.9 46.195 ;
    RECT 117.69 46.485 117.9 46.555 ;
    RECT 117.69 46.845 117.9 46.915 ;
    RECT 118.15 46.125 118.36 46.195 ;
    RECT 118.15 46.485 118.36 46.555 ;
    RECT 118.15 46.845 118.36 46.915 ;
    RECT 114.37 46.125 114.58 46.195 ;
    RECT 114.37 46.485 114.58 46.555 ;
    RECT 114.37 46.845 114.58 46.915 ;
    RECT 114.83 46.125 115.04 46.195 ;
    RECT 114.83 46.485 115.04 46.555 ;
    RECT 114.83 46.845 115.04 46.915 ;
    RECT 111.05 46.125 111.26 46.195 ;
    RECT 111.05 46.485 111.26 46.555 ;
    RECT 111.05 46.845 111.26 46.915 ;
    RECT 111.51 46.125 111.72 46.195 ;
    RECT 111.51 46.485 111.72 46.555 ;
    RECT 111.51 46.845 111.72 46.915 ;
    RECT 107.73 46.125 107.94 46.195 ;
    RECT 107.73 46.485 107.94 46.555 ;
    RECT 107.73 46.845 107.94 46.915 ;
    RECT 108.19 46.125 108.4 46.195 ;
    RECT 108.19 46.485 108.4 46.555 ;
    RECT 108.19 46.845 108.4 46.915 ;
    RECT 104.41 46.125 104.62 46.195 ;
    RECT 104.41 46.485 104.62 46.555 ;
    RECT 104.41 46.845 104.62 46.915 ;
    RECT 104.87 46.125 105.08 46.195 ;
    RECT 104.87 46.485 105.08 46.555 ;
    RECT 104.87 46.845 105.08 46.915 ;
    RECT 101.09 46.125 101.3 46.195 ;
    RECT 101.09 46.485 101.3 46.555 ;
    RECT 101.09 46.845 101.3 46.915 ;
    RECT 101.55 46.125 101.76 46.195 ;
    RECT 101.55 46.485 101.76 46.555 ;
    RECT 101.55 46.845 101.76 46.915 ;
    RECT 0.4 46.485 0.47 46.555 ;
    RECT 170.81 46.125 171.02 46.195 ;
    RECT 170.81 46.485 171.02 46.555 ;
    RECT 170.81 46.845 171.02 46.915 ;
    RECT 171.27 46.125 171.48 46.195 ;
    RECT 171.27 46.485 171.48 46.555 ;
    RECT 171.27 46.845 171.48 46.915 ;
    RECT 167.49 46.125 167.7 46.195 ;
    RECT 167.49 46.485 167.7 46.555 ;
    RECT 167.49 46.845 167.7 46.915 ;
    RECT 167.95 46.125 168.16 46.195 ;
    RECT 167.95 46.485 168.16 46.555 ;
    RECT 167.95 46.845 168.16 46.915 ;
    RECT 97.77 46.125 97.98 46.195 ;
    RECT 97.77 46.485 97.98 46.555 ;
    RECT 97.77 46.845 97.98 46.915 ;
    RECT 98.23 46.125 98.44 46.195 ;
    RECT 98.23 46.485 98.44 46.555 ;
    RECT 98.23 46.845 98.44 46.915 ;
    RECT 94.45 46.125 94.66 46.195 ;
    RECT 94.45 46.485 94.66 46.555 ;
    RECT 94.45 46.845 94.66 46.915 ;
    RECT 94.91 46.125 95.12 46.195 ;
    RECT 94.91 46.485 95.12 46.555 ;
    RECT 94.91 46.845 95.12 46.915 ;
    RECT 91.13 46.125 91.34 46.195 ;
    RECT 91.13 46.485 91.34 46.555 ;
    RECT 91.13 46.845 91.34 46.915 ;
    RECT 91.59 46.125 91.8 46.195 ;
    RECT 91.59 46.485 91.8 46.555 ;
    RECT 91.59 46.845 91.8 46.915 ;
    RECT 87.81 46.125 88.02 46.195 ;
    RECT 87.81 46.485 88.02 46.555 ;
    RECT 87.81 46.845 88.02 46.915 ;
    RECT 88.27 46.125 88.48 46.195 ;
    RECT 88.27 46.485 88.48 46.555 ;
    RECT 88.27 46.845 88.48 46.915 ;
    RECT 84.49 46.125 84.7 46.195 ;
    RECT 84.49 46.485 84.7 46.555 ;
    RECT 84.49 46.845 84.7 46.915 ;
    RECT 84.95 46.125 85.16 46.195 ;
    RECT 84.95 46.485 85.16 46.555 ;
    RECT 84.95 46.845 85.16 46.915 ;
    RECT 81.17 46.125 81.38 46.195 ;
    RECT 81.17 46.485 81.38 46.555 ;
    RECT 81.17 46.845 81.38 46.915 ;
    RECT 81.63 46.125 81.84 46.195 ;
    RECT 81.63 46.485 81.84 46.555 ;
    RECT 81.63 46.845 81.84 46.915 ;
    RECT 77.85 46.125 78.06 46.195 ;
    RECT 77.85 46.485 78.06 46.555 ;
    RECT 77.85 46.845 78.06 46.915 ;
    RECT 78.31 46.125 78.52 46.195 ;
    RECT 78.31 46.485 78.52 46.555 ;
    RECT 78.31 46.845 78.52 46.915 ;
    RECT 74.53 46.125 74.74 46.195 ;
    RECT 74.53 46.485 74.74 46.555 ;
    RECT 74.53 46.845 74.74 46.915 ;
    RECT 74.99 46.125 75.2 46.195 ;
    RECT 74.99 46.485 75.2 46.555 ;
    RECT 74.99 46.845 75.2 46.915 ;
    RECT 71.21 46.125 71.42 46.195 ;
    RECT 71.21 46.485 71.42 46.555 ;
    RECT 71.21 46.845 71.42 46.915 ;
    RECT 71.67 46.125 71.88 46.195 ;
    RECT 71.67 46.485 71.88 46.555 ;
    RECT 71.67 46.845 71.88 46.915 ;
    RECT 31.37 46.125 31.58 46.195 ;
    RECT 31.37 46.485 31.58 46.555 ;
    RECT 31.37 46.845 31.58 46.915 ;
    RECT 31.83 46.125 32.04 46.195 ;
    RECT 31.83 46.485 32.04 46.555 ;
    RECT 31.83 46.845 32.04 46.915 ;
    RECT 67.89 46.125 68.1 46.195 ;
    RECT 67.89 46.485 68.1 46.555 ;
    RECT 67.89 46.845 68.1 46.915 ;
    RECT 68.35 46.125 68.56 46.195 ;
    RECT 68.35 46.485 68.56 46.555 ;
    RECT 68.35 46.845 68.56 46.915 ;
    RECT 28.05 46.125 28.26 46.195 ;
    RECT 28.05 46.485 28.26 46.555 ;
    RECT 28.05 46.845 28.26 46.915 ;
    RECT 28.51 46.125 28.72 46.195 ;
    RECT 28.51 46.485 28.72 46.555 ;
    RECT 28.51 46.845 28.72 46.915 ;
    RECT 24.73 46.125 24.94 46.195 ;
    RECT 24.73 46.485 24.94 46.555 ;
    RECT 24.73 46.845 24.94 46.915 ;
    RECT 25.19 46.125 25.4 46.195 ;
    RECT 25.19 46.485 25.4 46.555 ;
    RECT 25.19 46.845 25.4 46.915 ;
    RECT 21.41 46.125 21.62 46.195 ;
    RECT 21.41 46.485 21.62 46.555 ;
    RECT 21.41 46.845 21.62 46.915 ;
    RECT 21.87 46.125 22.08 46.195 ;
    RECT 21.87 46.485 22.08 46.555 ;
    RECT 21.87 46.845 22.08 46.915 ;
    RECT 18.09 46.125 18.3 46.195 ;
    RECT 18.09 46.485 18.3 46.555 ;
    RECT 18.09 46.845 18.3 46.915 ;
    RECT 18.55 46.125 18.76 46.195 ;
    RECT 18.55 46.485 18.76 46.555 ;
    RECT 18.55 46.845 18.76 46.915 ;
    RECT 14.77 46.125 14.98 46.195 ;
    RECT 14.77 46.485 14.98 46.555 ;
    RECT 14.77 46.845 14.98 46.915 ;
    RECT 15.23 46.125 15.44 46.195 ;
    RECT 15.23 46.485 15.44 46.555 ;
    RECT 15.23 46.845 15.44 46.915 ;
    RECT 11.45 46.125 11.66 46.195 ;
    RECT 11.45 46.485 11.66 46.555 ;
    RECT 11.45 46.845 11.66 46.915 ;
    RECT 11.91 46.125 12.12 46.195 ;
    RECT 11.91 46.485 12.12 46.555 ;
    RECT 11.91 46.845 12.12 46.915 ;
    RECT 8.13 46.125 8.34 46.195 ;
    RECT 8.13 46.485 8.34 46.555 ;
    RECT 8.13 46.845 8.34 46.915 ;
    RECT 8.59 46.125 8.8 46.195 ;
    RECT 8.59 46.485 8.8 46.555 ;
    RECT 8.59 46.845 8.8 46.915 ;
    RECT 4.81 46.125 5.02 46.195 ;
    RECT 4.81 46.485 5.02 46.555 ;
    RECT 4.81 46.845 5.02 46.915 ;
    RECT 5.27 46.125 5.48 46.195 ;
    RECT 5.27 46.485 5.48 46.555 ;
    RECT 5.27 46.845 5.48 46.915 ;
    RECT 164.17 46.125 164.38 46.195 ;
    RECT 164.17 46.485 164.38 46.555 ;
    RECT 164.17 46.845 164.38 46.915 ;
    RECT 164.63 46.125 164.84 46.195 ;
    RECT 164.63 46.485 164.84 46.555 ;
    RECT 164.63 46.845 164.84 46.915 ;
    RECT 1.49 46.125 1.7 46.195 ;
    RECT 1.49 46.485 1.7 46.555 ;
    RECT 1.49 46.845 1.7 46.915 ;
    RECT 1.95 46.125 2.16 46.195 ;
    RECT 1.95 46.485 2.16 46.555 ;
    RECT 1.95 46.845 2.16 46.915 ;
    RECT 160.85 46.125 161.06 46.195 ;
    RECT 160.85 46.485 161.06 46.555 ;
    RECT 160.85 46.845 161.06 46.915 ;
    RECT 161.31 46.125 161.52 46.195 ;
    RECT 161.31 46.485 161.52 46.555 ;
    RECT 161.31 46.845 161.52 46.915 ;
    RECT 157.53 46.125 157.74 46.195 ;
    RECT 157.53 46.485 157.74 46.555 ;
    RECT 157.53 46.845 157.74 46.915 ;
    RECT 157.99 46.125 158.2 46.195 ;
    RECT 157.99 46.485 158.2 46.555 ;
    RECT 157.99 46.845 158.2 46.915 ;
    RECT 154.21 46.125 154.42 46.195 ;
    RECT 154.21 46.485 154.42 46.555 ;
    RECT 154.21 46.845 154.42 46.915 ;
    RECT 154.67 46.125 154.88 46.195 ;
    RECT 154.67 46.485 154.88 46.555 ;
    RECT 154.67 46.845 154.88 46.915 ;
    RECT 150.89 46.125 151.1 46.195 ;
    RECT 150.89 46.485 151.1 46.555 ;
    RECT 150.89 46.845 151.1 46.915 ;
    RECT 151.35 46.125 151.56 46.195 ;
    RECT 151.35 46.485 151.56 46.555 ;
    RECT 151.35 46.845 151.56 46.915 ;
    RECT 147.57 46.125 147.78 46.195 ;
    RECT 147.57 46.485 147.78 46.555 ;
    RECT 147.57 46.845 147.78 46.915 ;
    RECT 148.03 46.125 148.24 46.195 ;
    RECT 148.03 46.485 148.24 46.555 ;
    RECT 148.03 46.845 148.24 46.915 ;
    RECT 144.25 46.125 144.46 46.195 ;
    RECT 144.25 46.485 144.46 46.555 ;
    RECT 144.25 46.845 144.46 46.915 ;
    RECT 144.71 46.125 144.92 46.195 ;
    RECT 144.71 46.485 144.92 46.555 ;
    RECT 144.71 46.845 144.92 46.915 ;
    RECT 140.93 46.125 141.14 46.195 ;
    RECT 140.93 46.485 141.14 46.555 ;
    RECT 140.93 46.845 141.14 46.915 ;
    RECT 141.39 46.125 141.6 46.195 ;
    RECT 141.39 46.485 141.6 46.555 ;
    RECT 141.39 46.845 141.6 46.915 ;
    RECT 137.61 46.125 137.82 46.195 ;
    RECT 137.61 46.485 137.82 46.555 ;
    RECT 137.61 46.845 137.82 46.915 ;
    RECT 138.07 46.125 138.28 46.195 ;
    RECT 138.07 46.485 138.28 46.555 ;
    RECT 138.07 46.845 138.28 46.915 ;
    RECT 134.29 46.125 134.5 46.195 ;
    RECT 134.29 46.485 134.5 46.555 ;
    RECT 134.29 46.845 134.5 46.915 ;
    RECT 134.75 46.125 134.96 46.195 ;
    RECT 134.75 46.485 134.96 46.555 ;
    RECT 134.75 46.845 134.96 46.915 ;
    RECT 64.57 46.125 64.78 46.195 ;
    RECT 64.57 46.485 64.78 46.555 ;
    RECT 64.57 46.845 64.78 46.915 ;
    RECT 65.03 46.125 65.24 46.195 ;
    RECT 65.03 46.485 65.24 46.555 ;
    RECT 65.03 46.845 65.24 46.915 ;
    RECT 61.25 14.445 61.46 14.515 ;
    RECT 61.25 14.805 61.46 14.875 ;
    RECT 61.25 15.165 61.46 15.235 ;
    RECT 61.71 14.445 61.92 14.515 ;
    RECT 61.71 14.805 61.92 14.875 ;
    RECT 61.71 15.165 61.92 15.235 ;
    RECT 57.93 14.445 58.14 14.515 ;
    RECT 57.93 14.805 58.14 14.875 ;
    RECT 57.93 15.165 58.14 15.235 ;
    RECT 58.39 14.445 58.6 14.515 ;
    RECT 58.39 14.805 58.6 14.875 ;
    RECT 58.39 15.165 58.6 15.235 ;
    RECT 54.61 14.445 54.82 14.515 ;
    RECT 54.61 14.805 54.82 14.875 ;
    RECT 54.61 15.165 54.82 15.235 ;
    RECT 55.07 14.445 55.28 14.515 ;
    RECT 55.07 14.805 55.28 14.875 ;
    RECT 55.07 15.165 55.28 15.235 ;
    RECT 51.29 14.445 51.5 14.515 ;
    RECT 51.29 14.805 51.5 14.875 ;
    RECT 51.29 15.165 51.5 15.235 ;
    RECT 51.75 14.445 51.96 14.515 ;
    RECT 51.75 14.805 51.96 14.875 ;
    RECT 51.75 15.165 51.96 15.235 ;
    RECT 47.97 14.445 48.18 14.515 ;
    RECT 47.97 14.805 48.18 14.875 ;
    RECT 47.97 15.165 48.18 15.235 ;
    RECT 48.43 14.445 48.64 14.515 ;
    RECT 48.43 14.805 48.64 14.875 ;
    RECT 48.43 15.165 48.64 15.235 ;
    RECT 44.65 14.445 44.86 14.515 ;
    RECT 44.65 14.805 44.86 14.875 ;
    RECT 44.65 15.165 44.86 15.235 ;
    RECT 45.11 14.445 45.32 14.515 ;
    RECT 45.11 14.805 45.32 14.875 ;
    RECT 45.11 15.165 45.32 15.235 ;
    RECT 41.33 14.445 41.54 14.515 ;
    RECT 41.33 14.805 41.54 14.875 ;
    RECT 41.33 15.165 41.54 15.235 ;
    RECT 41.79 14.445 42.0 14.515 ;
    RECT 41.79 14.805 42.0 14.875 ;
    RECT 41.79 15.165 42.0 15.235 ;
    RECT 38.01 14.445 38.22 14.515 ;
    RECT 38.01 14.805 38.22 14.875 ;
    RECT 38.01 15.165 38.22 15.235 ;
    RECT 38.47 14.445 38.68 14.515 ;
    RECT 38.47 14.805 38.68 14.875 ;
    RECT 38.47 15.165 38.68 15.235 ;
    RECT 34.69 14.445 34.9 14.515 ;
    RECT 34.69 14.805 34.9 14.875 ;
    RECT 34.69 15.165 34.9 15.235 ;
    RECT 35.15 14.445 35.36 14.515 ;
    RECT 35.15 14.805 35.36 14.875 ;
    RECT 35.15 15.165 35.36 15.235 ;
    RECT 173.945 14.805 174.015 14.875 ;
    RECT 130.97 14.445 131.18 14.515 ;
    RECT 130.97 14.805 131.18 14.875 ;
    RECT 130.97 15.165 131.18 15.235 ;
    RECT 131.43 14.445 131.64 14.515 ;
    RECT 131.43 14.805 131.64 14.875 ;
    RECT 131.43 15.165 131.64 15.235 ;
    RECT 127.65 14.445 127.86 14.515 ;
    RECT 127.65 14.805 127.86 14.875 ;
    RECT 127.65 15.165 127.86 15.235 ;
    RECT 128.11 14.445 128.32 14.515 ;
    RECT 128.11 14.805 128.32 14.875 ;
    RECT 128.11 15.165 128.32 15.235 ;
    RECT 124.33 14.445 124.54 14.515 ;
    RECT 124.33 14.805 124.54 14.875 ;
    RECT 124.33 15.165 124.54 15.235 ;
    RECT 124.79 14.445 125.0 14.515 ;
    RECT 124.79 14.805 125.0 14.875 ;
    RECT 124.79 15.165 125.0 15.235 ;
    RECT 121.01 14.445 121.22 14.515 ;
    RECT 121.01 14.805 121.22 14.875 ;
    RECT 121.01 15.165 121.22 15.235 ;
    RECT 121.47 14.445 121.68 14.515 ;
    RECT 121.47 14.805 121.68 14.875 ;
    RECT 121.47 15.165 121.68 15.235 ;
    RECT 117.69 14.445 117.9 14.515 ;
    RECT 117.69 14.805 117.9 14.875 ;
    RECT 117.69 15.165 117.9 15.235 ;
    RECT 118.15 14.445 118.36 14.515 ;
    RECT 118.15 14.805 118.36 14.875 ;
    RECT 118.15 15.165 118.36 15.235 ;
    RECT 114.37 14.445 114.58 14.515 ;
    RECT 114.37 14.805 114.58 14.875 ;
    RECT 114.37 15.165 114.58 15.235 ;
    RECT 114.83 14.445 115.04 14.515 ;
    RECT 114.83 14.805 115.04 14.875 ;
    RECT 114.83 15.165 115.04 15.235 ;
    RECT 111.05 14.445 111.26 14.515 ;
    RECT 111.05 14.805 111.26 14.875 ;
    RECT 111.05 15.165 111.26 15.235 ;
    RECT 111.51 14.445 111.72 14.515 ;
    RECT 111.51 14.805 111.72 14.875 ;
    RECT 111.51 15.165 111.72 15.235 ;
    RECT 107.73 14.445 107.94 14.515 ;
    RECT 107.73 14.805 107.94 14.875 ;
    RECT 107.73 15.165 107.94 15.235 ;
    RECT 108.19 14.445 108.4 14.515 ;
    RECT 108.19 14.805 108.4 14.875 ;
    RECT 108.19 15.165 108.4 15.235 ;
    RECT 104.41 14.445 104.62 14.515 ;
    RECT 104.41 14.805 104.62 14.875 ;
    RECT 104.41 15.165 104.62 15.235 ;
    RECT 104.87 14.445 105.08 14.515 ;
    RECT 104.87 14.805 105.08 14.875 ;
    RECT 104.87 15.165 105.08 15.235 ;
    RECT 101.09 14.445 101.3 14.515 ;
    RECT 101.09 14.805 101.3 14.875 ;
    RECT 101.09 15.165 101.3 15.235 ;
    RECT 101.55 14.445 101.76 14.515 ;
    RECT 101.55 14.805 101.76 14.875 ;
    RECT 101.55 15.165 101.76 15.235 ;
    RECT 0.4 14.805 0.47 14.875 ;
    RECT 170.81 14.445 171.02 14.515 ;
    RECT 170.81 14.805 171.02 14.875 ;
    RECT 170.81 15.165 171.02 15.235 ;
    RECT 171.27 14.445 171.48 14.515 ;
    RECT 171.27 14.805 171.48 14.875 ;
    RECT 171.27 15.165 171.48 15.235 ;
    RECT 167.49 14.445 167.7 14.515 ;
    RECT 167.49 14.805 167.7 14.875 ;
    RECT 167.49 15.165 167.7 15.235 ;
    RECT 167.95 14.445 168.16 14.515 ;
    RECT 167.95 14.805 168.16 14.875 ;
    RECT 167.95 15.165 168.16 15.235 ;
    RECT 97.77 14.445 97.98 14.515 ;
    RECT 97.77 14.805 97.98 14.875 ;
    RECT 97.77 15.165 97.98 15.235 ;
    RECT 98.23 14.445 98.44 14.515 ;
    RECT 98.23 14.805 98.44 14.875 ;
    RECT 98.23 15.165 98.44 15.235 ;
    RECT 94.45 14.445 94.66 14.515 ;
    RECT 94.45 14.805 94.66 14.875 ;
    RECT 94.45 15.165 94.66 15.235 ;
    RECT 94.91 14.445 95.12 14.515 ;
    RECT 94.91 14.805 95.12 14.875 ;
    RECT 94.91 15.165 95.12 15.235 ;
    RECT 91.13 14.445 91.34 14.515 ;
    RECT 91.13 14.805 91.34 14.875 ;
    RECT 91.13 15.165 91.34 15.235 ;
    RECT 91.59 14.445 91.8 14.515 ;
    RECT 91.59 14.805 91.8 14.875 ;
    RECT 91.59 15.165 91.8 15.235 ;
    RECT 87.81 14.445 88.02 14.515 ;
    RECT 87.81 14.805 88.02 14.875 ;
    RECT 87.81 15.165 88.02 15.235 ;
    RECT 88.27 14.445 88.48 14.515 ;
    RECT 88.27 14.805 88.48 14.875 ;
    RECT 88.27 15.165 88.48 15.235 ;
    RECT 84.49 14.445 84.7 14.515 ;
    RECT 84.49 14.805 84.7 14.875 ;
    RECT 84.49 15.165 84.7 15.235 ;
    RECT 84.95 14.445 85.16 14.515 ;
    RECT 84.95 14.805 85.16 14.875 ;
    RECT 84.95 15.165 85.16 15.235 ;
    RECT 81.17 14.445 81.38 14.515 ;
    RECT 81.17 14.805 81.38 14.875 ;
    RECT 81.17 15.165 81.38 15.235 ;
    RECT 81.63 14.445 81.84 14.515 ;
    RECT 81.63 14.805 81.84 14.875 ;
    RECT 81.63 15.165 81.84 15.235 ;
    RECT 77.85 14.445 78.06 14.515 ;
    RECT 77.85 14.805 78.06 14.875 ;
    RECT 77.85 15.165 78.06 15.235 ;
    RECT 78.31 14.445 78.52 14.515 ;
    RECT 78.31 14.805 78.52 14.875 ;
    RECT 78.31 15.165 78.52 15.235 ;
    RECT 74.53 14.445 74.74 14.515 ;
    RECT 74.53 14.805 74.74 14.875 ;
    RECT 74.53 15.165 74.74 15.235 ;
    RECT 74.99 14.445 75.2 14.515 ;
    RECT 74.99 14.805 75.2 14.875 ;
    RECT 74.99 15.165 75.2 15.235 ;
    RECT 71.21 14.445 71.42 14.515 ;
    RECT 71.21 14.805 71.42 14.875 ;
    RECT 71.21 15.165 71.42 15.235 ;
    RECT 71.67 14.445 71.88 14.515 ;
    RECT 71.67 14.805 71.88 14.875 ;
    RECT 71.67 15.165 71.88 15.235 ;
    RECT 31.37 14.445 31.58 14.515 ;
    RECT 31.37 14.805 31.58 14.875 ;
    RECT 31.37 15.165 31.58 15.235 ;
    RECT 31.83 14.445 32.04 14.515 ;
    RECT 31.83 14.805 32.04 14.875 ;
    RECT 31.83 15.165 32.04 15.235 ;
    RECT 67.89 14.445 68.1 14.515 ;
    RECT 67.89 14.805 68.1 14.875 ;
    RECT 67.89 15.165 68.1 15.235 ;
    RECT 68.35 14.445 68.56 14.515 ;
    RECT 68.35 14.805 68.56 14.875 ;
    RECT 68.35 15.165 68.56 15.235 ;
    RECT 28.05 14.445 28.26 14.515 ;
    RECT 28.05 14.805 28.26 14.875 ;
    RECT 28.05 15.165 28.26 15.235 ;
    RECT 28.51 14.445 28.72 14.515 ;
    RECT 28.51 14.805 28.72 14.875 ;
    RECT 28.51 15.165 28.72 15.235 ;
    RECT 24.73 14.445 24.94 14.515 ;
    RECT 24.73 14.805 24.94 14.875 ;
    RECT 24.73 15.165 24.94 15.235 ;
    RECT 25.19 14.445 25.4 14.515 ;
    RECT 25.19 14.805 25.4 14.875 ;
    RECT 25.19 15.165 25.4 15.235 ;
    RECT 21.41 14.445 21.62 14.515 ;
    RECT 21.41 14.805 21.62 14.875 ;
    RECT 21.41 15.165 21.62 15.235 ;
    RECT 21.87 14.445 22.08 14.515 ;
    RECT 21.87 14.805 22.08 14.875 ;
    RECT 21.87 15.165 22.08 15.235 ;
    RECT 18.09 14.445 18.3 14.515 ;
    RECT 18.09 14.805 18.3 14.875 ;
    RECT 18.09 15.165 18.3 15.235 ;
    RECT 18.55 14.445 18.76 14.515 ;
    RECT 18.55 14.805 18.76 14.875 ;
    RECT 18.55 15.165 18.76 15.235 ;
    RECT 14.77 14.445 14.98 14.515 ;
    RECT 14.77 14.805 14.98 14.875 ;
    RECT 14.77 15.165 14.98 15.235 ;
    RECT 15.23 14.445 15.44 14.515 ;
    RECT 15.23 14.805 15.44 14.875 ;
    RECT 15.23 15.165 15.44 15.235 ;
    RECT 11.45 14.445 11.66 14.515 ;
    RECT 11.45 14.805 11.66 14.875 ;
    RECT 11.45 15.165 11.66 15.235 ;
    RECT 11.91 14.445 12.12 14.515 ;
    RECT 11.91 14.805 12.12 14.875 ;
    RECT 11.91 15.165 12.12 15.235 ;
    RECT 8.13 14.445 8.34 14.515 ;
    RECT 8.13 14.805 8.34 14.875 ;
    RECT 8.13 15.165 8.34 15.235 ;
    RECT 8.59 14.445 8.8 14.515 ;
    RECT 8.59 14.805 8.8 14.875 ;
    RECT 8.59 15.165 8.8 15.235 ;
    RECT 4.81 14.445 5.02 14.515 ;
    RECT 4.81 14.805 5.02 14.875 ;
    RECT 4.81 15.165 5.02 15.235 ;
    RECT 5.27 14.445 5.48 14.515 ;
    RECT 5.27 14.805 5.48 14.875 ;
    RECT 5.27 15.165 5.48 15.235 ;
    RECT 164.17 14.445 164.38 14.515 ;
    RECT 164.17 14.805 164.38 14.875 ;
    RECT 164.17 15.165 164.38 15.235 ;
    RECT 164.63 14.445 164.84 14.515 ;
    RECT 164.63 14.805 164.84 14.875 ;
    RECT 164.63 15.165 164.84 15.235 ;
    RECT 1.49 14.445 1.7 14.515 ;
    RECT 1.49 14.805 1.7 14.875 ;
    RECT 1.49 15.165 1.7 15.235 ;
    RECT 1.95 14.445 2.16 14.515 ;
    RECT 1.95 14.805 2.16 14.875 ;
    RECT 1.95 15.165 2.16 15.235 ;
    RECT 160.85 14.445 161.06 14.515 ;
    RECT 160.85 14.805 161.06 14.875 ;
    RECT 160.85 15.165 161.06 15.235 ;
    RECT 161.31 14.445 161.52 14.515 ;
    RECT 161.31 14.805 161.52 14.875 ;
    RECT 161.31 15.165 161.52 15.235 ;
    RECT 157.53 14.445 157.74 14.515 ;
    RECT 157.53 14.805 157.74 14.875 ;
    RECT 157.53 15.165 157.74 15.235 ;
    RECT 157.99 14.445 158.2 14.515 ;
    RECT 157.99 14.805 158.2 14.875 ;
    RECT 157.99 15.165 158.2 15.235 ;
    RECT 154.21 14.445 154.42 14.515 ;
    RECT 154.21 14.805 154.42 14.875 ;
    RECT 154.21 15.165 154.42 15.235 ;
    RECT 154.67 14.445 154.88 14.515 ;
    RECT 154.67 14.805 154.88 14.875 ;
    RECT 154.67 15.165 154.88 15.235 ;
    RECT 150.89 14.445 151.1 14.515 ;
    RECT 150.89 14.805 151.1 14.875 ;
    RECT 150.89 15.165 151.1 15.235 ;
    RECT 151.35 14.445 151.56 14.515 ;
    RECT 151.35 14.805 151.56 14.875 ;
    RECT 151.35 15.165 151.56 15.235 ;
    RECT 147.57 14.445 147.78 14.515 ;
    RECT 147.57 14.805 147.78 14.875 ;
    RECT 147.57 15.165 147.78 15.235 ;
    RECT 148.03 14.445 148.24 14.515 ;
    RECT 148.03 14.805 148.24 14.875 ;
    RECT 148.03 15.165 148.24 15.235 ;
    RECT 144.25 14.445 144.46 14.515 ;
    RECT 144.25 14.805 144.46 14.875 ;
    RECT 144.25 15.165 144.46 15.235 ;
    RECT 144.71 14.445 144.92 14.515 ;
    RECT 144.71 14.805 144.92 14.875 ;
    RECT 144.71 15.165 144.92 15.235 ;
    RECT 140.93 14.445 141.14 14.515 ;
    RECT 140.93 14.805 141.14 14.875 ;
    RECT 140.93 15.165 141.14 15.235 ;
    RECT 141.39 14.445 141.6 14.515 ;
    RECT 141.39 14.805 141.6 14.875 ;
    RECT 141.39 15.165 141.6 15.235 ;
    RECT 137.61 14.445 137.82 14.515 ;
    RECT 137.61 14.805 137.82 14.875 ;
    RECT 137.61 15.165 137.82 15.235 ;
    RECT 138.07 14.445 138.28 14.515 ;
    RECT 138.07 14.805 138.28 14.875 ;
    RECT 138.07 15.165 138.28 15.235 ;
    RECT 134.29 14.445 134.5 14.515 ;
    RECT 134.29 14.805 134.5 14.875 ;
    RECT 134.29 15.165 134.5 15.235 ;
    RECT 134.75 14.445 134.96 14.515 ;
    RECT 134.75 14.805 134.96 14.875 ;
    RECT 134.75 15.165 134.96 15.235 ;
    RECT 64.57 14.445 64.78 14.515 ;
    RECT 64.57 14.805 64.78 14.875 ;
    RECT 64.57 15.165 64.78 15.235 ;
    RECT 65.03 14.445 65.24 14.515 ;
    RECT 65.03 14.805 65.24 14.875 ;
    RECT 65.03 15.165 65.24 15.235 ;
    RECT 61.25 45.405 61.46 45.475 ;
    RECT 61.25 45.765 61.46 45.835 ;
    RECT 61.25 46.125 61.46 46.195 ;
    RECT 61.71 45.405 61.92 45.475 ;
    RECT 61.71 45.765 61.92 45.835 ;
    RECT 61.71 46.125 61.92 46.195 ;
    RECT 57.93 45.405 58.14 45.475 ;
    RECT 57.93 45.765 58.14 45.835 ;
    RECT 57.93 46.125 58.14 46.195 ;
    RECT 58.39 45.405 58.6 45.475 ;
    RECT 58.39 45.765 58.6 45.835 ;
    RECT 58.39 46.125 58.6 46.195 ;
    RECT 54.61 45.405 54.82 45.475 ;
    RECT 54.61 45.765 54.82 45.835 ;
    RECT 54.61 46.125 54.82 46.195 ;
    RECT 55.07 45.405 55.28 45.475 ;
    RECT 55.07 45.765 55.28 45.835 ;
    RECT 55.07 46.125 55.28 46.195 ;
    RECT 51.29 45.405 51.5 45.475 ;
    RECT 51.29 45.765 51.5 45.835 ;
    RECT 51.29 46.125 51.5 46.195 ;
    RECT 51.75 45.405 51.96 45.475 ;
    RECT 51.75 45.765 51.96 45.835 ;
    RECT 51.75 46.125 51.96 46.195 ;
    RECT 47.97 45.405 48.18 45.475 ;
    RECT 47.97 45.765 48.18 45.835 ;
    RECT 47.97 46.125 48.18 46.195 ;
    RECT 48.43 45.405 48.64 45.475 ;
    RECT 48.43 45.765 48.64 45.835 ;
    RECT 48.43 46.125 48.64 46.195 ;
    RECT 44.65 45.405 44.86 45.475 ;
    RECT 44.65 45.765 44.86 45.835 ;
    RECT 44.65 46.125 44.86 46.195 ;
    RECT 45.11 45.405 45.32 45.475 ;
    RECT 45.11 45.765 45.32 45.835 ;
    RECT 45.11 46.125 45.32 46.195 ;
    RECT 41.33 45.405 41.54 45.475 ;
    RECT 41.33 45.765 41.54 45.835 ;
    RECT 41.33 46.125 41.54 46.195 ;
    RECT 41.79 45.405 42.0 45.475 ;
    RECT 41.79 45.765 42.0 45.835 ;
    RECT 41.79 46.125 42.0 46.195 ;
    RECT 38.01 45.405 38.22 45.475 ;
    RECT 38.01 45.765 38.22 45.835 ;
    RECT 38.01 46.125 38.22 46.195 ;
    RECT 38.47 45.405 38.68 45.475 ;
    RECT 38.47 45.765 38.68 45.835 ;
    RECT 38.47 46.125 38.68 46.195 ;
    RECT 34.69 45.405 34.9 45.475 ;
    RECT 34.69 45.765 34.9 45.835 ;
    RECT 34.69 46.125 34.9 46.195 ;
    RECT 35.15 45.405 35.36 45.475 ;
    RECT 35.15 45.765 35.36 45.835 ;
    RECT 35.15 46.125 35.36 46.195 ;
    RECT 173.945 45.765 174.015 45.835 ;
    RECT 130.97 45.405 131.18 45.475 ;
    RECT 130.97 45.765 131.18 45.835 ;
    RECT 130.97 46.125 131.18 46.195 ;
    RECT 131.43 45.405 131.64 45.475 ;
    RECT 131.43 45.765 131.64 45.835 ;
    RECT 131.43 46.125 131.64 46.195 ;
    RECT 127.65 45.405 127.86 45.475 ;
    RECT 127.65 45.765 127.86 45.835 ;
    RECT 127.65 46.125 127.86 46.195 ;
    RECT 128.11 45.405 128.32 45.475 ;
    RECT 128.11 45.765 128.32 45.835 ;
    RECT 128.11 46.125 128.32 46.195 ;
    RECT 124.33 45.405 124.54 45.475 ;
    RECT 124.33 45.765 124.54 45.835 ;
    RECT 124.33 46.125 124.54 46.195 ;
    RECT 124.79 45.405 125.0 45.475 ;
    RECT 124.79 45.765 125.0 45.835 ;
    RECT 124.79 46.125 125.0 46.195 ;
    RECT 121.01 45.405 121.22 45.475 ;
    RECT 121.01 45.765 121.22 45.835 ;
    RECT 121.01 46.125 121.22 46.195 ;
    RECT 121.47 45.405 121.68 45.475 ;
    RECT 121.47 45.765 121.68 45.835 ;
    RECT 121.47 46.125 121.68 46.195 ;
    RECT 117.69 45.405 117.9 45.475 ;
    RECT 117.69 45.765 117.9 45.835 ;
    RECT 117.69 46.125 117.9 46.195 ;
    RECT 118.15 45.405 118.36 45.475 ;
    RECT 118.15 45.765 118.36 45.835 ;
    RECT 118.15 46.125 118.36 46.195 ;
    RECT 114.37 45.405 114.58 45.475 ;
    RECT 114.37 45.765 114.58 45.835 ;
    RECT 114.37 46.125 114.58 46.195 ;
    RECT 114.83 45.405 115.04 45.475 ;
    RECT 114.83 45.765 115.04 45.835 ;
    RECT 114.83 46.125 115.04 46.195 ;
    RECT 111.05 45.405 111.26 45.475 ;
    RECT 111.05 45.765 111.26 45.835 ;
    RECT 111.05 46.125 111.26 46.195 ;
    RECT 111.51 45.405 111.72 45.475 ;
    RECT 111.51 45.765 111.72 45.835 ;
    RECT 111.51 46.125 111.72 46.195 ;
    RECT 107.73 45.405 107.94 45.475 ;
    RECT 107.73 45.765 107.94 45.835 ;
    RECT 107.73 46.125 107.94 46.195 ;
    RECT 108.19 45.405 108.4 45.475 ;
    RECT 108.19 45.765 108.4 45.835 ;
    RECT 108.19 46.125 108.4 46.195 ;
    RECT 104.41 45.405 104.62 45.475 ;
    RECT 104.41 45.765 104.62 45.835 ;
    RECT 104.41 46.125 104.62 46.195 ;
    RECT 104.87 45.405 105.08 45.475 ;
    RECT 104.87 45.765 105.08 45.835 ;
    RECT 104.87 46.125 105.08 46.195 ;
    RECT 101.09 45.405 101.3 45.475 ;
    RECT 101.09 45.765 101.3 45.835 ;
    RECT 101.09 46.125 101.3 46.195 ;
    RECT 101.55 45.405 101.76 45.475 ;
    RECT 101.55 45.765 101.76 45.835 ;
    RECT 101.55 46.125 101.76 46.195 ;
    RECT 0.4 45.765 0.47 45.835 ;
    RECT 170.81 45.405 171.02 45.475 ;
    RECT 170.81 45.765 171.02 45.835 ;
    RECT 170.81 46.125 171.02 46.195 ;
    RECT 171.27 45.405 171.48 45.475 ;
    RECT 171.27 45.765 171.48 45.835 ;
    RECT 171.27 46.125 171.48 46.195 ;
    RECT 167.49 45.405 167.7 45.475 ;
    RECT 167.49 45.765 167.7 45.835 ;
    RECT 167.49 46.125 167.7 46.195 ;
    RECT 167.95 45.405 168.16 45.475 ;
    RECT 167.95 45.765 168.16 45.835 ;
    RECT 167.95 46.125 168.16 46.195 ;
    RECT 97.77 45.405 97.98 45.475 ;
    RECT 97.77 45.765 97.98 45.835 ;
    RECT 97.77 46.125 97.98 46.195 ;
    RECT 98.23 45.405 98.44 45.475 ;
    RECT 98.23 45.765 98.44 45.835 ;
    RECT 98.23 46.125 98.44 46.195 ;
    RECT 94.45 45.405 94.66 45.475 ;
    RECT 94.45 45.765 94.66 45.835 ;
    RECT 94.45 46.125 94.66 46.195 ;
    RECT 94.91 45.405 95.12 45.475 ;
    RECT 94.91 45.765 95.12 45.835 ;
    RECT 94.91 46.125 95.12 46.195 ;
    RECT 91.13 45.405 91.34 45.475 ;
    RECT 91.13 45.765 91.34 45.835 ;
    RECT 91.13 46.125 91.34 46.195 ;
    RECT 91.59 45.405 91.8 45.475 ;
    RECT 91.59 45.765 91.8 45.835 ;
    RECT 91.59 46.125 91.8 46.195 ;
    RECT 87.81 45.405 88.02 45.475 ;
    RECT 87.81 45.765 88.02 45.835 ;
    RECT 87.81 46.125 88.02 46.195 ;
    RECT 88.27 45.405 88.48 45.475 ;
    RECT 88.27 45.765 88.48 45.835 ;
    RECT 88.27 46.125 88.48 46.195 ;
    RECT 84.49 45.405 84.7 45.475 ;
    RECT 84.49 45.765 84.7 45.835 ;
    RECT 84.49 46.125 84.7 46.195 ;
    RECT 84.95 45.405 85.16 45.475 ;
    RECT 84.95 45.765 85.16 45.835 ;
    RECT 84.95 46.125 85.16 46.195 ;
    RECT 81.17 45.405 81.38 45.475 ;
    RECT 81.17 45.765 81.38 45.835 ;
    RECT 81.17 46.125 81.38 46.195 ;
    RECT 81.63 45.405 81.84 45.475 ;
    RECT 81.63 45.765 81.84 45.835 ;
    RECT 81.63 46.125 81.84 46.195 ;
    RECT 77.85 45.405 78.06 45.475 ;
    RECT 77.85 45.765 78.06 45.835 ;
    RECT 77.85 46.125 78.06 46.195 ;
    RECT 78.31 45.405 78.52 45.475 ;
    RECT 78.31 45.765 78.52 45.835 ;
    RECT 78.31 46.125 78.52 46.195 ;
    RECT 74.53 45.405 74.74 45.475 ;
    RECT 74.53 45.765 74.74 45.835 ;
    RECT 74.53 46.125 74.74 46.195 ;
    RECT 74.99 45.405 75.2 45.475 ;
    RECT 74.99 45.765 75.2 45.835 ;
    RECT 74.99 46.125 75.2 46.195 ;
    RECT 71.21 45.405 71.42 45.475 ;
    RECT 71.21 45.765 71.42 45.835 ;
    RECT 71.21 46.125 71.42 46.195 ;
    RECT 71.67 45.405 71.88 45.475 ;
    RECT 71.67 45.765 71.88 45.835 ;
    RECT 71.67 46.125 71.88 46.195 ;
    RECT 31.37 45.405 31.58 45.475 ;
    RECT 31.37 45.765 31.58 45.835 ;
    RECT 31.37 46.125 31.58 46.195 ;
    RECT 31.83 45.405 32.04 45.475 ;
    RECT 31.83 45.765 32.04 45.835 ;
    RECT 31.83 46.125 32.04 46.195 ;
    RECT 67.89 45.405 68.1 45.475 ;
    RECT 67.89 45.765 68.1 45.835 ;
    RECT 67.89 46.125 68.1 46.195 ;
    RECT 68.35 45.405 68.56 45.475 ;
    RECT 68.35 45.765 68.56 45.835 ;
    RECT 68.35 46.125 68.56 46.195 ;
    RECT 28.05 45.405 28.26 45.475 ;
    RECT 28.05 45.765 28.26 45.835 ;
    RECT 28.05 46.125 28.26 46.195 ;
    RECT 28.51 45.405 28.72 45.475 ;
    RECT 28.51 45.765 28.72 45.835 ;
    RECT 28.51 46.125 28.72 46.195 ;
    RECT 24.73 45.405 24.94 45.475 ;
    RECT 24.73 45.765 24.94 45.835 ;
    RECT 24.73 46.125 24.94 46.195 ;
    RECT 25.19 45.405 25.4 45.475 ;
    RECT 25.19 45.765 25.4 45.835 ;
    RECT 25.19 46.125 25.4 46.195 ;
    RECT 21.41 45.405 21.62 45.475 ;
    RECT 21.41 45.765 21.62 45.835 ;
    RECT 21.41 46.125 21.62 46.195 ;
    RECT 21.87 45.405 22.08 45.475 ;
    RECT 21.87 45.765 22.08 45.835 ;
    RECT 21.87 46.125 22.08 46.195 ;
    RECT 18.09 45.405 18.3 45.475 ;
    RECT 18.09 45.765 18.3 45.835 ;
    RECT 18.09 46.125 18.3 46.195 ;
    RECT 18.55 45.405 18.76 45.475 ;
    RECT 18.55 45.765 18.76 45.835 ;
    RECT 18.55 46.125 18.76 46.195 ;
    RECT 14.77 45.405 14.98 45.475 ;
    RECT 14.77 45.765 14.98 45.835 ;
    RECT 14.77 46.125 14.98 46.195 ;
    RECT 15.23 45.405 15.44 45.475 ;
    RECT 15.23 45.765 15.44 45.835 ;
    RECT 15.23 46.125 15.44 46.195 ;
    RECT 11.45 45.405 11.66 45.475 ;
    RECT 11.45 45.765 11.66 45.835 ;
    RECT 11.45 46.125 11.66 46.195 ;
    RECT 11.91 45.405 12.12 45.475 ;
    RECT 11.91 45.765 12.12 45.835 ;
    RECT 11.91 46.125 12.12 46.195 ;
    RECT 8.13 45.405 8.34 45.475 ;
    RECT 8.13 45.765 8.34 45.835 ;
    RECT 8.13 46.125 8.34 46.195 ;
    RECT 8.59 45.405 8.8 45.475 ;
    RECT 8.59 45.765 8.8 45.835 ;
    RECT 8.59 46.125 8.8 46.195 ;
    RECT 4.81 45.405 5.02 45.475 ;
    RECT 4.81 45.765 5.02 45.835 ;
    RECT 4.81 46.125 5.02 46.195 ;
    RECT 5.27 45.405 5.48 45.475 ;
    RECT 5.27 45.765 5.48 45.835 ;
    RECT 5.27 46.125 5.48 46.195 ;
    RECT 164.17 45.405 164.38 45.475 ;
    RECT 164.17 45.765 164.38 45.835 ;
    RECT 164.17 46.125 164.38 46.195 ;
    RECT 164.63 45.405 164.84 45.475 ;
    RECT 164.63 45.765 164.84 45.835 ;
    RECT 164.63 46.125 164.84 46.195 ;
    RECT 1.49 45.405 1.7 45.475 ;
    RECT 1.49 45.765 1.7 45.835 ;
    RECT 1.49 46.125 1.7 46.195 ;
    RECT 1.95 45.405 2.16 45.475 ;
    RECT 1.95 45.765 2.16 45.835 ;
    RECT 1.95 46.125 2.16 46.195 ;
    RECT 160.85 45.405 161.06 45.475 ;
    RECT 160.85 45.765 161.06 45.835 ;
    RECT 160.85 46.125 161.06 46.195 ;
    RECT 161.31 45.405 161.52 45.475 ;
    RECT 161.31 45.765 161.52 45.835 ;
    RECT 161.31 46.125 161.52 46.195 ;
    RECT 157.53 45.405 157.74 45.475 ;
    RECT 157.53 45.765 157.74 45.835 ;
    RECT 157.53 46.125 157.74 46.195 ;
    RECT 157.99 45.405 158.2 45.475 ;
    RECT 157.99 45.765 158.2 45.835 ;
    RECT 157.99 46.125 158.2 46.195 ;
    RECT 154.21 45.405 154.42 45.475 ;
    RECT 154.21 45.765 154.42 45.835 ;
    RECT 154.21 46.125 154.42 46.195 ;
    RECT 154.67 45.405 154.88 45.475 ;
    RECT 154.67 45.765 154.88 45.835 ;
    RECT 154.67 46.125 154.88 46.195 ;
    RECT 150.89 45.405 151.1 45.475 ;
    RECT 150.89 45.765 151.1 45.835 ;
    RECT 150.89 46.125 151.1 46.195 ;
    RECT 151.35 45.405 151.56 45.475 ;
    RECT 151.35 45.765 151.56 45.835 ;
    RECT 151.35 46.125 151.56 46.195 ;
    RECT 147.57 45.405 147.78 45.475 ;
    RECT 147.57 45.765 147.78 45.835 ;
    RECT 147.57 46.125 147.78 46.195 ;
    RECT 148.03 45.405 148.24 45.475 ;
    RECT 148.03 45.765 148.24 45.835 ;
    RECT 148.03 46.125 148.24 46.195 ;
    RECT 144.25 45.405 144.46 45.475 ;
    RECT 144.25 45.765 144.46 45.835 ;
    RECT 144.25 46.125 144.46 46.195 ;
    RECT 144.71 45.405 144.92 45.475 ;
    RECT 144.71 45.765 144.92 45.835 ;
    RECT 144.71 46.125 144.92 46.195 ;
    RECT 140.93 45.405 141.14 45.475 ;
    RECT 140.93 45.765 141.14 45.835 ;
    RECT 140.93 46.125 141.14 46.195 ;
    RECT 141.39 45.405 141.6 45.475 ;
    RECT 141.39 45.765 141.6 45.835 ;
    RECT 141.39 46.125 141.6 46.195 ;
    RECT 137.61 45.405 137.82 45.475 ;
    RECT 137.61 45.765 137.82 45.835 ;
    RECT 137.61 46.125 137.82 46.195 ;
    RECT 138.07 45.405 138.28 45.475 ;
    RECT 138.07 45.765 138.28 45.835 ;
    RECT 138.07 46.125 138.28 46.195 ;
    RECT 134.29 45.405 134.5 45.475 ;
    RECT 134.29 45.765 134.5 45.835 ;
    RECT 134.29 46.125 134.5 46.195 ;
    RECT 134.75 45.405 134.96 45.475 ;
    RECT 134.75 45.765 134.96 45.835 ;
    RECT 134.75 46.125 134.96 46.195 ;
    RECT 64.57 45.405 64.78 45.475 ;
    RECT 64.57 45.765 64.78 45.835 ;
    RECT 64.57 46.125 64.78 46.195 ;
    RECT 65.03 45.405 65.24 45.475 ;
    RECT 65.03 45.765 65.24 45.835 ;
    RECT 65.03 46.125 65.24 46.195 ;
    RECT 61.25 13.725 61.46 13.795 ;
    RECT 61.25 14.085 61.46 14.155 ;
    RECT 61.25 14.445 61.46 14.515 ;
    RECT 61.71 13.725 61.92 13.795 ;
    RECT 61.71 14.085 61.92 14.155 ;
    RECT 61.71 14.445 61.92 14.515 ;
    RECT 57.93 13.725 58.14 13.795 ;
    RECT 57.93 14.085 58.14 14.155 ;
    RECT 57.93 14.445 58.14 14.515 ;
    RECT 58.39 13.725 58.6 13.795 ;
    RECT 58.39 14.085 58.6 14.155 ;
    RECT 58.39 14.445 58.6 14.515 ;
    RECT 54.61 13.725 54.82 13.795 ;
    RECT 54.61 14.085 54.82 14.155 ;
    RECT 54.61 14.445 54.82 14.515 ;
    RECT 55.07 13.725 55.28 13.795 ;
    RECT 55.07 14.085 55.28 14.155 ;
    RECT 55.07 14.445 55.28 14.515 ;
    RECT 51.29 13.725 51.5 13.795 ;
    RECT 51.29 14.085 51.5 14.155 ;
    RECT 51.29 14.445 51.5 14.515 ;
    RECT 51.75 13.725 51.96 13.795 ;
    RECT 51.75 14.085 51.96 14.155 ;
    RECT 51.75 14.445 51.96 14.515 ;
    RECT 47.97 13.725 48.18 13.795 ;
    RECT 47.97 14.085 48.18 14.155 ;
    RECT 47.97 14.445 48.18 14.515 ;
    RECT 48.43 13.725 48.64 13.795 ;
    RECT 48.43 14.085 48.64 14.155 ;
    RECT 48.43 14.445 48.64 14.515 ;
    RECT 44.65 13.725 44.86 13.795 ;
    RECT 44.65 14.085 44.86 14.155 ;
    RECT 44.65 14.445 44.86 14.515 ;
    RECT 45.11 13.725 45.32 13.795 ;
    RECT 45.11 14.085 45.32 14.155 ;
    RECT 45.11 14.445 45.32 14.515 ;
    RECT 41.33 13.725 41.54 13.795 ;
    RECT 41.33 14.085 41.54 14.155 ;
    RECT 41.33 14.445 41.54 14.515 ;
    RECT 41.79 13.725 42.0 13.795 ;
    RECT 41.79 14.085 42.0 14.155 ;
    RECT 41.79 14.445 42.0 14.515 ;
    RECT 38.01 13.725 38.22 13.795 ;
    RECT 38.01 14.085 38.22 14.155 ;
    RECT 38.01 14.445 38.22 14.515 ;
    RECT 38.47 13.725 38.68 13.795 ;
    RECT 38.47 14.085 38.68 14.155 ;
    RECT 38.47 14.445 38.68 14.515 ;
    RECT 34.69 13.725 34.9 13.795 ;
    RECT 34.69 14.085 34.9 14.155 ;
    RECT 34.69 14.445 34.9 14.515 ;
    RECT 35.15 13.725 35.36 13.795 ;
    RECT 35.15 14.085 35.36 14.155 ;
    RECT 35.15 14.445 35.36 14.515 ;
    RECT 173.945 14.085 174.015 14.155 ;
    RECT 130.97 13.725 131.18 13.795 ;
    RECT 130.97 14.085 131.18 14.155 ;
    RECT 130.97 14.445 131.18 14.515 ;
    RECT 131.43 13.725 131.64 13.795 ;
    RECT 131.43 14.085 131.64 14.155 ;
    RECT 131.43 14.445 131.64 14.515 ;
    RECT 127.65 13.725 127.86 13.795 ;
    RECT 127.65 14.085 127.86 14.155 ;
    RECT 127.65 14.445 127.86 14.515 ;
    RECT 128.11 13.725 128.32 13.795 ;
    RECT 128.11 14.085 128.32 14.155 ;
    RECT 128.11 14.445 128.32 14.515 ;
    RECT 124.33 13.725 124.54 13.795 ;
    RECT 124.33 14.085 124.54 14.155 ;
    RECT 124.33 14.445 124.54 14.515 ;
    RECT 124.79 13.725 125.0 13.795 ;
    RECT 124.79 14.085 125.0 14.155 ;
    RECT 124.79 14.445 125.0 14.515 ;
    RECT 121.01 13.725 121.22 13.795 ;
    RECT 121.01 14.085 121.22 14.155 ;
    RECT 121.01 14.445 121.22 14.515 ;
    RECT 121.47 13.725 121.68 13.795 ;
    RECT 121.47 14.085 121.68 14.155 ;
    RECT 121.47 14.445 121.68 14.515 ;
    RECT 117.69 13.725 117.9 13.795 ;
    RECT 117.69 14.085 117.9 14.155 ;
    RECT 117.69 14.445 117.9 14.515 ;
    RECT 118.15 13.725 118.36 13.795 ;
    RECT 118.15 14.085 118.36 14.155 ;
    RECT 118.15 14.445 118.36 14.515 ;
    RECT 114.37 13.725 114.58 13.795 ;
    RECT 114.37 14.085 114.58 14.155 ;
    RECT 114.37 14.445 114.58 14.515 ;
    RECT 114.83 13.725 115.04 13.795 ;
    RECT 114.83 14.085 115.04 14.155 ;
    RECT 114.83 14.445 115.04 14.515 ;
    RECT 111.05 13.725 111.26 13.795 ;
    RECT 111.05 14.085 111.26 14.155 ;
    RECT 111.05 14.445 111.26 14.515 ;
    RECT 111.51 13.725 111.72 13.795 ;
    RECT 111.51 14.085 111.72 14.155 ;
    RECT 111.51 14.445 111.72 14.515 ;
    RECT 107.73 13.725 107.94 13.795 ;
    RECT 107.73 14.085 107.94 14.155 ;
    RECT 107.73 14.445 107.94 14.515 ;
    RECT 108.19 13.725 108.4 13.795 ;
    RECT 108.19 14.085 108.4 14.155 ;
    RECT 108.19 14.445 108.4 14.515 ;
    RECT 104.41 13.725 104.62 13.795 ;
    RECT 104.41 14.085 104.62 14.155 ;
    RECT 104.41 14.445 104.62 14.515 ;
    RECT 104.87 13.725 105.08 13.795 ;
    RECT 104.87 14.085 105.08 14.155 ;
    RECT 104.87 14.445 105.08 14.515 ;
    RECT 101.09 13.725 101.3 13.795 ;
    RECT 101.09 14.085 101.3 14.155 ;
    RECT 101.09 14.445 101.3 14.515 ;
    RECT 101.55 13.725 101.76 13.795 ;
    RECT 101.55 14.085 101.76 14.155 ;
    RECT 101.55 14.445 101.76 14.515 ;
    RECT 0.4 14.085 0.47 14.155 ;
    RECT 170.81 13.725 171.02 13.795 ;
    RECT 170.81 14.085 171.02 14.155 ;
    RECT 170.81 14.445 171.02 14.515 ;
    RECT 171.27 13.725 171.48 13.795 ;
    RECT 171.27 14.085 171.48 14.155 ;
    RECT 171.27 14.445 171.48 14.515 ;
    RECT 167.49 13.725 167.7 13.795 ;
    RECT 167.49 14.085 167.7 14.155 ;
    RECT 167.49 14.445 167.7 14.515 ;
    RECT 167.95 13.725 168.16 13.795 ;
    RECT 167.95 14.085 168.16 14.155 ;
    RECT 167.95 14.445 168.16 14.515 ;
    RECT 97.77 13.725 97.98 13.795 ;
    RECT 97.77 14.085 97.98 14.155 ;
    RECT 97.77 14.445 97.98 14.515 ;
    RECT 98.23 13.725 98.44 13.795 ;
    RECT 98.23 14.085 98.44 14.155 ;
    RECT 98.23 14.445 98.44 14.515 ;
    RECT 94.45 13.725 94.66 13.795 ;
    RECT 94.45 14.085 94.66 14.155 ;
    RECT 94.45 14.445 94.66 14.515 ;
    RECT 94.91 13.725 95.12 13.795 ;
    RECT 94.91 14.085 95.12 14.155 ;
    RECT 94.91 14.445 95.12 14.515 ;
    RECT 91.13 13.725 91.34 13.795 ;
    RECT 91.13 14.085 91.34 14.155 ;
    RECT 91.13 14.445 91.34 14.515 ;
    RECT 91.59 13.725 91.8 13.795 ;
    RECT 91.59 14.085 91.8 14.155 ;
    RECT 91.59 14.445 91.8 14.515 ;
    RECT 87.81 13.725 88.02 13.795 ;
    RECT 87.81 14.085 88.02 14.155 ;
    RECT 87.81 14.445 88.02 14.515 ;
    RECT 88.27 13.725 88.48 13.795 ;
    RECT 88.27 14.085 88.48 14.155 ;
    RECT 88.27 14.445 88.48 14.515 ;
    RECT 84.49 13.725 84.7 13.795 ;
    RECT 84.49 14.085 84.7 14.155 ;
    RECT 84.49 14.445 84.7 14.515 ;
    RECT 84.95 13.725 85.16 13.795 ;
    RECT 84.95 14.085 85.16 14.155 ;
    RECT 84.95 14.445 85.16 14.515 ;
    RECT 81.17 13.725 81.38 13.795 ;
    RECT 81.17 14.085 81.38 14.155 ;
    RECT 81.17 14.445 81.38 14.515 ;
    RECT 81.63 13.725 81.84 13.795 ;
    RECT 81.63 14.085 81.84 14.155 ;
    RECT 81.63 14.445 81.84 14.515 ;
    RECT 77.85 13.725 78.06 13.795 ;
    RECT 77.85 14.085 78.06 14.155 ;
    RECT 77.85 14.445 78.06 14.515 ;
    RECT 78.31 13.725 78.52 13.795 ;
    RECT 78.31 14.085 78.52 14.155 ;
    RECT 78.31 14.445 78.52 14.515 ;
    RECT 74.53 13.725 74.74 13.795 ;
    RECT 74.53 14.085 74.74 14.155 ;
    RECT 74.53 14.445 74.74 14.515 ;
    RECT 74.99 13.725 75.2 13.795 ;
    RECT 74.99 14.085 75.2 14.155 ;
    RECT 74.99 14.445 75.2 14.515 ;
    RECT 71.21 13.725 71.42 13.795 ;
    RECT 71.21 14.085 71.42 14.155 ;
    RECT 71.21 14.445 71.42 14.515 ;
    RECT 71.67 13.725 71.88 13.795 ;
    RECT 71.67 14.085 71.88 14.155 ;
    RECT 71.67 14.445 71.88 14.515 ;
    RECT 31.37 13.725 31.58 13.795 ;
    RECT 31.37 14.085 31.58 14.155 ;
    RECT 31.37 14.445 31.58 14.515 ;
    RECT 31.83 13.725 32.04 13.795 ;
    RECT 31.83 14.085 32.04 14.155 ;
    RECT 31.83 14.445 32.04 14.515 ;
    RECT 67.89 13.725 68.1 13.795 ;
    RECT 67.89 14.085 68.1 14.155 ;
    RECT 67.89 14.445 68.1 14.515 ;
    RECT 68.35 13.725 68.56 13.795 ;
    RECT 68.35 14.085 68.56 14.155 ;
    RECT 68.35 14.445 68.56 14.515 ;
    RECT 28.05 13.725 28.26 13.795 ;
    RECT 28.05 14.085 28.26 14.155 ;
    RECT 28.05 14.445 28.26 14.515 ;
    RECT 28.51 13.725 28.72 13.795 ;
    RECT 28.51 14.085 28.72 14.155 ;
    RECT 28.51 14.445 28.72 14.515 ;
    RECT 24.73 13.725 24.94 13.795 ;
    RECT 24.73 14.085 24.94 14.155 ;
    RECT 24.73 14.445 24.94 14.515 ;
    RECT 25.19 13.725 25.4 13.795 ;
    RECT 25.19 14.085 25.4 14.155 ;
    RECT 25.19 14.445 25.4 14.515 ;
    RECT 21.41 13.725 21.62 13.795 ;
    RECT 21.41 14.085 21.62 14.155 ;
    RECT 21.41 14.445 21.62 14.515 ;
    RECT 21.87 13.725 22.08 13.795 ;
    RECT 21.87 14.085 22.08 14.155 ;
    RECT 21.87 14.445 22.08 14.515 ;
    RECT 18.09 13.725 18.3 13.795 ;
    RECT 18.09 14.085 18.3 14.155 ;
    RECT 18.09 14.445 18.3 14.515 ;
    RECT 18.55 13.725 18.76 13.795 ;
    RECT 18.55 14.085 18.76 14.155 ;
    RECT 18.55 14.445 18.76 14.515 ;
    RECT 14.77 13.725 14.98 13.795 ;
    RECT 14.77 14.085 14.98 14.155 ;
    RECT 14.77 14.445 14.98 14.515 ;
    RECT 15.23 13.725 15.44 13.795 ;
    RECT 15.23 14.085 15.44 14.155 ;
    RECT 15.23 14.445 15.44 14.515 ;
    RECT 11.45 13.725 11.66 13.795 ;
    RECT 11.45 14.085 11.66 14.155 ;
    RECT 11.45 14.445 11.66 14.515 ;
    RECT 11.91 13.725 12.12 13.795 ;
    RECT 11.91 14.085 12.12 14.155 ;
    RECT 11.91 14.445 12.12 14.515 ;
    RECT 8.13 13.725 8.34 13.795 ;
    RECT 8.13 14.085 8.34 14.155 ;
    RECT 8.13 14.445 8.34 14.515 ;
    RECT 8.59 13.725 8.8 13.795 ;
    RECT 8.59 14.085 8.8 14.155 ;
    RECT 8.59 14.445 8.8 14.515 ;
    RECT 4.81 13.725 5.02 13.795 ;
    RECT 4.81 14.085 5.02 14.155 ;
    RECT 4.81 14.445 5.02 14.515 ;
    RECT 5.27 13.725 5.48 13.795 ;
    RECT 5.27 14.085 5.48 14.155 ;
    RECT 5.27 14.445 5.48 14.515 ;
    RECT 164.17 13.725 164.38 13.795 ;
    RECT 164.17 14.085 164.38 14.155 ;
    RECT 164.17 14.445 164.38 14.515 ;
    RECT 164.63 13.725 164.84 13.795 ;
    RECT 164.63 14.085 164.84 14.155 ;
    RECT 164.63 14.445 164.84 14.515 ;
    RECT 1.49 13.725 1.7 13.795 ;
    RECT 1.49 14.085 1.7 14.155 ;
    RECT 1.49 14.445 1.7 14.515 ;
    RECT 1.95 13.725 2.16 13.795 ;
    RECT 1.95 14.085 2.16 14.155 ;
    RECT 1.95 14.445 2.16 14.515 ;
    RECT 160.85 13.725 161.06 13.795 ;
    RECT 160.85 14.085 161.06 14.155 ;
    RECT 160.85 14.445 161.06 14.515 ;
    RECT 161.31 13.725 161.52 13.795 ;
    RECT 161.31 14.085 161.52 14.155 ;
    RECT 161.31 14.445 161.52 14.515 ;
    RECT 157.53 13.725 157.74 13.795 ;
    RECT 157.53 14.085 157.74 14.155 ;
    RECT 157.53 14.445 157.74 14.515 ;
    RECT 157.99 13.725 158.2 13.795 ;
    RECT 157.99 14.085 158.2 14.155 ;
    RECT 157.99 14.445 158.2 14.515 ;
    RECT 154.21 13.725 154.42 13.795 ;
    RECT 154.21 14.085 154.42 14.155 ;
    RECT 154.21 14.445 154.42 14.515 ;
    RECT 154.67 13.725 154.88 13.795 ;
    RECT 154.67 14.085 154.88 14.155 ;
    RECT 154.67 14.445 154.88 14.515 ;
    RECT 150.89 13.725 151.1 13.795 ;
    RECT 150.89 14.085 151.1 14.155 ;
    RECT 150.89 14.445 151.1 14.515 ;
    RECT 151.35 13.725 151.56 13.795 ;
    RECT 151.35 14.085 151.56 14.155 ;
    RECT 151.35 14.445 151.56 14.515 ;
    RECT 147.57 13.725 147.78 13.795 ;
    RECT 147.57 14.085 147.78 14.155 ;
    RECT 147.57 14.445 147.78 14.515 ;
    RECT 148.03 13.725 148.24 13.795 ;
    RECT 148.03 14.085 148.24 14.155 ;
    RECT 148.03 14.445 148.24 14.515 ;
    RECT 144.25 13.725 144.46 13.795 ;
    RECT 144.25 14.085 144.46 14.155 ;
    RECT 144.25 14.445 144.46 14.515 ;
    RECT 144.71 13.725 144.92 13.795 ;
    RECT 144.71 14.085 144.92 14.155 ;
    RECT 144.71 14.445 144.92 14.515 ;
    RECT 140.93 13.725 141.14 13.795 ;
    RECT 140.93 14.085 141.14 14.155 ;
    RECT 140.93 14.445 141.14 14.515 ;
    RECT 141.39 13.725 141.6 13.795 ;
    RECT 141.39 14.085 141.6 14.155 ;
    RECT 141.39 14.445 141.6 14.515 ;
    RECT 137.61 13.725 137.82 13.795 ;
    RECT 137.61 14.085 137.82 14.155 ;
    RECT 137.61 14.445 137.82 14.515 ;
    RECT 138.07 13.725 138.28 13.795 ;
    RECT 138.07 14.085 138.28 14.155 ;
    RECT 138.07 14.445 138.28 14.515 ;
    RECT 134.29 13.725 134.5 13.795 ;
    RECT 134.29 14.085 134.5 14.155 ;
    RECT 134.29 14.445 134.5 14.515 ;
    RECT 134.75 13.725 134.96 13.795 ;
    RECT 134.75 14.085 134.96 14.155 ;
    RECT 134.75 14.445 134.96 14.515 ;
    RECT 64.57 13.725 64.78 13.795 ;
    RECT 64.57 14.085 64.78 14.155 ;
    RECT 64.57 14.445 64.78 14.515 ;
    RECT 65.03 13.725 65.24 13.795 ;
    RECT 65.03 14.085 65.24 14.155 ;
    RECT 65.03 14.445 65.24 14.515 ;
    RECT 61.25 44.685 61.46 44.755 ;
    RECT 61.25 45.045 61.46 45.115 ;
    RECT 61.25 45.405 61.46 45.475 ;
    RECT 61.71 44.685 61.92 44.755 ;
    RECT 61.71 45.045 61.92 45.115 ;
    RECT 61.71 45.405 61.92 45.475 ;
    RECT 57.93 44.685 58.14 44.755 ;
    RECT 57.93 45.045 58.14 45.115 ;
    RECT 57.93 45.405 58.14 45.475 ;
    RECT 58.39 44.685 58.6 44.755 ;
    RECT 58.39 45.045 58.6 45.115 ;
    RECT 58.39 45.405 58.6 45.475 ;
    RECT 54.61 44.685 54.82 44.755 ;
    RECT 54.61 45.045 54.82 45.115 ;
    RECT 54.61 45.405 54.82 45.475 ;
    RECT 55.07 44.685 55.28 44.755 ;
    RECT 55.07 45.045 55.28 45.115 ;
    RECT 55.07 45.405 55.28 45.475 ;
    RECT 51.29 44.685 51.5 44.755 ;
    RECT 51.29 45.045 51.5 45.115 ;
    RECT 51.29 45.405 51.5 45.475 ;
    RECT 51.75 44.685 51.96 44.755 ;
    RECT 51.75 45.045 51.96 45.115 ;
    RECT 51.75 45.405 51.96 45.475 ;
    RECT 47.97 44.685 48.18 44.755 ;
    RECT 47.97 45.045 48.18 45.115 ;
    RECT 47.97 45.405 48.18 45.475 ;
    RECT 48.43 44.685 48.64 44.755 ;
    RECT 48.43 45.045 48.64 45.115 ;
    RECT 48.43 45.405 48.64 45.475 ;
    RECT 44.65 44.685 44.86 44.755 ;
    RECT 44.65 45.045 44.86 45.115 ;
    RECT 44.65 45.405 44.86 45.475 ;
    RECT 45.11 44.685 45.32 44.755 ;
    RECT 45.11 45.045 45.32 45.115 ;
    RECT 45.11 45.405 45.32 45.475 ;
    RECT 41.33 44.685 41.54 44.755 ;
    RECT 41.33 45.045 41.54 45.115 ;
    RECT 41.33 45.405 41.54 45.475 ;
    RECT 41.79 44.685 42.0 44.755 ;
    RECT 41.79 45.045 42.0 45.115 ;
    RECT 41.79 45.405 42.0 45.475 ;
    RECT 38.01 44.685 38.22 44.755 ;
    RECT 38.01 45.045 38.22 45.115 ;
    RECT 38.01 45.405 38.22 45.475 ;
    RECT 38.47 44.685 38.68 44.755 ;
    RECT 38.47 45.045 38.68 45.115 ;
    RECT 38.47 45.405 38.68 45.475 ;
    RECT 34.69 44.685 34.9 44.755 ;
    RECT 34.69 45.045 34.9 45.115 ;
    RECT 34.69 45.405 34.9 45.475 ;
    RECT 35.15 44.685 35.36 44.755 ;
    RECT 35.15 45.045 35.36 45.115 ;
    RECT 35.15 45.405 35.36 45.475 ;
    RECT 173.945 45.045 174.015 45.115 ;
    RECT 130.97 44.685 131.18 44.755 ;
    RECT 130.97 45.045 131.18 45.115 ;
    RECT 130.97 45.405 131.18 45.475 ;
    RECT 131.43 44.685 131.64 44.755 ;
    RECT 131.43 45.045 131.64 45.115 ;
    RECT 131.43 45.405 131.64 45.475 ;
    RECT 127.65 44.685 127.86 44.755 ;
    RECT 127.65 45.045 127.86 45.115 ;
    RECT 127.65 45.405 127.86 45.475 ;
    RECT 128.11 44.685 128.32 44.755 ;
    RECT 128.11 45.045 128.32 45.115 ;
    RECT 128.11 45.405 128.32 45.475 ;
    RECT 124.33 44.685 124.54 44.755 ;
    RECT 124.33 45.045 124.54 45.115 ;
    RECT 124.33 45.405 124.54 45.475 ;
    RECT 124.79 44.685 125.0 44.755 ;
    RECT 124.79 45.045 125.0 45.115 ;
    RECT 124.79 45.405 125.0 45.475 ;
    RECT 121.01 44.685 121.22 44.755 ;
    RECT 121.01 45.045 121.22 45.115 ;
    RECT 121.01 45.405 121.22 45.475 ;
    RECT 121.47 44.685 121.68 44.755 ;
    RECT 121.47 45.045 121.68 45.115 ;
    RECT 121.47 45.405 121.68 45.475 ;
    RECT 117.69 44.685 117.9 44.755 ;
    RECT 117.69 45.045 117.9 45.115 ;
    RECT 117.69 45.405 117.9 45.475 ;
    RECT 118.15 44.685 118.36 44.755 ;
    RECT 118.15 45.045 118.36 45.115 ;
    RECT 118.15 45.405 118.36 45.475 ;
    RECT 114.37 44.685 114.58 44.755 ;
    RECT 114.37 45.045 114.58 45.115 ;
    RECT 114.37 45.405 114.58 45.475 ;
    RECT 114.83 44.685 115.04 44.755 ;
    RECT 114.83 45.045 115.04 45.115 ;
    RECT 114.83 45.405 115.04 45.475 ;
    RECT 111.05 44.685 111.26 44.755 ;
    RECT 111.05 45.045 111.26 45.115 ;
    RECT 111.05 45.405 111.26 45.475 ;
    RECT 111.51 44.685 111.72 44.755 ;
    RECT 111.51 45.045 111.72 45.115 ;
    RECT 111.51 45.405 111.72 45.475 ;
    RECT 107.73 44.685 107.94 44.755 ;
    RECT 107.73 45.045 107.94 45.115 ;
    RECT 107.73 45.405 107.94 45.475 ;
    RECT 108.19 44.685 108.4 44.755 ;
    RECT 108.19 45.045 108.4 45.115 ;
    RECT 108.19 45.405 108.4 45.475 ;
    RECT 104.41 44.685 104.62 44.755 ;
    RECT 104.41 45.045 104.62 45.115 ;
    RECT 104.41 45.405 104.62 45.475 ;
    RECT 104.87 44.685 105.08 44.755 ;
    RECT 104.87 45.045 105.08 45.115 ;
    RECT 104.87 45.405 105.08 45.475 ;
    RECT 101.09 44.685 101.3 44.755 ;
    RECT 101.09 45.045 101.3 45.115 ;
    RECT 101.09 45.405 101.3 45.475 ;
    RECT 101.55 44.685 101.76 44.755 ;
    RECT 101.55 45.045 101.76 45.115 ;
    RECT 101.55 45.405 101.76 45.475 ;
    RECT 0.4 45.045 0.47 45.115 ;
    RECT 170.81 44.685 171.02 44.755 ;
    RECT 170.81 45.045 171.02 45.115 ;
    RECT 170.81 45.405 171.02 45.475 ;
    RECT 171.27 44.685 171.48 44.755 ;
    RECT 171.27 45.045 171.48 45.115 ;
    RECT 171.27 45.405 171.48 45.475 ;
    RECT 167.49 44.685 167.7 44.755 ;
    RECT 167.49 45.045 167.7 45.115 ;
    RECT 167.49 45.405 167.7 45.475 ;
    RECT 167.95 44.685 168.16 44.755 ;
    RECT 167.95 45.045 168.16 45.115 ;
    RECT 167.95 45.405 168.16 45.475 ;
    RECT 97.77 44.685 97.98 44.755 ;
    RECT 97.77 45.045 97.98 45.115 ;
    RECT 97.77 45.405 97.98 45.475 ;
    RECT 98.23 44.685 98.44 44.755 ;
    RECT 98.23 45.045 98.44 45.115 ;
    RECT 98.23 45.405 98.44 45.475 ;
    RECT 94.45 44.685 94.66 44.755 ;
    RECT 94.45 45.045 94.66 45.115 ;
    RECT 94.45 45.405 94.66 45.475 ;
    RECT 94.91 44.685 95.12 44.755 ;
    RECT 94.91 45.045 95.12 45.115 ;
    RECT 94.91 45.405 95.12 45.475 ;
    RECT 91.13 44.685 91.34 44.755 ;
    RECT 91.13 45.045 91.34 45.115 ;
    RECT 91.13 45.405 91.34 45.475 ;
    RECT 91.59 44.685 91.8 44.755 ;
    RECT 91.59 45.045 91.8 45.115 ;
    RECT 91.59 45.405 91.8 45.475 ;
    RECT 87.81 44.685 88.02 44.755 ;
    RECT 87.81 45.045 88.02 45.115 ;
    RECT 87.81 45.405 88.02 45.475 ;
    RECT 88.27 44.685 88.48 44.755 ;
    RECT 88.27 45.045 88.48 45.115 ;
    RECT 88.27 45.405 88.48 45.475 ;
    RECT 84.49 44.685 84.7 44.755 ;
    RECT 84.49 45.045 84.7 45.115 ;
    RECT 84.49 45.405 84.7 45.475 ;
    RECT 84.95 44.685 85.16 44.755 ;
    RECT 84.95 45.045 85.16 45.115 ;
    RECT 84.95 45.405 85.16 45.475 ;
    RECT 81.17 44.685 81.38 44.755 ;
    RECT 81.17 45.045 81.38 45.115 ;
    RECT 81.17 45.405 81.38 45.475 ;
    RECT 81.63 44.685 81.84 44.755 ;
    RECT 81.63 45.045 81.84 45.115 ;
    RECT 81.63 45.405 81.84 45.475 ;
    RECT 77.85 44.685 78.06 44.755 ;
    RECT 77.85 45.045 78.06 45.115 ;
    RECT 77.85 45.405 78.06 45.475 ;
    RECT 78.31 44.685 78.52 44.755 ;
    RECT 78.31 45.045 78.52 45.115 ;
    RECT 78.31 45.405 78.52 45.475 ;
    RECT 74.53 44.685 74.74 44.755 ;
    RECT 74.53 45.045 74.74 45.115 ;
    RECT 74.53 45.405 74.74 45.475 ;
    RECT 74.99 44.685 75.2 44.755 ;
    RECT 74.99 45.045 75.2 45.115 ;
    RECT 74.99 45.405 75.2 45.475 ;
    RECT 71.21 44.685 71.42 44.755 ;
    RECT 71.21 45.045 71.42 45.115 ;
    RECT 71.21 45.405 71.42 45.475 ;
    RECT 71.67 44.685 71.88 44.755 ;
    RECT 71.67 45.045 71.88 45.115 ;
    RECT 71.67 45.405 71.88 45.475 ;
    RECT 31.37 44.685 31.58 44.755 ;
    RECT 31.37 45.045 31.58 45.115 ;
    RECT 31.37 45.405 31.58 45.475 ;
    RECT 31.83 44.685 32.04 44.755 ;
    RECT 31.83 45.045 32.04 45.115 ;
    RECT 31.83 45.405 32.04 45.475 ;
    RECT 67.89 44.685 68.1 44.755 ;
    RECT 67.89 45.045 68.1 45.115 ;
    RECT 67.89 45.405 68.1 45.475 ;
    RECT 68.35 44.685 68.56 44.755 ;
    RECT 68.35 45.045 68.56 45.115 ;
    RECT 68.35 45.405 68.56 45.475 ;
    RECT 28.05 44.685 28.26 44.755 ;
    RECT 28.05 45.045 28.26 45.115 ;
    RECT 28.05 45.405 28.26 45.475 ;
    RECT 28.51 44.685 28.72 44.755 ;
    RECT 28.51 45.045 28.72 45.115 ;
    RECT 28.51 45.405 28.72 45.475 ;
    RECT 24.73 44.685 24.94 44.755 ;
    RECT 24.73 45.045 24.94 45.115 ;
    RECT 24.73 45.405 24.94 45.475 ;
    RECT 25.19 44.685 25.4 44.755 ;
    RECT 25.19 45.045 25.4 45.115 ;
    RECT 25.19 45.405 25.4 45.475 ;
    RECT 21.41 44.685 21.62 44.755 ;
    RECT 21.41 45.045 21.62 45.115 ;
    RECT 21.41 45.405 21.62 45.475 ;
    RECT 21.87 44.685 22.08 44.755 ;
    RECT 21.87 45.045 22.08 45.115 ;
    RECT 21.87 45.405 22.08 45.475 ;
    RECT 18.09 44.685 18.3 44.755 ;
    RECT 18.09 45.045 18.3 45.115 ;
    RECT 18.09 45.405 18.3 45.475 ;
    RECT 18.55 44.685 18.76 44.755 ;
    RECT 18.55 45.045 18.76 45.115 ;
    RECT 18.55 45.405 18.76 45.475 ;
    RECT 14.77 44.685 14.98 44.755 ;
    RECT 14.77 45.045 14.98 45.115 ;
    RECT 14.77 45.405 14.98 45.475 ;
    RECT 15.23 44.685 15.44 44.755 ;
    RECT 15.23 45.045 15.44 45.115 ;
    RECT 15.23 45.405 15.44 45.475 ;
    RECT 11.45 44.685 11.66 44.755 ;
    RECT 11.45 45.045 11.66 45.115 ;
    RECT 11.45 45.405 11.66 45.475 ;
    RECT 11.91 44.685 12.12 44.755 ;
    RECT 11.91 45.045 12.12 45.115 ;
    RECT 11.91 45.405 12.12 45.475 ;
    RECT 8.13 44.685 8.34 44.755 ;
    RECT 8.13 45.045 8.34 45.115 ;
    RECT 8.13 45.405 8.34 45.475 ;
    RECT 8.59 44.685 8.8 44.755 ;
    RECT 8.59 45.045 8.8 45.115 ;
    RECT 8.59 45.405 8.8 45.475 ;
    RECT 4.81 44.685 5.02 44.755 ;
    RECT 4.81 45.045 5.02 45.115 ;
    RECT 4.81 45.405 5.02 45.475 ;
    RECT 5.27 44.685 5.48 44.755 ;
    RECT 5.27 45.045 5.48 45.115 ;
    RECT 5.27 45.405 5.48 45.475 ;
    RECT 164.17 44.685 164.38 44.755 ;
    RECT 164.17 45.045 164.38 45.115 ;
    RECT 164.17 45.405 164.38 45.475 ;
    RECT 164.63 44.685 164.84 44.755 ;
    RECT 164.63 45.045 164.84 45.115 ;
    RECT 164.63 45.405 164.84 45.475 ;
    RECT 1.49 44.685 1.7 44.755 ;
    RECT 1.49 45.045 1.7 45.115 ;
    RECT 1.49 45.405 1.7 45.475 ;
    RECT 1.95 44.685 2.16 44.755 ;
    RECT 1.95 45.045 2.16 45.115 ;
    RECT 1.95 45.405 2.16 45.475 ;
    RECT 160.85 44.685 161.06 44.755 ;
    RECT 160.85 45.045 161.06 45.115 ;
    RECT 160.85 45.405 161.06 45.475 ;
    RECT 161.31 44.685 161.52 44.755 ;
    RECT 161.31 45.045 161.52 45.115 ;
    RECT 161.31 45.405 161.52 45.475 ;
    RECT 157.53 44.685 157.74 44.755 ;
    RECT 157.53 45.045 157.74 45.115 ;
    RECT 157.53 45.405 157.74 45.475 ;
    RECT 157.99 44.685 158.2 44.755 ;
    RECT 157.99 45.045 158.2 45.115 ;
    RECT 157.99 45.405 158.2 45.475 ;
    RECT 154.21 44.685 154.42 44.755 ;
    RECT 154.21 45.045 154.42 45.115 ;
    RECT 154.21 45.405 154.42 45.475 ;
    RECT 154.67 44.685 154.88 44.755 ;
    RECT 154.67 45.045 154.88 45.115 ;
    RECT 154.67 45.405 154.88 45.475 ;
    RECT 150.89 44.685 151.1 44.755 ;
    RECT 150.89 45.045 151.1 45.115 ;
    RECT 150.89 45.405 151.1 45.475 ;
    RECT 151.35 44.685 151.56 44.755 ;
    RECT 151.35 45.045 151.56 45.115 ;
    RECT 151.35 45.405 151.56 45.475 ;
    RECT 147.57 44.685 147.78 44.755 ;
    RECT 147.57 45.045 147.78 45.115 ;
    RECT 147.57 45.405 147.78 45.475 ;
    RECT 148.03 44.685 148.24 44.755 ;
    RECT 148.03 45.045 148.24 45.115 ;
    RECT 148.03 45.405 148.24 45.475 ;
    RECT 144.25 44.685 144.46 44.755 ;
    RECT 144.25 45.045 144.46 45.115 ;
    RECT 144.25 45.405 144.46 45.475 ;
    RECT 144.71 44.685 144.92 44.755 ;
    RECT 144.71 45.045 144.92 45.115 ;
    RECT 144.71 45.405 144.92 45.475 ;
    RECT 140.93 44.685 141.14 44.755 ;
    RECT 140.93 45.045 141.14 45.115 ;
    RECT 140.93 45.405 141.14 45.475 ;
    RECT 141.39 44.685 141.6 44.755 ;
    RECT 141.39 45.045 141.6 45.115 ;
    RECT 141.39 45.405 141.6 45.475 ;
    RECT 137.61 44.685 137.82 44.755 ;
    RECT 137.61 45.045 137.82 45.115 ;
    RECT 137.61 45.405 137.82 45.475 ;
    RECT 138.07 44.685 138.28 44.755 ;
    RECT 138.07 45.045 138.28 45.115 ;
    RECT 138.07 45.405 138.28 45.475 ;
    RECT 134.29 44.685 134.5 44.755 ;
    RECT 134.29 45.045 134.5 45.115 ;
    RECT 134.29 45.405 134.5 45.475 ;
    RECT 134.75 44.685 134.96 44.755 ;
    RECT 134.75 45.045 134.96 45.115 ;
    RECT 134.75 45.405 134.96 45.475 ;
    RECT 64.57 44.685 64.78 44.755 ;
    RECT 64.57 45.045 64.78 45.115 ;
    RECT 64.57 45.405 64.78 45.475 ;
    RECT 65.03 44.685 65.24 44.755 ;
    RECT 65.03 45.045 65.24 45.115 ;
    RECT 65.03 45.405 65.24 45.475 ;
    RECT 61.25 13.005 61.46 13.075 ;
    RECT 61.25 13.365 61.46 13.435 ;
    RECT 61.25 13.725 61.46 13.795 ;
    RECT 61.71 13.005 61.92 13.075 ;
    RECT 61.71 13.365 61.92 13.435 ;
    RECT 61.71 13.725 61.92 13.795 ;
    RECT 57.93 13.005 58.14 13.075 ;
    RECT 57.93 13.365 58.14 13.435 ;
    RECT 57.93 13.725 58.14 13.795 ;
    RECT 58.39 13.005 58.6 13.075 ;
    RECT 58.39 13.365 58.6 13.435 ;
    RECT 58.39 13.725 58.6 13.795 ;
    RECT 54.61 13.005 54.82 13.075 ;
    RECT 54.61 13.365 54.82 13.435 ;
    RECT 54.61 13.725 54.82 13.795 ;
    RECT 55.07 13.005 55.28 13.075 ;
    RECT 55.07 13.365 55.28 13.435 ;
    RECT 55.07 13.725 55.28 13.795 ;
    RECT 51.29 13.005 51.5 13.075 ;
    RECT 51.29 13.365 51.5 13.435 ;
    RECT 51.29 13.725 51.5 13.795 ;
    RECT 51.75 13.005 51.96 13.075 ;
    RECT 51.75 13.365 51.96 13.435 ;
    RECT 51.75 13.725 51.96 13.795 ;
    RECT 47.97 13.005 48.18 13.075 ;
    RECT 47.97 13.365 48.18 13.435 ;
    RECT 47.97 13.725 48.18 13.795 ;
    RECT 48.43 13.005 48.64 13.075 ;
    RECT 48.43 13.365 48.64 13.435 ;
    RECT 48.43 13.725 48.64 13.795 ;
    RECT 44.65 13.005 44.86 13.075 ;
    RECT 44.65 13.365 44.86 13.435 ;
    RECT 44.65 13.725 44.86 13.795 ;
    RECT 45.11 13.005 45.32 13.075 ;
    RECT 45.11 13.365 45.32 13.435 ;
    RECT 45.11 13.725 45.32 13.795 ;
    RECT 41.33 13.005 41.54 13.075 ;
    RECT 41.33 13.365 41.54 13.435 ;
    RECT 41.33 13.725 41.54 13.795 ;
    RECT 41.79 13.005 42.0 13.075 ;
    RECT 41.79 13.365 42.0 13.435 ;
    RECT 41.79 13.725 42.0 13.795 ;
    RECT 38.01 13.005 38.22 13.075 ;
    RECT 38.01 13.365 38.22 13.435 ;
    RECT 38.01 13.725 38.22 13.795 ;
    RECT 38.47 13.005 38.68 13.075 ;
    RECT 38.47 13.365 38.68 13.435 ;
    RECT 38.47 13.725 38.68 13.795 ;
    RECT 34.69 13.005 34.9 13.075 ;
    RECT 34.69 13.365 34.9 13.435 ;
    RECT 34.69 13.725 34.9 13.795 ;
    RECT 35.15 13.005 35.36 13.075 ;
    RECT 35.15 13.365 35.36 13.435 ;
    RECT 35.15 13.725 35.36 13.795 ;
    RECT 173.945 13.365 174.015 13.435 ;
    RECT 130.97 13.005 131.18 13.075 ;
    RECT 130.97 13.365 131.18 13.435 ;
    RECT 130.97 13.725 131.18 13.795 ;
    RECT 131.43 13.005 131.64 13.075 ;
    RECT 131.43 13.365 131.64 13.435 ;
    RECT 131.43 13.725 131.64 13.795 ;
    RECT 127.65 13.005 127.86 13.075 ;
    RECT 127.65 13.365 127.86 13.435 ;
    RECT 127.65 13.725 127.86 13.795 ;
    RECT 128.11 13.005 128.32 13.075 ;
    RECT 128.11 13.365 128.32 13.435 ;
    RECT 128.11 13.725 128.32 13.795 ;
    RECT 124.33 13.005 124.54 13.075 ;
    RECT 124.33 13.365 124.54 13.435 ;
    RECT 124.33 13.725 124.54 13.795 ;
    RECT 124.79 13.005 125.0 13.075 ;
    RECT 124.79 13.365 125.0 13.435 ;
    RECT 124.79 13.725 125.0 13.795 ;
    RECT 121.01 13.005 121.22 13.075 ;
    RECT 121.01 13.365 121.22 13.435 ;
    RECT 121.01 13.725 121.22 13.795 ;
    RECT 121.47 13.005 121.68 13.075 ;
    RECT 121.47 13.365 121.68 13.435 ;
    RECT 121.47 13.725 121.68 13.795 ;
    RECT 117.69 13.005 117.9 13.075 ;
    RECT 117.69 13.365 117.9 13.435 ;
    RECT 117.69 13.725 117.9 13.795 ;
    RECT 118.15 13.005 118.36 13.075 ;
    RECT 118.15 13.365 118.36 13.435 ;
    RECT 118.15 13.725 118.36 13.795 ;
    RECT 114.37 13.005 114.58 13.075 ;
    RECT 114.37 13.365 114.58 13.435 ;
    RECT 114.37 13.725 114.58 13.795 ;
    RECT 114.83 13.005 115.04 13.075 ;
    RECT 114.83 13.365 115.04 13.435 ;
    RECT 114.83 13.725 115.04 13.795 ;
    RECT 111.05 13.005 111.26 13.075 ;
    RECT 111.05 13.365 111.26 13.435 ;
    RECT 111.05 13.725 111.26 13.795 ;
    RECT 111.51 13.005 111.72 13.075 ;
    RECT 111.51 13.365 111.72 13.435 ;
    RECT 111.51 13.725 111.72 13.795 ;
    RECT 107.73 13.005 107.94 13.075 ;
    RECT 107.73 13.365 107.94 13.435 ;
    RECT 107.73 13.725 107.94 13.795 ;
    RECT 108.19 13.005 108.4 13.075 ;
    RECT 108.19 13.365 108.4 13.435 ;
    RECT 108.19 13.725 108.4 13.795 ;
    RECT 104.41 13.005 104.62 13.075 ;
    RECT 104.41 13.365 104.62 13.435 ;
    RECT 104.41 13.725 104.62 13.795 ;
    RECT 104.87 13.005 105.08 13.075 ;
    RECT 104.87 13.365 105.08 13.435 ;
    RECT 104.87 13.725 105.08 13.795 ;
    RECT 101.09 13.005 101.3 13.075 ;
    RECT 101.09 13.365 101.3 13.435 ;
    RECT 101.09 13.725 101.3 13.795 ;
    RECT 101.55 13.005 101.76 13.075 ;
    RECT 101.55 13.365 101.76 13.435 ;
    RECT 101.55 13.725 101.76 13.795 ;
    RECT 0.4 13.365 0.47 13.435 ;
    RECT 170.81 13.005 171.02 13.075 ;
    RECT 170.81 13.365 171.02 13.435 ;
    RECT 170.81 13.725 171.02 13.795 ;
    RECT 171.27 13.005 171.48 13.075 ;
    RECT 171.27 13.365 171.48 13.435 ;
    RECT 171.27 13.725 171.48 13.795 ;
    RECT 167.49 13.005 167.7 13.075 ;
    RECT 167.49 13.365 167.7 13.435 ;
    RECT 167.49 13.725 167.7 13.795 ;
    RECT 167.95 13.005 168.16 13.075 ;
    RECT 167.95 13.365 168.16 13.435 ;
    RECT 167.95 13.725 168.16 13.795 ;
    RECT 97.77 13.005 97.98 13.075 ;
    RECT 97.77 13.365 97.98 13.435 ;
    RECT 97.77 13.725 97.98 13.795 ;
    RECT 98.23 13.005 98.44 13.075 ;
    RECT 98.23 13.365 98.44 13.435 ;
    RECT 98.23 13.725 98.44 13.795 ;
    RECT 94.45 13.005 94.66 13.075 ;
    RECT 94.45 13.365 94.66 13.435 ;
    RECT 94.45 13.725 94.66 13.795 ;
    RECT 94.91 13.005 95.12 13.075 ;
    RECT 94.91 13.365 95.12 13.435 ;
    RECT 94.91 13.725 95.12 13.795 ;
    RECT 91.13 13.005 91.34 13.075 ;
    RECT 91.13 13.365 91.34 13.435 ;
    RECT 91.13 13.725 91.34 13.795 ;
    RECT 91.59 13.005 91.8 13.075 ;
    RECT 91.59 13.365 91.8 13.435 ;
    RECT 91.59 13.725 91.8 13.795 ;
    RECT 87.81 13.005 88.02 13.075 ;
    RECT 87.81 13.365 88.02 13.435 ;
    RECT 87.81 13.725 88.02 13.795 ;
    RECT 88.27 13.005 88.48 13.075 ;
    RECT 88.27 13.365 88.48 13.435 ;
    RECT 88.27 13.725 88.48 13.795 ;
    RECT 84.49 13.005 84.7 13.075 ;
    RECT 84.49 13.365 84.7 13.435 ;
    RECT 84.49 13.725 84.7 13.795 ;
    RECT 84.95 13.005 85.16 13.075 ;
    RECT 84.95 13.365 85.16 13.435 ;
    RECT 84.95 13.725 85.16 13.795 ;
    RECT 81.17 13.005 81.38 13.075 ;
    RECT 81.17 13.365 81.38 13.435 ;
    RECT 81.17 13.725 81.38 13.795 ;
    RECT 81.63 13.005 81.84 13.075 ;
    RECT 81.63 13.365 81.84 13.435 ;
    RECT 81.63 13.725 81.84 13.795 ;
    RECT 77.85 13.005 78.06 13.075 ;
    RECT 77.85 13.365 78.06 13.435 ;
    RECT 77.85 13.725 78.06 13.795 ;
    RECT 78.31 13.005 78.52 13.075 ;
    RECT 78.31 13.365 78.52 13.435 ;
    RECT 78.31 13.725 78.52 13.795 ;
    RECT 74.53 13.005 74.74 13.075 ;
    RECT 74.53 13.365 74.74 13.435 ;
    RECT 74.53 13.725 74.74 13.795 ;
    RECT 74.99 13.005 75.2 13.075 ;
    RECT 74.99 13.365 75.2 13.435 ;
    RECT 74.99 13.725 75.2 13.795 ;
    RECT 71.21 13.005 71.42 13.075 ;
    RECT 71.21 13.365 71.42 13.435 ;
    RECT 71.21 13.725 71.42 13.795 ;
    RECT 71.67 13.005 71.88 13.075 ;
    RECT 71.67 13.365 71.88 13.435 ;
    RECT 71.67 13.725 71.88 13.795 ;
    RECT 31.37 13.005 31.58 13.075 ;
    RECT 31.37 13.365 31.58 13.435 ;
    RECT 31.37 13.725 31.58 13.795 ;
    RECT 31.83 13.005 32.04 13.075 ;
    RECT 31.83 13.365 32.04 13.435 ;
    RECT 31.83 13.725 32.04 13.795 ;
    RECT 67.89 13.005 68.1 13.075 ;
    RECT 67.89 13.365 68.1 13.435 ;
    RECT 67.89 13.725 68.1 13.795 ;
    RECT 68.35 13.005 68.56 13.075 ;
    RECT 68.35 13.365 68.56 13.435 ;
    RECT 68.35 13.725 68.56 13.795 ;
    RECT 28.05 13.005 28.26 13.075 ;
    RECT 28.05 13.365 28.26 13.435 ;
    RECT 28.05 13.725 28.26 13.795 ;
    RECT 28.51 13.005 28.72 13.075 ;
    RECT 28.51 13.365 28.72 13.435 ;
    RECT 28.51 13.725 28.72 13.795 ;
    RECT 24.73 13.005 24.94 13.075 ;
    RECT 24.73 13.365 24.94 13.435 ;
    RECT 24.73 13.725 24.94 13.795 ;
    RECT 25.19 13.005 25.4 13.075 ;
    RECT 25.19 13.365 25.4 13.435 ;
    RECT 25.19 13.725 25.4 13.795 ;
    RECT 21.41 13.005 21.62 13.075 ;
    RECT 21.41 13.365 21.62 13.435 ;
    RECT 21.41 13.725 21.62 13.795 ;
    RECT 21.87 13.005 22.08 13.075 ;
    RECT 21.87 13.365 22.08 13.435 ;
    RECT 21.87 13.725 22.08 13.795 ;
    RECT 18.09 13.005 18.3 13.075 ;
    RECT 18.09 13.365 18.3 13.435 ;
    RECT 18.09 13.725 18.3 13.795 ;
    RECT 18.55 13.005 18.76 13.075 ;
    RECT 18.55 13.365 18.76 13.435 ;
    RECT 18.55 13.725 18.76 13.795 ;
    RECT 14.77 13.005 14.98 13.075 ;
    RECT 14.77 13.365 14.98 13.435 ;
    RECT 14.77 13.725 14.98 13.795 ;
    RECT 15.23 13.005 15.44 13.075 ;
    RECT 15.23 13.365 15.44 13.435 ;
    RECT 15.23 13.725 15.44 13.795 ;
    RECT 11.45 13.005 11.66 13.075 ;
    RECT 11.45 13.365 11.66 13.435 ;
    RECT 11.45 13.725 11.66 13.795 ;
    RECT 11.91 13.005 12.12 13.075 ;
    RECT 11.91 13.365 12.12 13.435 ;
    RECT 11.91 13.725 12.12 13.795 ;
    RECT 8.13 13.005 8.34 13.075 ;
    RECT 8.13 13.365 8.34 13.435 ;
    RECT 8.13 13.725 8.34 13.795 ;
    RECT 8.59 13.005 8.8 13.075 ;
    RECT 8.59 13.365 8.8 13.435 ;
    RECT 8.59 13.725 8.8 13.795 ;
    RECT 4.81 13.005 5.02 13.075 ;
    RECT 4.81 13.365 5.02 13.435 ;
    RECT 4.81 13.725 5.02 13.795 ;
    RECT 5.27 13.005 5.48 13.075 ;
    RECT 5.27 13.365 5.48 13.435 ;
    RECT 5.27 13.725 5.48 13.795 ;
    RECT 164.17 13.005 164.38 13.075 ;
    RECT 164.17 13.365 164.38 13.435 ;
    RECT 164.17 13.725 164.38 13.795 ;
    RECT 164.63 13.005 164.84 13.075 ;
    RECT 164.63 13.365 164.84 13.435 ;
    RECT 164.63 13.725 164.84 13.795 ;
    RECT 1.49 13.005 1.7 13.075 ;
    RECT 1.49 13.365 1.7 13.435 ;
    RECT 1.49 13.725 1.7 13.795 ;
    RECT 1.95 13.005 2.16 13.075 ;
    RECT 1.95 13.365 2.16 13.435 ;
    RECT 1.95 13.725 2.16 13.795 ;
    RECT 160.85 13.005 161.06 13.075 ;
    RECT 160.85 13.365 161.06 13.435 ;
    RECT 160.85 13.725 161.06 13.795 ;
    RECT 161.31 13.005 161.52 13.075 ;
    RECT 161.31 13.365 161.52 13.435 ;
    RECT 161.31 13.725 161.52 13.795 ;
    RECT 157.53 13.005 157.74 13.075 ;
    RECT 157.53 13.365 157.74 13.435 ;
    RECT 157.53 13.725 157.74 13.795 ;
    RECT 157.99 13.005 158.2 13.075 ;
    RECT 157.99 13.365 158.2 13.435 ;
    RECT 157.99 13.725 158.2 13.795 ;
    RECT 154.21 13.005 154.42 13.075 ;
    RECT 154.21 13.365 154.42 13.435 ;
    RECT 154.21 13.725 154.42 13.795 ;
    RECT 154.67 13.005 154.88 13.075 ;
    RECT 154.67 13.365 154.88 13.435 ;
    RECT 154.67 13.725 154.88 13.795 ;
    RECT 150.89 13.005 151.1 13.075 ;
    RECT 150.89 13.365 151.1 13.435 ;
    RECT 150.89 13.725 151.1 13.795 ;
    RECT 151.35 13.005 151.56 13.075 ;
    RECT 151.35 13.365 151.56 13.435 ;
    RECT 151.35 13.725 151.56 13.795 ;
    RECT 147.57 13.005 147.78 13.075 ;
    RECT 147.57 13.365 147.78 13.435 ;
    RECT 147.57 13.725 147.78 13.795 ;
    RECT 148.03 13.005 148.24 13.075 ;
    RECT 148.03 13.365 148.24 13.435 ;
    RECT 148.03 13.725 148.24 13.795 ;
    RECT 144.25 13.005 144.46 13.075 ;
    RECT 144.25 13.365 144.46 13.435 ;
    RECT 144.25 13.725 144.46 13.795 ;
    RECT 144.71 13.005 144.92 13.075 ;
    RECT 144.71 13.365 144.92 13.435 ;
    RECT 144.71 13.725 144.92 13.795 ;
    RECT 140.93 13.005 141.14 13.075 ;
    RECT 140.93 13.365 141.14 13.435 ;
    RECT 140.93 13.725 141.14 13.795 ;
    RECT 141.39 13.005 141.6 13.075 ;
    RECT 141.39 13.365 141.6 13.435 ;
    RECT 141.39 13.725 141.6 13.795 ;
    RECT 137.61 13.005 137.82 13.075 ;
    RECT 137.61 13.365 137.82 13.435 ;
    RECT 137.61 13.725 137.82 13.795 ;
    RECT 138.07 13.005 138.28 13.075 ;
    RECT 138.07 13.365 138.28 13.435 ;
    RECT 138.07 13.725 138.28 13.795 ;
    RECT 134.29 13.005 134.5 13.075 ;
    RECT 134.29 13.365 134.5 13.435 ;
    RECT 134.29 13.725 134.5 13.795 ;
    RECT 134.75 13.005 134.96 13.075 ;
    RECT 134.75 13.365 134.96 13.435 ;
    RECT 134.75 13.725 134.96 13.795 ;
    RECT 64.57 13.005 64.78 13.075 ;
    RECT 64.57 13.365 64.78 13.435 ;
    RECT 64.57 13.725 64.78 13.795 ;
    RECT 65.03 13.005 65.24 13.075 ;
    RECT 65.03 13.365 65.24 13.435 ;
    RECT 65.03 13.725 65.24 13.795 ;
    RECT 61.25 43.965 61.46 44.035 ;
    RECT 61.25 44.325 61.46 44.395 ;
    RECT 61.25 44.685 61.46 44.755 ;
    RECT 61.71 43.965 61.92 44.035 ;
    RECT 61.71 44.325 61.92 44.395 ;
    RECT 61.71 44.685 61.92 44.755 ;
    RECT 57.93 43.965 58.14 44.035 ;
    RECT 57.93 44.325 58.14 44.395 ;
    RECT 57.93 44.685 58.14 44.755 ;
    RECT 58.39 43.965 58.6 44.035 ;
    RECT 58.39 44.325 58.6 44.395 ;
    RECT 58.39 44.685 58.6 44.755 ;
    RECT 54.61 43.965 54.82 44.035 ;
    RECT 54.61 44.325 54.82 44.395 ;
    RECT 54.61 44.685 54.82 44.755 ;
    RECT 55.07 43.965 55.28 44.035 ;
    RECT 55.07 44.325 55.28 44.395 ;
    RECT 55.07 44.685 55.28 44.755 ;
    RECT 51.29 43.965 51.5 44.035 ;
    RECT 51.29 44.325 51.5 44.395 ;
    RECT 51.29 44.685 51.5 44.755 ;
    RECT 51.75 43.965 51.96 44.035 ;
    RECT 51.75 44.325 51.96 44.395 ;
    RECT 51.75 44.685 51.96 44.755 ;
    RECT 47.97 43.965 48.18 44.035 ;
    RECT 47.97 44.325 48.18 44.395 ;
    RECT 47.97 44.685 48.18 44.755 ;
    RECT 48.43 43.965 48.64 44.035 ;
    RECT 48.43 44.325 48.64 44.395 ;
    RECT 48.43 44.685 48.64 44.755 ;
    RECT 44.65 43.965 44.86 44.035 ;
    RECT 44.65 44.325 44.86 44.395 ;
    RECT 44.65 44.685 44.86 44.755 ;
    RECT 45.11 43.965 45.32 44.035 ;
    RECT 45.11 44.325 45.32 44.395 ;
    RECT 45.11 44.685 45.32 44.755 ;
    RECT 41.33 43.965 41.54 44.035 ;
    RECT 41.33 44.325 41.54 44.395 ;
    RECT 41.33 44.685 41.54 44.755 ;
    RECT 41.79 43.965 42.0 44.035 ;
    RECT 41.79 44.325 42.0 44.395 ;
    RECT 41.79 44.685 42.0 44.755 ;
    RECT 38.01 43.965 38.22 44.035 ;
    RECT 38.01 44.325 38.22 44.395 ;
    RECT 38.01 44.685 38.22 44.755 ;
    RECT 38.47 43.965 38.68 44.035 ;
    RECT 38.47 44.325 38.68 44.395 ;
    RECT 38.47 44.685 38.68 44.755 ;
    RECT 34.69 43.965 34.9 44.035 ;
    RECT 34.69 44.325 34.9 44.395 ;
    RECT 34.69 44.685 34.9 44.755 ;
    RECT 35.15 43.965 35.36 44.035 ;
    RECT 35.15 44.325 35.36 44.395 ;
    RECT 35.15 44.685 35.36 44.755 ;
    RECT 173.945 44.325 174.015 44.395 ;
    RECT 130.97 43.965 131.18 44.035 ;
    RECT 130.97 44.325 131.18 44.395 ;
    RECT 130.97 44.685 131.18 44.755 ;
    RECT 131.43 43.965 131.64 44.035 ;
    RECT 131.43 44.325 131.64 44.395 ;
    RECT 131.43 44.685 131.64 44.755 ;
    RECT 127.65 43.965 127.86 44.035 ;
    RECT 127.65 44.325 127.86 44.395 ;
    RECT 127.65 44.685 127.86 44.755 ;
    RECT 128.11 43.965 128.32 44.035 ;
    RECT 128.11 44.325 128.32 44.395 ;
    RECT 128.11 44.685 128.32 44.755 ;
    RECT 124.33 43.965 124.54 44.035 ;
    RECT 124.33 44.325 124.54 44.395 ;
    RECT 124.33 44.685 124.54 44.755 ;
    RECT 124.79 43.965 125.0 44.035 ;
    RECT 124.79 44.325 125.0 44.395 ;
    RECT 124.79 44.685 125.0 44.755 ;
    RECT 121.01 43.965 121.22 44.035 ;
    RECT 121.01 44.325 121.22 44.395 ;
    RECT 121.01 44.685 121.22 44.755 ;
    RECT 121.47 43.965 121.68 44.035 ;
    RECT 121.47 44.325 121.68 44.395 ;
    RECT 121.47 44.685 121.68 44.755 ;
    RECT 117.69 43.965 117.9 44.035 ;
    RECT 117.69 44.325 117.9 44.395 ;
    RECT 117.69 44.685 117.9 44.755 ;
    RECT 118.15 43.965 118.36 44.035 ;
    RECT 118.15 44.325 118.36 44.395 ;
    RECT 118.15 44.685 118.36 44.755 ;
    RECT 114.37 43.965 114.58 44.035 ;
    RECT 114.37 44.325 114.58 44.395 ;
    RECT 114.37 44.685 114.58 44.755 ;
    RECT 114.83 43.965 115.04 44.035 ;
    RECT 114.83 44.325 115.04 44.395 ;
    RECT 114.83 44.685 115.04 44.755 ;
    RECT 111.05 43.965 111.26 44.035 ;
    RECT 111.05 44.325 111.26 44.395 ;
    RECT 111.05 44.685 111.26 44.755 ;
    RECT 111.51 43.965 111.72 44.035 ;
    RECT 111.51 44.325 111.72 44.395 ;
    RECT 111.51 44.685 111.72 44.755 ;
    RECT 107.73 43.965 107.94 44.035 ;
    RECT 107.73 44.325 107.94 44.395 ;
    RECT 107.73 44.685 107.94 44.755 ;
    RECT 108.19 43.965 108.4 44.035 ;
    RECT 108.19 44.325 108.4 44.395 ;
    RECT 108.19 44.685 108.4 44.755 ;
    RECT 104.41 43.965 104.62 44.035 ;
    RECT 104.41 44.325 104.62 44.395 ;
    RECT 104.41 44.685 104.62 44.755 ;
    RECT 104.87 43.965 105.08 44.035 ;
    RECT 104.87 44.325 105.08 44.395 ;
    RECT 104.87 44.685 105.08 44.755 ;
    RECT 101.09 43.965 101.3 44.035 ;
    RECT 101.09 44.325 101.3 44.395 ;
    RECT 101.09 44.685 101.3 44.755 ;
    RECT 101.55 43.965 101.76 44.035 ;
    RECT 101.55 44.325 101.76 44.395 ;
    RECT 101.55 44.685 101.76 44.755 ;
    RECT 0.4 44.325 0.47 44.395 ;
    RECT 170.81 43.965 171.02 44.035 ;
    RECT 170.81 44.325 171.02 44.395 ;
    RECT 170.81 44.685 171.02 44.755 ;
    RECT 171.27 43.965 171.48 44.035 ;
    RECT 171.27 44.325 171.48 44.395 ;
    RECT 171.27 44.685 171.48 44.755 ;
    RECT 167.49 43.965 167.7 44.035 ;
    RECT 167.49 44.325 167.7 44.395 ;
    RECT 167.49 44.685 167.7 44.755 ;
    RECT 167.95 43.965 168.16 44.035 ;
    RECT 167.95 44.325 168.16 44.395 ;
    RECT 167.95 44.685 168.16 44.755 ;
    RECT 97.77 43.965 97.98 44.035 ;
    RECT 97.77 44.325 97.98 44.395 ;
    RECT 97.77 44.685 97.98 44.755 ;
    RECT 98.23 43.965 98.44 44.035 ;
    RECT 98.23 44.325 98.44 44.395 ;
    RECT 98.23 44.685 98.44 44.755 ;
    RECT 94.45 43.965 94.66 44.035 ;
    RECT 94.45 44.325 94.66 44.395 ;
    RECT 94.45 44.685 94.66 44.755 ;
    RECT 94.91 43.965 95.12 44.035 ;
    RECT 94.91 44.325 95.12 44.395 ;
    RECT 94.91 44.685 95.12 44.755 ;
    RECT 91.13 43.965 91.34 44.035 ;
    RECT 91.13 44.325 91.34 44.395 ;
    RECT 91.13 44.685 91.34 44.755 ;
    RECT 91.59 43.965 91.8 44.035 ;
    RECT 91.59 44.325 91.8 44.395 ;
    RECT 91.59 44.685 91.8 44.755 ;
    RECT 87.81 43.965 88.02 44.035 ;
    RECT 87.81 44.325 88.02 44.395 ;
    RECT 87.81 44.685 88.02 44.755 ;
    RECT 88.27 43.965 88.48 44.035 ;
    RECT 88.27 44.325 88.48 44.395 ;
    RECT 88.27 44.685 88.48 44.755 ;
    RECT 84.49 43.965 84.7 44.035 ;
    RECT 84.49 44.325 84.7 44.395 ;
    RECT 84.49 44.685 84.7 44.755 ;
    RECT 84.95 43.965 85.16 44.035 ;
    RECT 84.95 44.325 85.16 44.395 ;
    RECT 84.95 44.685 85.16 44.755 ;
    RECT 81.17 43.965 81.38 44.035 ;
    RECT 81.17 44.325 81.38 44.395 ;
    RECT 81.17 44.685 81.38 44.755 ;
    RECT 81.63 43.965 81.84 44.035 ;
    RECT 81.63 44.325 81.84 44.395 ;
    RECT 81.63 44.685 81.84 44.755 ;
    RECT 77.85 43.965 78.06 44.035 ;
    RECT 77.85 44.325 78.06 44.395 ;
    RECT 77.85 44.685 78.06 44.755 ;
    RECT 78.31 43.965 78.52 44.035 ;
    RECT 78.31 44.325 78.52 44.395 ;
    RECT 78.31 44.685 78.52 44.755 ;
    RECT 74.53 43.965 74.74 44.035 ;
    RECT 74.53 44.325 74.74 44.395 ;
    RECT 74.53 44.685 74.74 44.755 ;
    RECT 74.99 43.965 75.2 44.035 ;
    RECT 74.99 44.325 75.2 44.395 ;
    RECT 74.99 44.685 75.2 44.755 ;
    RECT 71.21 43.965 71.42 44.035 ;
    RECT 71.21 44.325 71.42 44.395 ;
    RECT 71.21 44.685 71.42 44.755 ;
    RECT 71.67 43.965 71.88 44.035 ;
    RECT 71.67 44.325 71.88 44.395 ;
    RECT 71.67 44.685 71.88 44.755 ;
    RECT 31.37 43.965 31.58 44.035 ;
    RECT 31.37 44.325 31.58 44.395 ;
    RECT 31.37 44.685 31.58 44.755 ;
    RECT 31.83 43.965 32.04 44.035 ;
    RECT 31.83 44.325 32.04 44.395 ;
    RECT 31.83 44.685 32.04 44.755 ;
    RECT 67.89 43.965 68.1 44.035 ;
    RECT 67.89 44.325 68.1 44.395 ;
    RECT 67.89 44.685 68.1 44.755 ;
    RECT 68.35 43.965 68.56 44.035 ;
    RECT 68.35 44.325 68.56 44.395 ;
    RECT 68.35 44.685 68.56 44.755 ;
    RECT 28.05 43.965 28.26 44.035 ;
    RECT 28.05 44.325 28.26 44.395 ;
    RECT 28.05 44.685 28.26 44.755 ;
    RECT 28.51 43.965 28.72 44.035 ;
    RECT 28.51 44.325 28.72 44.395 ;
    RECT 28.51 44.685 28.72 44.755 ;
    RECT 24.73 43.965 24.94 44.035 ;
    RECT 24.73 44.325 24.94 44.395 ;
    RECT 24.73 44.685 24.94 44.755 ;
    RECT 25.19 43.965 25.4 44.035 ;
    RECT 25.19 44.325 25.4 44.395 ;
    RECT 25.19 44.685 25.4 44.755 ;
    RECT 21.41 43.965 21.62 44.035 ;
    RECT 21.41 44.325 21.62 44.395 ;
    RECT 21.41 44.685 21.62 44.755 ;
    RECT 21.87 43.965 22.08 44.035 ;
    RECT 21.87 44.325 22.08 44.395 ;
    RECT 21.87 44.685 22.08 44.755 ;
    RECT 18.09 43.965 18.3 44.035 ;
    RECT 18.09 44.325 18.3 44.395 ;
    RECT 18.09 44.685 18.3 44.755 ;
    RECT 18.55 43.965 18.76 44.035 ;
    RECT 18.55 44.325 18.76 44.395 ;
    RECT 18.55 44.685 18.76 44.755 ;
    RECT 14.77 43.965 14.98 44.035 ;
    RECT 14.77 44.325 14.98 44.395 ;
    RECT 14.77 44.685 14.98 44.755 ;
    RECT 15.23 43.965 15.44 44.035 ;
    RECT 15.23 44.325 15.44 44.395 ;
    RECT 15.23 44.685 15.44 44.755 ;
    RECT 11.45 43.965 11.66 44.035 ;
    RECT 11.45 44.325 11.66 44.395 ;
    RECT 11.45 44.685 11.66 44.755 ;
    RECT 11.91 43.965 12.12 44.035 ;
    RECT 11.91 44.325 12.12 44.395 ;
    RECT 11.91 44.685 12.12 44.755 ;
    RECT 8.13 43.965 8.34 44.035 ;
    RECT 8.13 44.325 8.34 44.395 ;
    RECT 8.13 44.685 8.34 44.755 ;
    RECT 8.59 43.965 8.8 44.035 ;
    RECT 8.59 44.325 8.8 44.395 ;
    RECT 8.59 44.685 8.8 44.755 ;
    RECT 4.81 43.965 5.02 44.035 ;
    RECT 4.81 44.325 5.02 44.395 ;
    RECT 4.81 44.685 5.02 44.755 ;
    RECT 5.27 43.965 5.48 44.035 ;
    RECT 5.27 44.325 5.48 44.395 ;
    RECT 5.27 44.685 5.48 44.755 ;
    RECT 164.17 43.965 164.38 44.035 ;
    RECT 164.17 44.325 164.38 44.395 ;
    RECT 164.17 44.685 164.38 44.755 ;
    RECT 164.63 43.965 164.84 44.035 ;
    RECT 164.63 44.325 164.84 44.395 ;
    RECT 164.63 44.685 164.84 44.755 ;
    RECT 1.49 43.965 1.7 44.035 ;
    RECT 1.49 44.325 1.7 44.395 ;
    RECT 1.49 44.685 1.7 44.755 ;
    RECT 1.95 43.965 2.16 44.035 ;
    RECT 1.95 44.325 2.16 44.395 ;
    RECT 1.95 44.685 2.16 44.755 ;
    RECT 160.85 43.965 161.06 44.035 ;
    RECT 160.85 44.325 161.06 44.395 ;
    RECT 160.85 44.685 161.06 44.755 ;
    RECT 161.31 43.965 161.52 44.035 ;
    RECT 161.31 44.325 161.52 44.395 ;
    RECT 161.31 44.685 161.52 44.755 ;
    RECT 157.53 43.965 157.74 44.035 ;
    RECT 157.53 44.325 157.74 44.395 ;
    RECT 157.53 44.685 157.74 44.755 ;
    RECT 157.99 43.965 158.2 44.035 ;
    RECT 157.99 44.325 158.2 44.395 ;
    RECT 157.99 44.685 158.2 44.755 ;
    RECT 154.21 43.965 154.42 44.035 ;
    RECT 154.21 44.325 154.42 44.395 ;
    RECT 154.21 44.685 154.42 44.755 ;
    RECT 154.67 43.965 154.88 44.035 ;
    RECT 154.67 44.325 154.88 44.395 ;
    RECT 154.67 44.685 154.88 44.755 ;
    RECT 150.89 43.965 151.1 44.035 ;
    RECT 150.89 44.325 151.1 44.395 ;
    RECT 150.89 44.685 151.1 44.755 ;
    RECT 151.35 43.965 151.56 44.035 ;
    RECT 151.35 44.325 151.56 44.395 ;
    RECT 151.35 44.685 151.56 44.755 ;
    RECT 147.57 43.965 147.78 44.035 ;
    RECT 147.57 44.325 147.78 44.395 ;
    RECT 147.57 44.685 147.78 44.755 ;
    RECT 148.03 43.965 148.24 44.035 ;
    RECT 148.03 44.325 148.24 44.395 ;
    RECT 148.03 44.685 148.24 44.755 ;
    RECT 144.25 43.965 144.46 44.035 ;
    RECT 144.25 44.325 144.46 44.395 ;
    RECT 144.25 44.685 144.46 44.755 ;
    RECT 144.71 43.965 144.92 44.035 ;
    RECT 144.71 44.325 144.92 44.395 ;
    RECT 144.71 44.685 144.92 44.755 ;
    RECT 140.93 43.965 141.14 44.035 ;
    RECT 140.93 44.325 141.14 44.395 ;
    RECT 140.93 44.685 141.14 44.755 ;
    RECT 141.39 43.965 141.6 44.035 ;
    RECT 141.39 44.325 141.6 44.395 ;
    RECT 141.39 44.685 141.6 44.755 ;
    RECT 137.61 43.965 137.82 44.035 ;
    RECT 137.61 44.325 137.82 44.395 ;
    RECT 137.61 44.685 137.82 44.755 ;
    RECT 138.07 43.965 138.28 44.035 ;
    RECT 138.07 44.325 138.28 44.395 ;
    RECT 138.07 44.685 138.28 44.755 ;
    RECT 134.29 43.965 134.5 44.035 ;
    RECT 134.29 44.325 134.5 44.395 ;
    RECT 134.29 44.685 134.5 44.755 ;
    RECT 134.75 43.965 134.96 44.035 ;
    RECT 134.75 44.325 134.96 44.395 ;
    RECT 134.75 44.685 134.96 44.755 ;
    RECT 64.57 43.965 64.78 44.035 ;
    RECT 64.57 44.325 64.78 44.395 ;
    RECT 64.57 44.685 64.78 44.755 ;
    RECT 65.03 43.965 65.24 44.035 ;
    RECT 65.03 44.325 65.24 44.395 ;
    RECT 65.03 44.685 65.24 44.755 ;
    RECT 61.25 12.285 61.46 12.355 ;
    RECT 61.25 12.645 61.46 12.715 ;
    RECT 61.25 13.005 61.46 13.075 ;
    RECT 61.71 12.285 61.92 12.355 ;
    RECT 61.71 12.645 61.92 12.715 ;
    RECT 61.71 13.005 61.92 13.075 ;
    RECT 57.93 12.285 58.14 12.355 ;
    RECT 57.93 12.645 58.14 12.715 ;
    RECT 57.93 13.005 58.14 13.075 ;
    RECT 58.39 12.285 58.6 12.355 ;
    RECT 58.39 12.645 58.6 12.715 ;
    RECT 58.39 13.005 58.6 13.075 ;
    RECT 54.61 12.285 54.82 12.355 ;
    RECT 54.61 12.645 54.82 12.715 ;
    RECT 54.61 13.005 54.82 13.075 ;
    RECT 55.07 12.285 55.28 12.355 ;
    RECT 55.07 12.645 55.28 12.715 ;
    RECT 55.07 13.005 55.28 13.075 ;
    RECT 51.29 12.285 51.5 12.355 ;
    RECT 51.29 12.645 51.5 12.715 ;
    RECT 51.29 13.005 51.5 13.075 ;
    RECT 51.75 12.285 51.96 12.355 ;
    RECT 51.75 12.645 51.96 12.715 ;
    RECT 51.75 13.005 51.96 13.075 ;
    RECT 47.97 12.285 48.18 12.355 ;
    RECT 47.97 12.645 48.18 12.715 ;
    RECT 47.97 13.005 48.18 13.075 ;
    RECT 48.43 12.285 48.64 12.355 ;
    RECT 48.43 12.645 48.64 12.715 ;
    RECT 48.43 13.005 48.64 13.075 ;
    RECT 44.65 12.285 44.86 12.355 ;
    RECT 44.65 12.645 44.86 12.715 ;
    RECT 44.65 13.005 44.86 13.075 ;
    RECT 45.11 12.285 45.32 12.355 ;
    RECT 45.11 12.645 45.32 12.715 ;
    RECT 45.11 13.005 45.32 13.075 ;
    RECT 41.33 12.285 41.54 12.355 ;
    RECT 41.33 12.645 41.54 12.715 ;
    RECT 41.33 13.005 41.54 13.075 ;
    RECT 41.79 12.285 42.0 12.355 ;
    RECT 41.79 12.645 42.0 12.715 ;
    RECT 41.79 13.005 42.0 13.075 ;
    RECT 38.01 12.285 38.22 12.355 ;
    RECT 38.01 12.645 38.22 12.715 ;
    RECT 38.01 13.005 38.22 13.075 ;
    RECT 38.47 12.285 38.68 12.355 ;
    RECT 38.47 12.645 38.68 12.715 ;
    RECT 38.47 13.005 38.68 13.075 ;
    RECT 34.69 12.285 34.9 12.355 ;
    RECT 34.69 12.645 34.9 12.715 ;
    RECT 34.69 13.005 34.9 13.075 ;
    RECT 35.15 12.285 35.36 12.355 ;
    RECT 35.15 12.645 35.36 12.715 ;
    RECT 35.15 13.005 35.36 13.075 ;
    RECT 173.945 12.645 174.015 12.715 ;
    RECT 130.97 12.285 131.18 12.355 ;
    RECT 130.97 12.645 131.18 12.715 ;
    RECT 130.97 13.005 131.18 13.075 ;
    RECT 131.43 12.285 131.64 12.355 ;
    RECT 131.43 12.645 131.64 12.715 ;
    RECT 131.43 13.005 131.64 13.075 ;
    RECT 127.65 12.285 127.86 12.355 ;
    RECT 127.65 12.645 127.86 12.715 ;
    RECT 127.65 13.005 127.86 13.075 ;
    RECT 128.11 12.285 128.32 12.355 ;
    RECT 128.11 12.645 128.32 12.715 ;
    RECT 128.11 13.005 128.32 13.075 ;
    RECT 124.33 12.285 124.54 12.355 ;
    RECT 124.33 12.645 124.54 12.715 ;
    RECT 124.33 13.005 124.54 13.075 ;
    RECT 124.79 12.285 125.0 12.355 ;
    RECT 124.79 12.645 125.0 12.715 ;
    RECT 124.79 13.005 125.0 13.075 ;
    RECT 121.01 12.285 121.22 12.355 ;
    RECT 121.01 12.645 121.22 12.715 ;
    RECT 121.01 13.005 121.22 13.075 ;
    RECT 121.47 12.285 121.68 12.355 ;
    RECT 121.47 12.645 121.68 12.715 ;
    RECT 121.47 13.005 121.68 13.075 ;
    RECT 117.69 12.285 117.9 12.355 ;
    RECT 117.69 12.645 117.9 12.715 ;
    RECT 117.69 13.005 117.9 13.075 ;
    RECT 118.15 12.285 118.36 12.355 ;
    RECT 118.15 12.645 118.36 12.715 ;
    RECT 118.15 13.005 118.36 13.075 ;
    RECT 114.37 12.285 114.58 12.355 ;
    RECT 114.37 12.645 114.58 12.715 ;
    RECT 114.37 13.005 114.58 13.075 ;
    RECT 114.83 12.285 115.04 12.355 ;
    RECT 114.83 12.645 115.04 12.715 ;
    RECT 114.83 13.005 115.04 13.075 ;
    RECT 111.05 12.285 111.26 12.355 ;
    RECT 111.05 12.645 111.26 12.715 ;
    RECT 111.05 13.005 111.26 13.075 ;
    RECT 111.51 12.285 111.72 12.355 ;
    RECT 111.51 12.645 111.72 12.715 ;
    RECT 111.51 13.005 111.72 13.075 ;
    RECT 107.73 12.285 107.94 12.355 ;
    RECT 107.73 12.645 107.94 12.715 ;
    RECT 107.73 13.005 107.94 13.075 ;
    RECT 108.19 12.285 108.4 12.355 ;
    RECT 108.19 12.645 108.4 12.715 ;
    RECT 108.19 13.005 108.4 13.075 ;
    RECT 104.41 12.285 104.62 12.355 ;
    RECT 104.41 12.645 104.62 12.715 ;
    RECT 104.41 13.005 104.62 13.075 ;
    RECT 104.87 12.285 105.08 12.355 ;
    RECT 104.87 12.645 105.08 12.715 ;
    RECT 104.87 13.005 105.08 13.075 ;
    RECT 101.09 12.285 101.3 12.355 ;
    RECT 101.09 12.645 101.3 12.715 ;
    RECT 101.09 13.005 101.3 13.075 ;
    RECT 101.55 12.285 101.76 12.355 ;
    RECT 101.55 12.645 101.76 12.715 ;
    RECT 101.55 13.005 101.76 13.075 ;
    RECT 0.4 12.645 0.47 12.715 ;
    RECT 170.81 12.285 171.02 12.355 ;
    RECT 170.81 12.645 171.02 12.715 ;
    RECT 170.81 13.005 171.02 13.075 ;
    RECT 171.27 12.285 171.48 12.355 ;
    RECT 171.27 12.645 171.48 12.715 ;
    RECT 171.27 13.005 171.48 13.075 ;
    RECT 167.49 12.285 167.7 12.355 ;
    RECT 167.49 12.645 167.7 12.715 ;
    RECT 167.49 13.005 167.7 13.075 ;
    RECT 167.95 12.285 168.16 12.355 ;
    RECT 167.95 12.645 168.16 12.715 ;
    RECT 167.95 13.005 168.16 13.075 ;
    RECT 97.77 12.285 97.98 12.355 ;
    RECT 97.77 12.645 97.98 12.715 ;
    RECT 97.77 13.005 97.98 13.075 ;
    RECT 98.23 12.285 98.44 12.355 ;
    RECT 98.23 12.645 98.44 12.715 ;
    RECT 98.23 13.005 98.44 13.075 ;
    RECT 94.45 12.285 94.66 12.355 ;
    RECT 94.45 12.645 94.66 12.715 ;
    RECT 94.45 13.005 94.66 13.075 ;
    RECT 94.91 12.285 95.12 12.355 ;
    RECT 94.91 12.645 95.12 12.715 ;
    RECT 94.91 13.005 95.12 13.075 ;
    RECT 91.13 12.285 91.34 12.355 ;
    RECT 91.13 12.645 91.34 12.715 ;
    RECT 91.13 13.005 91.34 13.075 ;
    RECT 91.59 12.285 91.8 12.355 ;
    RECT 91.59 12.645 91.8 12.715 ;
    RECT 91.59 13.005 91.8 13.075 ;
    RECT 87.81 12.285 88.02 12.355 ;
    RECT 87.81 12.645 88.02 12.715 ;
    RECT 87.81 13.005 88.02 13.075 ;
    RECT 88.27 12.285 88.48 12.355 ;
    RECT 88.27 12.645 88.48 12.715 ;
    RECT 88.27 13.005 88.48 13.075 ;
    RECT 84.49 12.285 84.7 12.355 ;
    RECT 84.49 12.645 84.7 12.715 ;
    RECT 84.49 13.005 84.7 13.075 ;
    RECT 84.95 12.285 85.16 12.355 ;
    RECT 84.95 12.645 85.16 12.715 ;
    RECT 84.95 13.005 85.16 13.075 ;
    RECT 81.17 12.285 81.38 12.355 ;
    RECT 81.17 12.645 81.38 12.715 ;
    RECT 81.17 13.005 81.38 13.075 ;
    RECT 81.63 12.285 81.84 12.355 ;
    RECT 81.63 12.645 81.84 12.715 ;
    RECT 81.63 13.005 81.84 13.075 ;
    RECT 77.85 12.285 78.06 12.355 ;
    RECT 77.85 12.645 78.06 12.715 ;
    RECT 77.85 13.005 78.06 13.075 ;
    RECT 78.31 12.285 78.52 12.355 ;
    RECT 78.31 12.645 78.52 12.715 ;
    RECT 78.31 13.005 78.52 13.075 ;
    RECT 74.53 12.285 74.74 12.355 ;
    RECT 74.53 12.645 74.74 12.715 ;
    RECT 74.53 13.005 74.74 13.075 ;
    RECT 74.99 12.285 75.2 12.355 ;
    RECT 74.99 12.645 75.2 12.715 ;
    RECT 74.99 13.005 75.2 13.075 ;
    RECT 71.21 12.285 71.42 12.355 ;
    RECT 71.21 12.645 71.42 12.715 ;
    RECT 71.21 13.005 71.42 13.075 ;
    RECT 71.67 12.285 71.88 12.355 ;
    RECT 71.67 12.645 71.88 12.715 ;
    RECT 71.67 13.005 71.88 13.075 ;
    RECT 31.37 12.285 31.58 12.355 ;
    RECT 31.37 12.645 31.58 12.715 ;
    RECT 31.37 13.005 31.58 13.075 ;
    RECT 31.83 12.285 32.04 12.355 ;
    RECT 31.83 12.645 32.04 12.715 ;
    RECT 31.83 13.005 32.04 13.075 ;
    RECT 67.89 12.285 68.1 12.355 ;
    RECT 67.89 12.645 68.1 12.715 ;
    RECT 67.89 13.005 68.1 13.075 ;
    RECT 68.35 12.285 68.56 12.355 ;
    RECT 68.35 12.645 68.56 12.715 ;
    RECT 68.35 13.005 68.56 13.075 ;
    RECT 28.05 12.285 28.26 12.355 ;
    RECT 28.05 12.645 28.26 12.715 ;
    RECT 28.05 13.005 28.26 13.075 ;
    RECT 28.51 12.285 28.72 12.355 ;
    RECT 28.51 12.645 28.72 12.715 ;
    RECT 28.51 13.005 28.72 13.075 ;
    RECT 24.73 12.285 24.94 12.355 ;
    RECT 24.73 12.645 24.94 12.715 ;
    RECT 24.73 13.005 24.94 13.075 ;
    RECT 25.19 12.285 25.4 12.355 ;
    RECT 25.19 12.645 25.4 12.715 ;
    RECT 25.19 13.005 25.4 13.075 ;
    RECT 21.41 12.285 21.62 12.355 ;
    RECT 21.41 12.645 21.62 12.715 ;
    RECT 21.41 13.005 21.62 13.075 ;
    RECT 21.87 12.285 22.08 12.355 ;
    RECT 21.87 12.645 22.08 12.715 ;
    RECT 21.87 13.005 22.08 13.075 ;
    RECT 18.09 12.285 18.3 12.355 ;
    RECT 18.09 12.645 18.3 12.715 ;
    RECT 18.09 13.005 18.3 13.075 ;
    RECT 18.55 12.285 18.76 12.355 ;
    RECT 18.55 12.645 18.76 12.715 ;
    RECT 18.55 13.005 18.76 13.075 ;
    RECT 14.77 12.285 14.98 12.355 ;
    RECT 14.77 12.645 14.98 12.715 ;
    RECT 14.77 13.005 14.98 13.075 ;
    RECT 15.23 12.285 15.44 12.355 ;
    RECT 15.23 12.645 15.44 12.715 ;
    RECT 15.23 13.005 15.44 13.075 ;
    RECT 11.45 12.285 11.66 12.355 ;
    RECT 11.45 12.645 11.66 12.715 ;
    RECT 11.45 13.005 11.66 13.075 ;
    RECT 11.91 12.285 12.12 12.355 ;
    RECT 11.91 12.645 12.12 12.715 ;
    RECT 11.91 13.005 12.12 13.075 ;
    RECT 8.13 12.285 8.34 12.355 ;
    RECT 8.13 12.645 8.34 12.715 ;
    RECT 8.13 13.005 8.34 13.075 ;
    RECT 8.59 12.285 8.8 12.355 ;
    RECT 8.59 12.645 8.8 12.715 ;
    RECT 8.59 13.005 8.8 13.075 ;
    RECT 4.81 12.285 5.02 12.355 ;
    RECT 4.81 12.645 5.02 12.715 ;
    RECT 4.81 13.005 5.02 13.075 ;
    RECT 5.27 12.285 5.48 12.355 ;
    RECT 5.27 12.645 5.48 12.715 ;
    RECT 5.27 13.005 5.48 13.075 ;
    RECT 164.17 12.285 164.38 12.355 ;
    RECT 164.17 12.645 164.38 12.715 ;
    RECT 164.17 13.005 164.38 13.075 ;
    RECT 164.63 12.285 164.84 12.355 ;
    RECT 164.63 12.645 164.84 12.715 ;
    RECT 164.63 13.005 164.84 13.075 ;
    RECT 1.49 12.285 1.7 12.355 ;
    RECT 1.49 12.645 1.7 12.715 ;
    RECT 1.49 13.005 1.7 13.075 ;
    RECT 1.95 12.285 2.16 12.355 ;
    RECT 1.95 12.645 2.16 12.715 ;
    RECT 1.95 13.005 2.16 13.075 ;
    RECT 160.85 12.285 161.06 12.355 ;
    RECT 160.85 12.645 161.06 12.715 ;
    RECT 160.85 13.005 161.06 13.075 ;
    RECT 161.31 12.285 161.52 12.355 ;
    RECT 161.31 12.645 161.52 12.715 ;
    RECT 161.31 13.005 161.52 13.075 ;
    RECT 157.53 12.285 157.74 12.355 ;
    RECT 157.53 12.645 157.74 12.715 ;
    RECT 157.53 13.005 157.74 13.075 ;
    RECT 157.99 12.285 158.2 12.355 ;
    RECT 157.99 12.645 158.2 12.715 ;
    RECT 157.99 13.005 158.2 13.075 ;
    RECT 154.21 12.285 154.42 12.355 ;
    RECT 154.21 12.645 154.42 12.715 ;
    RECT 154.21 13.005 154.42 13.075 ;
    RECT 154.67 12.285 154.88 12.355 ;
    RECT 154.67 12.645 154.88 12.715 ;
    RECT 154.67 13.005 154.88 13.075 ;
    RECT 150.89 12.285 151.1 12.355 ;
    RECT 150.89 12.645 151.1 12.715 ;
    RECT 150.89 13.005 151.1 13.075 ;
    RECT 151.35 12.285 151.56 12.355 ;
    RECT 151.35 12.645 151.56 12.715 ;
    RECT 151.35 13.005 151.56 13.075 ;
    RECT 147.57 12.285 147.78 12.355 ;
    RECT 147.57 12.645 147.78 12.715 ;
    RECT 147.57 13.005 147.78 13.075 ;
    RECT 148.03 12.285 148.24 12.355 ;
    RECT 148.03 12.645 148.24 12.715 ;
    RECT 148.03 13.005 148.24 13.075 ;
    RECT 144.25 12.285 144.46 12.355 ;
    RECT 144.25 12.645 144.46 12.715 ;
    RECT 144.25 13.005 144.46 13.075 ;
    RECT 144.71 12.285 144.92 12.355 ;
    RECT 144.71 12.645 144.92 12.715 ;
    RECT 144.71 13.005 144.92 13.075 ;
    RECT 140.93 12.285 141.14 12.355 ;
    RECT 140.93 12.645 141.14 12.715 ;
    RECT 140.93 13.005 141.14 13.075 ;
    RECT 141.39 12.285 141.6 12.355 ;
    RECT 141.39 12.645 141.6 12.715 ;
    RECT 141.39 13.005 141.6 13.075 ;
    RECT 137.61 12.285 137.82 12.355 ;
    RECT 137.61 12.645 137.82 12.715 ;
    RECT 137.61 13.005 137.82 13.075 ;
    RECT 138.07 12.285 138.28 12.355 ;
    RECT 138.07 12.645 138.28 12.715 ;
    RECT 138.07 13.005 138.28 13.075 ;
    RECT 134.29 12.285 134.5 12.355 ;
    RECT 134.29 12.645 134.5 12.715 ;
    RECT 134.29 13.005 134.5 13.075 ;
    RECT 134.75 12.285 134.96 12.355 ;
    RECT 134.75 12.645 134.96 12.715 ;
    RECT 134.75 13.005 134.96 13.075 ;
    RECT 64.57 12.285 64.78 12.355 ;
    RECT 64.57 12.645 64.78 12.715 ;
    RECT 64.57 13.005 64.78 13.075 ;
    RECT 65.03 12.285 65.24 12.355 ;
    RECT 65.03 12.645 65.24 12.715 ;
    RECT 65.03 13.005 65.24 13.075 ;
    RECT 61.25 43.245 61.46 43.315 ;
    RECT 61.25 43.605 61.46 43.675 ;
    RECT 61.25 43.965 61.46 44.035 ;
    RECT 61.71 43.245 61.92 43.315 ;
    RECT 61.71 43.605 61.92 43.675 ;
    RECT 61.71 43.965 61.92 44.035 ;
    RECT 57.93 43.245 58.14 43.315 ;
    RECT 57.93 43.605 58.14 43.675 ;
    RECT 57.93 43.965 58.14 44.035 ;
    RECT 58.39 43.245 58.6 43.315 ;
    RECT 58.39 43.605 58.6 43.675 ;
    RECT 58.39 43.965 58.6 44.035 ;
    RECT 54.61 43.245 54.82 43.315 ;
    RECT 54.61 43.605 54.82 43.675 ;
    RECT 54.61 43.965 54.82 44.035 ;
    RECT 55.07 43.245 55.28 43.315 ;
    RECT 55.07 43.605 55.28 43.675 ;
    RECT 55.07 43.965 55.28 44.035 ;
    RECT 51.29 43.245 51.5 43.315 ;
    RECT 51.29 43.605 51.5 43.675 ;
    RECT 51.29 43.965 51.5 44.035 ;
    RECT 51.75 43.245 51.96 43.315 ;
    RECT 51.75 43.605 51.96 43.675 ;
    RECT 51.75 43.965 51.96 44.035 ;
    RECT 47.97 43.245 48.18 43.315 ;
    RECT 47.97 43.605 48.18 43.675 ;
    RECT 47.97 43.965 48.18 44.035 ;
    RECT 48.43 43.245 48.64 43.315 ;
    RECT 48.43 43.605 48.64 43.675 ;
    RECT 48.43 43.965 48.64 44.035 ;
    RECT 44.65 43.245 44.86 43.315 ;
    RECT 44.65 43.605 44.86 43.675 ;
    RECT 44.65 43.965 44.86 44.035 ;
    RECT 45.11 43.245 45.32 43.315 ;
    RECT 45.11 43.605 45.32 43.675 ;
    RECT 45.11 43.965 45.32 44.035 ;
    RECT 41.33 43.245 41.54 43.315 ;
    RECT 41.33 43.605 41.54 43.675 ;
    RECT 41.33 43.965 41.54 44.035 ;
    RECT 41.79 43.245 42.0 43.315 ;
    RECT 41.79 43.605 42.0 43.675 ;
    RECT 41.79 43.965 42.0 44.035 ;
    RECT 38.01 43.245 38.22 43.315 ;
    RECT 38.01 43.605 38.22 43.675 ;
    RECT 38.01 43.965 38.22 44.035 ;
    RECT 38.47 43.245 38.68 43.315 ;
    RECT 38.47 43.605 38.68 43.675 ;
    RECT 38.47 43.965 38.68 44.035 ;
    RECT 34.69 43.245 34.9 43.315 ;
    RECT 34.69 43.605 34.9 43.675 ;
    RECT 34.69 43.965 34.9 44.035 ;
    RECT 35.15 43.245 35.36 43.315 ;
    RECT 35.15 43.605 35.36 43.675 ;
    RECT 35.15 43.965 35.36 44.035 ;
    RECT 173.945 43.605 174.015 43.675 ;
    RECT 130.97 43.245 131.18 43.315 ;
    RECT 130.97 43.605 131.18 43.675 ;
    RECT 130.97 43.965 131.18 44.035 ;
    RECT 131.43 43.245 131.64 43.315 ;
    RECT 131.43 43.605 131.64 43.675 ;
    RECT 131.43 43.965 131.64 44.035 ;
    RECT 127.65 43.245 127.86 43.315 ;
    RECT 127.65 43.605 127.86 43.675 ;
    RECT 127.65 43.965 127.86 44.035 ;
    RECT 128.11 43.245 128.32 43.315 ;
    RECT 128.11 43.605 128.32 43.675 ;
    RECT 128.11 43.965 128.32 44.035 ;
    RECT 124.33 43.245 124.54 43.315 ;
    RECT 124.33 43.605 124.54 43.675 ;
    RECT 124.33 43.965 124.54 44.035 ;
    RECT 124.79 43.245 125.0 43.315 ;
    RECT 124.79 43.605 125.0 43.675 ;
    RECT 124.79 43.965 125.0 44.035 ;
    RECT 121.01 43.245 121.22 43.315 ;
    RECT 121.01 43.605 121.22 43.675 ;
    RECT 121.01 43.965 121.22 44.035 ;
    RECT 121.47 43.245 121.68 43.315 ;
    RECT 121.47 43.605 121.68 43.675 ;
    RECT 121.47 43.965 121.68 44.035 ;
    RECT 117.69 43.245 117.9 43.315 ;
    RECT 117.69 43.605 117.9 43.675 ;
    RECT 117.69 43.965 117.9 44.035 ;
    RECT 118.15 43.245 118.36 43.315 ;
    RECT 118.15 43.605 118.36 43.675 ;
    RECT 118.15 43.965 118.36 44.035 ;
    RECT 114.37 43.245 114.58 43.315 ;
    RECT 114.37 43.605 114.58 43.675 ;
    RECT 114.37 43.965 114.58 44.035 ;
    RECT 114.83 43.245 115.04 43.315 ;
    RECT 114.83 43.605 115.04 43.675 ;
    RECT 114.83 43.965 115.04 44.035 ;
    RECT 111.05 43.245 111.26 43.315 ;
    RECT 111.05 43.605 111.26 43.675 ;
    RECT 111.05 43.965 111.26 44.035 ;
    RECT 111.51 43.245 111.72 43.315 ;
    RECT 111.51 43.605 111.72 43.675 ;
    RECT 111.51 43.965 111.72 44.035 ;
    RECT 107.73 43.245 107.94 43.315 ;
    RECT 107.73 43.605 107.94 43.675 ;
    RECT 107.73 43.965 107.94 44.035 ;
    RECT 108.19 43.245 108.4 43.315 ;
    RECT 108.19 43.605 108.4 43.675 ;
    RECT 108.19 43.965 108.4 44.035 ;
    RECT 104.41 43.245 104.62 43.315 ;
    RECT 104.41 43.605 104.62 43.675 ;
    RECT 104.41 43.965 104.62 44.035 ;
    RECT 104.87 43.245 105.08 43.315 ;
    RECT 104.87 43.605 105.08 43.675 ;
    RECT 104.87 43.965 105.08 44.035 ;
    RECT 101.09 43.245 101.3 43.315 ;
    RECT 101.09 43.605 101.3 43.675 ;
    RECT 101.09 43.965 101.3 44.035 ;
    RECT 101.55 43.245 101.76 43.315 ;
    RECT 101.55 43.605 101.76 43.675 ;
    RECT 101.55 43.965 101.76 44.035 ;
    RECT 0.4 43.605 0.47 43.675 ;
    RECT 170.81 43.245 171.02 43.315 ;
    RECT 170.81 43.605 171.02 43.675 ;
    RECT 170.81 43.965 171.02 44.035 ;
    RECT 171.27 43.245 171.48 43.315 ;
    RECT 171.27 43.605 171.48 43.675 ;
    RECT 171.27 43.965 171.48 44.035 ;
    RECT 167.49 43.245 167.7 43.315 ;
    RECT 167.49 43.605 167.7 43.675 ;
    RECT 167.49 43.965 167.7 44.035 ;
    RECT 167.95 43.245 168.16 43.315 ;
    RECT 167.95 43.605 168.16 43.675 ;
    RECT 167.95 43.965 168.16 44.035 ;
    RECT 97.77 43.245 97.98 43.315 ;
    RECT 97.77 43.605 97.98 43.675 ;
    RECT 97.77 43.965 97.98 44.035 ;
    RECT 98.23 43.245 98.44 43.315 ;
    RECT 98.23 43.605 98.44 43.675 ;
    RECT 98.23 43.965 98.44 44.035 ;
    RECT 94.45 43.245 94.66 43.315 ;
    RECT 94.45 43.605 94.66 43.675 ;
    RECT 94.45 43.965 94.66 44.035 ;
    RECT 94.91 43.245 95.12 43.315 ;
    RECT 94.91 43.605 95.12 43.675 ;
    RECT 94.91 43.965 95.12 44.035 ;
    RECT 91.13 43.245 91.34 43.315 ;
    RECT 91.13 43.605 91.34 43.675 ;
    RECT 91.13 43.965 91.34 44.035 ;
    RECT 91.59 43.245 91.8 43.315 ;
    RECT 91.59 43.605 91.8 43.675 ;
    RECT 91.59 43.965 91.8 44.035 ;
    RECT 87.81 43.245 88.02 43.315 ;
    RECT 87.81 43.605 88.02 43.675 ;
    RECT 87.81 43.965 88.02 44.035 ;
    RECT 88.27 43.245 88.48 43.315 ;
    RECT 88.27 43.605 88.48 43.675 ;
    RECT 88.27 43.965 88.48 44.035 ;
    RECT 84.49 43.245 84.7 43.315 ;
    RECT 84.49 43.605 84.7 43.675 ;
    RECT 84.49 43.965 84.7 44.035 ;
    RECT 84.95 43.245 85.16 43.315 ;
    RECT 84.95 43.605 85.16 43.675 ;
    RECT 84.95 43.965 85.16 44.035 ;
    RECT 81.17 43.245 81.38 43.315 ;
    RECT 81.17 43.605 81.38 43.675 ;
    RECT 81.17 43.965 81.38 44.035 ;
    RECT 81.63 43.245 81.84 43.315 ;
    RECT 81.63 43.605 81.84 43.675 ;
    RECT 81.63 43.965 81.84 44.035 ;
    RECT 77.85 43.245 78.06 43.315 ;
    RECT 77.85 43.605 78.06 43.675 ;
    RECT 77.85 43.965 78.06 44.035 ;
    RECT 78.31 43.245 78.52 43.315 ;
    RECT 78.31 43.605 78.52 43.675 ;
    RECT 78.31 43.965 78.52 44.035 ;
    RECT 74.53 43.245 74.74 43.315 ;
    RECT 74.53 43.605 74.74 43.675 ;
    RECT 74.53 43.965 74.74 44.035 ;
    RECT 74.99 43.245 75.2 43.315 ;
    RECT 74.99 43.605 75.2 43.675 ;
    RECT 74.99 43.965 75.2 44.035 ;
    RECT 71.21 43.245 71.42 43.315 ;
    RECT 71.21 43.605 71.42 43.675 ;
    RECT 71.21 43.965 71.42 44.035 ;
    RECT 71.67 43.245 71.88 43.315 ;
    RECT 71.67 43.605 71.88 43.675 ;
    RECT 71.67 43.965 71.88 44.035 ;
    RECT 31.37 43.245 31.58 43.315 ;
    RECT 31.37 43.605 31.58 43.675 ;
    RECT 31.37 43.965 31.58 44.035 ;
    RECT 31.83 43.245 32.04 43.315 ;
    RECT 31.83 43.605 32.04 43.675 ;
    RECT 31.83 43.965 32.04 44.035 ;
    RECT 67.89 43.245 68.1 43.315 ;
    RECT 67.89 43.605 68.1 43.675 ;
    RECT 67.89 43.965 68.1 44.035 ;
    RECT 68.35 43.245 68.56 43.315 ;
    RECT 68.35 43.605 68.56 43.675 ;
    RECT 68.35 43.965 68.56 44.035 ;
    RECT 28.05 43.245 28.26 43.315 ;
    RECT 28.05 43.605 28.26 43.675 ;
    RECT 28.05 43.965 28.26 44.035 ;
    RECT 28.51 43.245 28.72 43.315 ;
    RECT 28.51 43.605 28.72 43.675 ;
    RECT 28.51 43.965 28.72 44.035 ;
    RECT 24.73 43.245 24.94 43.315 ;
    RECT 24.73 43.605 24.94 43.675 ;
    RECT 24.73 43.965 24.94 44.035 ;
    RECT 25.19 43.245 25.4 43.315 ;
    RECT 25.19 43.605 25.4 43.675 ;
    RECT 25.19 43.965 25.4 44.035 ;
    RECT 21.41 43.245 21.62 43.315 ;
    RECT 21.41 43.605 21.62 43.675 ;
    RECT 21.41 43.965 21.62 44.035 ;
    RECT 21.87 43.245 22.08 43.315 ;
    RECT 21.87 43.605 22.08 43.675 ;
    RECT 21.87 43.965 22.08 44.035 ;
    RECT 18.09 43.245 18.3 43.315 ;
    RECT 18.09 43.605 18.3 43.675 ;
    RECT 18.09 43.965 18.3 44.035 ;
    RECT 18.55 43.245 18.76 43.315 ;
    RECT 18.55 43.605 18.76 43.675 ;
    RECT 18.55 43.965 18.76 44.035 ;
    RECT 14.77 43.245 14.98 43.315 ;
    RECT 14.77 43.605 14.98 43.675 ;
    RECT 14.77 43.965 14.98 44.035 ;
    RECT 15.23 43.245 15.44 43.315 ;
    RECT 15.23 43.605 15.44 43.675 ;
    RECT 15.23 43.965 15.44 44.035 ;
    RECT 11.45 43.245 11.66 43.315 ;
    RECT 11.45 43.605 11.66 43.675 ;
    RECT 11.45 43.965 11.66 44.035 ;
    RECT 11.91 43.245 12.12 43.315 ;
    RECT 11.91 43.605 12.12 43.675 ;
    RECT 11.91 43.965 12.12 44.035 ;
    RECT 8.13 43.245 8.34 43.315 ;
    RECT 8.13 43.605 8.34 43.675 ;
    RECT 8.13 43.965 8.34 44.035 ;
    RECT 8.59 43.245 8.8 43.315 ;
    RECT 8.59 43.605 8.8 43.675 ;
    RECT 8.59 43.965 8.8 44.035 ;
    RECT 4.81 43.245 5.02 43.315 ;
    RECT 4.81 43.605 5.02 43.675 ;
    RECT 4.81 43.965 5.02 44.035 ;
    RECT 5.27 43.245 5.48 43.315 ;
    RECT 5.27 43.605 5.48 43.675 ;
    RECT 5.27 43.965 5.48 44.035 ;
    RECT 164.17 43.245 164.38 43.315 ;
    RECT 164.17 43.605 164.38 43.675 ;
    RECT 164.17 43.965 164.38 44.035 ;
    RECT 164.63 43.245 164.84 43.315 ;
    RECT 164.63 43.605 164.84 43.675 ;
    RECT 164.63 43.965 164.84 44.035 ;
    RECT 1.49 43.245 1.7 43.315 ;
    RECT 1.49 43.605 1.7 43.675 ;
    RECT 1.49 43.965 1.7 44.035 ;
    RECT 1.95 43.245 2.16 43.315 ;
    RECT 1.95 43.605 2.16 43.675 ;
    RECT 1.95 43.965 2.16 44.035 ;
    RECT 160.85 43.245 161.06 43.315 ;
    RECT 160.85 43.605 161.06 43.675 ;
    RECT 160.85 43.965 161.06 44.035 ;
    RECT 161.31 43.245 161.52 43.315 ;
    RECT 161.31 43.605 161.52 43.675 ;
    RECT 161.31 43.965 161.52 44.035 ;
    RECT 157.53 43.245 157.74 43.315 ;
    RECT 157.53 43.605 157.74 43.675 ;
    RECT 157.53 43.965 157.74 44.035 ;
    RECT 157.99 43.245 158.2 43.315 ;
    RECT 157.99 43.605 158.2 43.675 ;
    RECT 157.99 43.965 158.2 44.035 ;
    RECT 154.21 43.245 154.42 43.315 ;
    RECT 154.21 43.605 154.42 43.675 ;
    RECT 154.21 43.965 154.42 44.035 ;
    RECT 154.67 43.245 154.88 43.315 ;
    RECT 154.67 43.605 154.88 43.675 ;
    RECT 154.67 43.965 154.88 44.035 ;
    RECT 150.89 43.245 151.1 43.315 ;
    RECT 150.89 43.605 151.1 43.675 ;
    RECT 150.89 43.965 151.1 44.035 ;
    RECT 151.35 43.245 151.56 43.315 ;
    RECT 151.35 43.605 151.56 43.675 ;
    RECT 151.35 43.965 151.56 44.035 ;
    RECT 147.57 43.245 147.78 43.315 ;
    RECT 147.57 43.605 147.78 43.675 ;
    RECT 147.57 43.965 147.78 44.035 ;
    RECT 148.03 43.245 148.24 43.315 ;
    RECT 148.03 43.605 148.24 43.675 ;
    RECT 148.03 43.965 148.24 44.035 ;
    RECT 144.25 43.245 144.46 43.315 ;
    RECT 144.25 43.605 144.46 43.675 ;
    RECT 144.25 43.965 144.46 44.035 ;
    RECT 144.71 43.245 144.92 43.315 ;
    RECT 144.71 43.605 144.92 43.675 ;
    RECT 144.71 43.965 144.92 44.035 ;
    RECT 140.93 43.245 141.14 43.315 ;
    RECT 140.93 43.605 141.14 43.675 ;
    RECT 140.93 43.965 141.14 44.035 ;
    RECT 141.39 43.245 141.6 43.315 ;
    RECT 141.39 43.605 141.6 43.675 ;
    RECT 141.39 43.965 141.6 44.035 ;
    RECT 137.61 43.245 137.82 43.315 ;
    RECT 137.61 43.605 137.82 43.675 ;
    RECT 137.61 43.965 137.82 44.035 ;
    RECT 138.07 43.245 138.28 43.315 ;
    RECT 138.07 43.605 138.28 43.675 ;
    RECT 138.07 43.965 138.28 44.035 ;
    RECT 134.29 43.245 134.5 43.315 ;
    RECT 134.29 43.605 134.5 43.675 ;
    RECT 134.29 43.965 134.5 44.035 ;
    RECT 134.75 43.245 134.96 43.315 ;
    RECT 134.75 43.605 134.96 43.675 ;
    RECT 134.75 43.965 134.96 44.035 ;
    RECT 64.57 43.245 64.78 43.315 ;
    RECT 64.57 43.605 64.78 43.675 ;
    RECT 64.57 43.965 64.78 44.035 ;
    RECT 65.03 43.245 65.24 43.315 ;
    RECT 65.03 43.605 65.24 43.675 ;
    RECT 65.03 43.965 65.24 44.035 ;
    RECT 61.25 42.525 61.46 42.595 ;
    RECT 61.25 42.885 61.46 42.955 ;
    RECT 61.25 43.245 61.46 43.315 ;
    RECT 61.71 42.525 61.92 42.595 ;
    RECT 61.71 42.885 61.92 42.955 ;
    RECT 61.71 43.245 61.92 43.315 ;
    RECT 57.93 42.525 58.14 42.595 ;
    RECT 57.93 42.885 58.14 42.955 ;
    RECT 57.93 43.245 58.14 43.315 ;
    RECT 58.39 42.525 58.6 42.595 ;
    RECT 58.39 42.885 58.6 42.955 ;
    RECT 58.39 43.245 58.6 43.315 ;
    RECT 54.61 42.525 54.82 42.595 ;
    RECT 54.61 42.885 54.82 42.955 ;
    RECT 54.61 43.245 54.82 43.315 ;
    RECT 55.07 42.525 55.28 42.595 ;
    RECT 55.07 42.885 55.28 42.955 ;
    RECT 55.07 43.245 55.28 43.315 ;
    RECT 51.29 42.525 51.5 42.595 ;
    RECT 51.29 42.885 51.5 42.955 ;
    RECT 51.29 43.245 51.5 43.315 ;
    RECT 51.75 42.525 51.96 42.595 ;
    RECT 51.75 42.885 51.96 42.955 ;
    RECT 51.75 43.245 51.96 43.315 ;
    RECT 47.97 42.525 48.18 42.595 ;
    RECT 47.97 42.885 48.18 42.955 ;
    RECT 47.97 43.245 48.18 43.315 ;
    RECT 48.43 42.525 48.64 42.595 ;
    RECT 48.43 42.885 48.64 42.955 ;
    RECT 48.43 43.245 48.64 43.315 ;
    RECT 44.65 42.525 44.86 42.595 ;
    RECT 44.65 42.885 44.86 42.955 ;
    RECT 44.65 43.245 44.86 43.315 ;
    RECT 45.11 42.525 45.32 42.595 ;
    RECT 45.11 42.885 45.32 42.955 ;
    RECT 45.11 43.245 45.32 43.315 ;
    RECT 41.33 42.525 41.54 42.595 ;
    RECT 41.33 42.885 41.54 42.955 ;
    RECT 41.33 43.245 41.54 43.315 ;
    RECT 41.79 42.525 42.0 42.595 ;
    RECT 41.79 42.885 42.0 42.955 ;
    RECT 41.79 43.245 42.0 43.315 ;
    RECT 38.01 42.525 38.22 42.595 ;
    RECT 38.01 42.885 38.22 42.955 ;
    RECT 38.01 43.245 38.22 43.315 ;
    RECT 38.47 42.525 38.68 42.595 ;
    RECT 38.47 42.885 38.68 42.955 ;
    RECT 38.47 43.245 38.68 43.315 ;
    RECT 34.69 42.525 34.9 42.595 ;
    RECT 34.69 42.885 34.9 42.955 ;
    RECT 34.69 43.245 34.9 43.315 ;
    RECT 35.15 42.525 35.36 42.595 ;
    RECT 35.15 42.885 35.36 42.955 ;
    RECT 35.15 43.245 35.36 43.315 ;
    RECT 173.945 42.885 174.015 42.955 ;
    RECT 130.97 42.525 131.18 42.595 ;
    RECT 130.97 42.885 131.18 42.955 ;
    RECT 130.97 43.245 131.18 43.315 ;
    RECT 131.43 42.525 131.64 42.595 ;
    RECT 131.43 42.885 131.64 42.955 ;
    RECT 131.43 43.245 131.64 43.315 ;
    RECT 127.65 42.525 127.86 42.595 ;
    RECT 127.65 42.885 127.86 42.955 ;
    RECT 127.65 43.245 127.86 43.315 ;
    RECT 128.11 42.525 128.32 42.595 ;
    RECT 128.11 42.885 128.32 42.955 ;
    RECT 128.11 43.245 128.32 43.315 ;
    RECT 124.33 42.525 124.54 42.595 ;
    RECT 124.33 42.885 124.54 42.955 ;
    RECT 124.33 43.245 124.54 43.315 ;
    RECT 124.79 42.525 125.0 42.595 ;
    RECT 124.79 42.885 125.0 42.955 ;
    RECT 124.79 43.245 125.0 43.315 ;
    RECT 121.01 42.525 121.22 42.595 ;
    RECT 121.01 42.885 121.22 42.955 ;
    RECT 121.01 43.245 121.22 43.315 ;
    RECT 121.47 42.525 121.68 42.595 ;
    RECT 121.47 42.885 121.68 42.955 ;
    RECT 121.47 43.245 121.68 43.315 ;
    RECT 117.69 42.525 117.9 42.595 ;
    RECT 117.69 42.885 117.9 42.955 ;
    RECT 117.69 43.245 117.9 43.315 ;
    RECT 118.15 42.525 118.36 42.595 ;
    RECT 118.15 42.885 118.36 42.955 ;
    RECT 118.15 43.245 118.36 43.315 ;
    RECT 114.37 42.525 114.58 42.595 ;
    RECT 114.37 42.885 114.58 42.955 ;
    RECT 114.37 43.245 114.58 43.315 ;
    RECT 114.83 42.525 115.04 42.595 ;
    RECT 114.83 42.885 115.04 42.955 ;
    RECT 114.83 43.245 115.04 43.315 ;
    RECT 111.05 42.525 111.26 42.595 ;
    RECT 111.05 42.885 111.26 42.955 ;
    RECT 111.05 43.245 111.26 43.315 ;
    RECT 111.51 42.525 111.72 42.595 ;
    RECT 111.51 42.885 111.72 42.955 ;
    RECT 111.51 43.245 111.72 43.315 ;
    RECT 107.73 42.525 107.94 42.595 ;
    RECT 107.73 42.885 107.94 42.955 ;
    RECT 107.73 43.245 107.94 43.315 ;
    RECT 108.19 42.525 108.4 42.595 ;
    RECT 108.19 42.885 108.4 42.955 ;
    RECT 108.19 43.245 108.4 43.315 ;
    RECT 104.41 42.525 104.62 42.595 ;
    RECT 104.41 42.885 104.62 42.955 ;
    RECT 104.41 43.245 104.62 43.315 ;
    RECT 104.87 42.525 105.08 42.595 ;
    RECT 104.87 42.885 105.08 42.955 ;
    RECT 104.87 43.245 105.08 43.315 ;
    RECT 101.09 42.525 101.3 42.595 ;
    RECT 101.09 42.885 101.3 42.955 ;
    RECT 101.09 43.245 101.3 43.315 ;
    RECT 101.55 42.525 101.76 42.595 ;
    RECT 101.55 42.885 101.76 42.955 ;
    RECT 101.55 43.245 101.76 43.315 ;
    RECT 0.4 42.885 0.47 42.955 ;
    RECT 170.81 42.525 171.02 42.595 ;
    RECT 170.81 42.885 171.02 42.955 ;
    RECT 170.81 43.245 171.02 43.315 ;
    RECT 171.27 42.525 171.48 42.595 ;
    RECT 171.27 42.885 171.48 42.955 ;
    RECT 171.27 43.245 171.48 43.315 ;
    RECT 167.49 42.525 167.7 42.595 ;
    RECT 167.49 42.885 167.7 42.955 ;
    RECT 167.49 43.245 167.7 43.315 ;
    RECT 167.95 42.525 168.16 42.595 ;
    RECT 167.95 42.885 168.16 42.955 ;
    RECT 167.95 43.245 168.16 43.315 ;
    RECT 97.77 42.525 97.98 42.595 ;
    RECT 97.77 42.885 97.98 42.955 ;
    RECT 97.77 43.245 97.98 43.315 ;
    RECT 98.23 42.525 98.44 42.595 ;
    RECT 98.23 42.885 98.44 42.955 ;
    RECT 98.23 43.245 98.44 43.315 ;
    RECT 94.45 42.525 94.66 42.595 ;
    RECT 94.45 42.885 94.66 42.955 ;
    RECT 94.45 43.245 94.66 43.315 ;
    RECT 94.91 42.525 95.12 42.595 ;
    RECT 94.91 42.885 95.12 42.955 ;
    RECT 94.91 43.245 95.12 43.315 ;
    RECT 91.13 42.525 91.34 42.595 ;
    RECT 91.13 42.885 91.34 42.955 ;
    RECT 91.13 43.245 91.34 43.315 ;
    RECT 91.59 42.525 91.8 42.595 ;
    RECT 91.59 42.885 91.8 42.955 ;
    RECT 91.59 43.245 91.8 43.315 ;
    RECT 87.81 42.525 88.02 42.595 ;
    RECT 87.81 42.885 88.02 42.955 ;
    RECT 87.81 43.245 88.02 43.315 ;
    RECT 88.27 42.525 88.48 42.595 ;
    RECT 88.27 42.885 88.48 42.955 ;
    RECT 88.27 43.245 88.48 43.315 ;
    RECT 84.49 42.525 84.7 42.595 ;
    RECT 84.49 42.885 84.7 42.955 ;
    RECT 84.49 43.245 84.7 43.315 ;
    RECT 84.95 42.525 85.16 42.595 ;
    RECT 84.95 42.885 85.16 42.955 ;
    RECT 84.95 43.245 85.16 43.315 ;
    RECT 81.17 42.525 81.38 42.595 ;
    RECT 81.17 42.885 81.38 42.955 ;
    RECT 81.17 43.245 81.38 43.315 ;
    RECT 81.63 42.525 81.84 42.595 ;
    RECT 81.63 42.885 81.84 42.955 ;
    RECT 81.63 43.245 81.84 43.315 ;
    RECT 77.85 42.525 78.06 42.595 ;
    RECT 77.85 42.885 78.06 42.955 ;
    RECT 77.85 43.245 78.06 43.315 ;
    RECT 78.31 42.525 78.52 42.595 ;
    RECT 78.31 42.885 78.52 42.955 ;
    RECT 78.31 43.245 78.52 43.315 ;
    RECT 74.53 42.525 74.74 42.595 ;
    RECT 74.53 42.885 74.74 42.955 ;
    RECT 74.53 43.245 74.74 43.315 ;
    RECT 74.99 42.525 75.2 42.595 ;
    RECT 74.99 42.885 75.2 42.955 ;
    RECT 74.99 43.245 75.2 43.315 ;
    RECT 71.21 42.525 71.42 42.595 ;
    RECT 71.21 42.885 71.42 42.955 ;
    RECT 71.21 43.245 71.42 43.315 ;
    RECT 71.67 42.525 71.88 42.595 ;
    RECT 71.67 42.885 71.88 42.955 ;
    RECT 71.67 43.245 71.88 43.315 ;
    RECT 31.37 42.525 31.58 42.595 ;
    RECT 31.37 42.885 31.58 42.955 ;
    RECT 31.37 43.245 31.58 43.315 ;
    RECT 31.83 42.525 32.04 42.595 ;
    RECT 31.83 42.885 32.04 42.955 ;
    RECT 31.83 43.245 32.04 43.315 ;
    RECT 67.89 42.525 68.1 42.595 ;
    RECT 67.89 42.885 68.1 42.955 ;
    RECT 67.89 43.245 68.1 43.315 ;
    RECT 68.35 42.525 68.56 42.595 ;
    RECT 68.35 42.885 68.56 42.955 ;
    RECT 68.35 43.245 68.56 43.315 ;
    RECT 28.05 42.525 28.26 42.595 ;
    RECT 28.05 42.885 28.26 42.955 ;
    RECT 28.05 43.245 28.26 43.315 ;
    RECT 28.51 42.525 28.72 42.595 ;
    RECT 28.51 42.885 28.72 42.955 ;
    RECT 28.51 43.245 28.72 43.315 ;
    RECT 24.73 42.525 24.94 42.595 ;
    RECT 24.73 42.885 24.94 42.955 ;
    RECT 24.73 43.245 24.94 43.315 ;
    RECT 25.19 42.525 25.4 42.595 ;
    RECT 25.19 42.885 25.4 42.955 ;
    RECT 25.19 43.245 25.4 43.315 ;
    RECT 21.41 42.525 21.62 42.595 ;
    RECT 21.41 42.885 21.62 42.955 ;
    RECT 21.41 43.245 21.62 43.315 ;
    RECT 21.87 42.525 22.08 42.595 ;
    RECT 21.87 42.885 22.08 42.955 ;
    RECT 21.87 43.245 22.08 43.315 ;
    RECT 18.09 42.525 18.3 42.595 ;
    RECT 18.09 42.885 18.3 42.955 ;
    RECT 18.09 43.245 18.3 43.315 ;
    RECT 18.55 42.525 18.76 42.595 ;
    RECT 18.55 42.885 18.76 42.955 ;
    RECT 18.55 43.245 18.76 43.315 ;
    RECT 14.77 42.525 14.98 42.595 ;
    RECT 14.77 42.885 14.98 42.955 ;
    RECT 14.77 43.245 14.98 43.315 ;
    RECT 15.23 42.525 15.44 42.595 ;
    RECT 15.23 42.885 15.44 42.955 ;
    RECT 15.23 43.245 15.44 43.315 ;
    RECT 11.45 42.525 11.66 42.595 ;
    RECT 11.45 42.885 11.66 42.955 ;
    RECT 11.45 43.245 11.66 43.315 ;
    RECT 11.91 42.525 12.12 42.595 ;
    RECT 11.91 42.885 12.12 42.955 ;
    RECT 11.91 43.245 12.12 43.315 ;
    RECT 8.13 42.525 8.34 42.595 ;
    RECT 8.13 42.885 8.34 42.955 ;
    RECT 8.13 43.245 8.34 43.315 ;
    RECT 8.59 42.525 8.8 42.595 ;
    RECT 8.59 42.885 8.8 42.955 ;
    RECT 8.59 43.245 8.8 43.315 ;
    RECT 4.81 42.525 5.02 42.595 ;
    RECT 4.81 42.885 5.02 42.955 ;
    RECT 4.81 43.245 5.02 43.315 ;
    RECT 5.27 42.525 5.48 42.595 ;
    RECT 5.27 42.885 5.48 42.955 ;
    RECT 5.27 43.245 5.48 43.315 ;
    RECT 164.17 42.525 164.38 42.595 ;
    RECT 164.17 42.885 164.38 42.955 ;
    RECT 164.17 43.245 164.38 43.315 ;
    RECT 164.63 42.525 164.84 42.595 ;
    RECT 164.63 42.885 164.84 42.955 ;
    RECT 164.63 43.245 164.84 43.315 ;
    RECT 1.49 42.525 1.7 42.595 ;
    RECT 1.49 42.885 1.7 42.955 ;
    RECT 1.49 43.245 1.7 43.315 ;
    RECT 1.95 42.525 2.16 42.595 ;
    RECT 1.95 42.885 2.16 42.955 ;
    RECT 1.95 43.245 2.16 43.315 ;
    RECT 160.85 42.525 161.06 42.595 ;
    RECT 160.85 42.885 161.06 42.955 ;
    RECT 160.85 43.245 161.06 43.315 ;
    RECT 161.31 42.525 161.52 42.595 ;
    RECT 161.31 42.885 161.52 42.955 ;
    RECT 161.31 43.245 161.52 43.315 ;
    RECT 157.53 42.525 157.74 42.595 ;
    RECT 157.53 42.885 157.74 42.955 ;
    RECT 157.53 43.245 157.74 43.315 ;
    RECT 157.99 42.525 158.2 42.595 ;
    RECT 157.99 42.885 158.2 42.955 ;
    RECT 157.99 43.245 158.2 43.315 ;
    RECT 154.21 42.525 154.42 42.595 ;
    RECT 154.21 42.885 154.42 42.955 ;
    RECT 154.21 43.245 154.42 43.315 ;
    RECT 154.67 42.525 154.88 42.595 ;
    RECT 154.67 42.885 154.88 42.955 ;
    RECT 154.67 43.245 154.88 43.315 ;
    RECT 150.89 42.525 151.1 42.595 ;
    RECT 150.89 42.885 151.1 42.955 ;
    RECT 150.89 43.245 151.1 43.315 ;
    RECT 151.35 42.525 151.56 42.595 ;
    RECT 151.35 42.885 151.56 42.955 ;
    RECT 151.35 43.245 151.56 43.315 ;
    RECT 147.57 42.525 147.78 42.595 ;
    RECT 147.57 42.885 147.78 42.955 ;
    RECT 147.57 43.245 147.78 43.315 ;
    RECT 148.03 42.525 148.24 42.595 ;
    RECT 148.03 42.885 148.24 42.955 ;
    RECT 148.03 43.245 148.24 43.315 ;
    RECT 144.25 42.525 144.46 42.595 ;
    RECT 144.25 42.885 144.46 42.955 ;
    RECT 144.25 43.245 144.46 43.315 ;
    RECT 144.71 42.525 144.92 42.595 ;
    RECT 144.71 42.885 144.92 42.955 ;
    RECT 144.71 43.245 144.92 43.315 ;
    RECT 140.93 42.525 141.14 42.595 ;
    RECT 140.93 42.885 141.14 42.955 ;
    RECT 140.93 43.245 141.14 43.315 ;
    RECT 141.39 42.525 141.6 42.595 ;
    RECT 141.39 42.885 141.6 42.955 ;
    RECT 141.39 43.245 141.6 43.315 ;
    RECT 137.61 42.525 137.82 42.595 ;
    RECT 137.61 42.885 137.82 42.955 ;
    RECT 137.61 43.245 137.82 43.315 ;
    RECT 138.07 42.525 138.28 42.595 ;
    RECT 138.07 42.885 138.28 42.955 ;
    RECT 138.07 43.245 138.28 43.315 ;
    RECT 134.29 42.525 134.5 42.595 ;
    RECT 134.29 42.885 134.5 42.955 ;
    RECT 134.29 43.245 134.5 43.315 ;
    RECT 134.75 42.525 134.96 42.595 ;
    RECT 134.75 42.885 134.96 42.955 ;
    RECT 134.75 43.245 134.96 43.315 ;
    RECT 64.57 42.525 64.78 42.595 ;
    RECT 64.57 42.885 64.78 42.955 ;
    RECT 64.57 43.245 64.78 43.315 ;
    RECT 65.03 42.525 65.24 42.595 ;
    RECT 65.03 42.885 65.24 42.955 ;
    RECT 65.03 43.245 65.24 43.315 ;
    RECT 61.25 41.805 61.46 41.875 ;
    RECT 61.25 42.165 61.46 42.235 ;
    RECT 61.25 42.525 61.46 42.595 ;
    RECT 61.71 41.805 61.92 41.875 ;
    RECT 61.71 42.165 61.92 42.235 ;
    RECT 61.71 42.525 61.92 42.595 ;
    RECT 57.93 41.805 58.14 41.875 ;
    RECT 57.93 42.165 58.14 42.235 ;
    RECT 57.93 42.525 58.14 42.595 ;
    RECT 58.39 41.805 58.6 41.875 ;
    RECT 58.39 42.165 58.6 42.235 ;
    RECT 58.39 42.525 58.6 42.595 ;
    RECT 54.61 41.805 54.82 41.875 ;
    RECT 54.61 42.165 54.82 42.235 ;
    RECT 54.61 42.525 54.82 42.595 ;
    RECT 55.07 41.805 55.28 41.875 ;
    RECT 55.07 42.165 55.28 42.235 ;
    RECT 55.07 42.525 55.28 42.595 ;
    RECT 51.29 41.805 51.5 41.875 ;
    RECT 51.29 42.165 51.5 42.235 ;
    RECT 51.29 42.525 51.5 42.595 ;
    RECT 51.75 41.805 51.96 41.875 ;
    RECT 51.75 42.165 51.96 42.235 ;
    RECT 51.75 42.525 51.96 42.595 ;
    RECT 47.97 41.805 48.18 41.875 ;
    RECT 47.97 42.165 48.18 42.235 ;
    RECT 47.97 42.525 48.18 42.595 ;
    RECT 48.43 41.805 48.64 41.875 ;
    RECT 48.43 42.165 48.64 42.235 ;
    RECT 48.43 42.525 48.64 42.595 ;
    RECT 44.65 41.805 44.86 41.875 ;
    RECT 44.65 42.165 44.86 42.235 ;
    RECT 44.65 42.525 44.86 42.595 ;
    RECT 45.11 41.805 45.32 41.875 ;
    RECT 45.11 42.165 45.32 42.235 ;
    RECT 45.11 42.525 45.32 42.595 ;
    RECT 41.33 41.805 41.54 41.875 ;
    RECT 41.33 42.165 41.54 42.235 ;
    RECT 41.33 42.525 41.54 42.595 ;
    RECT 41.79 41.805 42.0 41.875 ;
    RECT 41.79 42.165 42.0 42.235 ;
    RECT 41.79 42.525 42.0 42.595 ;
    RECT 38.01 41.805 38.22 41.875 ;
    RECT 38.01 42.165 38.22 42.235 ;
    RECT 38.01 42.525 38.22 42.595 ;
    RECT 38.47 41.805 38.68 41.875 ;
    RECT 38.47 42.165 38.68 42.235 ;
    RECT 38.47 42.525 38.68 42.595 ;
    RECT 34.69 41.805 34.9 41.875 ;
    RECT 34.69 42.165 34.9 42.235 ;
    RECT 34.69 42.525 34.9 42.595 ;
    RECT 35.15 41.805 35.36 41.875 ;
    RECT 35.15 42.165 35.36 42.235 ;
    RECT 35.15 42.525 35.36 42.595 ;
    RECT 173.945 42.165 174.015 42.235 ;
    RECT 130.97 41.805 131.18 41.875 ;
    RECT 130.97 42.165 131.18 42.235 ;
    RECT 130.97 42.525 131.18 42.595 ;
    RECT 131.43 41.805 131.64 41.875 ;
    RECT 131.43 42.165 131.64 42.235 ;
    RECT 131.43 42.525 131.64 42.595 ;
    RECT 127.65 41.805 127.86 41.875 ;
    RECT 127.65 42.165 127.86 42.235 ;
    RECT 127.65 42.525 127.86 42.595 ;
    RECT 128.11 41.805 128.32 41.875 ;
    RECT 128.11 42.165 128.32 42.235 ;
    RECT 128.11 42.525 128.32 42.595 ;
    RECT 124.33 41.805 124.54 41.875 ;
    RECT 124.33 42.165 124.54 42.235 ;
    RECT 124.33 42.525 124.54 42.595 ;
    RECT 124.79 41.805 125.0 41.875 ;
    RECT 124.79 42.165 125.0 42.235 ;
    RECT 124.79 42.525 125.0 42.595 ;
    RECT 121.01 41.805 121.22 41.875 ;
    RECT 121.01 42.165 121.22 42.235 ;
    RECT 121.01 42.525 121.22 42.595 ;
    RECT 121.47 41.805 121.68 41.875 ;
    RECT 121.47 42.165 121.68 42.235 ;
    RECT 121.47 42.525 121.68 42.595 ;
    RECT 117.69 41.805 117.9 41.875 ;
    RECT 117.69 42.165 117.9 42.235 ;
    RECT 117.69 42.525 117.9 42.595 ;
    RECT 118.15 41.805 118.36 41.875 ;
    RECT 118.15 42.165 118.36 42.235 ;
    RECT 118.15 42.525 118.36 42.595 ;
    RECT 114.37 41.805 114.58 41.875 ;
    RECT 114.37 42.165 114.58 42.235 ;
    RECT 114.37 42.525 114.58 42.595 ;
    RECT 114.83 41.805 115.04 41.875 ;
    RECT 114.83 42.165 115.04 42.235 ;
    RECT 114.83 42.525 115.04 42.595 ;
    RECT 111.05 41.805 111.26 41.875 ;
    RECT 111.05 42.165 111.26 42.235 ;
    RECT 111.05 42.525 111.26 42.595 ;
    RECT 111.51 41.805 111.72 41.875 ;
    RECT 111.51 42.165 111.72 42.235 ;
    RECT 111.51 42.525 111.72 42.595 ;
    RECT 107.73 41.805 107.94 41.875 ;
    RECT 107.73 42.165 107.94 42.235 ;
    RECT 107.73 42.525 107.94 42.595 ;
    RECT 108.19 41.805 108.4 41.875 ;
    RECT 108.19 42.165 108.4 42.235 ;
    RECT 108.19 42.525 108.4 42.595 ;
    RECT 104.41 41.805 104.62 41.875 ;
    RECT 104.41 42.165 104.62 42.235 ;
    RECT 104.41 42.525 104.62 42.595 ;
    RECT 104.87 41.805 105.08 41.875 ;
    RECT 104.87 42.165 105.08 42.235 ;
    RECT 104.87 42.525 105.08 42.595 ;
    RECT 101.09 41.805 101.3 41.875 ;
    RECT 101.09 42.165 101.3 42.235 ;
    RECT 101.09 42.525 101.3 42.595 ;
    RECT 101.55 41.805 101.76 41.875 ;
    RECT 101.55 42.165 101.76 42.235 ;
    RECT 101.55 42.525 101.76 42.595 ;
    RECT 0.4 42.165 0.47 42.235 ;
    RECT 170.81 41.805 171.02 41.875 ;
    RECT 170.81 42.165 171.02 42.235 ;
    RECT 170.81 42.525 171.02 42.595 ;
    RECT 171.27 41.805 171.48 41.875 ;
    RECT 171.27 42.165 171.48 42.235 ;
    RECT 171.27 42.525 171.48 42.595 ;
    RECT 167.49 41.805 167.7 41.875 ;
    RECT 167.49 42.165 167.7 42.235 ;
    RECT 167.49 42.525 167.7 42.595 ;
    RECT 167.95 41.805 168.16 41.875 ;
    RECT 167.95 42.165 168.16 42.235 ;
    RECT 167.95 42.525 168.16 42.595 ;
    RECT 97.77 41.805 97.98 41.875 ;
    RECT 97.77 42.165 97.98 42.235 ;
    RECT 97.77 42.525 97.98 42.595 ;
    RECT 98.23 41.805 98.44 41.875 ;
    RECT 98.23 42.165 98.44 42.235 ;
    RECT 98.23 42.525 98.44 42.595 ;
    RECT 94.45 41.805 94.66 41.875 ;
    RECT 94.45 42.165 94.66 42.235 ;
    RECT 94.45 42.525 94.66 42.595 ;
    RECT 94.91 41.805 95.12 41.875 ;
    RECT 94.91 42.165 95.12 42.235 ;
    RECT 94.91 42.525 95.12 42.595 ;
    RECT 91.13 41.805 91.34 41.875 ;
    RECT 91.13 42.165 91.34 42.235 ;
    RECT 91.13 42.525 91.34 42.595 ;
    RECT 91.59 41.805 91.8 41.875 ;
    RECT 91.59 42.165 91.8 42.235 ;
    RECT 91.59 42.525 91.8 42.595 ;
    RECT 87.81 41.805 88.02 41.875 ;
    RECT 87.81 42.165 88.02 42.235 ;
    RECT 87.81 42.525 88.02 42.595 ;
    RECT 88.27 41.805 88.48 41.875 ;
    RECT 88.27 42.165 88.48 42.235 ;
    RECT 88.27 42.525 88.48 42.595 ;
    RECT 84.49 41.805 84.7 41.875 ;
    RECT 84.49 42.165 84.7 42.235 ;
    RECT 84.49 42.525 84.7 42.595 ;
    RECT 84.95 41.805 85.16 41.875 ;
    RECT 84.95 42.165 85.16 42.235 ;
    RECT 84.95 42.525 85.16 42.595 ;
    RECT 81.17 41.805 81.38 41.875 ;
    RECT 81.17 42.165 81.38 42.235 ;
    RECT 81.17 42.525 81.38 42.595 ;
    RECT 81.63 41.805 81.84 41.875 ;
    RECT 81.63 42.165 81.84 42.235 ;
    RECT 81.63 42.525 81.84 42.595 ;
    RECT 77.85 41.805 78.06 41.875 ;
    RECT 77.85 42.165 78.06 42.235 ;
    RECT 77.85 42.525 78.06 42.595 ;
    RECT 78.31 41.805 78.52 41.875 ;
    RECT 78.31 42.165 78.52 42.235 ;
    RECT 78.31 42.525 78.52 42.595 ;
    RECT 74.53 41.805 74.74 41.875 ;
    RECT 74.53 42.165 74.74 42.235 ;
    RECT 74.53 42.525 74.74 42.595 ;
    RECT 74.99 41.805 75.2 41.875 ;
    RECT 74.99 42.165 75.2 42.235 ;
    RECT 74.99 42.525 75.2 42.595 ;
    RECT 71.21 41.805 71.42 41.875 ;
    RECT 71.21 42.165 71.42 42.235 ;
    RECT 71.21 42.525 71.42 42.595 ;
    RECT 71.67 41.805 71.88 41.875 ;
    RECT 71.67 42.165 71.88 42.235 ;
    RECT 71.67 42.525 71.88 42.595 ;
    RECT 31.37 41.805 31.58 41.875 ;
    RECT 31.37 42.165 31.58 42.235 ;
    RECT 31.37 42.525 31.58 42.595 ;
    RECT 31.83 41.805 32.04 41.875 ;
    RECT 31.83 42.165 32.04 42.235 ;
    RECT 31.83 42.525 32.04 42.595 ;
    RECT 67.89 41.805 68.1 41.875 ;
    RECT 67.89 42.165 68.1 42.235 ;
    RECT 67.89 42.525 68.1 42.595 ;
    RECT 68.35 41.805 68.56 41.875 ;
    RECT 68.35 42.165 68.56 42.235 ;
    RECT 68.35 42.525 68.56 42.595 ;
    RECT 28.05 41.805 28.26 41.875 ;
    RECT 28.05 42.165 28.26 42.235 ;
    RECT 28.05 42.525 28.26 42.595 ;
    RECT 28.51 41.805 28.72 41.875 ;
    RECT 28.51 42.165 28.72 42.235 ;
    RECT 28.51 42.525 28.72 42.595 ;
    RECT 24.73 41.805 24.94 41.875 ;
    RECT 24.73 42.165 24.94 42.235 ;
    RECT 24.73 42.525 24.94 42.595 ;
    RECT 25.19 41.805 25.4 41.875 ;
    RECT 25.19 42.165 25.4 42.235 ;
    RECT 25.19 42.525 25.4 42.595 ;
    RECT 21.41 41.805 21.62 41.875 ;
    RECT 21.41 42.165 21.62 42.235 ;
    RECT 21.41 42.525 21.62 42.595 ;
    RECT 21.87 41.805 22.08 41.875 ;
    RECT 21.87 42.165 22.08 42.235 ;
    RECT 21.87 42.525 22.08 42.595 ;
    RECT 18.09 41.805 18.3 41.875 ;
    RECT 18.09 42.165 18.3 42.235 ;
    RECT 18.09 42.525 18.3 42.595 ;
    RECT 18.55 41.805 18.76 41.875 ;
    RECT 18.55 42.165 18.76 42.235 ;
    RECT 18.55 42.525 18.76 42.595 ;
    RECT 14.77 41.805 14.98 41.875 ;
    RECT 14.77 42.165 14.98 42.235 ;
    RECT 14.77 42.525 14.98 42.595 ;
    RECT 15.23 41.805 15.44 41.875 ;
    RECT 15.23 42.165 15.44 42.235 ;
    RECT 15.23 42.525 15.44 42.595 ;
    RECT 11.45 41.805 11.66 41.875 ;
    RECT 11.45 42.165 11.66 42.235 ;
    RECT 11.45 42.525 11.66 42.595 ;
    RECT 11.91 41.805 12.12 41.875 ;
    RECT 11.91 42.165 12.12 42.235 ;
    RECT 11.91 42.525 12.12 42.595 ;
    RECT 8.13 41.805 8.34 41.875 ;
    RECT 8.13 42.165 8.34 42.235 ;
    RECT 8.13 42.525 8.34 42.595 ;
    RECT 8.59 41.805 8.8 41.875 ;
    RECT 8.59 42.165 8.8 42.235 ;
    RECT 8.59 42.525 8.8 42.595 ;
    RECT 4.81 41.805 5.02 41.875 ;
    RECT 4.81 42.165 5.02 42.235 ;
    RECT 4.81 42.525 5.02 42.595 ;
    RECT 5.27 41.805 5.48 41.875 ;
    RECT 5.27 42.165 5.48 42.235 ;
    RECT 5.27 42.525 5.48 42.595 ;
    RECT 164.17 41.805 164.38 41.875 ;
    RECT 164.17 42.165 164.38 42.235 ;
    RECT 164.17 42.525 164.38 42.595 ;
    RECT 164.63 41.805 164.84 41.875 ;
    RECT 164.63 42.165 164.84 42.235 ;
    RECT 164.63 42.525 164.84 42.595 ;
    RECT 1.49 41.805 1.7 41.875 ;
    RECT 1.49 42.165 1.7 42.235 ;
    RECT 1.49 42.525 1.7 42.595 ;
    RECT 1.95 41.805 2.16 41.875 ;
    RECT 1.95 42.165 2.16 42.235 ;
    RECT 1.95 42.525 2.16 42.595 ;
    RECT 160.85 41.805 161.06 41.875 ;
    RECT 160.85 42.165 161.06 42.235 ;
    RECT 160.85 42.525 161.06 42.595 ;
    RECT 161.31 41.805 161.52 41.875 ;
    RECT 161.31 42.165 161.52 42.235 ;
    RECT 161.31 42.525 161.52 42.595 ;
    RECT 157.53 41.805 157.74 41.875 ;
    RECT 157.53 42.165 157.74 42.235 ;
    RECT 157.53 42.525 157.74 42.595 ;
    RECT 157.99 41.805 158.2 41.875 ;
    RECT 157.99 42.165 158.2 42.235 ;
    RECT 157.99 42.525 158.2 42.595 ;
    RECT 154.21 41.805 154.42 41.875 ;
    RECT 154.21 42.165 154.42 42.235 ;
    RECT 154.21 42.525 154.42 42.595 ;
    RECT 154.67 41.805 154.88 41.875 ;
    RECT 154.67 42.165 154.88 42.235 ;
    RECT 154.67 42.525 154.88 42.595 ;
    RECT 150.89 41.805 151.1 41.875 ;
    RECT 150.89 42.165 151.1 42.235 ;
    RECT 150.89 42.525 151.1 42.595 ;
    RECT 151.35 41.805 151.56 41.875 ;
    RECT 151.35 42.165 151.56 42.235 ;
    RECT 151.35 42.525 151.56 42.595 ;
    RECT 147.57 41.805 147.78 41.875 ;
    RECT 147.57 42.165 147.78 42.235 ;
    RECT 147.57 42.525 147.78 42.595 ;
    RECT 148.03 41.805 148.24 41.875 ;
    RECT 148.03 42.165 148.24 42.235 ;
    RECT 148.03 42.525 148.24 42.595 ;
    RECT 144.25 41.805 144.46 41.875 ;
    RECT 144.25 42.165 144.46 42.235 ;
    RECT 144.25 42.525 144.46 42.595 ;
    RECT 144.71 41.805 144.92 41.875 ;
    RECT 144.71 42.165 144.92 42.235 ;
    RECT 144.71 42.525 144.92 42.595 ;
    RECT 140.93 41.805 141.14 41.875 ;
    RECT 140.93 42.165 141.14 42.235 ;
    RECT 140.93 42.525 141.14 42.595 ;
    RECT 141.39 41.805 141.6 41.875 ;
    RECT 141.39 42.165 141.6 42.235 ;
    RECT 141.39 42.525 141.6 42.595 ;
    RECT 137.61 41.805 137.82 41.875 ;
    RECT 137.61 42.165 137.82 42.235 ;
    RECT 137.61 42.525 137.82 42.595 ;
    RECT 138.07 41.805 138.28 41.875 ;
    RECT 138.07 42.165 138.28 42.235 ;
    RECT 138.07 42.525 138.28 42.595 ;
    RECT 134.29 41.805 134.5 41.875 ;
    RECT 134.29 42.165 134.5 42.235 ;
    RECT 134.29 42.525 134.5 42.595 ;
    RECT 134.75 41.805 134.96 41.875 ;
    RECT 134.75 42.165 134.96 42.235 ;
    RECT 134.75 42.525 134.96 42.595 ;
    RECT 64.57 41.805 64.78 41.875 ;
    RECT 64.57 42.165 64.78 42.235 ;
    RECT 64.57 42.525 64.78 42.595 ;
    RECT 65.03 41.805 65.24 41.875 ;
    RECT 65.03 42.165 65.24 42.235 ;
    RECT 65.03 42.525 65.24 42.595 ;
    RECT 61.25 41.085 61.46 41.155 ;
    RECT 61.25 41.445 61.46 41.515 ;
    RECT 61.25 41.805 61.46 41.875 ;
    RECT 61.71 41.085 61.92 41.155 ;
    RECT 61.71 41.445 61.92 41.515 ;
    RECT 61.71 41.805 61.92 41.875 ;
    RECT 57.93 41.085 58.14 41.155 ;
    RECT 57.93 41.445 58.14 41.515 ;
    RECT 57.93 41.805 58.14 41.875 ;
    RECT 58.39 41.085 58.6 41.155 ;
    RECT 58.39 41.445 58.6 41.515 ;
    RECT 58.39 41.805 58.6 41.875 ;
    RECT 54.61 41.085 54.82 41.155 ;
    RECT 54.61 41.445 54.82 41.515 ;
    RECT 54.61 41.805 54.82 41.875 ;
    RECT 55.07 41.085 55.28 41.155 ;
    RECT 55.07 41.445 55.28 41.515 ;
    RECT 55.07 41.805 55.28 41.875 ;
    RECT 51.29 41.085 51.5 41.155 ;
    RECT 51.29 41.445 51.5 41.515 ;
    RECT 51.29 41.805 51.5 41.875 ;
    RECT 51.75 41.085 51.96 41.155 ;
    RECT 51.75 41.445 51.96 41.515 ;
    RECT 51.75 41.805 51.96 41.875 ;
    RECT 47.97 41.085 48.18 41.155 ;
    RECT 47.97 41.445 48.18 41.515 ;
    RECT 47.97 41.805 48.18 41.875 ;
    RECT 48.43 41.085 48.64 41.155 ;
    RECT 48.43 41.445 48.64 41.515 ;
    RECT 48.43 41.805 48.64 41.875 ;
    RECT 44.65 41.085 44.86 41.155 ;
    RECT 44.65 41.445 44.86 41.515 ;
    RECT 44.65 41.805 44.86 41.875 ;
    RECT 45.11 41.085 45.32 41.155 ;
    RECT 45.11 41.445 45.32 41.515 ;
    RECT 45.11 41.805 45.32 41.875 ;
    RECT 41.33 41.085 41.54 41.155 ;
    RECT 41.33 41.445 41.54 41.515 ;
    RECT 41.33 41.805 41.54 41.875 ;
    RECT 41.79 41.085 42.0 41.155 ;
    RECT 41.79 41.445 42.0 41.515 ;
    RECT 41.79 41.805 42.0 41.875 ;
    RECT 38.01 41.085 38.22 41.155 ;
    RECT 38.01 41.445 38.22 41.515 ;
    RECT 38.01 41.805 38.22 41.875 ;
    RECT 38.47 41.085 38.68 41.155 ;
    RECT 38.47 41.445 38.68 41.515 ;
    RECT 38.47 41.805 38.68 41.875 ;
    RECT 34.69 41.085 34.9 41.155 ;
    RECT 34.69 41.445 34.9 41.515 ;
    RECT 34.69 41.805 34.9 41.875 ;
    RECT 35.15 41.085 35.36 41.155 ;
    RECT 35.15 41.445 35.36 41.515 ;
    RECT 35.15 41.805 35.36 41.875 ;
    RECT 173.945 41.445 174.015 41.515 ;
    RECT 130.97 41.085 131.18 41.155 ;
    RECT 130.97 41.445 131.18 41.515 ;
    RECT 130.97 41.805 131.18 41.875 ;
    RECT 131.43 41.085 131.64 41.155 ;
    RECT 131.43 41.445 131.64 41.515 ;
    RECT 131.43 41.805 131.64 41.875 ;
    RECT 127.65 41.085 127.86 41.155 ;
    RECT 127.65 41.445 127.86 41.515 ;
    RECT 127.65 41.805 127.86 41.875 ;
    RECT 128.11 41.085 128.32 41.155 ;
    RECT 128.11 41.445 128.32 41.515 ;
    RECT 128.11 41.805 128.32 41.875 ;
    RECT 124.33 41.085 124.54 41.155 ;
    RECT 124.33 41.445 124.54 41.515 ;
    RECT 124.33 41.805 124.54 41.875 ;
    RECT 124.79 41.085 125.0 41.155 ;
    RECT 124.79 41.445 125.0 41.515 ;
    RECT 124.79 41.805 125.0 41.875 ;
    RECT 121.01 41.085 121.22 41.155 ;
    RECT 121.01 41.445 121.22 41.515 ;
    RECT 121.01 41.805 121.22 41.875 ;
    RECT 121.47 41.085 121.68 41.155 ;
    RECT 121.47 41.445 121.68 41.515 ;
    RECT 121.47 41.805 121.68 41.875 ;
    RECT 117.69 41.085 117.9 41.155 ;
    RECT 117.69 41.445 117.9 41.515 ;
    RECT 117.69 41.805 117.9 41.875 ;
    RECT 118.15 41.085 118.36 41.155 ;
    RECT 118.15 41.445 118.36 41.515 ;
    RECT 118.15 41.805 118.36 41.875 ;
    RECT 114.37 41.085 114.58 41.155 ;
    RECT 114.37 41.445 114.58 41.515 ;
    RECT 114.37 41.805 114.58 41.875 ;
    RECT 114.83 41.085 115.04 41.155 ;
    RECT 114.83 41.445 115.04 41.515 ;
    RECT 114.83 41.805 115.04 41.875 ;
    RECT 111.05 41.085 111.26 41.155 ;
    RECT 111.05 41.445 111.26 41.515 ;
    RECT 111.05 41.805 111.26 41.875 ;
    RECT 111.51 41.085 111.72 41.155 ;
    RECT 111.51 41.445 111.72 41.515 ;
    RECT 111.51 41.805 111.72 41.875 ;
    RECT 107.73 41.085 107.94 41.155 ;
    RECT 107.73 41.445 107.94 41.515 ;
    RECT 107.73 41.805 107.94 41.875 ;
    RECT 108.19 41.085 108.4 41.155 ;
    RECT 108.19 41.445 108.4 41.515 ;
    RECT 108.19 41.805 108.4 41.875 ;
    RECT 104.41 41.085 104.62 41.155 ;
    RECT 104.41 41.445 104.62 41.515 ;
    RECT 104.41 41.805 104.62 41.875 ;
    RECT 104.87 41.085 105.08 41.155 ;
    RECT 104.87 41.445 105.08 41.515 ;
    RECT 104.87 41.805 105.08 41.875 ;
    RECT 101.09 41.085 101.3 41.155 ;
    RECT 101.09 41.445 101.3 41.515 ;
    RECT 101.09 41.805 101.3 41.875 ;
    RECT 101.55 41.085 101.76 41.155 ;
    RECT 101.55 41.445 101.76 41.515 ;
    RECT 101.55 41.805 101.76 41.875 ;
    RECT 0.4 41.445 0.47 41.515 ;
    RECT 170.81 41.085 171.02 41.155 ;
    RECT 170.81 41.445 171.02 41.515 ;
    RECT 170.81 41.805 171.02 41.875 ;
    RECT 171.27 41.085 171.48 41.155 ;
    RECT 171.27 41.445 171.48 41.515 ;
    RECT 171.27 41.805 171.48 41.875 ;
    RECT 167.49 41.085 167.7 41.155 ;
    RECT 167.49 41.445 167.7 41.515 ;
    RECT 167.49 41.805 167.7 41.875 ;
    RECT 167.95 41.085 168.16 41.155 ;
    RECT 167.95 41.445 168.16 41.515 ;
    RECT 167.95 41.805 168.16 41.875 ;
    RECT 97.77 41.085 97.98 41.155 ;
    RECT 97.77 41.445 97.98 41.515 ;
    RECT 97.77 41.805 97.98 41.875 ;
    RECT 98.23 41.085 98.44 41.155 ;
    RECT 98.23 41.445 98.44 41.515 ;
    RECT 98.23 41.805 98.44 41.875 ;
    RECT 94.45 41.085 94.66 41.155 ;
    RECT 94.45 41.445 94.66 41.515 ;
    RECT 94.45 41.805 94.66 41.875 ;
    RECT 94.91 41.085 95.12 41.155 ;
    RECT 94.91 41.445 95.12 41.515 ;
    RECT 94.91 41.805 95.12 41.875 ;
    RECT 91.13 41.085 91.34 41.155 ;
    RECT 91.13 41.445 91.34 41.515 ;
    RECT 91.13 41.805 91.34 41.875 ;
    RECT 91.59 41.085 91.8 41.155 ;
    RECT 91.59 41.445 91.8 41.515 ;
    RECT 91.59 41.805 91.8 41.875 ;
    RECT 87.81 41.085 88.02 41.155 ;
    RECT 87.81 41.445 88.02 41.515 ;
    RECT 87.81 41.805 88.02 41.875 ;
    RECT 88.27 41.085 88.48 41.155 ;
    RECT 88.27 41.445 88.48 41.515 ;
    RECT 88.27 41.805 88.48 41.875 ;
    RECT 84.49 41.085 84.7 41.155 ;
    RECT 84.49 41.445 84.7 41.515 ;
    RECT 84.49 41.805 84.7 41.875 ;
    RECT 84.95 41.085 85.16 41.155 ;
    RECT 84.95 41.445 85.16 41.515 ;
    RECT 84.95 41.805 85.16 41.875 ;
    RECT 81.17 41.085 81.38 41.155 ;
    RECT 81.17 41.445 81.38 41.515 ;
    RECT 81.17 41.805 81.38 41.875 ;
    RECT 81.63 41.085 81.84 41.155 ;
    RECT 81.63 41.445 81.84 41.515 ;
    RECT 81.63 41.805 81.84 41.875 ;
    RECT 77.85 41.085 78.06 41.155 ;
    RECT 77.85 41.445 78.06 41.515 ;
    RECT 77.85 41.805 78.06 41.875 ;
    RECT 78.31 41.085 78.52 41.155 ;
    RECT 78.31 41.445 78.52 41.515 ;
    RECT 78.31 41.805 78.52 41.875 ;
    RECT 74.53 41.085 74.74 41.155 ;
    RECT 74.53 41.445 74.74 41.515 ;
    RECT 74.53 41.805 74.74 41.875 ;
    RECT 74.99 41.085 75.2 41.155 ;
    RECT 74.99 41.445 75.2 41.515 ;
    RECT 74.99 41.805 75.2 41.875 ;
    RECT 71.21 41.085 71.42 41.155 ;
    RECT 71.21 41.445 71.42 41.515 ;
    RECT 71.21 41.805 71.42 41.875 ;
    RECT 71.67 41.085 71.88 41.155 ;
    RECT 71.67 41.445 71.88 41.515 ;
    RECT 71.67 41.805 71.88 41.875 ;
    RECT 31.37 41.085 31.58 41.155 ;
    RECT 31.37 41.445 31.58 41.515 ;
    RECT 31.37 41.805 31.58 41.875 ;
    RECT 31.83 41.085 32.04 41.155 ;
    RECT 31.83 41.445 32.04 41.515 ;
    RECT 31.83 41.805 32.04 41.875 ;
    RECT 67.89 41.085 68.1 41.155 ;
    RECT 67.89 41.445 68.1 41.515 ;
    RECT 67.89 41.805 68.1 41.875 ;
    RECT 68.35 41.085 68.56 41.155 ;
    RECT 68.35 41.445 68.56 41.515 ;
    RECT 68.35 41.805 68.56 41.875 ;
    RECT 28.05 41.085 28.26 41.155 ;
    RECT 28.05 41.445 28.26 41.515 ;
    RECT 28.05 41.805 28.26 41.875 ;
    RECT 28.51 41.085 28.72 41.155 ;
    RECT 28.51 41.445 28.72 41.515 ;
    RECT 28.51 41.805 28.72 41.875 ;
    RECT 24.73 41.085 24.94 41.155 ;
    RECT 24.73 41.445 24.94 41.515 ;
    RECT 24.73 41.805 24.94 41.875 ;
    RECT 25.19 41.085 25.4 41.155 ;
    RECT 25.19 41.445 25.4 41.515 ;
    RECT 25.19 41.805 25.4 41.875 ;
    RECT 21.41 41.085 21.62 41.155 ;
    RECT 21.41 41.445 21.62 41.515 ;
    RECT 21.41 41.805 21.62 41.875 ;
    RECT 21.87 41.085 22.08 41.155 ;
    RECT 21.87 41.445 22.08 41.515 ;
    RECT 21.87 41.805 22.08 41.875 ;
    RECT 18.09 41.085 18.3 41.155 ;
    RECT 18.09 41.445 18.3 41.515 ;
    RECT 18.09 41.805 18.3 41.875 ;
    RECT 18.55 41.085 18.76 41.155 ;
    RECT 18.55 41.445 18.76 41.515 ;
    RECT 18.55 41.805 18.76 41.875 ;
    RECT 14.77 41.085 14.98 41.155 ;
    RECT 14.77 41.445 14.98 41.515 ;
    RECT 14.77 41.805 14.98 41.875 ;
    RECT 15.23 41.085 15.44 41.155 ;
    RECT 15.23 41.445 15.44 41.515 ;
    RECT 15.23 41.805 15.44 41.875 ;
    RECT 11.45 41.085 11.66 41.155 ;
    RECT 11.45 41.445 11.66 41.515 ;
    RECT 11.45 41.805 11.66 41.875 ;
    RECT 11.91 41.085 12.12 41.155 ;
    RECT 11.91 41.445 12.12 41.515 ;
    RECT 11.91 41.805 12.12 41.875 ;
    RECT 8.13 41.085 8.34 41.155 ;
    RECT 8.13 41.445 8.34 41.515 ;
    RECT 8.13 41.805 8.34 41.875 ;
    RECT 8.59 41.085 8.8 41.155 ;
    RECT 8.59 41.445 8.8 41.515 ;
    RECT 8.59 41.805 8.8 41.875 ;
    RECT 4.81 41.085 5.02 41.155 ;
    RECT 4.81 41.445 5.02 41.515 ;
    RECT 4.81 41.805 5.02 41.875 ;
    RECT 5.27 41.085 5.48 41.155 ;
    RECT 5.27 41.445 5.48 41.515 ;
    RECT 5.27 41.805 5.48 41.875 ;
    RECT 164.17 41.085 164.38 41.155 ;
    RECT 164.17 41.445 164.38 41.515 ;
    RECT 164.17 41.805 164.38 41.875 ;
    RECT 164.63 41.085 164.84 41.155 ;
    RECT 164.63 41.445 164.84 41.515 ;
    RECT 164.63 41.805 164.84 41.875 ;
    RECT 1.49 41.085 1.7 41.155 ;
    RECT 1.49 41.445 1.7 41.515 ;
    RECT 1.49 41.805 1.7 41.875 ;
    RECT 1.95 41.085 2.16 41.155 ;
    RECT 1.95 41.445 2.16 41.515 ;
    RECT 1.95 41.805 2.16 41.875 ;
    RECT 160.85 41.085 161.06 41.155 ;
    RECT 160.85 41.445 161.06 41.515 ;
    RECT 160.85 41.805 161.06 41.875 ;
    RECT 161.31 41.085 161.52 41.155 ;
    RECT 161.31 41.445 161.52 41.515 ;
    RECT 161.31 41.805 161.52 41.875 ;
    RECT 157.53 41.085 157.74 41.155 ;
    RECT 157.53 41.445 157.74 41.515 ;
    RECT 157.53 41.805 157.74 41.875 ;
    RECT 157.99 41.085 158.2 41.155 ;
    RECT 157.99 41.445 158.2 41.515 ;
    RECT 157.99 41.805 158.2 41.875 ;
    RECT 154.21 41.085 154.42 41.155 ;
    RECT 154.21 41.445 154.42 41.515 ;
    RECT 154.21 41.805 154.42 41.875 ;
    RECT 154.67 41.085 154.88 41.155 ;
    RECT 154.67 41.445 154.88 41.515 ;
    RECT 154.67 41.805 154.88 41.875 ;
    RECT 150.89 41.085 151.1 41.155 ;
    RECT 150.89 41.445 151.1 41.515 ;
    RECT 150.89 41.805 151.1 41.875 ;
    RECT 151.35 41.085 151.56 41.155 ;
    RECT 151.35 41.445 151.56 41.515 ;
    RECT 151.35 41.805 151.56 41.875 ;
    RECT 147.57 41.085 147.78 41.155 ;
    RECT 147.57 41.445 147.78 41.515 ;
    RECT 147.57 41.805 147.78 41.875 ;
    RECT 148.03 41.085 148.24 41.155 ;
    RECT 148.03 41.445 148.24 41.515 ;
    RECT 148.03 41.805 148.24 41.875 ;
    RECT 144.25 41.085 144.46 41.155 ;
    RECT 144.25 41.445 144.46 41.515 ;
    RECT 144.25 41.805 144.46 41.875 ;
    RECT 144.71 41.085 144.92 41.155 ;
    RECT 144.71 41.445 144.92 41.515 ;
    RECT 144.71 41.805 144.92 41.875 ;
    RECT 140.93 41.085 141.14 41.155 ;
    RECT 140.93 41.445 141.14 41.515 ;
    RECT 140.93 41.805 141.14 41.875 ;
    RECT 141.39 41.085 141.6 41.155 ;
    RECT 141.39 41.445 141.6 41.515 ;
    RECT 141.39 41.805 141.6 41.875 ;
    RECT 137.61 41.085 137.82 41.155 ;
    RECT 137.61 41.445 137.82 41.515 ;
    RECT 137.61 41.805 137.82 41.875 ;
    RECT 138.07 41.085 138.28 41.155 ;
    RECT 138.07 41.445 138.28 41.515 ;
    RECT 138.07 41.805 138.28 41.875 ;
    RECT 134.29 41.085 134.5 41.155 ;
    RECT 134.29 41.445 134.5 41.515 ;
    RECT 134.29 41.805 134.5 41.875 ;
    RECT 134.75 41.085 134.96 41.155 ;
    RECT 134.75 41.445 134.96 41.515 ;
    RECT 134.75 41.805 134.96 41.875 ;
    RECT 64.57 41.085 64.78 41.155 ;
    RECT 64.57 41.445 64.78 41.515 ;
    RECT 64.57 41.805 64.78 41.875 ;
    RECT 65.03 41.085 65.24 41.155 ;
    RECT 65.03 41.445 65.24 41.515 ;
    RECT 65.03 41.805 65.24 41.875 ;
    RECT 61.25 40.365 61.46 40.435 ;
    RECT 61.25 40.725 61.46 40.795 ;
    RECT 61.25 41.085 61.46 41.155 ;
    RECT 61.71 40.365 61.92 40.435 ;
    RECT 61.71 40.725 61.92 40.795 ;
    RECT 61.71 41.085 61.92 41.155 ;
    RECT 57.93 40.365 58.14 40.435 ;
    RECT 57.93 40.725 58.14 40.795 ;
    RECT 57.93 41.085 58.14 41.155 ;
    RECT 58.39 40.365 58.6 40.435 ;
    RECT 58.39 40.725 58.6 40.795 ;
    RECT 58.39 41.085 58.6 41.155 ;
    RECT 54.61 40.365 54.82 40.435 ;
    RECT 54.61 40.725 54.82 40.795 ;
    RECT 54.61 41.085 54.82 41.155 ;
    RECT 55.07 40.365 55.28 40.435 ;
    RECT 55.07 40.725 55.28 40.795 ;
    RECT 55.07 41.085 55.28 41.155 ;
    RECT 51.29 40.365 51.5 40.435 ;
    RECT 51.29 40.725 51.5 40.795 ;
    RECT 51.29 41.085 51.5 41.155 ;
    RECT 51.75 40.365 51.96 40.435 ;
    RECT 51.75 40.725 51.96 40.795 ;
    RECT 51.75 41.085 51.96 41.155 ;
    RECT 47.97 40.365 48.18 40.435 ;
    RECT 47.97 40.725 48.18 40.795 ;
    RECT 47.97 41.085 48.18 41.155 ;
    RECT 48.43 40.365 48.64 40.435 ;
    RECT 48.43 40.725 48.64 40.795 ;
    RECT 48.43 41.085 48.64 41.155 ;
    RECT 44.65 40.365 44.86 40.435 ;
    RECT 44.65 40.725 44.86 40.795 ;
    RECT 44.65 41.085 44.86 41.155 ;
    RECT 45.11 40.365 45.32 40.435 ;
    RECT 45.11 40.725 45.32 40.795 ;
    RECT 45.11 41.085 45.32 41.155 ;
    RECT 41.33 40.365 41.54 40.435 ;
    RECT 41.33 40.725 41.54 40.795 ;
    RECT 41.33 41.085 41.54 41.155 ;
    RECT 41.79 40.365 42.0 40.435 ;
    RECT 41.79 40.725 42.0 40.795 ;
    RECT 41.79 41.085 42.0 41.155 ;
    RECT 38.01 40.365 38.22 40.435 ;
    RECT 38.01 40.725 38.22 40.795 ;
    RECT 38.01 41.085 38.22 41.155 ;
    RECT 38.47 40.365 38.68 40.435 ;
    RECT 38.47 40.725 38.68 40.795 ;
    RECT 38.47 41.085 38.68 41.155 ;
    RECT 34.69 40.365 34.9 40.435 ;
    RECT 34.69 40.725 34.9 40.795 ;
    RECT 34.69 41.085 34.9 41.155 ;
    RECT 35.15 40.365 35.36 40.435 ;
    RECT 35.15 40.725 35.36 40.795 ;
    RECT 35.15 41.085 35.36 41.155 ;
    RECT 173.945 40.725 174.015 40.795 ;
    RECT 130.97 40.365 131.18 40.435 ;
    RECT 130.97 40.725 131.18 40.795 ;
    RECT 130.97 41.085 131.18 41.155 ;
    RECT 131.43 40.365 131.64 40.435 ;
    RECT 131.43 40.725 131.64 40.795 ;
    RECT 131.43 41.085 131.64 41.155 ;
    RECT 127.65 40.365 127.86 40.435 ;
    RECT 127.65 40.725 127.86 40.795 ;
    RECT 127.65 41.085 127.86 41.155 ;
    RECT 128.11 40.365 128.32 40.435 ;
    RECT 128.11 40.725 128.32 40.795 ;
    RECT 128.11 41.085 128.32 41.155 ;
    RECT 124.33 40.365 124.54 40.435 ;
    RECT 124.33 40.725 124.54 40.795 ;
    RECT 124.33 41.085 124.54 41.155 ;
    RECT 124.79 40.365 125.0 40.435 ;
    RECT 124.79 40.725 125.0 40.795 ;
    RECT 124.79 41.085 125.0 41.155 ;
    RECT 121.01 40.365 121.22 40.435 ;
    RECT 121.01 40.725 121.22 40.795 ;
    RECT 121.01 41.085 121.22 41.155 ;
    RECT 121.47 40.365 121.68 40.435 ;
    RECT 121.47 40.725 121.68 40.795 ;
    RECT 121.47 41.085 121.68 41.155 ;
    RECT 117.69 40.365 117.9 40.435 ;
    RECT 117.69 40.725 117.9 40.795 ;
    RECT 117.69 41.085 117.9 41.155 ;
    RECT 118.15 40.365 118.36 40.435 ;
    RECT 118.15 40.725 118.36 40.795 ;
    RECT 118.15 41.085 118.36 41.155 ;
    RECT 114.37 40.365 114.58 40.435 ;
    RECT 114.37 40.725 114.58 40.795 ;
    RECT 114.37 41.085 114.58 41.155 ;
    RECT 114.83 40.365 115.04 40.435 ;
    RECT 114.83 40.725 115.04 40.795 ;
    RECT 114.83 41.085 115.04 41.155 ;
    RECT 111.05 40.365 111.26 40.435 ;
    RECT 111.05 40.725 111.26 40.795 ;
    RECT 111.05 41.085 111.26 41.155 ;
    RECT 111.51 40.365 111.72 40.435 ;
    RECT 111.51 40.725 111.72 40.795 ;
    RECT 111.51 41.085 111.72 41.155 ;
    RECT 107.73 40.365 107.94 40.435 ;
    RECT 107.73 40.725 107.94 40.795 ;
    RECT 107.73 41.085 107.94 41.155 ;
    RECT 108.19 40.365 108.4 40.435 ;
    RECT 108.19 40.725 108.4 40.795 ;
    RECT 108.19 41.085 108.4 41.155 ;
    RECT 104.41 40.365 104.62 40.435 ;
    RECT 104.41 40.725 104.62 40.795 ;
    RECT 104.41 41.085 104.62 41.155 ;
    RECT 104.87 40.365 105.08 40.435 ;
    RECT 104.87 40.725 105.08 40.795 ;
    RECT 104.87 41.085 105.08 41.155 ;
    RECT 101.09 40.365 101.3 40.435 ;
    RECT 101.09 40.725 101.3 40.795 ;
    RECT 101.09 41.085 101.3 41.155 ;
    RECT 101.55 40.365 101.76 40.435 ;
    RECT 101.55 40.725 101.76 40.795 ;
    RECT 101.55 41.085 101.76 41.155 ;
    RECT 0.4 40.725 0.47 40.795 ;
    RECT 170.81 40.365 171.02 40.435 ;
    RECT 170.81 40.725 171.02 40.795 ;
    RECT 170.81 41.085 171.02 41.155 ;
    RECT 171.27 40.365 171.48 40.435 ;
    RECT 171.27 40.725 171.48 40.795 ;
    RECT 171.27 41.085 171.48 41.155 ;
    RECT 167.49 40.365 167.7 40.435 ;
    RECT 167.49 40.725 167.7 40.795 ;
    RECT 167.49 41.085 167.7 41.155 ;
    RECT 167.95 40.365 168.16 40.435 ;
    RECT 167.95 40.725 168.16 40.795 ;
    RECT 167.95 41.085 168.16 41.155 ;
    RECT 97.77 40.365 97.98 40.435 ;
    RECT 97.77 40.725 97.98 40.795 ;
    RECT 97.77 41.085 97.98 41.155 ;
    RECT 98.23 40.365 98.44 40.435 ;
    RECT 98.23 40.725 98.44 40.795 ;
    RECT 98.23 41.085 98.44 41.155 ;
    RECT 94.45 40.365 94.66 40.435 ;
    RECT 94.45 40.725 94.66 40.795 ;
    RECT 94.45 41.085 94.66 41.155 ;
    RECT 94.91 40.365 95.12 40.435 ;
    RECT 94.91 40.725 95.12 40.795 ;
    RECT 94.91 41.085 95.12 41.155 ;
    RECT 91.13 40.365 91.34 40.435 ;
    RECT 91.13 40.725 91.34 40.795 ;
    RECT 91.13 41.085 91.34 41.155 ;
    RECT 91.59 40.365 91.8 40.435 ;
    RECT 91.59 40.725 91.8 40.795 ;
    RECT 91.59 41.085 91.8 41.155 ;
    RECT 87.81 40.365 88.02 40.435 ;
    RECT 87.81 40.725 88.02 40.795 ;
    RECT 87.81 41.085 88.02 41.155 ;
    RECT 88.27 40.365 88.48 40.435 ;
    RECT 88.27 40.725 88.48 40.795 ;
    RECT 88.27 41.085 88.48 41.155 ;
    RECT 84.49 40.365 84.7 40.435 ;
    RECT 84.49 40.725 84.7 40.795 ;
    RECT 84.49 41.085 84.7 41.155 ;
    RECT 84.95 40.365 85.16 40.435 ;
    RECT 84.95 40.725 85.16 40.795 ;
    RECT 84.95 41.085 85.16 41.155 ;
    RECT 81.17 40.365 81.38 40.435 ;
    RECT 81.17 40.725 81.38 40.795 ;
    RECT 81.17 41.085 81.38 41.155 ;
    RECT 81.63 40.365 81.84 40.435 ;
    RECT 81.63 40.725 81.84 40.795 ;
    RECT 81.63 41.085 81.84 41.155 ;
    RECT 77.85 40.365 78.06 40.435 ;
    RECT 77.85 40.725 78.06 40.795 ;
    RECT 77.85 41.085 78.06 41.155 ;
    RECT 78.31 40.365 78.52 40.435 ;
    RECT 78.31 40.725 78.52 40.795 ;
    RECT 78.31 41.085 78.52 41.155 ;
    RECT 74.53 40.365 74.74 40.435 ;
    RECT 74.53 40.725 74.74 40.795 ;
    RECT 74.53 41.085 74.74 41.155 ;
    RECT 74.99 40.365 75.2 40.435 ;
    RECT 74.99 40.725 75.2 40.795 ;
    RECT 74.99 41.085 75.2 41.155 ;
    RECT 71.21 40.365 71.42 40.435 ;
    RECT 71.21 40.725 71.42 40.795 ;
    RECT 71.21 41.085 71.42 41.155 ;
    RECT 71.67 40.365 71.88 40.435 ;
    RECT 71.67 40.725 71.88 40.795 ;
    RECT 71.67 41.085 71.88 41.155 ;
    RECT 31.37 40.365 31.58 40.435 ;
    RECT 31.37 40.725 31.58 40.795 ;
    RECT 31.37 41.085 31.58 41.155 ;
    RECT 31.83 40.365 32.04 40.435 ;
    RECT 31.83 40.725 32.04 40.795 ;
    RECT 31.83 41.085 32.04 41.155 ;
    RECT 67.89 40.365 68.1 40.435 ;
    RECT 67.89 40.725 68.1 40.795 ;
    RECT 67.89 41.085 68.1 41.155 ;
    RECT 68.35 40.365 68.56 40.435 ;
    RECT 68.35 40.725 68.56 40.795 ;
    RECT 68.35 41.085 68.56 41.155 ;
    RECT 28.05 40.365 28.26 40.435 ;
    RECT 28.05 40.725 28.26 40.795 ;
    RECT 28.05 41.085 28.26 41.155 ;
    RECT 28.51 40.365 28.72 40.435 ;
    RECT 28.51 40.725 28.72 40.795 ;
    RECT 28.51 41.085 28.72 41.155 ;
    RECT 24.73 40.365 24.94 40.435 ;
    RECT 24.73 40.725 24.94 40.795 ;
    RECT 24.73 41.085 24.94 41.155 ;
    RECT 25.19 40.365 25.4 40.435 ;
    RECT 25.19 40.725 25.4 40.795 ;
    RECT 25.19 41.085 25.4 41.155 ;
    RECT 21.41 40.365 21.62 40.435 ;
    RECT 21.41 40.725 21.62 40.795 ;
    RECT 21.41 41.085 21.62 41.155 ;
    RECT 21.87 40.365 22.08 40.435 ;
    RECT 21.87 40.725 22.08 40.795 ;
    RECT 21.87 41.085 22.08 41.155 ;
    RECT 18.09 40.365 18.3 40.435 ;
    RECT 18.09 40.725 18.3 40.795 ;
    RECT 18.09 41.085 18.3 41.155 ;
    RECT 18.55 40.365 18.76 40.435 ;
    RECT 18.55 40.725 18.76 40.795 ;
    RECT 18.55 41.085 18.76 41.155 ;
    RECT 14.77 40.365 14.98 40.435 ;
    RECT 14.77 40.725 14.98 40.795 ;
    RECT 14.77 41.085 14.98 41.155 ;
    RECT 15.23 40.365 15.44 40.435 ;
    RECT 15.23 40.725 15.44 40.795 ;
    RECT 15.23 41.085 15.44 41.155 ;
    RECT 11.45 40.365 11.66 40.435 ;
    RECT 11.45 40.725 11.66 40.795 ;
    RECT 11.45 41.085 11.66 41.155 ;
    RECT 11.91 40.365 12.12 40.435 ;
    RECT 11.91 40.725 12.12 40.795 ;
    RECT 11.91 41.085 12.12 41.155 ;
    RECT 8.13 40.365 8.34 40.435 ;
    RECT 8.13 40.725 8.34 40.795 ;
    RECT 8.13 41.085 8.34 41.155 ;
    RECT 8.59 40.365 8.8 40.435 ;
    RECT 8.59 40.725 8.8 40.795 ;
    RECT 8.59 41.085 8.8 41.155 ;
    RECT 4.81 40.365 5.02 40.435 ;
    RECT 4.81 40.725 5.02 40.795 ;
    RECT 4.81 41.085 5.02 41.155 ;
    RECT 5.27 40.365 5.48 40.435 ;
    RECT 5.27 40.725 5.48 40.795 ;
    RECT 5.27 41.085 5.48 41.155 ;
    RECT 164.17 40.365 164.38 40.435 ;
    RECT 164.17 40.725 164.38 40.795 ;
    RECT 164.17 41.085 164.38 41.155 ;
    RECT 164.63 40.365 164.84 40.435 ;
    RECT 164.63 40.725 164.84 40.795 ;
    RECT 164.63 41.085 164.84 41.155 ;
    RECT 1.49 40.365 1.7 40.435 ;
    RECT 1.49 40.725 1.7 40.795 ;
    RECT 1.49 41.085 1.7 41.155 ;
    RECT 1.95 40.365 2.16 40.435 ;
    RECT 1.95 40.725 2.16 40.795 ;
    RECT 1.95 41.085 2.16 41.155 ;
    RECT 160.85 40.365 161.06 40.435 ;
    RECT 160.85 40.725 161.06 40.795 ;
    RECT 160.85 41.085 161.06 41.155 ;
    RECT 161.31 40.365 161.52 40.435 ;
    RECT 161.31 40.725 161.52 40.795 ;
    RECT 161.31 41.085 161.52 41.155 ;
    RECT 157.53 40.365 157.74 40.435 ;
    RECT 157.53 40.725 157.74 40.795 ;
    RECT 157.53 41.085 157.74 41.155 ;
    RECT 157.99 40.365 158.2 40.435 ;
    RECT 157.99 40.725 158.2 40.795 ;
    RECT 157.99 41.085 158.2 41.155 ;
    RECT 154.21 40.365 154.42 40.435 ;
    RECT 154.21 40.725 154.42 40.795 ;
    RECT 154.21 41.085 154.42 41.155 ;
    RECT 154.67 40.365 154.88 40.435 ;
    RECT 154.67 40.725 154.88 40.795 ;
    RECT 154.67 41.085 154.88 41.155 ;
    RECT 150.89 40.365 151.1 40.435 ;
    RECT 150.89 40.725 151.1 40.795 ;
    RECT 150.89 41.085 151.1 41.155 ;
    RECT 151.35 40.365 151.56 40.435 ;
    RECT 151.35 40.725 151.56 40.795 ;
    RECT 151.35 41.085 151.56 41.155 ;
    RECT 147.57 40.365 147.78 40.435 ;
    RECT 147.57 40.725 147.78 40.795 ;
    RECT 147.57 41.085 147.78 41.155 ;
    RECT 148.03 40.365 148.24 40.435 ;
    RECT 148.03 40.725 148.24 40.795 ;
    RECT 148.03 41.085 148.24 41.155 ;
    RECT 144.25 40.365 144.46 40.435 ;
    RECT 144.25 40.725 144.46 40.795 ;
    RECT 144.25 41.085 144.46 41.155 ;
    RECT 144.71 40.365 144.92 40.435 ;
    RECT 144.71 40.725 144.92 40.795 ;
    RECT 144.71 41.085 144.92 41.155 ;
    RECT 140.93 40.365 141.14 40.435 ;
    RECT 140.93 40.725 141.14 40.795 ;
    RECT 140.93 41.085 141.14 41.155 ;
    RECT 141.39 40.365 141.6 40.435 ;
    RECT 141.39 40.725 141.6 40.795 ;
    RECT 141.39 41.085 141.6 41.155 ;
    RECT 137.61 40.365 137.82 40.435 ;
    RECT 137.61 40.725 137.82 40.795 ;
    RECT 137.61 41.085 137.82 41.155 ;
    RECT 138.07 40.365 138.28 40.435 ;
    RECT 138.07 40.725 138.28 40.795 ;
    RECT 138.07 41.085 138.28 41.155 ;
    RECT 134.29 40.365 134.5 40.435 ;
    RECT 134.29 40.725 134.5 40.795 ;
    RECT 134.29 41.085 134.5 41.155 ;
    RECT 134.75 40.365 134.96 40.435 ;
    RECT 134.75 40.725 134.96 40.795 ;
    RECT 134.75 41.085 134.96 41.155 ;
    RECT 64.57 40.365 64.78 40.435 ;
    RECT 64.57 40.725 64.78 40.795 ;
    RECT 64.57 41.085 64.78 41.155 ;
    RECT 65.03 40.365 65.24 40.435 ;
    RECT 65.03 40.725 65.24 40.795 ;
    RECT 65.03 41.085 65.24 41.155 ;
    RECT 61.25 39.645 61.46 39.715 ;
    RECT 61.25 40.005 61.46 40.075 ;
    RECT 61.25 40.365 61.46 40.435 ;
    RECT 61.71 39.645 61.92 39.715 ;
    RECT 61.71 40.005 61.92 40.075 ;
    RECT 61.71 40.365 61.92 40.435 ;
    RECT 57.93 39.645 58.14 39.715 ;
    RECT 57.93 40.005 58.14 40.075 ;
    RECT 57.93 40.365 58.14 40.435 ;
    RECT 58.39 39.645 58.6 39.715 ;
    RECT 58.39 40.005 58.6 40.075 ;
    RECT 58.39 40.365 58.6 40.435 ;
    RECT 54.61 39.645 54.82 39.715 ;
    RECT 54.61 40.005 54.82 40.075 ;
    RECT 54.61 40.365 54.82 40.435 ;
    RECT 55.07 39.645 55.28 39.715 ;
    RECT 55.07 40.005 55.28 40.075 ;
    RECT 55.07 40.365 55.28 40.435 ;
    RECT 51.29 39.645 51.5 39.715 ;
    RECT 51.29 40.005 51.5 40.075 ;
    RECT 51.29 40.365 51.5 40.435 ;
    RECT 51.75 39.645 51.96 39.715 ;
    RECT 51.75 40.005 51.96 40.075 ;
    RECT 51.75 40.365 51.96 40.435 ;
    RECT 47.97 39.645 48.18 39.715 ;
    RECT 47.97 40.005 48.18 40.075 ;
    RECT 47.97 40.365 48.18 40.435 ;
    RECT 48.43 39.645 48.64 39.715 ;
    RECT 48.43 40.005 48.64 40.075 ;
    RECT 48.43 40.365 48.64 40.435 ;
    RECT 44.65 39.645 44.86 39.715 ;
    RECT 44.65 40.005 44.86 40.075 ;
    RECT 44.65 40.365 44.86 40.435 ;
    RECT 45.11 39.645 45.32 39.715 ;
    RECT 45.11 40.005 45.32 40.075 ;
    RECT 45.11 40.365 45.32 40.435 ;
    RECT 41.33 39.645 41.54 39.715 ;
    RECT 41.33 40.005 41.54 40.075 ;
    RECT 41.33 40.365 41.54 40.435 ;
    RECT 41.79 39.645 42.0 39.715 ;
    RECT 41.79 40.005 42.0 40.075 ;
    RECT 41.79 40.365 42.0 40.435 ;
    RECT 38.01 39.645 38.22 39.715 ;
    RECT 38.01 40.005 38.22 40.075 ;
    RECT 38.01 40.365 38.22 40.435 ;
    RECT 38.47 39.645 38.68 39.715 ;
    RECT 38.47 40.005 38.68 40.075 ;
    RECT 38.47 40.365 38.68 40.435 ;
    RECT 34.69 39.645 34.9 39.715 ;
    RECT 34.69 40.005 34.9 40.075 ;
    RECT 34.69 40.365 34.9 40.435 ;
    RECT 35.15 39.645 35.36 39.715 ;
    RECT 35.15 40.005 35.36 40.075 ;
    RECT 35.15 40.365 35.36 40.435 ;
    RECT 173.945 40.005 174.015 40.075 ;
    RECT 130.97 39.645 131.18 39.715 ;
    RECT 130.97 40.005 131.18 40.075 ;
    RECT 130.97 40.365 131.18 40.435 ;
    RECT 131.43 39.645 131.64 39.715 ;
    RECT 131.43 40.005 131.64 40.075 ;
    RECT 131.43 40.365 131.64 40.435 ;
    RECT 127.65 39.645 127.86 39.715 ;
    RECT 127.65 40.005 127.86 40.075 ;
    RECT 127.65 40.365 127.86 40.435 ;
    RECT 128.11 39.645 128.32 39.715 ;
    RECT 128.11 40.005 128.32 40.075 ;
    RECT 128.11 40.365 128.32 40.435 ;
    RECT 124.33 39.645 124.54 39.715 ;
    RECT 124.33 40.005 124.54 40.075 ;
    RECT 124.33 40.365 124.54 40.435 ;
    RECT 124.79 39.645 125.0 39.715 ;
    RECT 124.79 40.005 125.0 40.075 ;
    RECT 124.79 40.365 125.0 40.435 ;
    RECT 121.01 39.645 121.22 39.715 ;
    RECT 121.01 40.005 121.22 40.075 ;
    RECT 121.01 40.365 121.22 40.435 ;
    RECT 121.47 39.645 121.68 39.715 ;
    RECT 121.47 40.005 121.68 40.075 ;
    RECT 121.47 40.365 121.68 40.435 ;
    RECT 117.69 39.645 117.9 39.715 ;
    RECT 117.69 40.005 117.9 40.075 ;
    RECT 117.69 40.365 117.9 40.435 ;
    RECT 118.15 39.645 118.36 39.715 ;
    RECT 118.15 40.005 118.36 40.075 ;
    RECT 118.15 40.365 118.36 40.435 ;
    RECT 114.37 39.645 114.58 39.715 ;
    RECT 114.37 40.005 114.58 40.075 ;
    RECT 114.37 40.365 114.58 40.435 ;
    RECT 114.83 39.645 115.04 39.715 ;
    RECT 114.83 40.005 115.04 40.075 ;
    RECT 114.83 40.365 115.04 40.435 ;
    RECT 111.05 39.645 111.26 39.715 ;
    RECT 111.05 40.005 111.26 40.075 ;
    RECT 111.05 40.365 111.26 40.435 ;
    RECT 111.51 39.645 111.72 39.715 ;
    RECT 111.51 40.005 111.72 40.075 ;
    RECT 111.51 40.365 111.72 40.435 ;
    RECT 107.73 39.645 107.94 39.715 ;
    RECT 107.73 40.005 107.94 40.075 ;
    RECT 107.73 40.365 107.94 40.435 ;
    RECT 108.19 39.645 108.4 39.715 ;
    RECT 108.19 40.005 108.4 40.075 ;
    RECT 108.19 40.365 108.4 40.435 ;
    RECT 104.41 39.645 104.62 39.715 ;
    RECT 104.41 40.005 104.62 40.075 ;
    RECT 104.41 40.365 104.62 40.435 ;
    RECT 104.87 39.645 105.08 39.715 ;
    RECT 104.87 40.005 105.08 40.075 ;
    RECT 104.87 40.365 105.08 40.435 ;
    RECT 101.09 39.645 101.3 39.715 ;
    RECT 101.09 40.005 101.3 40.075 ;
    RECT 101.09 40.365 101.3 40.435 ;
    RECT 101.55 39.645 101.76 39.715 ;
    RECT 101.55 40.005 101.76 40.075 ;
    RECT 101.55 40.365 101.76 40.435 ;
    RECT 0.4 40.005 0.47 40.075 ;
    RECT 170.81 39.645 171.02 39.715 ;
    RECT 170.81 40.005 171.02 40.075 ;
    RECT 170.81 40.365 171.02 40.435 ;
    RECT 171.27 39.645 171.48 39.715 ;
    RECT 171.27 40.005 171.48 40.075 ;
    RECT 171.27 40.365 171.48 40.435 ;
    RECT 167.49 39.645 167.7 39.715 ;
    RECT 167.49 40.005 167.7 40.075 ;
    RECT 167.49 40.365 167.7 40.435 ;
    RECT 167.95 39.645 168.16 39.715 ;
    RECT 167.95 40.005 168.16 40.075 ;
    RECT 167.95 40.365 168.16 40.435 ;
    RECT 97.77 39.645 97.98 39.715 ;
    RECT 97.77 40.005 97.98 40.075 ;
    RECT 97.77 40.365 97.98 40.435 ;
    RECT 98.23 39.645 98.44 39.715 ;
    RECT 98.23 40.005 98.44 40.075 ;
    RECT 98.23 40.365 98.44 40.435 ;
    RECT 94.45 39.645 94.66 39.715 ;
    RECT 94.45 40.005 94.66 40.075 ;
    RECT 94.45 40.365 94.66 40.435 ;
    RECT 94.91 39.645 95.12 39.715 ;
    RECT 94.91 40.005 95.12 40.075 ;
    RECT 94.91 40.365 95.12 40.435 ;
    RECT 91.13 39.645 91.34 39.715 ;
    RECT 91.13 40.005 91.34 40.075 ;
    RECT 91.13 40.365 91.34 40.435 ;
    RECT 91.59 39.645 91.8 39.715 ;
    RECT 91.59 40.005 91.8 40.075 ;
    RECT 91.59 40.365 91.8 40.435 ;
    RECT 87.81 39.645 88.02 39.715 ;
    RECT 87.81 40.005 88.02 40.075 ;
    RECT 87.81 40.365 88.02 40.435 ;
    RECT 88.27 39.645 88.48 39.715 ;
    RECT 88.27 40.005 88.48 40.075 ;
    RECT 88.27 40.365 88.48 40.435 ;
    RECT 84.49 39.645 84.7 39.715 ;
    RECT 84.49 40.005 84.7 40.075 ;
    RECT 84.49 40.365 84.7 40.435 ;
    RECT 84.95 39.645 85.16 39.715 ;
    RECT 84.95 40.005 85.16 40.075 ;
    RECT 84.95 40.365 85.16 40.435 ;
    RECT 81.17 39.645 81.38 39.715 ;
    RECT 81.17 40.005 81.38 40.075 ;
    RECT 81.17 40.365 81.38 40.435 ;
    RECT 81.63 39.645 81.84 39.715 ;
    RECT 81.63 40.005 81.84 40.075 ;
    RECT 81.63 40.365 81.84 40.435 ;
    RECT 77.85 39.645 78.06 39.715 ;
    RECT 77.85 40.005 78.06 40.075 ;
    RECT 77.85 40.365 78.06 40.435 ;
    RECT 78.31 39.645 78.52 39.715 ;
    RECT 78.31 40.005 78.52 40.075 ;
    RECT 78.31 40.365 78.52 40.435 ;
    RECT 74.53 39.645 74.74 39.715 ;
    RECT 74.53 40.005 74.74 40.075 ;
    RECT 74.53 40.365 74.74 40.435 ;
    RECT 74.99 39.645 75.2 39.715 ;
    RECT 74.99 40.005 75.2 40.075 ;
    RECT 74.99 40.365 75.2 40.435 ;
    RECT 71.21 39.645 71.42 39.715 ;
    RECT 71.21 40.005 71.42 40.075 ;
    RECT 71.21 40.365 71.42 40.435 ;
    RECT 71.67 39.645 71.88 39.715 ;
    RECT 71.67 40.005 71.88 40.075 ;
    RECT 71.67 40.365 71.88 40.435 ;
    RECT 31.37 39.645 31.58 39.715 ;
    RECT 31.37 40.005 31.58 40.075 ;
    RECT 31.37 40.365 31.58 40.435 ;
    RECT 31.83 39.645 32.04 39.715 ;
    RECT 31.83 40.005 32.04 40.075 ;
    RECT 31.83 40.365 32.04 40.435 ;
    RECT 67.89 39.645 68.1 39.715 ;
    RECT 67.89 40.005 68.1 40.075 ;
    RECT 67.89 40.365 68.1 40.435 ;
    RECT 68.35 39.645 68.56 39.715 ;
    RECT 68.35 40.005 68.56 40.075 ;
    RECT 68.35 40.365 68.56 40.435 ;
    RECT 28.05 39.645 28.26 39.715 ;
    RECT 28.05 40.005 28.26 40.075 ;
    RECT 28.05 40.365 28.26 40.435 ;
    RECT 28.51 39.645 28.72 39.715 ;
    RECT 28.51 40.005 28.72 40.075 ;
    RECT 28.51 40.365 28.72 40.435 ;
    RECT 24.73 39.645 24.94 39.715 ;
    RECT 24.73 40.005 24.94 40.075 ;
    RECT 24.73 40.365 24.94 40.435 ;
    RECT 25.19 39.645 25.4 39.715 ;
    RECT 25.19 40.005 25.4 40.075 ;
    RECT 25.19 40.365 25.4 40.435 ;
    RECT 21.41 39.645 21.62 39.715 ;
    RECT 21.41 40.005 21.62 40.075 ;
    RECT 21.41 40.365 21.62 40.435 ;
    RECT 21.87 39.645 22.08 39.715 ;
    RECT 21.87 40.005 22.08 40.075 ;
    RECT 21.87 40.365 22.08 40.435 ;
    RECT 18.09 39.645 18.3 39.715 ;
    RECT 18.09 40.005 18.3 40.075 ;
    RECT 18.09 40.365 18.3 40.435 ;
    RECT 18.55 39.645 18.76 39.715 ;
    RECT 18.55 40.005 18.76 40.075 ;
    RECT 18.55 40.365 18.76 40.435 ;
    RECT 14.77 39.645 14.98 39.715 ;
    RECT 14.77 40.005 14.98 40.075 ;
    RECT 14.77 40.365 14.98 40.435 ;
    RECT 15.23 39.645 15.44 39.715 ;
    RECT 15.23 40.005 15.44 40.075 ;
    RECT 15.23 40.365 15.44 40.435 ;
    RECT 11.45 39.645 11.66 39.715 ;
    RECT 11.45 40.005 11.66 40.075 ;
    RECT 11.45 40.365 11.66 40.435 ;
    RECT 11.91 39.645 12.12 39.715 ;
    RECT 11.91 40.005 12.12 40.075 ;
    RECT 11.91 40.365 12.12 40.435 ;
    RECT 8.13 39.645 8.34 39.715 ;
    RECT 8.13 40.005 8.34 40.075 ;
    RECT 8.13 40.365 8.34 40.435 ;
    RECT 8.59 39.645 8.8 39.715 ;
    RECT 8.59 40.005 8.8 40.075 ;
    RECT 8.59 40.365 8.8 40.435 ;
    RECT 4.81 39.645 5.02 39.715 ;
    RECT 4.81 40.005 5.02 40.075 ;
    RECT 4.81 40.365 5.02 40.435 ;
    RECT 5.27 39.645 5.48 39.715 ;
    RECT 5.27 40.005 5.48 40.075 ;
    RECT 5.27 40.365 5.48 40.435 ;
    RECT 164.17 39.645 164.38 39.715 ;
    RECT 164.17 40.005 164.38 40.075 ;
    RECT 164.17 40.365 164.38 40.435 ;
    RECT 164.63 39.645 164.84 39.715 ;
    RECT 164.63 40.005 164.84 40.075 ;
    RECT 164.63 40.365 164.84 40.435 ;
    RECT 1.49 39.645 1.7 39.715 ;
    RECT 1.49 40.005 1.7 40.075 ;
    RECT 1.49 40.365 1.7 40.435 ;
    RECT 1.95 39.645 2.16 39.715 ;
    RECT 1.95 40.005 2.16 40.075 ;
    RECT 1.95 40.365 2.16 40.435 ;
    RECT 160.85 39.645 161.06 39.715 ;
    RECT 160.85 40.005 161.06 40.075 ;
    RECT 160.85 40.365 161.06 40.435 ;
    RECT 161.31 39.645 161.52 39.715 ;
    RECT 161.31 40.005 161.52 40.075 ;
    RECT 161.31 40.365 161.52 40.435 ;
    RECT 157.53 39.645 157.74 39.715 ;
    RECT 157.53 40.005 157.74 40.075 ;
    RECT 157.53 40.365 157.74 40.435 ;
    RECT 157.99 39.645 158.2 39.715 ;
    RECT 157.99 40.005 158.2 40.075 ;
    RECT 157.99 40.365 158.2 40.435 ;
    RECT 154.21 39.645 154.42 39.715 ;
    RECT 154.21 40.005 154.42 40.075 ;
    RECT 154.21 40.365 154.42 40.435 ;
    RECT 154.67 39.645 154.88 39.715 ;
    RECT 154.67 40.005 154.88 40.075 ;
    RECT 154.67 40.365 154.88 40.435 ;
    RECT 150.89 39.645 151.1 39.715 ;
    RECT 150.89 40.005 151.1 40.075 ;
    RECT 150.89 40.365 151.1 40.435 ;
    RECT 151.35 39.645 151.56 39.715 ;
    RECT 151.35 40.005 151.56 40.075 ;
    RECT 151.35 40.365 151.56 40.435 ;
    RECT 147.57 39.645 147.78 39.715 ;
    RECT 147.57 40.005 147.78 40.075 ;
    RECT 147.57 40.365 147.78 40.435 ;
    RECT 148.03 39.645 148.24 39.715 ;
    RECT 148.03 40.005 148.24 40.075 ;
    RECT 148.03 40.365 148.24 40.435 ;
    RECT 144.25 39.645 144.46 39.715 ;
    RECT 144.25 40.005 144.46 40.075 ;
    RECT 144.25 40.365 144.46 40.435 ;
    RECT 144.71 39.645 144.92 39.715 ;
    RECT 144.71 40.005 144.92 40.075 ;
    RECT 144.71 40.365 144.92 40.435 ;
    RECT 140.93 39.645 141.14 39.715 ;
    RECT 140.93 40.005 141.14 40.075 ;
    RECT 140.93 40.365 141.14 40.435 ;
    RECT 141.39 39.645 141.6 39.715 ;
    RECT 141.39 40.005 141.6 40.075 ;
    RECT 141.39 40.365 141.6 40.435 ;
    RECT 137.61 39.645 137.82 39.715 ;
    RECT 137.61 40.005 137.82 40.075 ;
    RECT 137.61 40.365 137.82 40.435 ;
    RECT 138.07 39.645 138.28 39.715 ;
    RECT 138.07 40.005 138.28 40.075 ;
    RECT 138.07 40.365 138.28 40.435 ;
    RECT 134.29 39.645 134.5 39.715 ;
    RECT 134.29 40.005 134.5 40.075 ;
    RECT 134.29 40.365 134.5 40.435 ;
    RECT 134.75 39.645 134.96 39.715 ;
    RECT 134.75 40.005 134.96 40.075 ;
    RECT 134.75 40.365 134.96 40.435 ;
    RECT 64.57 39.645 64.78 39.715 ;
    RECT 64.57 40.005 64.78 40.075 ;
    RECT 64.57 40.365 64.78 40.435 ;
    RECT 65.03 39.645 65.24 39.715 ;
    RECT 65.03 40.005 65.24 40.075 ;
    RECT 65.03 40.365 65.24 40.435 ;
    RECT 61.25 58.385 61.46 58.455 ;
    RECT 61.25 58.745 61.46 58.815 ;
    RECT 61.25 59.105 61.46 59.175 ;
    RECT 61.71 58.385 61.92 58.455 ;
    RECT 61.71 58.745 61.92 58.815 ;
    RECT 61.71 59.105 61.92 59.175 ;
    RECT 57.93 58.385 58.14 58.455 ;
    RECT 57.93 58.745 58.14 58.815 ;
    RECT 57.93 59.105 58.14 59.175 ;
    RECT 58.39 58.385 58.6 58.455 ;
    RECT 58.39 58.745 58.6 58.815 ;
    RECT 58.39 59.105 58.6 59.175 ;
    RECT 54.61 58.385 54.82 58.455 ;
    RECT 54.61 58.745 54.82 58.815 ;
    RECT 54.61 59.105 54.82 59.175 ;
    RECT 55.07 58.385 55.28 58.455 ;
    RECT 55.07 58.745 55.28 58.815 ;
    RECT 55.07 59.105 55.28 59.175 ;
    RECT 170.81 58.385 171.02 58.455 ;
    RECT 170.81 58.745 171.02 58.815 ;
    RECT 170.81 59.105 171.02 59.175 ;
    RECT 171.27 58.385 171.48 58.455 ;
    RECT 171.27 58.745 171.48 58.815 ;
    RECT 171.27 59.105 171.48 59.175 ;
    RECT 51.29 58.385 51.5 58.455 ;
    RECT 51.29 58.745 51.5 58.815 ;
    RECT 51.29 59.105 51.5 59.175 ;
    RECT 51.75 58.385 51.96 58.455 ;
    RECT 51.75 58.745 51.96 58.815 ;
    RECT 51.75 59.105 51.96 59.175 ;
    RECT 47.97 58.385 48.18 58.455 ;
    RECT 47.97 58.745 48.18 58.815 ;
    RECT 47.97 59.105 48.18 59.175 ;
    RECT 48.43 58.385 48.64 58.455 ;
    RECT 48.43 58.745 48.64 58.815 ;
    RECT 48.43 59.105 48.64 59.175 ;
    RECT 44.65 58.385 44.86 58.455 ;
    RECT 44.65 58.745 44.86 58.815 ;
    RECT 44.65 59.105 44.86 59.175 ;
    RECT 45.11 58.385 45.32 58.455 ;
    RECT 45.11 58.745 45.32 58.815 ;
    RECT 45.11 59.105 45.32 59.175 ;
    RECT 41.33 58.385 41.54 58.455 ;
    RECT 41.33 58.745 41.54 58.815 ;
    RECT 41.33 59.105 41.54 59.175 ;
    RECT 41.79 58.385 42.0 58.455 ;
    RECT 41.79 58.745 42.0 58.815 ;
    RECT 41.79 59.105 42.0 59.175 ;
    RECT 38.01 58.385 38.22 58.455 ;
    RECT 38.01 58.745 38.22 58.815 ;
    RECT 38.01 59.105 38.22 59.175 ;
    RECT 38.47 58.385 38.68 58.455 ;
    RECT 38.47 58.745 38.68 58.815 ;
    RECT 38.47 59.105 38.68 59.175 ;
    RECT 34.69 58.385 34.9 58.455 ;
    RECT 34.69 58.745 34.9 58.815 ;
    RECT 34.69 59.105 34.9 59.175 ;
    RECT 35.15 58.385 35.36 58.455 ;
    RECT 35.15 58.745 35.36 58.815 ;
    RECT 35.15 59.105 35.36 59.175 ;
    RECT 1.49 58.385 1.7 58.455 ;
    RECT 1.49 58.745 1.7 58.815 ;
    RECT 1.49 59.105 1.7 59.175 ;
    RECT 1.95 58.385 2.16 58.455 ;
    RECT 1.95 58.745 2.16 58.815 ;
    RECT 1.95 59.105 2.16 59.175 ;
    RECT 130.97 58.385 131.18 58.455 ;
    RECT 130.97 58.745 131.18 58.815 ;
    RECT 130.97 59.105 131.18 59.175 ;
    RECT 131.43 58.385 131.64 58.455 ;
    RECT 131.43 58.745 131.64 58.815 ;
    RECT 131.43 59.105 131.64 59.175 ;
    RECT 127.65 58.385 127.86 58.455 ;
    RECT 127.65 58.745 127.86 58.815 ;
    RECT 127.65 59.105 127.86 59.175 ;
    RECT 128.11 58.385 128.32 58.455 ;
    RECT 128.11 58.745 128.32 58.815 ;
    RECT 128.11 59.105 128.32 59.175 ;
    RECT 124.33 58.385 124.54 58.455 ;
    RECT 124.33 58.745 124.54 58.815 ;
    RECT 124.33 59.105 124.54 59.175 ;
    RECT 124.79 58.385 125.0 58.455 ;
    RECT 124.79 58.745 125.0 58.815 ;
    RECT 124.79 59.105 125.0 59.175 ;
    RECT 121.01 58.385 121.22 58.455 ;
    RECT 121.01 58.745 121.22 58.815 ;
    RECT 121.01 59.105 121.22 59.175 ;
    RECT 121.47 58.385 121.68 58.455 ;
    RECT 121.47 58.745 121.68 58.815 ;
    RECT 121.47 59.105 121.68 59.175 ;
    RECT 117.69 58.385 117.9 58.455 ;
    RECT 117.69 58.745 117.9 58.815 ;
    RECT 117.69 59.105 117.9 59.175 ;
    RECT 118.15 58.385 118.36 58.455 ;
    RECT 118.15 58.745 118.36 58.815 ;
    RECT 118.15 59.105 118.36 59.175 ;
    RECT 114.37 58.385 114.58 58.455 ;
    RECT 114.37 58.745 114.58 58.815 ;
    RECT 114.37 59.105 114.58 59.175 ;
    RECT 114.83 58.385 115.04 58.455 ;
    RECT 114.83 58.745 115.04 58.815 ;
    RECT 114.83 59.105 115.04 59.175 ;
    RECT 111.05 58.385 111.26 58.455 ;
    RECT 111.05 58.745 111.26 58.815 ;
    RECT 111.05 59.105 111.26 59.175 ;
    RECT 111.51 58.385 111.72 58.455 ;
    RECT 111.51 58.745 111.72 58.815 ;
    RECT 111.51 59.105 111.72 59.175 ;
    RECT 107.73 58.385 107.94 58.455 ;
    RECT 107.73 58.745 107.94 58.815 ;
    RECT 107.73 59.105 107.94 59.175 ;
    RECT 108.19 58.385 108.4 58.455 ;
    RECT 108.19 58.745 108.4 58.815 ;
    RECT 108.19 59.105 108.4 59.175 ;
    RECT 104.41 58.385 104.62 58.455 ;
    RECT 104.41 58.745 104.62 58.815 ;
    RECT 104.41 59.105 104.62 59.175 ;
    RECT 104.87 58.385 105.08 58.455 ;
    RECT 104.87 58.745 105.08 58.815 ;
    RECT 104.87 59.105 105.08 59.175 ;
    RECT 101.09 58.385 101.3 58.455 ;
    RECT 101.09 58.745 101.3 58.815 ;
    RECT 101.09 59.105 101.3 59.175 ;
    RECT 101.55 58.385 101.76 58.455 ;
    RECT 101.55 58.745 101.76 58.815 ;
    RECT 101.55 59.105 101.76 59.175 ;
    RECT 167.49 58.385 167.7 58.455 ;
    RECT 167.49 58.745 167.7 58.815 ;
    RECT 167.49 59.105 167.7 59.175 ;
    RECT 167.95 58.385 168.16 58.455 ;
    RECT 167.95 58.745 168.16 58.815 ;
    RECT 167.95 59.105 168.16 59.175 ;
    RECT 173.945 58.745 174.015 58.815 ;
    RECT 97.77 58.385 97.98 58.455 ;
    RECT 97.77 58.745 97.98 58.815 ;
    RECT 97.77 59.105 97.98 59.175 ;
    RECT 98.23 58.385 98.44 58.455 ;
    RECT 98.23 58.745 98.44 58.815 ;
    RECT 98.23 59.105 98.44 59.175 ;
    RECT 94.45 58.385 94.66 58.455 ;
    RECT 94.45 58.745 94.66 58.815 ;
    RECT 94.45 59.105 94.66 59.175 ;
    RECT 94.91 58.385 95.12 58.455 ;
    RECT 94.91 58.745 95.12 58.815 ;
    RECT 94.91 59.105 95.12 59.175 ;
    RECT 91.13 58.385 91.34 58.455 ;
    RECT 91.13 58.745 91.34 58.815 ;
    RECT 91.13 59.105 91.34 59.175 ;
    RECT 91.59 58.385 91.8 58.455 ;
    RECT 91.59 58.745 91.8 58.815 ;
    RECT 91.59 59.105 91.8 59.175 ;
    RECT 87.81 58.385 88.02 58.455 ;
    RECT 87.81 58.745 88.02 58.815 ;
    RECT 87.81 59.105 88.02 59.175 ;
    RECT 88.27 58.385 88.48 58.455 ;
    RECT 88.27 58.745 88.48 58.815 ;
    RECT 88.27 59.105 88.48 59.175 ;
    RECT 84.49 58.385 84.7 58.455 ;
    RECT 84.49 58.745 84.7 58.815 ;
    RECT 84.49 59.105 84.7 59.175 ;
    RECT 84.95 58.385 85.16 58.455 ;
    RECT 84.95 58.745 85.16 58.815 ;
    RECT 84.95 59.105 85.16 59.175 ;
    RECT 81.17 58.385 81.38 58.455 ;
    RECT 81.17 58.745 81.38 58.815 ;
    RECT 81.17 59.105 81.38 59.175 ;
    RECT 81.63 58.385 81.84 58.455 ;
    RECT 81.63 58.745 81.84 58.815 ;
    RECT 81.63 59.105 81.84 59.175 ;
    RECT 77.85 58.385 78.06 58.455 ;
    RECT 77.85 58.745 78.06 58.815 ;
    RECT 77.85 59.105 78.06 59.175 ;
    RECT 78.31 58.385 78.52 58.455 ;
    RECT 78.31 58.745 78.52 58.815 ;
    RECT 78.31 59.105 78.52 59.175 ;
    RECT 74.53 58.385 74.74 58.455 ;
    RECT 74.53 58.745 74.74 58.815 ;
    RECT 74.53 59.105 74.74 59.175 ;
    RECT 74.99 58.385 75.2 58.455 ;
    RECT 74.99 58.745 75.2 58.815 ;
    RECT 74.99 59.105 75.2 59.175 ;
    RECT 71.21 58.385 71.42 58.455 ;
    RECT 71.21 58.745 71.42 58.815 ;
    RECT 71.21 59.105 71.42 59.175 ;
    RECT 71.67 58.385 71.88 58.455 ;
    RECT 71.67 58.745 71.88 58.815 ;
    RECT 71.67 59.105 71.88 59.175 ;
    RECT 31.37 58.385 31.58 58.455 ;
    RECT 31.37 58.745 31.58 58.815 ;
    RECT 31.37 59.105 31.58 59.175 ;
    RECT 31.83 58.385 32.04 58.455 ;
    RECT 31.83 58.745 32.04 58.815 ;
    RECT 31.83 59.105 32.04 59.175 ;
    RECT 67.89 58.385 68.1 58.455 ;
    RECT 67.89 58.745 68.1 58.815 ;
    RECT 67.89 59.105 68.1 59.175 ;
    RECT 68.35 58.385 68.56 58.455 ;
    RECT 68.35 58.745 68.56 58.815 ;
    RECT 68.35 59.105 68.56 59.175 ;
    RECT 28.05 58.385 28.26 58.455 ;
    RECT 28.05 58.745 28.26 58.815 ;
    RECT 28.05 59.105 28.26 59.175 ;
    RECT 28.51 58.385 28.72 58.455 ;
    RECT 28.51 58.745 28.72 58.815 ;
    RECT 28.51 59.105 28.72 59.175 ;
    RECT 24.73 58.385 24.94 58.455 ;
    RECT 24.73 58.745 24.94 58.815 ;
    RECT 24.73 59.105 24.94 59.175 ;
    RECT 25.19 58.385 25.4 58.455 ;
    RECT 25.19 58.745 25.4 58.815 ;
    RECT 25.19 59.105 25.4 59.175 ;
    RECT 21.41 58.385 21.62 58.455 ;
    RECT 21.41 58.745 21.62 58.815 ;
    RECT 21.41 59.105 21.62 59.175 ;
    RECT 21.87 58.385 22.08 58.455 ;
    RECT 21.87 58.745 22.08 58.815 ;
    RECT 21.87 59.105 22.08 59.175 ;
    RECT 18.09 58.385 18.3 58.455 ;
    RECT 18.09 58.745 18.3 58.815 ;
    RECT 18.09 59.105 18.3 59.175 ;
    RECT 18.55 58.385 18.76 58.455 ;
    RECT 18.55 58.745 18.76 58.815 ;
    RECT 18.55 59.105 18.76 59.175 ;
    RECT 14.77 58.385 14.98 58.455 ;
    RECT 14.77 58.745 14.98 58.815 ;
    RECT 14.77 59.105 14.98 59.175 ;
    RECT 15.23 58.385 15.44 58.455 ;
    RECT 15.23 58.745 15.44 58.815 ;
    RECT 15.23 59.105 15.44 59.175 ;
    RECT 11.45 58.385 11.66 58.455 ;
    RECT 11.45 58.745 11.66 58.815 ;
    RECT 11.45 59.105 11.66 59.175 ;
    RECT 11.91 58.385 12.12 58.455 ;
    RECT 11.91 58.745 12.12 58.815 ;
    RECT 11.91 59.105 12.12 59.175 ;
    RECT 8.13 58.385 8.34 58.455 ;
    RECT 8.13 58.745 8.34 58.815 ;
    RECT 8.13 59.105 8.34 59.175 ;
    RECT 8.59 58.385 8.8 58.455 ;
    RECT 8.59 58.745 8.8 58.815 ;
    RECT 8.59 59.105 8.8 59.175 ;
    RECT 4.81 58.385 5.02 58.455 ;
    RECT 4.81 58.745 5.02 58.815 ;
    RECT 4.81 59.105 5.02 59.175 ;
    RECT 5.27 58.385 5.48 58.455 ;
    RECT 5.27 58.745 5.48 58.815 ;
    RECT 5.27 59.105 5.48 59.175 ;
    RECT 164.17 58.385 164.38 58.455 ;
    RECT 164.17 58.745 164.38 58.815 ;
    RECT 164.17 59.105 164.38 59.175 ;
    RECT 164.63 58.385 164.84 58.455 ;
    RECT 164.63 58.745 164.84 58.815 ;
    RECT 164.63 59.105 164.84 59.175 ;
    RECT 160.85 58.385 161.06 58.455 ;
    RECT 160.85 58.745 161.06 58.815 ;
    RECT 160.85 59.105 161.06 59.175 ;
    RECT 161.31 58.385 161.52 58.455 ;
    RECT 161.31 58.745 161.52 58.815 ;
    RECT 161.31 59.105 161.52 59.175 ;
    RECT 157.53 58.385 157.74 58.455 ;
    RECT 157.53 58.745 157.74 58.815 ;
    RECT 157.53 59.105 157.74 59.175 ;
    RECT 157.99 58.385 158.2 58.455 ;
    RECT 157.99 58.745 158.2 58.815 ;
    RECT 157.99 59.105 158.2 59.175 ;
    RECT 154.21 58.385 154.42 58.455 ;
    RECT 154.21 58.745 154.42 58.815 ;
    RECT 154.21 59.105 154.42 59.175 ;
    RECT 154.67 58.385 154.88 58.455 ;
    RECT 154.67 58.745 154.88 58.815 ;
    RECT 154.67 59.105 154.88 59.175 ;
    RECT 150.89 58.385 151.1 58.455 ;
    RECT 150.89 58.745 151.1 58.815 ;
    RECT 150.89 59.105 151.1 59.175 ;
    RECT 151.35 58.385 151.56 58.455 ;
    RECT 151.35 58.745 151.56 58.815 ;
    RECT 151.35 59.105 151.56 59.175 ;
    RECT 147.57 58.385 147.78 58.455 ;
    RECT 147.57 58.745 147.78 58.815 ;
    RECT 147.57 59.105 147.78 59.175 ;
    RECT 148.03 58.385 148.24 58.455 ;
    RECT 148.03 58.745 148.24 58.815 ;
    RECT 148.03 59.105 148.24 59.175 ;
    RECT 144.25 58.385 144.46 58.455 ;
    RECT 144.25 58.745 144.46 58.815 ;
    RECT 144.25 59.105 144.46 59.175 ;
    RECT 144.71 58.385 144.92 58.455 ;
    RECT 144.71 58.745 144.92 58.815 ;
    RECT 144.71 59.105 144.92 59.175 ;
    RECT 0.4 58.745 0.47 58.815 ;
    RECT 140.93 58.385 141.14 58.455 ;
    RECT 140.93 58.745 141.14 58.815 ;
    RECT 140.93 59.105 141.14 59.175 ;
    RECT 141.39 58.385 141.6 58.455 ;
    RECT 141.39 58.745 141.6 58.815 ;
    RECT 141.39 59.105 141.6 59.175 ;
    RECT 137.61 58.385 137.82 58.455 ;
    RECT 137.61 58.745 137.82 58.815 ;
    RECT 137.61 59.105 137.82 59.175 ;
    RECT 138.07 58.385 138.28 58.455 ;
    RECT 138.07 58.745 138.28 58.815 ;
    RECT 138.07 59.105 138.28 59.175 ;
    RECT 134.29 58.385 134.5 58.455 ;
    RECT 134.29 58.745 134.5 58.815 ;
    RECT 134.29 59.105 134.5 59.175 ;
    RECT 134.75 58.385 134.96 58.455 ;
    RECT 134.75 58.745 134.96 58.815 ;
    RECT 134.75 59.105 134.96 59.175 ;
    RECT 64.57 58.385 64.78 58.455 ;
    RECT 64.57 58.745 64.78 58.815 ;
    RECT 64.57 59.105 64.78 59.175 ;
    RECT 65.03 58.385 65.24 58.455 ;
    RECT 65.03 58.745 65.24 58.815 ;
    RECT 65.03 59.105 65.24 59.175 ;
    RECT 61.25 38.925 61.46 38.995 ;
    RECT 61.25 39.285 61.46 39.355 ;
    RECT 61.25 39.645 61.46 39.715 ;
    RECT 61.71 38.925 61.92 38.995 ;
    RECT 61.71 39.285 61.92 39.355 ;
    RECT 61.71 39.645 61.92 39.715 ;
    RECT 57.93 38.925 58.14 38.995 ;
    RECT 57.93 39.285 58.14 39.355 ;
    RECT 57.93 39.645 58.14 39.715 ;
    RECT 58.39 38.925 58.6 38.995 ;
    RECT 58.39 39.285 58.6 39.355 ;
    RECT 58.39 39.645 58.6 39.715 ;
    RECT 54.61 38.925 54.82 38.995 ;
    RECT 54.61 39.285 54.82 39.355 ;
    RECT 54.61 39.645 54.82 39.715 ;
    RECT 55.07 38.925 55.28 38.995 ;
    RECT 55.07 39.285 55.28 39.355 ;
    RECT 55.07 39.645 55.28 39.715 ;
    RECT 51.29 38.925 51.5 38.995 ;
    RECT 51.29 39.285 51.5 39.355 ;
    RECT 51.29 39.645 51.5 39.715 ;
    RECT 51.75 38.925 51.96 38.995 ;
    RECT 51.75 39.285 51.96 39.355 ;
    RECT 51.75 39.645 51.96 39.715 ;
    RECT 47.97 38.925 48.18 38.995 ;
    RECT 47.97 39.285 48.18 39.355 ;
    RECT 47.97 39.645 48.18 39.715 ;
    RECT 48.43 38.925 48.64 38.995 ;
    RECT 48.43 39.285 48.64 39.355 ;
    RECT 48.43 39.645 48.64 39.715 ;
    RECT 44.65 38.925 44.86 38.995 ;
    RECT 44.65 39.285 44.86 39.355 ;
    RECT 44.65 39.645 44.86 39.715 ;
    RECT 45.11 38.925 45.32 38.995 ;
    RECT 45.11 39.285 45.32 39.355 ;
    RECT 45.11 39.645 45.32 39.715 ;
    RECT 41.33 38.925 41.54 38.995 ;
    RECT 41.33 39.285 41.54 39.355 ;
    RECT 41.33 39.645 41.54 39.715 ;
    RECT 41.79 38.925 42.0 38.995 ;
    RECT 41.79 39.285 42.0 39.355 ;
    RECT 41.79 39.645 42.0 39.715 ;
    RECT 38.01 38.925 38.22 38.995 ;
    RECT 38.01 39.285 38.22 39.355 ;
    RECT 38.01 39.645 38.22 39.715 ;
    RECT 38.47 38.925 38.68 38.995 ;
    RECT 38.47 39.285 38.68 39.355 ;
    RECT 38.47 39.645 38.68 39.715 ;
    RECT 34.69 38.925 34.9 38.995 ;
    RECT 34.69 39.285 34.9 39.355 ;
    RECT 34.69 39.645 34.9 39.715 ;
    RECT 35.15 38.925 35.36 38.995 ;
    RECT 35.15 39.285 35.36 39.355 ;
    RECT 35.15 39.645 35.36 39.715 ;
    RECT 173.945 39.285 174.015 39.355 ;
    RECT 130.97 38.925 131.18 38.995 ;
    RECT 130.97 39.285 131.18 39.355 ;
    RECT 130.97 39.645 131.18 39.715 ;
    RECT 131.43 38.925 131.64 38.995 ;
    RECT 131.43 39.285 131.64 39.355 ;
    RECT 131.43 39.645 131.64 39.715 ;
    RECT 127.65 38.925 127.86 38.995 ;
    RECT 127.65 39.285 127.86 39.355 ;
    RECT 127.65 39.645 127.86 39.715 ;
    RECT 128.11 38.925 128.32 38.995 ;
    RECT 128.11 39.285 128.32 39.355 ;
    RECT 128.11 39.645 128.32 39.715 ;
    RECT 124.33 38.925 124.54 38.995 ;
    RECT 124.33 39.285 124.54 39.355 ;
    RECT 124.33 39.645 124.54 39.715 ;
    RECT 124.79 38.925 125.0 38.995 ;
    RECT 124.79 39.285 125.0 39.355 ;
    RECT 124.79 39.645 125.0 39.715 ;
    RECT 121.01 38.925 121.22 38.995 ;
    RECT 121.01 39.285 121.22 39.355 ;
    RECT 121.01 39.645 121.22 39.715 ;
    RECT 121.47 38.925 121.68 38.995 ;
    RECT 121.47 39.285 121.68 39.355 ;
    RECT 121.47 39.645 121.68 39.715 ;
    RECT 117.69 38.925 117.9 38.995 ;
    RECT 117.69 39.285 117.9 39.355 ;
    RECT 117.69 39.645 117.9 39.715 ;
    RECT 118.15 38.925 118.36 38.995 ;
    RECT 118.15 39.285 118.36 39.355 ;
    RECT 118.15 39.645 118.36 39.715 ;
    RECT 114.37 38.925 114.58 38.995 ;
    RECT 114.37 39.285 114.58 39.355 ;
    RECT 114.37 39.645 114.58 39.715 ;
    RECT 114.83 38.925 115.04 38.995 ;
    RECT 114.83 39.285 115.04 39.355 ;
    RECT 114.83 39.645 115.04 39.715 ;
    RECT 111.05 38.925 111.26 38.995 ;
    RECT 111.05 39.285 111.26 39.355 ;
    RECT 111.05 39.645 111.26 39.715 ;
    RECT 111.51 38.925 111.72 38.995 ;
    RECT 111.51 39.285 111.72 39.355 ;
    RECT 111.51 39.645 111.72 39.715 ;
    RECT 107.73 38.925 107.94 38.995 ;
    RECT 107.73 39.285 107.94 39.355 ;
    RECT 107.73 39.645 107.94 39.715 ;
    RECT 108.19 38.925 108.4 38.995 ;
    RECT 108.19 39.285 108.4 39.355 ;
    RECT 108.19 39.645 108.4 39.715 ;
    RECT 104.41 38.925 104.62 38.995 ;
    RECT 104.41 39.285 104.62 39.355 ;
    RECT 104.41 39.645 104.62 39.715 ;
    RECT 104.87 38.925 105.08 38.995 ;
    RECT 104.87 39.285 105.08 39.355 ;
    RECT 104.87 39.645 105.08 39.715 ;
    RECT 101.09 38.925 101.3 38.995 ;
    RECT 101.09 39.285 101.3 39.355 ;
    RECT 101.09 39.645 101.3 39.715 ;
    RECT 101.55 38.925 101.76 38.995 ;
    RECT 101.55 39.285 101.76 39.355 ;
    RECT 101.55 39.645 101.76 39.715 ;
    RECT 0.4 39.285 0.47 39.355 ;
    RECT 170.81 38.925 171.02 38.995 ;
    RECT 170.81 39.285 171.02 39.355 ;
    RECT 170.81 39.645 171.02 39.715 ;
    RECT 171.27 38.925 171.48 38.995 ;
    RECT 171.27 39.285 171.48 39.355 ;
    RECT 171.27 39.645 171.48 39.715 ;
    RECT 167.49 38.925 167.7 38.995 ;
    RECT 167.49 39.285 167.7 39.355 ;
    RECT 167.49 39.645 167.7 39.715 ;
    RECT 167.95 38.925 168.16 38.995 ;
    RECT 167.95 39.285 168.16 39.355 ;
    RECT 167.95 39.645 168.16 39.715 ;
    RECT 97.77 38.925 97.98 38.995 ;
    RECT 97.77 39.285 97.98 39.355 ;
    RECT 97.77 39.645 97.98 39.715 ;
    RECT 98.23 38.925 98.44 38.995 ;
    RECT 98.23 39.285 98.44 39.355 ;
    RECT 98.23 39.645 98.44 39.715 ;
    RECT 94.45 38.925 94.66 38.995 ;
    RECT 94.45 39.285 94.66 39.355 ;
    RECT 94.45 39.645 94.66 39.715 ;
    RECT 94.91 38.925 95.12 38.995 ;
    RECT 94.91 39.285 95.12 39.355 ;
    RECT 94.91 39.645 95.12 39.715 ;
    RECT 91.13 38.925 91.34 38.995 ;
    RECT 91.13 39.285 91.34 39.355 ;
    RECT 91.13 39.645 91.34 39.715 ;
    RECT 91.59 38.925 91.8 38.995 ;
    RECT 91.59 39.285 91.8 39.355 ;
    RECT 91.59 39.645 91.8 39.715 ;
    RECT 87.81 38.925 88.02 38.995 ;
    RECT 87.81 39.285 88.02 39.355 ;
    RECT 87.81 39.645 88.02 39.715 ;
    RECT 88.27 38.925 88.48 38.995 ;
    RECT 88.27 39.285 88.48 39.355 ;
    RECT 88.27 39.645 88.48 39.715 ;
    RECT 84.49 38.925 84.7 38.995 ;
    RECT 84.49 39.285 84.7 39.355 ;
    RECT 84.49 39.645 84.7 39.715 ;
    RECT 84.95 38.925 85.16 38.995 ;
    RECT 84.95 39.285 85.16 39.355 ;
    RECT 84.95 39.645 85.16 39.715 ;
    RECT 81.17 38.925 81.38 38.995 ;
    RECT 81.17 39.285 81.38 39.355 ;
    RECT 81.17 39.645 81.38 39.715 ;
    RECT 81.63 38.925 81.84 38.995 ;
    RECT 81.63 39.285 81.84 39.355 ;
    RECT 81.63 39.645 81.84 39.715 ;
    RECT 77.85 38.925 78.06 38.995 ;
    RECT 77.85 39.285 78.06 39.355 ;
    RECT 77.85 39.645 78.06 39.715 ;
    RECT 78.31 38.925 78.52 38.995 ;
    RECT 78.31 39.285 78.52 39.355 ;
    RECT 78.31 39.645 78.52 39.715 ;
    RECT 74.53 38.925 74.74 38.995 ;
    RECT 74.53 39.285 74.74 39.355 ;
    RECT 74.53 39.645 74.74 39.715 ;
    RECT 74.99 38.925 75.2 38.995 ;
    RECT 74.99 39.285 75.2 39.355 ;
    RECT 74.99 39.645 75.2 39.715 ;
    RECT 71.21 38.925 71.42 38.995 ;
    RECT 71.21 39.285 71.42 39.355 ;
    RECT 71.21 39.645 71.42 39.715 ;
    RECT 71.67 38.925 71.88 38.995 ;
    RECT 71.67 39.285 71.88 39.355 ;
    RECT 71.67 39.645 71.88 39.715 ;
    RECT 31.37 38.925 31.58 38.995 ;
    RECT 31.37 39.285 31.58 39.355 ;
    RECT 31.37 39.645 31.58 39.715 ;
    RECT 31.83 38.925 32.04 38.995 ;
    RECT 31.83 39.285 32.04 39.355 ;
    RECT 31.83 39.645 32.04 39.715 ;
    RECT 67.89 38.925 68.1 38.995 ;
    RECT 67.89 39.285 68.1 39.355 ;
    RECT 67.89 39.645 68.1 39.715 ;
    RECT 68.35 38.925 68.56 38.995 ;
    RECT 68.35 39.285 68.56 39.355 ;
    RECT 68.35 39.645 68.56 39.715 ;
    RECT 28.05 38.925 28.26 38.995 ;
    RECT 28.05 39.285 28.26 39.355 ;
    RECT 28.05 39.645 28.26 39.715 ;
    RECT 28.51 38.925 28.72 38.995 ;
    RECT 28.51 39.285 28.72 39.355 ;
    RECT 28.51 39.645 28.72 39.715 ;
    RECT 24.73 38.925 24.94 38.995 ;
    RECT 24.73 39.285 24.94 39.355 ;
    RECT 24.73 39.645 24.94 39.715 ;
    RECT 25.19 38.925 25.4 38.995 ;
    RECT 25.19 39.285 25.4 39.355 ;
    RECT 25.19 39.645 25.4 39.715 ;
    RECT 21.41 38.925 21.62 38.995 ;
    RECT 21.41 39.285 21.62 39.355 ;
    RECT 21.41 39.645 21.62 39.715 ;
    RECT 21.87 38.925 22.08 38.995 ;
    RECT 21.87 39.285 22.08 39.355 ;
    RECT 21.87 39.645 22.08 39.715 ;
    RECT 18.09 38.925 18.3 38.995 ;
    RECT 18.09 39.285 18.3 39.355 ;
    RECT 18.09 39.645 18.3 39.715 ;
    RECT 18.55 38.925 18.76 38.995 ;
    RECT 18.55 39.285 18.76 39.355 ;
    RECT 18.55 39.645 18.76 39.715 ;
    RECT 14.77 38.925 14.98 38.995 ;
    RECT 14.77 39.285 14.98 39.355 ;
    RECT 14.77 39.645 14.98 39.715 ;
    RECT 15.23 38.925 15.44 38.995 ;
    RECT 15.23 39.285 15.44 39.355 ;
    RECT 15.23 39.645 15.44 39.715 ;
    RECT 11.45 38.925 11.66 38.995 ;
    RECT 11.45 39.285 11.66 39.355 ;
    RECT 11.45 39.645 11.66 39.715 ;
    RECT 11.91 38.925 12.12 38.995 ;
    RECT 11.91 39.285 12.12 39.355 ;
    RECT 11.91 39.645 12.12 39.715 ;
    RECT 8.13 38.925 8.34 38.995 ;
    RECT 8.13 39.285 8.34 39.355 ;
    RECT 8.13 39.645 8.34 39.715 ;
    RECT 8.59 38.925 8.8 38.995 ;
    RECT 8.59 39.285 8.8 39.355 ;
    RECT 8.59 39.645 8.8 39.715 ;
    RECT 4.81 38.925 5.02 38.995 ;
    RECT 4.81 39.285 5.02 39.355 ;
    RECT 4.81 39.645 5.02 39.715 ;
    RECT 5.27 38.925 5.48 38.995 ;
    RECT 5.27 39.285 5.48 39.355 ;
    RECT 5.27 39.645 5.48 39.715 ;
    RECT 164.17 38.925 164.38 38.995 ;
    RECT 164.17 39.285 164.38 39.355 ;
    RECT 164.17 39.645 164.38 39.715 ;
    RECT 164.63 38.925 164.84 38.995 ;
    RECT 164.63 39.285 164.84 39.355 ;
    RECT 164.63 39.645 164.84 39.715 ;
    RECT 1.49 38.925 1.7 38.995 ;
    RECT 1.49 39.285 1.7 39.355 ;
    RECT 1.49 39.645 1.7 39.715 ;
    RECT 1.95 38.925 2.16 38.995 ;
    RECT 1.95 39.285 2.16 39.355 ;
    RECT 1.95 39.645 2.16 39.715 ;
    RECT 160.85 38.925 161.06 38.995 ;
    RECT 160.85 39.285 161.06 39.355 ;
    RECT 160.85 39.645 161.06 39.715 ;
    RECT 161.31 38.925 161.52 38.995 ;
    RECT 161.31 39.285 161.52 39.355 ;
    RECT 161.31 39.645 161.52 39.715 ;
    RECT 157.53 38.925 157.74 38.995 ;
    RECT 157.53 39.285 157.74 39.355 ;
    RECT 157.53 39.645 157.74 39.715 ;
    RECT 157.99 38.925 158.2 38.995 ;
    RECT 157.99 39.285 158.2 39.355 ;
    RECT 157.99 39.645 158.2 39.715 ;
    RECT 154.21 38.925 154.42 38.995 ;
    RECT 154.21 39.285 154.42 39.355 ;
    RECT 154.21 39.645 154.42 39.715 ;
    RECT 154.67 38.925 154.88 38.995 ;
    RECT 154.67 39.285 154.88 39.355 ;
    RECT 154.67 39.645 154.88 39.715 ;
    RECT 150.89 38.925 151.1 38.995 ;
    RECT 150.89 39.285 151.1 39.355 ;
    RECT 150.89 39.645 151.1 39.715 ;
    RECT 151.35 38.925 151.56 38.995 ;
    RECT 151.35 39.285 151.56 39.355 ;
    RECT 151.35 39.645 151.56 39.715 ;
    RECT 147.57 38.925 147.78 38.995 ;
    RECT 147.57 39.285 147.78 39.355 ;
    RECT 147.57 39.645 147.78 39.715 ;
    RECT 148.03 38.925 148.24 38.995 ;
    RECT 148.03 39.285 148.24 39.355 ;
    RECT 148.03 39.645 148.24 39.715 ;
    RECT 144.25 38.925 144.46 38.995 ;
    RECT 144.25 39.285 144.46 39.355 ;
    RECT 144.25 39.645 144.46 39.715 ;
    RECT 144.71 38.925 144.92 38.995 ;
    RECT 144.71 39.285 144.92 39.355 ;
    RECT 144.71 39.645 144.92 39.715 ;
    RECT 140.93 38.925 141.14 38.995 ;
    RECT 140.93 39.285 141.14 39.355 ;
    RECT 140.93 39.645 141.14 39.715 ;
    RECT 141.39 38.925 141.6 38.995 ;
    RECT 141.39 39.285 141.6 39.355 ;
    RECT 141.39 39.645 141.6 39.715 ;
    RECT 137.61 38.925 137.82 38.995 ;
    RECT 137.61 39.285 137.82 39.355 ;
    RECT 137.61 39.645 137.82 39.715 ;
    RECT 138.07 38.925 138.28 38.995 ;
    RECT 138.07 39.285 138.28 39.355 ;
    RECT 138.07 39.645 138.28 39.715 ;
    RECT 134.29 38.925 134.5 38.995 ;
    RECT 134.29 39.285 134.5 39.355 ;
    RECT 134.29 39.645 134.5 39.715 ;
    RECT 134.75 38.925 134.96 38.995 ;
    RECT 134.75 39.285 134.96 39.355 ;
    RECT 134.75 39.645 134.96 39.715 ;
    RECT 64.57 38.925 64.78 38.995 ;
    RECT 64.57 39.285 64.78 39.355 ;
    RECT 64.57 39.645 64.78 39.715 ;
    RECT 65.03 38.925 65.24 38.995 ;
    RECT 65.03 39.285 65.24 39.355 ;
    RECT 65.03 39.645 65.24 39.715 ;
    RECT 61.25 38.205 61.46 38.275 ;
    RECT 61.25 38.565 61.46 38.635 ;
    RECT 61.25 38.925 61.46 38.995 ;
    RECT 61.71 38.205 61.92 38.275 ;
    RECT 61.71 38.565 61.92 38.635 ;
    RECT 61.71 38.925 61.92 38.995 ;
    RECT 57.93 38.205 58.14 38.275 ;
    RECT 57.93 38.565 58.14 38.635 ;
    RECT 57.93 38.925 58.14 38.995 ;
    RECT 58.39 38.205 58.6 38.275 ;
    RECT 58.39 38.565 58.6 38.635 ;
    RECT 58.39 38.925 58.6 38.995 ;
    RECT 54.61 38.205 54.82 38.275 ;
    RECT 54.61 38.565 54.82 38.635 ;
    RECT 54.61 38.925 54.82 38.995 ;
    RECT 55.07 38.205 55.28 38.275 ;
    RECT 55.07 38.565 55.28 38.635 ;
    RECT 55.07 38.925 55.28 38.995 ;
    RECT 51.29 38.205 51.5 38.275 ;
    RECT 51.29 38.565 51.5 38.635 ;
    RECT 51.29 38.925 51.5 38.995 ;
    RECT 51.75 38.205 51.96 38.275 ;
    RECT 51.75 38.565 51.96 38.635 ;
    RECT 51.75 38.925 51.96 38.995 ;
    RECT 47.97 38.205 48.18 38.275 ;
    RECT 47.97 38.565 48.18 38.635 ;
    RECT 47.97 38.925 48.18 38.995 ;
    RECT 48.43 38.205 48.64 38.275 ;
    RECT 48.43 38.565 48.64 38.635 ;
    RECT 48.43 38.925 48.64 38.995 ;
    RECT 44.65 38.205 44.86 38.275 ;
    RECT 44.65 38.565 44.86 38.635 ;
    RECT 44.65 38.925 44.86 38.995 ;
    RECT 45.11 38.205 45.32 38.275 ;
    RECT 45.11 38.565 45.32 38.635 ;
    RECT 45.11 38.925 45.32 38.995 ;
    RECT 41.33 38.205 41.54 38.275 ;
    RECT 41.33 38.565 41.54 38.635 ;
    RECT 41.33 38.925 41.54 38.995 ;
    RECT 41.79 38.205 42.0 38.275 ;
    RECT 41.79 38.565 42.0 38.635 ;
    RECT 41.79 38.925 42.0 38.995 ;
    RECT 38.01 38.205 38.22 38.275 ;
    RECT 38.01 38.565 38.22 38.635 ;
    RECT 38.01 38.925 38.22 38.995 ;
    RECT 38.47 38.205 38.68 38.275 ;
    RECT 38.47 38.565 38.68 38.635 ;
    RECT 38.47 38.925 38.68 38.995 ;
    RECT 34.69 38.205 34.9 38.275 ;
    RECT 34.69 38.565 34.9 38.635 ;
    RECT 34.69 38.925 34.9 38.995 ;
    RECT 35.15 38.205 35.36 38.275 ;
    RECT 35.15 38.565 35.36 38.635 ;
    RECT 35.15 38.925 35.36 38.995 ;
    RECT 173.945 38.565 174.015 38.635 ;
    RECT 130.97 38.205 131.18 38.275 ;
    RECT 130.97 38.565 131.18 38.635 ;
    RECT 130.97 38.925 131.18 38.995 ;
    RECT 131.43 38.205 131.64 38.275 ;
    RECT 131.43 38.565 131.64 38.635 ;
    RECT 131.43 38.925 131.64 38.995 ;
    RECT 127.65 38.205 127.86 38.275 ;
    RECT 127.65 38.565 127.86 38.635 ;
    RECT 127.65 38.925 127.86 38.995 ;
    RECT 128.11 38.205 128.32 38.275 ;
    RECT 128.11 38.565 128.32 38.635 ;
    RECT 128.11 38.925 128.32 38.995 ;
    RECT 124.33 38.205 124.54 38.275 ;
    RECT 124.33 38.565 124.54 38.635 ;
    RECT 124.33 38.925 124.54 38.995 ;
    RECT 124.79 38.205 125.0 38.275 ;
    RECT 124.79 38.565 125.0 38.635 ;
    RECT 124.79 38.925 125.0 38.995 ;
    RECT 121.01 38.205 121.22 38.275 ;
    RECT 121.01 38.565 121.22 38.635 ;
    RECT 121.01 38.925 121.22 38.995 ;
    RECT 121.47 38.205 121.68 38.275 ;
    RECT 121.47 38.565 121.68 38.635 ;
    RECT 121.47 38.925 121.68 38.995 ;
    RECT 117.69 38.205 117.9 38.275 ;
    RECT 117.69 38.565 117.9 38.635 ;
    RECT 117.69 38.925 117.9 38.995 ;
    RECT 118.15 38.205 118.36 38.275 ;
    RECT 118.15 38.565 118.36 38.635 ;
    RECT 118.15 38.925 118.36 38.995 ;
    RECT 114.37 38.205 114.58 38.275 ;
    RECT 114.37 38.565 114.58 38.635 ;
    RECT 114.37 38.925 114.58 38.995 ;
    RECT 114.83 38.205 115.04 38.275 ;
    RECT 114.83 38.565 115.04 38.635 ;
    RECT 114.83 38.925 115.04 38.995 ;
    RECT 111.05 38.205 111.26 38.275 ;
    RECT 111.05 38.565 111.26 38.635 ;
    RECT 111.05 38.925 111.26 38.995 ;
    RECT 111.51 38.205 111.72 38.275 ;
    RECT 111.51 38.565 111.72 38.635 ;
    RECT 111.51 38.925 111.72 38.995 ;
    RECT 107.73 38.205 107.94 38.275 ;
    RECT 107.73 38.565 107.94 38.635 ;
    RECT 107.73 38.925 107.94 38.995 ;
    RECT 108.19 38.205 108.4 38.275 ;
    RECT 108.19 38.565 108.4 38.635 ;
    RECT 108.19 38.925 108.4 38.995 ;
    RECT 104.41 38.205 104.62 38.275 ;
    RECT 104.41 38.565 104.62 38.635 ;
    RECT 104.41 38.925 104.62 38.995 ;
    RECT 104.87 38.205 105.08 38.275 ;
    RECT 104.87 38.565 105.08 38.635 ;
    RECT 104.87 38.925 105.08 38.995 ;
    RECT 101.09 38.205 101.3 38.275 ;
    RECT 101.09 38.565 101.3 38.635 ;
    RECT 101.09 38.925 101.3 38.995 ;
    RECT 101.55 38.205 101.76 38.275 ;
    RECT 101.55 38.565 101.76 38.635 ;
    RECT 101.55 38.925 101.76 38.995 ;
    RECT 0.4 38.565 0.47 38.635 ;
    RECT 170.81 38.205 171.02 38.275 ;
    RECT 170.81 38.565 171.02 38.635 ;
    RECT 170.81 38.925 171.02 38.995 ;
    RECT 171.27 38.205 171.48 38.275 ;
    RECT 171.27 38.565 171.48 38.635 ;
    RECT 171.27 38.925 171.48 38.995 ;
    RECT 167.49 38.205 167.7 38.275 ;
    RECT 167.49 38.565 167.7 38.635 ;
    RECT 167.49 38.925 167.7 38.995 ;
    RECT 167.95 38.205 168.16 38.275 ;
    RECT 167.95 38.565 168.16 38.635 ;
    RECT 167.95 38.925 168.16 38.995 ;
    RECT 97.77 38.205 97.98 38.275 ;
    RECT 97.77 38.565 97.98 38.635 ;
    RECT 97.77 38.925 97.98 38.995 ;
    RECT 98.23 38.205 98.44 38.275 ;
    RECT 98.23 38.565 98.44 38.635 ;
    RECT 98.23 38.925 98.44 38.995 ;
    RECT 94.45 38.205 94.66 38.275 ;
    RECT 94.45 38.565 94.66 38.635 ;
    RECT 94.45 38.925 94.66 38.995 ;
    RECT 94.91 38.205 95.12 38.275 ;
    RECT 94.91 38.565 95.12 38.635 ;
    RECT 94.91 38.925 95.12 38.995 ;
    RECT 91.13 38.205 91.34 38.275 ;
    RECT 91.13 38.565 91.34 38.635 ;
    RECT 91.13 38.925 91.34 38.995 ;
    RECT 91.59 38.205 91.8 38.275 ;
    RECT 91.59 38.565 91.8 38.635 ;
    RECT 91.59 38.925 91.8 38.995 ;
    RECT 87.81 38.205 88.02 38.275 ;
    RECT 87.81 38.565 88.02 38.635 ;
    RECT 87.81 38.925 88.02 38.995 ;
    RECT 88.27 38.205 88.48 38.275 ;
    RECT 88.27 38.565 88.48 38.635 ;
    RECT 88.27 38.925 88.48 38.995 ;
    RECT 84.49 38.205 84.7 38.275 ;
    RECT 84.49 38.565 84.7 38.635 ;
    RECT 84.49 38.925 84.7 38.995 ;
    RECT 84.95 38.205 85.16 38.275 ;
    RECT 84.95 38.565 85.16 38.635 ;
    RECT 84.95 38.925 85.16 38.995 ;
    RECT 81.17 38.205 81.38 38.275 ;
    RECT 81.17 38.565 81.38 38.635 ;
    RECT 81.17 38.925 81.38 38.995 ;
    RECT 81.63 38.205 81.84 38.275 ;
    RECT 81.63 38.565 81.84 38.635 ;
    RECT 81.63 38.925 81.84 38.995 ;
    RECT 77.85 38.205 78.06 38.275 ;
    RECT 77.85 38.565 78.06 38.635 ;
    RECT 77.85 38.925 78.06 38.995 ;
    RECT 78.31 38.205 78.52 38.275 ;
    RECT 78.31 38.565 78.52 38.635 ;
    RECT 78.31 38.925 78.52 38.995 ;
    RECT 74.53 38.205 74.74 38.275 ;
    RECT 74.53 38.565 74.74 38.635 ;
    RECT 74.53 38.925 74.74 38.995 ;
    RECT 74.99 38.205 75.2 38.275 ;
    RECT 74.99 38.565 75.2 38.635 ;
    RECT 74.99 38.925 75.2 38.995 ;
    RECT 71.21 38.205 71.42 38.275 ;
    RECT 71.21 38.565 71.42 38.635 ;
    RECT 71.21 38.925 71.42 38.995 ;
    RECT 71.67 38.205 71.88 38.275 ;
    RECT 71.67 38.565 71.88 38.635 ;
    RECT 71.67 38.925 71.88 38.995 ;
    RECT 31.37 38.205 31.58 38.275 ;
    RECT 31.37 38.565 31.58 38.635 ;
    RECT 31.37 38.925 31.58 38.995 ;
    RECT 31.83 38.205 32.04 38.275 ;
    RECT 31.83 38.565 32.04 38.635 ;
    RECT 31.83 38.925 32.04 38.995 ;
    RECT 67.89 38.205 68.1 38.275 ;
    RECT 67.89 38.565 68.1 38.635 ;
    RECT 67.89 38.925 68.1 38.995 ;
    RECT 68.35 38.205 68.56 38.275 ;
    RECT 68.35 38.565 68.56 38.635 ;
    RECT 68.35 38.925 68.56 38.995 ;
    RECT 28.05 38.205 28.26 38.275 ;
    RECT 28.05 38.565 28.26 38.635 ;
    RECT 28.05 38.925 28.26 38.995 ;
    RECT 28.51 38.205 28.72 38.275 ;
    RECT 28.51 38.565 28.72 38.635 ;
    RECT 28.51 38.925 28.72 38.995 ;
    RECT 24.73 38.205 24.94 38.275 ;
    RECT 24.73 38.565 24.94 38.635 ;
    RECT 24.73 38.925 24.94 38.995 ;
    RECT 25.19 38.205 25.4 38.275 ;
    RECT 25.19 38.565 25.4 38.635 ;
    RECT 25.19 38.925 25.4 38.995 ;
    RECT 21.41 38.205 21.62 38.275 ;
    RECT 21.41 38.565 21.62 38.635 ;
    RECT 21.41 38.925 21.62 38.995 ;
    RECT 21.87 38.205 22.08 38.275 ;
    RECT 21.87 38.565 22.08 38.635 ;
    RECT 21.87 38.925 22.08 38.995 ;
    RECT 18.09 38.205 18.3 38.275 ;
    RECT 18.09 38.565 18.3 38.635 ;
    RECT 18.09 38.925 18.3 38.995 ;
    RECT 18.55 38.205 18.76 38.275 ;
    RECT 18.55 38.565 18.76 38.635 ;
    RECT 18.55 38.925 18.76 38.995 ;
    RECT 14.77 38.205 14.98 38.275 ;
    RECT 14.77 38.565 14.98 38.635 ;
    RECT 14.77 38.925 14.98 38.995 ;
    RECT 15.23 38.205 15.44 38.275 ;
    RECT 15.23 38.565 15.44 38.635 ;
    RECT 15.23 38.925 15.44 38.995 ;
    RECT 11.45 38.205 11.66 38.275 ;
    RECT 11.45 38.565 11.66 38.635 ;
    RECT 11.45 38.925 11.66 38.995 ;
    RECT 11.91 38.205 12.12 38.275 ;
    RECT 11.91 38.565 12.12 38.635 ;
    RECT 11.91 38.925 12.12 38.995 ;
    RECT 8.13 38.205 8.34 38.275 ;
    RECT 8.13 38.565 8.34 38.635 ;
    RECT 8.13 38.925 8.34 38.995 ;
    RECT 8.59 38.205 8.8 38.275 ;
    RECT 8.59 38.565 8.8 38.635 ;
    RECT 8.59 38.925 8.8 38.995 ;
    RECT 4.81 38.205 5.02 38.275 ;
    RECT 4.81 38.565 5.02 38.635 ;
    RECT 4.81 38.925 5.02 38.995 ;
    RECT 5.27 38.205 5.48 38.275 ;
    RECT 5.27 38.565 5.48 38.635 ;
    RECT 5.27 38.925 5.48 38.995 ;
    RECT 164.17 38.205 164.38 38.275 ;
    RECT 164.17 38.565 164.38 38.635 ;
    RECT 164.17 38.925 164.38 38.995 ;
    RECT 164.63 38.205 164.84 38.275 ;
    RECT 164.63 38.565 164.84 38.635 ;
    RECT 164.63 38.925 164.84 38.995 ;
    RECT 1.49 38.205 1.7 38.275 ;
    RECT 1.49 38.565 1.7 38.635 ;
    RECT 1.49 38.925 1.7 38.995 ;
    RECT 1.95 38.205 2.16 38.275 ;
    RECT 1.95 38.565 2.16 38.635 ;
    RECT 1.95 38.925 2.16 38.995 ;
    RECT 160.85 38.205 161.06 38.275 ;
    RECT 160.85 38.565 161.06 38.635 ;
    RECT 160.85 38.925 161.06 38.995 ;
    RECT 161.31 38.205 161.52 38.275 ;
    RECT 161.31 38.565 161.52 38.635 ;
    RECT 161.31 38.925 161.52 38.995 ;
    RECT 157.53 38.205 157.74 38.275 ;
    RECT 157.53 38.565 157.74 38.635 ;
    RECT 157.53 38.925 157.74 38.995 ;
    RECT 157.99 38.205 158.2 38.275 ;
    RECT 157.99 38.565 158.2 38.635 ;
    RECT 157.99 38.925 158.2 38.995 ;
    RECT 154.21 38.205 154.42 38.275 ;
    RECT 154.21 38.565 154.42 38.635 ;
    RECT 154.21 38.925 154.42 38.995 ;
    RECT 154.67 38.205 154.88 38.275 ;
    RECT 154.67 38.565 154.88 38.635 ;
    RECT 154.67 38.925 154.88 38.995 ;
    RECT 150.89 38.205 151.1 38.275 ;
    RECT 150.89 38.565 151.1 38.635 ;
    RECT 150.89 38.925 151.1 38.995 ;
    RECT 151.35 38.205 151.56 38.275 ;
    RECT 151.35 38.565 151.56 38.635 ;
    RECT 151.35 38.925 151.56 38.995 ;
    RECT 147.57 38.205 147.78 38.275 ;
    RECT 147.57 38.565 147.78 38.635 ;
    RECT 147.57 38.925 147.78 38.995 ;
    RECT 148.03 38.205 148.24 38.275 ;
    RECT 148.03 38.565 148.24 38.635 ;
    RECT 148.03 38.925 148.24 38.995 ;
    RECT 144.25 38.205 144.46 38.275 ;
    RECT 144.25 38.565 144.46 38.635 ;
    RECT 144.25 38.925 144.46 38.995 ;
    RECT 144.71 38.205 144.92 38.275 ;
    RECT 144.71 38.565 144.92 38.635 ;
    RECT 144.71 38.925 144.92 38.995 ;
    RECT 140.93 38.205 141.14 38.275 ;
    RECT 140.93 38.565 141.14 38.635 ;
    RECT 140.93 38.925 141.14 38.995 ;
    RECT 141.39 38.205 141.6 38.275 ;
    RECT 141.39 38.565 141.6 38.635 ;
    RECT 141.39 38.925 141.6 38.995 ;
    RECT 137.61 38.205 137.82 38.275 ;
    RECT 137.61 38.565 137.82 38.635 ;
    RECT 137.61 38.925 137.82 38.995 ;
    RECT 138.07 38.205 138.28 38.275 ;
    RECT 138.07 38.565 138.28 38.635 ;
    RECT 138.07 38.925 138.28 38.995 ;
    RECT 134.29 38.205 134.5 38.275 ;
    RECT 134.29 38.565 134.5 38.635 ;
    RECT 134.29 38.925 134.5 38.995 ;
    RECT 134.75 38.205 134.96 38.275 ;
    RECT 134.75 38.565 134.96 38.635 ;
    RECT 134.75 38.925 134.96 38.995 ;
    RECT 64.57 38.205 64.78 38.275 ;
    RECT 64.57 38.565 64.78 38.635 ;
    RECT 64.57 38.925 64.78 38.995 ;
    RECT 65.03 38.205 65.24 38.275 ;
    RECT 65.03 38.565 65.24 38.635 ;
    RECT 65.03 38.925 65.24 38.995 ;
    RECT 61.25 37.485 61.46 37.555 ;
    RECT 61.25 37.845 61.46 37.915 ;
    RECT 61.25 38.205 61.46 38.275 ;
    RECT 61.71 37.485 61.92 37.555 ;
    RECT 61.71 37.845 61.92 37.915 ;
    RECT 61.71 38.205 61.92 38.275 ;
    RECT 57.93 37.485 58.14 37.555 ;
    RECT 57.93 37.845 58.14 37.915 ;
    RECT 57.93 38.205 58.14 38.275 ;
    RECT 58.39 37.485 58.6 37.555 ;
    RECT 58.39 37.845 58.6 37.915 ;
    RECT 58.39 38.205 58.6 38.275 ;
    RECT 54.61 37.485 54.82 37.555 ;
    RECT 54.61 37.845 54.82 37.915 ;
    RECT 54.61 38.205 54.82 38.275 ;
    RECT 55.07 37.485 55.28 37.555 ;
    RECT 55.07 37.845 55.28 37.915 ;
    RECT 55.07 38.205 55.28 38.275 ;
    RECT 51.29 37.485 51.5 37.555 ;
    RECT 51.29 37.845 51.5 37.915 ;
    RECT 51.29 38.205 51.5 38.275 ;
    RECT 51.75 37.485 51.96 37.555 ;
    RECT 51.75 37.845 51.96 37.915 ;
    RECT 51.75 38.205 51.96 38.275 ;
    RECT 47.97 37.485 48.18 37.555 ;
    RECT 47.97 37.845 48.18 37.915 ;
    RECT 47.97 38.205 48.18 38.275 ;
    RECT 48.43 37.485 48.64 37.555 ;
    RECT 48.43 37.845 48.64 37.915 ;
    RECT 48.43 38.205 48.64 38.275 ;
    RECT 44.65 37.485 44.86 37.555 ;
    RECT 44.65 37.845 44.86 37.915 ;
    RECT 44.65 38.205 44.86 38.275 ;
    RECT 45.11 37.485 45.32 37.555 ;
    RECT 45.11 37.845 45.32 37.915 ;
    RECT 45.11 38.205 45.32 38.275 ;
    RECT 41.33 37.485 41.54 37.555 ;
    RECT 41.33 37.845 41.54 37.915 ;
    RECT 41.33 38.205 41.54 38.275 ;
    RECT 41.79 37.485 42.0 37.555 ;
    RECT 41.79 37.845 42.0 37.915 ;
    RECT 41.79 38.205 42.0 38.275 ;
    RECT 38.01 37.485 38.22 37.555 ;
    RECT 38.01 37.845 38.22 37.915 ;
    RECT 38.01 38.205 38.22 38.275 ;
    RECT 38.47 37.485 38.68 37.555 ;
    RECT 38.47 37.845 38.68 37.915 ;
    RECT 38.47 38.205 38.68 38.275 ;
    RECT 34.69 37.485 34.9 37.555 ;
    RECT 34.69 37.845 34.9 37.915 ;
    RECT 34.69 38.205 34.9 38.275 ;
    RECT 35.15 37.485 35.36 37.555 ;
    RECT 35.15 37.845 35.36 37.915 ;
    RECT 35.15 38.205 35.36 38.275 ;
    RECT 173.945 37.845 174.015 37.915 ;
    RECT 130.97 37.485 131.18 37.555 ;
    RECT 130.97 37.845 131.18 37.915 ;
    RECT 130.97 38.205 131.18 38.275 ;
    RECT 131.43 37.485 131.64 37.555 ;
    RECT 131.43 37.845 131.64 37.915 ;
    RECT 131.43 38.205 131.64 38.275 ;
    RECT 127.65 37.485 127.86 37.555 ;
    RECT 127.65 37.845 127.86 37.915 ;
    RECT 127.65 38.205 127.86 38.275 ;
    RECT 128.11 37.485 128.32 37.555 ;
    RECT 128.11 37.845 128.32 37.915 ;
    RECT 128.11 38.205 128.32 38.275 ;
    RECT 124.33 37.485 124.54 37.555 ;
    RECT 124.33 37.845 124.54 37.915 ;
    RECT 124.33 38.205 124.54 38.275 ;
    RECT 124.79 37.485 125.0 37.555 ;
    RECT 124.79 37.845 125.0 37.915 ;
    RECT 124.79 38.205 125.0 38.275 ;
    RECT 121.01 37.485 121.22 37.555 ;
    RECT 121.01 37.845 121.22 37.915 ;
    RECT 121.01 38.205 121.22 38.275 ;
    RECT 121.47 37.485 121.68 37.555 ;
    RECT 121.47 37.845 121.68 37.915 ;
    RECT 121.47 38.205 121.68 38.275 ;
    RECT 117.69 37.485 117.9 37.555 ;
    RECT 117.69 37.845 117.9 37.915 ;
    RECT 117.69 38.205 117.9 38.275 ;
    RECT 118.15 37.485 118.36 37.555 ;
    RECT 118.15 37.845 118.36 37.915 ;
    RECT 118.15 38.205 118.36 38.275 ;
    RECT 114.37 37.485 114.58 37.555 ;
    RECT 114.37 37.845 114.58 37.915 ;
    RECT 114.37 38.205 114.58 38.275 ;
    RECT 114.83 37.485 115.04 37.555 ;
    RECT 114.83 37.845 115.04 37.915 ;
    RECT 114.83 38.205 115.04 38.275 ;
    RECT 111.05 37.485 111.26 37.555 ;
    RECT 111.05 37.845 111.26 37.915 ;
    RECT 111.05 38.205 111.26 38.275 ;
    RECT 111.51 37.485 111.72 37.555 ;
    RECT 111.51 37.845 111.72 37.915 ;
    RECT 111.51 38.205 111.72 38.275 ;
    RECT 107.73 37.485 107.94 37.555 ;
    RECT 107.73 37.845 107.94 37.915 ;
    RECT 107.73 38.205 107.94 38.275 ;
    RECT 108.19 37.485 108.4 37.555 ;
    RECT 108.19 37.845 108.4 37.915 ;
    RECT 108.19 38.205 108.4 38.275 ;
    RECT 104.41 37.485 104.62 37.555 ;
    RECT 104.41 37.845 104.62 37.915 ;
    RECT 104.41 38.205 104.62 38.275 ;
    RECT 104.87 37.485 105.08 37.555 ;
    RECT 104.87 37.845 105.08 37.915 ;
    RECT 104.87 38.205 105.08 38.275 ;
    RECT 101.09 37.485 101.3 37.555 ;
    RECT 101.09 37.845 101.3 37.915 ;
    RECT 101.09 38.205 101.3 38.275 ;
    RECT 101.55 37.485 101.76 37.555 ;
    RECT 101.55 37.845 101.76 37.915 ;
    RECT 101.55 38.205 101.76 38.275 ;
    RECT 0.4 37.845 0.47 37.915 ;
    RECT 170.81 37.485 171.02 37.555 ;
    RECT 170.81 37.845 171.02 37.915 ;
    RECT 170.81 38.205 171.02 38.275 ;
    RECT 171.27 37.485 171.48 37.555 ;
    RECT 171.27 37.845 171.48 37.915 ;
    RECT 171.27 38.205 171.48 38.275 ;
    RECT 167.49 37.485 167.7 37.555 ;
    RECT 167.49 37.845 167.7 37.915 ;
    RECT 167.49 38.205 167.7 38.275 ;
    RECT 167.95 37.485 168.16 37.555 ;
    RECT 167.95 37.845 168.16 37.915 ;
    RECT 167.95 38.205 168.16 38.275 ;
    RECT 97.77 37.485 97.98 37.555 ;
    RECT 97.77 37.845 97.98 37.915 ;
    RECT 97.77 38.205 97.98 38.275 ;
    RECT 98.23 37.485 98.44 37.555 ;
    RECT 98.23 37.845 98.44 37.915 ;
    RECT 98.23 38.205 98.44 38.275 ;
    RECT 94.45 37.485 94.66 37.555 ;
    RECT 94.45 37.845 94.66 37.915 ;
    RECT 94.45 38.205 94.66 38.275 ;
    RECT 94.91 37.485 95.12 37.555 ;
    RECT 94.91 37.845 95.12 37.915 ;
    RECT 94.91 38.205 95.12 38.275 ;
    RECT 91.13 37.485 91.34 37.555 ;
    RECT 91.13 37.845 91.34 37.915 ;
    RECT 91.13 38.205 91.34 38.275 ;
    RECT 91.59 37.485 91.8 37.555 ;
    RECT 91.59 37.845 91.8 37.915 ;
    RECT 91.59 38.205 91.8 38.275 ;
    RECT 87.81 37.485 88.02 37.555 ;
    RECT 87.81 37.845 88.02 37.915 ;
    RECT 87.81 38.205 88.02 38.275 ;
    RECT 88.27 37.485 88.48 37.555 ;
    RECT 88.27 37.845 88.48 37.915 ;
    RECT 88.27 38.205 88.48 38.275 ;
    RECT 84.49 37.485 84.7 37.555 ;
    RECT 84.49 37.845 84.7 37.915 ;
    RECT 84.49 38.205 84.7 38.275 ;
    RECT 84.95 37.485 85.16 37.555 ;
    RECT 84.95 37.845 85.16 37.915 ;
    RECT 84.95 38.205 85.16 38.275 ;
    RECT 81.17 37.485 81.38 37.555 ;
    RECT 81.17 37.845 81.38 37.915 ;
    RECT 81.17 38.205 81.38 38.275 ;
    RECT 81.63 37.485 81.84 37.555 ;
    RECT 81.63 37.845 81.84 37.915 ;
    RECT 81.63 38.205 81.84 38.275 ;
    RECT 77.85 37.485 78.06 37.555 ;
    RECT 77.85 37.845 78.06 37.915 ;
    RECT 77.85 38.205 78.06 38.275 ;
    RECT 78.31 37.485 78.52 37.555 ;
    RECT 78.31 37.845 78.52 37.915 ;
    RECT 78.31 38.205 78.52 38.275 ;
    RECT 74.53 37.485 74.74 37.555 ;
    RECT 74.53 37.845 74.74 37.915 ;
    RECT 74.53 38.205 74.74 38.275 ;
    RECT 74.99 37.485 75.2 37.555 ;
    RECT 74.99 37.845 75.2 37.915 ;
    RECT 74.99 38.205 75.2 38.275 ;
    RECT 71.21 37.485 71.42 37.555 ;
    RECT 71.21 37.845 71.42 37.915 ;
    RECT 71.21 38.205 71.42 38.275 ;
    RECT 71.67 37.485 71.88 37.555 ;
    RECT 71.67 37.845 71.88 37.915 ;
    RECT 71.67 38.205 71.88 38.275 ;
    RECT 31.37 37.485 31.58 37.555 ;
    RECT 31.37 37.845 31.58 37.915 ;
    RECT 31.37 38.205 31.58 38.275 ;
    RECT 31.83 37.485 32.04 37.555 ;
    RECT 31.83 37.845 32.04 37.915 ;
    RECT 31.83 38.205 32.04 38.275 ;
    RECT 67.89 37.485 68.1 37.555 ;
    RECT 67.89 37.845 68.1 37.915 ;
    RECT 67.89 38.205 68.1 38.275 ;
    RECT 68.35 37.485 68.56 37.555 ;
    RECT 68.35 37.845 68.56 37.915 ;
    RECT 68.35 38.205 68.56 38.275 ;
    RECT 28.05 37.485 28.26 37.555 ;
    RECT 28.05 37.845 28.26 37.915 ;
    RECT 28.05 38.205 28.26 38.275 ;
    RECT 28.51 37.485 28.72 37.555 ;
    RECT 28.51 37.845 28.72 37.915 ;
    RECT 28.51 38.205 28.72 38.275 ;
    RECT 24.73 37.485 24.94 37.555 ;
    RECT 24.73 37.845 24.94 37.915 ;
    RECT 24.73 38.205 24.94 38.275 ;
    RECT 25.19 37.485 25.4 37.555 ;
    RECT 25.19 37.845 25.4 37.915 ;
    RECT 25.19 38.205 25.4 38.275 ;
    RECT 21.41 37.485 21.62 37.555 ;
    RECT 21.41 37.845 21.62 37.915 ;
    RECT 21.41 38.205 21.62 38.275 ;
    RECT 21.87 37.485 22.08 37.555 ;
    RECT 21.87 37.845 22.08 37.915 ;
    RECT 21.87 38.205 22.08 38.275 ;
    RECT 18.09 37.485 18.3 37.555 ;
    RECT 18.09 37.845 18.3 37.915 ;
    RECT 18.09 38.205 18.3 38.275 ;
    RECT 18.55 37.485 18.76 37.555 ;
    RECT 18.55 37.845 18.76 37.915 ;
    RECT 18.55 38.205 18.76 38.275 ;
    RECT 14.77 37.485 14.98 37.555 ;
    RECT 14.77 37.845 14.98 37.915 ;
    RECT 14.77 38.205 14.98 38.275 ;
    RECT 15.23 37.485 15.44 37.555 ;
    RECT 15.23 37.845 15.44 37.915 ;
    RECT 15.23 38.205 15.44 38.275 ;
    RECT 11.45 37.485 11.66 37.555 ;
    RECT 11.45 37.845 11.66 37.915 ;
    RECT 11.45 38.205 11.66 38.275 ;
    RECT 11.91 37.485 12.12 37.555 ;
    RECT 11.91 37.845 12.12 37.915 ;
    RECT 11.91 38.205 12.12 38.275 ;
    RECT 8.13 37.485 8.34 37.555 ;
    RECT 8.13 37.845 8.34 37.915 ;
    RECT 8.13 38.205 8.34 38.275 ;
    RECT 8.59 37.485 8.8 37.555 ;
    RECT 8.59 37.845 8.8 37.915 ;
    RECT 8.59 38.205 8.8 38.275 ;
    RECT 4.81 37.485 5.02 37.555 ;
    RECT 4.81 37.845 5.02 37.915 ;
    RECT 4.81 38.205 5.02 38.275 ;
    RECT 5.27 37.485 5.48 37.555 ;
    RECT 5.27 37.845 5.48 37.915 ;
    RECT 5.27 38.205 5.48 38.275 ;
    RECT 164.17 37.485 164.38 37.555 ;
    RECT 164.17 37.845 164.38 37.915 ;
    RECT 164.17 38.205 164.38 38.275 ;
    RECT 164.63 37.485 164.84 37.555 ;
    RECT 164.63 37.845 164.84 37.915 ;
    RECT 164.63 38.205 164.84 38.275 ;
    RECT 1.49 37.485 1.7 37.555 ;
    RECT 1.49 37.845 1.7 37.915 ;
    RECT 1.49 38.205 1.7 38.275 ;
    RECT 1.95 37.485 2.16 37.555 ;
    RECT 1.95 37.845 2.16 37.915 ;
    RECT 1.95 38.205 2.16 38.275 ;
    RECT 160.85 37.485 161.06 37.555 ;
    RECT 160.85 37.845 161.06 37.915 ;
    RECT 160.85 38.205 161.06 38.275 ;
    RECT 161.31 37.485 161.52 37.555 ;
    RECT 161.31 37.845 161.52 37.915 ;
    RECT 161.31 38.205 161.52 38.275 ;
    RECT 157.53 37.485 157.74 37.555 ;
    RECT 157.53 37.845 157.74 37.915 ;
    RECT 157.53 38.205 157.74 38.275 ;
    RECT 157.99 37.485 158.2 37.555 ;
    RECT 157.99 37.845 158.2 37.915 ;
    RECT 157.99 38.205 158.2 38.275 ;
    RECT 154.21 37.485 154.42 37.555 ;
    RECT 154.21 37.845 154.42 37.915 ;
    RECT 154.21 38.205 154.42 38.275 ;
    RECT 154.67 37.485 154.88 37.555 ;
    RECT 154.67 37.845 154.88 37.915 ;
    RECT 154.67 38.205 154.88 38.275 ;
    RECT 150.89 37.485 151.1 37.555 ;
    RECT 150.89 37.845 151.1 37.915 ;
    RECT 150.89 38.205 151.1 38.275 ;
    RECT 151.35 37.485 151.56 37.555 ;
    RECT 151.35 37.845 151.56 37.915 ;
    RECT 151.35 38.205 151.56 38.275 ;
    RECT 147.57 37.485 147.78 37.555 ;
    RECT 147.57 37.845 147.78 37.915 ;
    RECT 147.57 38.205 147.78 38.275 ;
    RECT 148.03 37.485 148.24 37.555 ;
    RECT 148.03 37.845 148.24 37.915 ;
    RECT 148.03 38.205 148.24 38.275 ;
    RECT 144.25 37.485 144.46 37.555 ;
    RECT 144.25 37.845 144.46 37.915 ;
    RECT 144.25 38.205 144.46 38.275 ;
    RECT 144.71 37.485 144.92 37.555 ;
    RECT 144.71 37.845 144.92 37.915 ;
    RECT 144.71 38.205 144.92 38.275 ;
    RECT 140.93 37.485 141.14 37.555 ;
    RECT 140.93 37.845 141.14 37.915 ;
    RECT 140.93 38.205 141.14 38.275 ;
    RECT 141.39 37.485 141.6 37.555 ;
    RECT 141.39 37.845 141.6 37.915 ;
    RECT 141.39 38.205 141.6 38.275 ;
    RECT 137.61 37.485 137.82 37.555 ;
    RECT 137.61 37.845 137.82 37.915 ;
    RECT 137.61 38.205 137.82 38.275 ;
    RECT 138.07 37.485 138.28 37.555 ;
    RECT 138.07 37.845 138.28 37.915 ;
    RECT 138.07 38.205 138.28 38.275 ;
    RECT 134.29 37.485 134.5 37.555 ;
    RECT 134.29 37.845 134.5 37.915 ;
    RECT 134.29 38.205 134.5 38.275 ;
    RECT 134.75 37.485 134.96 37.555 ;
    RECT 134.75 37.845 134.96 37.915 ;
    RECT 134.75 38.205 134.96 38.275 ;
    RECT 64.57 37.485 64.78 37.555 ;
    RECT 64.57 37.845 64.78 37.915 ;
    RECT 64.57 38.205 64.78 38.275 ;
    RECT 65.03 37.485 65.24 37.555 ;
    RECT 65.03 37.845 65.24 37.915 ;
    RECT 65.03 38.205 65.24 38.275 ;
    RECT 61.25 36.765 61.46 36.835 ;
    RECT 61.25 37.125 61.46 37.195 ;
    RECT 61.25 37.485 61.46 37.555 ;
    RECT 61.71 36.765 61.92 36.835 ;
    RECT 61.71 37.125 61.92 37.195 ;
    RECT 61.71 37.485 61.92 37.555 ;
    RECT 57.93 36.765 58.14 36.835 ;
    RECT 57.93 37.125 58.14 37.195 ;
    RECT 57.93 37.485 58.14 37.555 ;
    RECT 58.39 36.765 58.6 36.835 ;
    RECT 58.39 37.125 58.6 37.195 ;
    RECT 58.39 37.485 58.6 37.555 ;
    RECT 54.61 36.765 54.82 36.835 ;
    RECT 54.61 37.125 54.82 37.195 ;
    RECT 54.61 37.485 54.82 37.555 ;
    RECT 55.07 36.765 55.28 36.835 ;
    RECT 55.07 37.125 55.28 37.195 ;
    RECT 55.07 37.485 55.28 37.555 ;
    RECT 51.29 36.765 51.5 36.835 ;
    RECT 51.29 37.125 51.5 37.195 ;
    RECT 51.29 37.485 51.5 37.555 ;
    RECT 51.75 36.765 51.96 36.835 ;
    RECT 51.75 37.125 51.96 37.195 ;
    RECT 51.75 37.485 51.96 37.555 ;
    RECT 47.97 36.765 48.18 36.835 ;
    RECT 47.97 37.125 48.18 37.195 ;
    RECT 47.97 37.485 48.18 37.555 ;
    RECT 48.43 36.765 48.64 36.835 ;
    RECT 48.43 37.125 48.64 37.195 ;
    RECT 48.43 37.485 48.64 37.555 ;
    RECT 44.65 36.765 44.86 36.835 ;
    RECT 44.65 37.125 44.86 37.195 ;
    RECT 44.65 37.485 44.86 37.555 ;
    RECT 45.11 36.765 45.32 36.835 ;
    RECT 45.11 37.125 45.32 37.195 ;
    RECT 45.11 37.485 45.32 37.555 ;
    RECT 41.33 36.765 41.54 36.835 ;
    RECT 41.33 37.125 41.54 37.195 ;
    RECT 41.33 37.485 41.54 37.555 ;
    RECT 41.79 36.765 42.0 36.835 ;
    RECT 41.79 37.125 42.0 37.195 ;
    RECT 41.79 37.485 42.0 37.555 ;
    RECT 38.01 36.765 38.22 36.835 ;
    RECT 38.01 37.125 38.22 37.195 ;
    RECT 38.01 37.485 38.22 37.555 ;
    RECT 38.47 36.765 38.68 36.835 ;
    RECT 38.47 37.125 38.68 37.195 ;
    RECT 38.47 37.485 38.68 37.555 ;
    RECT 34.69 36.765 34.9 36.835 ;
    RECT 34.69 37.125 34.9 37.195 ;
    RECT 34.69 37.485 34.9 37.555 ;
    RECT 35.15 36.765 35.36 36.835 ;
    RECT 35.15 37.125 35.36 37.195 ;
    RECT 35.15 37.485 35.36 37.555 ;
    RECT 173.945 37.125 174.015 37.195 ;
    RECT 130.97 36.765 131.18 36.835 ;
    RECT 130.97 37.125 131.18 37.195 ;
    RECT 130.97 37.485 131.18 37.555 ;
    RECT 131.43 36.765 131.64 36.835 ;
    RECT 131.43 37.125 131.64 37.195 ;
    RECT 131.43 37.485 131.64 37.555 ;
    RECT 127.65 36.765 127.86 36.835 ;
    RECT 127.65 37.125 127.86 37.195 ;
    RECT 127.65 37.485 127.86 37.555 ;
    RECT 128.11 36.765 128.32 36.835 ;
    RECT 128.11 37.125 128.32 37.195 ;
    RECT 128.11 37.485 128.32 37.555 ;
    RECT 124.33 36.765 124.54 36.835 ;
    RECT 124.33 37.125 124.54 37.195 ;
    RECT 124.33 37.485 124.54 37.555 ;
    RECT 124.79 36.765 125.0 36.835 ;
    RECT 124.79 37.125 125.0 37.195 ;
    RECT 124.79 37.485 125.0 37.555 ;
    RECT 121.01 36.765 121.22 36.835 ;
    RECT 121.01 37.125 121.22 37.195 ;
    RECT 121.01 37.485 121.22 37.555 ;
    RECT 121.47 36.765 121.68 36.835 ;
    RECT 121.47 37.125 121.68 37.195 ;
    RECT 121.47 37.485 121.68 37.555 ;
    RECT 117.69 36.765 117.9 36.835 ;
    RECT 117.69 37.125 117.9 37.195 ;
    RECT 117.69 37.485 117.9 37.555 ;
    RECT 118.15 36.765 118.36 36.835 ;
    RECT 118.15 37.125 118.36 37.195 ;
    RECT 118.15 37.485 118.36 37.555 ;
    RECT 114.37 36.765 114.58 36.835 ;
    RECT 114.37 37.125 114.58 37.195 ;
    RECT 114.37 37.485 114.58 37.555 ;
    RECT 114.83 36.765 115.04 36.835 ;
    RECT 114.83 37.125 115.04 37.195 ;
    RECT 114.83 37.485 115.04 37.555 ;
    RECT 111.05 36.765 111.26 36.835 ;
    RECT 111.05 37.125 111.26 37.195 ;
    RECT 111.05 37.485 111.26 37.555 ;
    RECT 111.51 36.765 111.72 36.835 ;
    RECT 111.51 37.125 111.72 37.195 ;
    RECT 111.51 37.485 111.72 37.555 ;
    RECT 107.73 36.765 107.94 36.835 ;
    RECT 107.73 37.125 107.94 37.195 ;
    RECT 107.73 37.485 107.94 37.555 ;
    RECT 108.19 36.765 108.4 36.835 ;
    RECT 108.19 37.125 108.4 37.195 ;
    RECT 108.19 37.485 108.4 37.555 ;
    RECT 104.41 36.765 104.62 36.835 ;
    RECT 104.41 37.125 104.62 37.195 ;
    RECT 104.41 37.485 104.62 37.555 ;
    RECT 104.87 36.765 105.08 36.835 ;
    RECT 104.87 37.125 105.08 37.195 ;
    RECT 104.87 37.485 105.08 37.555 ;
    RECT 101.09 36.765 101.3 36.835 ;
    RECT 101.09 37.125 101.3 37.195 ;
    RECT 101.09 37.485 101.3 37.555 ;
    RECT 101.55 36.765 101.76 36.835 ;
    RECT 101.55 37.125 101.76 37.195 ;
    RECT 101.55 37.485 101.76 37.555 ;
    RECT 0.4 37.125 0.47 37.195 ;
    RECT 170.81 36.765 171.02 36.835 ;
    RECT 170.81 37.125 171.02 37.195 ;
    RECT 170.81 37.485 171.02 37.555 ;
    RECT 171.27 36.765 171.48 36.835 ;
    RECT 171.27 37.125 171.48 37.195 ;
    RECT 171.27 37.485 171.48 37.555 ;
    RECT 167.49 36.765 167.7 36.835 ;
    RECT 167.49 37.125 167.7 37.195 ;
    RECT 167.49 37.485 167.7 37.555 ;
    RECT 167.95 36.765 168.16 36.835 ;
    RECT 167.95 37.125 168.16 37.195 ;
    RECT 167.95 37.485 168.16 37.555 ;
    RECT 97.77 36.765 97.98 36.835 ;
    RECT 97.77 37.125 97.98 37.195 ;
    RECT 97.77 37.485 97.98 37.555 ;
    RECT 98.23 36.765 98.44 36.835 ;
    RECT 98.23 37.125 98.44 37.195 ;
    RECT 98.23 37.485 98.44 37.555 ;
    RECT 94.45 36.765 94.66 36.835 ;
    RECT 94.45 37.125 94.66 37.195 ;
    RECT 94.45 37.485 94.66 37.555 ;
    RECT 94.91 36.765 95.12 36.835 ;
    RECT 94.91 37.125 95.12 37.195 ;
    RECT 94.91 37.485 95.12 37.555 ;
    RECT 91.13 36.765 91.34 36.835 ;
    RECT 91.13 37.125 91.34 37.195 ;
    RECT 91.13 37.485 91.34 37.555 ;
    RECT 91.59 36.765 91.8 36.835 ;
    RECT 91.59 37.125 91.8 37.195 ;
    RECT 91.59 37.485 91.8 37.555 ;
    RECT 87.81 36.765 88.02 36.835 ;
    RECT 87.81 37.125 88.02 37.195 ;
    RECT 87.81 37.485 88.02 37.555 ;
    RECT 88.27 36.765 88.48 36.835 ;
    RECT 88.27 37.125 88.48 37.195 ;
    RECT 88.27 37.485 88.48 37.555 ;
    RECT 84.49 36.765 84.7 36.835 ;
    RECT 84.49 37.125 84.7 37.195 ;
    RECT 84.49 37.485 84.7 37.555 ;
    RECT 84.95 36.765 85.16 36.835 ;
    RECT 84.95 37.125 85.16 37.195 ;
    RECT 84.95 37.485 85.16 37.555 ;
    RECT 81.17 36.765 81.38 36.835 ;
    RECT 81.17 37.125 81.38 37.195 ;
    RECT 81.17 37.485 81.38 37.555 ;
    RECT 81.63 36.765 81.84 36.835 ;
    RECT 81.63 37.125 81.84 37.195 ;
    RECT 81.63 37.485 81.84 37.555 ;
    RECT 77.85 36.765 78.06 36.835 ;
    RECT 77.85 37.125 78.06 37.195 ;
    RECT 77.85 37.485 78.06 37.555 ;
    RECT 78.31 36.765 78.52 36.835 ;
    RECT 78.31 37.125 78.52 37.195 ;
    RECT 78.31 37.485 78.52 37.555 ;
    RECT 74.53 36.765 74.74 36.835 ;
    RECT 74.53 37.125 74.74 37.195 ;
    RECT 74.53 37.485 74.74 37.555 ;
    RECT 74.99 36.765 75.2 36.835 ;
    RECT 74.99 37.125 75.2 37.195 ;
    RECT 74.99 37.485 75.2 37.555 ;
    RECT 71.21 36.765 71.42 36.835 ;
    RECT 71.21 37.125 71.42 37.195 ;
    RECT 71.21 37.485 71.42 37.555 ;
    RECT 71.67 36.765 71.88 36.835 ;
    RECT 71.67 37.125 71.88 37.195 ;
    RECT 71.67 37.485 71.88 37.555 ;
    RECT 31.37 36.765 31.58 36.835 ;
    RECT 31.37 37.125 31.58 37.195 ;
    RECT 31.37 37.485 31.58 37.555 ;
    RECT 31.83 36.765 32.04 36.835 ;
    RECT 31.83 37.125 32.04 37.195 ;
    RECT 31.83 37.485 32.04 37.555 ;
    RECT 67.89 36.765 68.1 36.835 ;
    RECT 67.89 37.125 68.1 37.195 ;
    RECT 67.89 37.485 68.1 37.555 ;
    RECT 68.35 36.765 68.56 36.835 ;
    RECT 68.35 37.125 68.56 37.195 ;
    RECT 68.35 37.485 68.56 37.555 ;
    RECT 28.05 36.765 28.26 36.835 ;
    RECT 28.05 37.125 28.26 37.195 ;
    RECT 28.05 37.485 28.26 37.555 ;
    RECT 28.51 36.765 28.72 36.835 ;
    RECT 28.51 37.125 28.72 37.195 ;
    RECT 28.51 37.485 28.72 37.555 ;
    RECT 24.73 36.765 24.94 36.835 ;
    RECT 24.73 37.125 24.94 37.195 ;
    RECT 24.73 37.485 24.94 37.555 ;
    RECT 25.19 36.765 25.4 36.835 ;
    RECT 25.19 37.125 25.4 37.195 ;
    RECT 25.19 37.485 25.4 37.555 ;
    RECT 21.41 36.765 21.62 36.835 ;
    RECT 21.41 37.125 21.62 37.195 ;
    RECT 21.41 37.485 21.62 37.555 ;
    RECT 21.87 36.765 22.08 36.835 ;
    RECT 21.87 37.125 22.08 37.195 ;
    RECT 21.87 37.485 22.08 37.555 ;
    RECT 18.09 36.765 18.3 36.835 ;
    RECT 18.09 37.125 18.3 37.195 ;
    RECT 18.09 37.485 18.3 37.555 ;
    RECT 18.55 36.765 18.76 36.835 ;
    RECT 18.55 37.125 18.76 37.195 ;
    RECT 18.55 37.485 18.76 37.555 ;
    RECT 14.77 36.765 14.98 36.835 ;
    RECT 14.77 37.125 14.98 37.195 ;
    RECT 14.77 37.485 14.98 37.555 ;
    RECT 15.23 36.765 15.44 36.835 ;
    RECT 15.23 37.125 15.44 37.195 ;
    RECT 15.23 37.485 15.44 37.555 ;
    RECT 11.45 36.765 11.66 36.835 ;
    RECT 11.45 37.125 11.66 37.195 ;
    RECT 11.45 37.485 11.66 37.555 ;
    RECT 11.91 36.765 12.12 36.835 ;
    RECT 11.91 37.125 12.12 37.195 ;
    RECT 11.91 37.485 12.12 37.555 ;
    RECT 8.13 36.765 8.34 36.835 ;
    RECT 8.13 37.125 8.34 37.195 ;
    RECT 8.13 37.485 8.34 37.555 ;
    RECT 8.59 36.765 8.8 36.835 ;
    RECT 8.59 37.125 8.8 37.195 ;
    RECT 8.59 37.485 8.8 37.555 ;
    RECT 4.81 36.765 5.02 36.835 ;
    RECT 4.81 37.125 5.02 37.195 ;
    RECT 4.81 37.485 5.02 37.555 ;
    RECT 5.27 36.765 5.48 36.835 ;
    RECT 5.27 37.125 5.48 37.195 ;
    RECT 5.27 37.485 5.48 37.555 ;
    RECT 164.17 36.765 164.38 36.835 ;
    RECT 164.17 37.125 164.38 37.195 ;
    RECT 164.17 37.485 164.38 37.555 ;
    RECT 164.63 36.765 164.84 36.835 ;
    RECT 164.63 37.125 164.84 37.195 ;
    RECT 164.63 37.485 164.84 37.555 ;
    RECT 1.49 36.765 1.7 36.835 ;
    RECT 1.49 37.125 1.7 37.195 ;
    RECT 1.49 37.485 1.7 37.555 ;
    RECT 1.95 36.765 2.16 36.835 ;
    RECT 1.95 37.125 2.16 37.195 ;
    RECT 1.95 37.485 2.16 37.555 ;
    RECT 160.85 36.765 161.06 36.835 ;
    RECT 160.85 37.125 161.06 37.195 ;
    RECT 160.85 37.485 161.06 37.555 ;
    RECT 161.31 36.765 161.52 36.835 ;
    RECT 161.31 37.125 161.52 37.195 ;
    RECT 161.31 37.485 161.52 37.555 ;
    RECT 157.53 36.765 157.74 36.835 ;
    RECT 157.53 37.125 157.74 37.195 ;
    RECT 157.53 37.485 157.74 37.555 ;
    RECT 157.99 36.765 158.2 36.835 ;
    RECT 157.99 37.125 158.2 37.195 ;
    RECT 157.99 37.485 158.2 37.555 ;
    RECT 154.21 36.765 154.42 36.835 ;
    RECT 154.21 37.125 154.42 37.195 ;
    RECT 154.21 37.485 154.42 37.555 ;
    RECT 154.67 36.765 154.88 36.835 ;
    RECT 154.67 37.125 154.88 37.195 ;
    RECT 154.67 37.485 154.88 37.555 ;
    RECT 150.89 36.765 151.1 36.835 ;
    RECT 150.89 37.125 151.1 37.195 ;
    RECT 150.89 37.485 151.1 37.555 ;
    RECT 151.35 36.765 151.56 36.835 ;
    RECT 151.35 37.125 151.56 37.195 ;
    RECT 151.35 37.485 151.56 37.555 ;
    RECT 147.57 36.765 147.78 36.835 ;
    RECT 147.57 37.125 147.78 37.195 ;
    RECT 147.57 37.485 147.78 37.555 ;
    RECT 148.03 36.765 148.24 36.835 ;
    RECT 148.03 37.125 148.24 37.195 ;
    RECT 148.03 37.485 148.24 37.555 ;
    RECT 144.25 36.765 144.46 36.835 ;
    RECT 144.25 37.125 144.46 37.195 ;
    RECT 144.25 37.485 144.46 37.555 ;
    RECT 144.71 36.765 144.92 36.835 ;
    RECT 144.71 37.125 144.92 37.195 ;
    RECT 144.71 37.485 144.92 37.555 ;
    RECT 140.93 36.765 141.14 36.835 ;
    RECT 140.93 37.125 141.14 37.195 ;
    RECT 140.93 37.485 141.14 37.555 ;
    RECT 141.39 36.765 141.6 36.835 ;
    RECT 141.39 37.125 141.6 37.195 ;
    RECT 141.39 37.485 141.6 37.555 ;
    RECT 137.61 36.765 137.82 36.835 ;
    RECT 137.61 37.125 137.82 37.195 ;
    RECT 137.61 37.485 137.82 37.555 ;
    RECT 138.07 36.765 138.28 36.835 ;
    RECT 138.07 37.125 138.28 37.195 ;
    RECT 138.07 37.485 138.28 37.555 ;
    RECT 134.29 36.765 134.5 36.835 ;
    RECT 134.29 37.125 134.5 37.195 ;
    RECT 134.29 37.485 134.5 37.555 ;
    RECT 134.75 36.765 134.96 36.835 ;
    RECT 134.75 37.125 134.96 37.195 ;
    RECT 134.75 37.485 134.96 37.555 ;
    RECT 64.57 36.765 64.78 36.835 ;
    RECT 64.57 37.125 64.78 37.195 ;
    RECT 64.57 37.485 64.78 37.555 ;
    RECT 65.03 36.765 65.24 36.835 ;
    RECT 65.03 37.125 65.24 37.195 ;
    RECT 65.03 37.485 65.24 37.555 ;
    RECT 61.25 36.045 61.46 36.115 ;
    RECT 61.25 36.405 61.46 36.475 ;
    RECT 61.25 36.765 61.46 36.835 ;
    RECT 61.71 36.045 61.92 36.115 ;
    RECT 61.71 36.405 61.92 36.475 ;
    RECT 61.71 36.765 61.92 36.835 ;
    RECT 57.93 36.045 58.14 36.115 ;
    RECT 57.93 36.405 58.14 36.475 ;
    RECT 57.93 36.765 58.14 36.835 ;
    RECT 58.39 36.045 58.6 36.115 ;
    RECT 58.39 36.405 58.6 36.475 ;
    RECT 58.39 36.765 58.6 36.835 ;
    RECT 54.61 36.045 54.82 36.115 ;
    RECT 54.61 36.405 54.82 36.475 ;
    RECT 54.61 36.765 54.82 36.835 ;
    RECT 55.07 36.045 55.28 36.115 ;
    RECT 55.07 36.405 55.28 36.475 ;
    RECT 55.07 36.765 55.28 36.835 ;
    RECT 51.29 36.045 51.5 36.115 ;
    RECT 51.29 36.405 51.5 36.475 ;
    RECT 51.29 36.765 51.5 36.835 ;
    RECT 51.75 36.045 51.96 36.115 ;
    RECT 51.75 36.405 51.96 36.475 ;
    RECT 51.75 36.765 51.96 36.835 ;
    RECT 47.97 36.045 48.18 36.115 ;
    RECT 47.97 36.405 48.18 36.475 ;
    RECT 47.97 36.765 48.18 36.835 ;
    RECT 48.43 36.045 48.64 36.115 ;
    RECT 48.43 36.405 48.64 36.475 ;
    RECT 48.43 36.765 48.64 36.835 ;
    RECT 44.65 36.045 44.86 36.115 ;
    RECT 44.65 36.405 44.86 36.475 ;
    RECT 44.65 36.765 44.86 36.835 ;
    RECT 45.11 36.045 45.32 36.115 ;
    RECT 45.11 36.405 45.32 36.475 ;
    RECT 45.11 36.765 45.32 36.835 ;
    RECT 41.33 36.045 41.54 36.115 ;
    RECT 41.33 36.405 41.54 36.475 ;
    RECT 41.33 36.765 41.54 36.835 ;
    RECT 41.79 36.045 42.0 36.115 ;
    RECT 41.79 36.405 42.0 36.475 ;
    RECT 41.79 36.765 42.0 36.835 ;
    RECT 38.01 36.045 38.22 36.115 ;
    RECT 38.01 36.405 38.22 36.475 ;
    RECT 38.01 36.765 38.22 36.835 ;
    RECT 38.47 36.045 38.68 36.115 ;
    RECT 38.47 36.405 38.68 36.475 ;
    RECT 38.47 36.765 38.68 36.835 ;
    RECT 34.69 36.045 34.9 36.115 ;
    RECT 34.69 36.405 34.9 36.475 ;
    RECT 34.69 36.765 34.9 36.835 ;
    RECT 35.15 36.045 35.36 36.115 ;
    RECT 35.15 36.405 35.36 36.475 ;
    RECT 35.15 36.765 35.36 36.835 ;
    RECT 173.945 36.405 174.015 36.475 ;
    RECT 130.97 36.045 131.18 36.115 ;
    RECT 130.97 36.405 131.18 36.475 ;
    RECT 130.97 36.765 131.18 36.835 ;
    RECT 131.43 36.045 131.64 36.115 ;
    RECT 131.43 36.405 131.64 36.475 ;
    RECT 131.43 36.765 131.64 36.835 ;
    RECT 127.65 36.045 127.86 36.115 ;
    RECT 127.65 36.405 127.86 36.475 ;
    RECT 127.65 36.765 127.86 36.835 ;
    RECT 128.11 36.045 128.32 36.115 ;
    RECT 128.11 36.405 128.32 36.475 ;
    RECT 128.11 36.765 128.32 36.835 ;
    RECT 124.33 36.045 124.54 36.115 ;
    RECT 124.33 36.405 124.54 36.475 ;
    RECT 124.33 36.765 124.54 36.835 ;
    RECT 124.79 36.045 125.0 36.115 ;
    RECT 124.79 36.405 125.0 36.475 ;
    RECT 124.79 36.765 125.0 36.835 ;
    RECT 121.01 36.045 121.22 36.115 ;
    RECT 121.01 36.405 121.22 36.475 ;
    RECT 121.01 36.765 121.22 36.835 ;
    RECT 121.47 36.045 121.68 36.115 ;
    RECT 121.47 36.405 121.68 36.475 ;
    RECT 121.47 36.765 121.68 36.835 ;
    RECT 117.69 36.045 117.9 36.115 ;
    RECT 117.69 36.405 117.9 36.475 ;
    RECT 117.69 36.765 117.9 36.835 ;
    RECT 118.15 36.045 118.36 36.115 ;
    RECT 118.15 36.405 118.36 36.475 ;
    RECT 118.15 36.765 118.36 36.835 ;
    RECT 114.37 36.045 114.58 36.115 ;
    RECT 114.37 36.405 114.58 36.475 ;
    RECT 114.37 36.765 114.58 36.835 ;
    RECT 114.83 36.045 115.04 36.115 ;
    RECT 114.83 36.405 115.04 36.475 ;
    RECT 114.83 36.765 115.04 36.835 ;
    RECT 111.05 36.045 111.26 36.115 ;
    RECT 111.05 36.405 111.26 36.475 ;
    RECT 111.05 36.765 111.26 36.835 ;
    RECT 111.51 36.045 111.72 36.115 ;
    RECT 111.51 36.405 111.72 36.475 ;
    RECT 111.51 36.765 111.72 36.835 ;
    RECT 107.73 36.045 107.94 36.115 ;
    RECT 107.73 36.405 107.94 36.475 ;
    RECT 107.73 36.765 107.94 36.835 ;
    RECT 108.19 36.045 108.4 36.115 ;
    RECT 108.19 36.405 108.4 36.475 ;
    RECT 108.19 36.765 108.4 36.835 ;
    RECT 104.41 36.045 104.62 36.115 ;
    RECT 104.41 36.405 104.62 36.475 ;
    RECT 104.41 36.765 104.62 36.835 ;
    RECT 104.87 36.045 105.08 36.115 ;
    RECT 104.87 36.405 105.08 36.475 ;
    RECT 104.87 36.765 105.08 36.835 ;
    RECT 101.09 36.045 101.3 36.115 ;
    RECT 101.09 36.405 101.3 36.475 ;
    RECT 101.09 36.765 101.3 36.835 ;
    RECT 101.55 36.045 101.76 36.115 ;
    RECT 101.55 36.405 101.76 36.475 ;
    RECT 101.55 36.765 101.76 36.835 ;
    RECT 0.4 36.405 0.47 36.475 ;
    RECT 170.81 36.045 171.02 36.115 ;
    RECT 170.81 36.405 171.02 36.475 ;
    RECT 170.81 36.765 171.02 36.835 ;
    RECT 171.27 36.045 171.48 36.115 ;
    RECT 171.27 36.405 171.48 36.475 ;
    RECT 171.27 36.765 171.48 36.835 ;
    RECT 167.49 36.045 167.7 36.115 ;
    RECT 167.49 36.405 167.7 36.475 ;
    RECT 167.49 36.765 167.7 36.835 ;
    RECT 167.95 36.045 168.16 36.115 ;
    RECT 167.95 36.405 168.16 36.475 ;
    RECT 167.95 36.765 168.16 36.835 ;
    RECT 97.77 36.045 97.98 36.115 ;
    RECT 97.77 36.405 97.98 36.475 ;
    RECT 97.77 36.765 97.98 36.835 ;
    RECT 98.23 36.045 98.44 36.115 ;
    RECT 98.23 36.405 98.44 36.475 ;
    RECT 98.23 36.765 98.44 36.835 ;
    RECT 94.45 36.045 94.66 36.115 ;
    RECT 94.45 36.405 94.66 36.475 ;
    RECT 94.45 36.765 94.66 36.835 ;
    RECT 94.91 36.045 95.12 36.115 ;
    RECT 94.91 36.405 95.12 36.475 ;
    RECT 94.91 36.765 95.12 36.835 ;
    RECT 91.13 36.045 91.34 36.115 ;
    RECT 91.13 36.405 91.34 36.475 ;
    RECT 91.13 36.765 91.34 36.835 ;
    RECT 91.59 36.045 91.8 36.115 ;
    RECT 91.59 36.405 91.8 36.475 ;
    RECT 91.59 36.765 91.8 36.835 ;
    RECT 87.81 36.045 88.02 36.115 ;
    RECT 87.81 36.405 88.02 36.475 ;
    RECT 87.81 36.765 88.02 36.835 ;
    RECT 88.27 36.045 88.48 36.115 ;
    RECT 88.27 36.405 88.48 36.475 ;
    RECT 88.27 36.765 88.48 36.835 ;
    RECT 84.49 36.045 84.7 36.115 ;
    RECT 84.49 36.405 84.7 36.475 ;
    RECT 84.49 36.765 84.7 36.835 ;
    RECT 84.95 36.045 85.16 36.115 ;
    RECT 84.95 36.405 85.16 36.475 ;
    RECT 84.95 36.765 85.16 36.835 ;
    RECT 81.17 36.045 81.38 36.115 ;
    RECT 81.17 36.405 81.38 36.475 ;
    RECT 81.17 36.765 81.38 36.835 ;
    RECT 81.63 36.045 81.84 36.115 ;
    RECT 81.63 36.405 81.84 36.475 ;
    RECT 81.63 36.765 81.84 36.835 ;
    RECT 77.85 36.045 78.06 36.115 ;
    RECT 77.85 36.405 78.06 36.475 ;
    RECT 77.85 36.765 78.06 36.835 ;
    RECT 78.31 36.045 78.52 36.115 ;
    RECT 78.31 36.405 78.52 36.475 ;
    RECT 78.31 36.765 78.52 36.835 ;
    RECT 74.53 36.045 74.74 36.115 ;
    RECT 74.53 36.405 74.74 36.475 ;
    RECT 74.53 36.765 74.74 36.835 ;
    RECT 74.99 36.045 75.2 36.115 ;
    RECT 74.99 36.405 75.2 36.475 ;
    RECT 74.99 36.765 75.2 36.835 ;
    RECT 71.21 36.045 71.42 36.115 ;
    RECT 71.21 36.405 71.42 36.475 ;
    RECT 71.21 36.765 71.42 36.835 ;
    RECT 71.67 36.045 71.88 36.115 ;
    RECT 71.67 36.405 71.88 36.475 ;
    RECT 71.67 36.765 71.88 36.835 ;
    RECT 31.37 36.045 31.58 36.115 ;
    RECT 31.37 36.405 31.58 36.475 ;
    RECT 31.37 36.765 31.58 36.835 ;
    RECT 31.83 36.045 32.04 36.115 ;
    RECT 31.83 36.405 32.04 36.475 ;
    RECT 31.83 36.765 32.04 36.835 ;
    RECT 67.89 36.045 68.1 36.115 ;
    RECT 67.89 36.405 68.1 36.475 ;
    RECT 67.89 36.765 68.1 36.835 ;
    RECT 68.35 36.045 68.56 36.115 ;
    RECT 68.35 36.405 68.56 36.475 ;
    RECT 68.35 36.765 68.56 36.835 ;
    RECT 28.05 36.045 28.26 36.115 ;
    RECT 28.05 36.405 28.26 36.475 ;
    RECT 28.05 36.765 28.26 36.835 ;
    RECT 28.51 36.045 28.72 36.115 ;
    RECT 28.51 36.405 28.72 36.475 ;
    RECT 28.51 36.765 28.72 36.835 ;
    RECT 24.73 36.045 24.94 36.115 ;
    RECT 24.73 36.405 24.94 36.475 ;
    RECT 24.73 36.765 24.94 36.835 ;
    RECT 25.19 36.045 25.4 36.115 ;
    RECT 25.19 36.405 25.4 36.475 ;
    RECT 25.19 36.765 25.4 36.835 ;
    RECT 21.41 36.045 21.62 36.115 ;
    RECT 21.41 36.405 21.62 36.475 ;
    RECT 21.41 36.765 21.62 36.835 ;
    RECT 21.87 36.045 22.08 36.115 ;
    RECT 21.87 36.405 22.08 36.475 ;
    RECT 21.87 36.765 22.08 36.835 ;
    RECT 18.09 36.045 18.3 36.115 ;
    RECT 18.09 36.405 18.3 36.475 ;
    RECT 18.09 36.765 18.3 36.835 ;
    RECT 18.55 36.045 18.76 36.115 ;
    RECT 18.55 36.405 18.76 36.475 ;
    RECT 18.55 36.765 18.76 36.835 ;
    RECT 14.77 36.045 14.98 36.115 ;
    RECT 14.77 36.405 14.98 36.475 ;
    RECT 14.77 36.765 14.98 36.835 ;
    RECT 15.23 36.045 15.44 36.115 ;
    RECT 15.23 36.405 15.44 36.475 ;
    RECT 15.23 36.765 15.44 36.835 ;
    RECT 11.45 36.045 11.66 36.115 ;
    RECT 11.45 36.405 11.66 36.475 ;
    RECT 11.45 36.765 11.66 36.835 ;
    RECT 11.91 36.045 12.12 36.115 ;
    RECT 11.91 36.405 12.12 36.475 ;
    RECT 11.91 36.765 12.12 36.835 ;
    RECT 8.13 36.045 8.34 36.115 ;
    RECT 8.13 36.405 8.34 36.475 ;
    RECT 8.13 36.765 8.34 36.835 ;
    RECT 8.59 36.045 8.8 36.115 ;
    RECT 8.59 36.405 8.8 36.475 ;
    RECT 8.59 36.765 8.8 36.835 ;
    RECT 4.81 36.045 5.02 36.115 ;
    RECT 4.81 36.405 5.02 36.475 ;
    RECT 4.81 36.765 5.02 36.835 ;
    RECT 5.27 36.045 5.48 36.115 ;
    RECT 5.27 36.405 5.48 36.475 ;
    RECT 5.27 36.765 5.48 36.835 ;
    RECT 164.17 36.045 164.38 36.115 ;
    RECT 164.17 36.405 164.38 36.475 ;
    RECT 164.17 36.765 164.38 36.835 ;
    RECT 164.63 36.045 164.84 36.115 ;
    RECT 164.63 36.405 164.84 36.475 ;
    RECT 164.63 36.765 164.84 36.835 ;
    RECT 1.49 36.045 1.7 36.115 ;
    RECT 1.49 36.405 1.7 36.475 ;
    RECT 1.49 36.765 1.7 36.835 ;
    RECT 1.95 36.045 2.16 36.115 ;
    RECT 1.95 36.405 2.16 36.475 ;
    RECT 1.95 36.765 2.16 36.835 ;
    RECT 160.85 36.045 161.06 36.115 ;
    RECT 160.85 36.405 161.06 36.475 ;
    RECT 160.85 36.765 161.06 36.835 ;
    RECT 161.31 36.045 161.52 36.115 ;
    RECT 161.31 36.405 161.52 36.475 ;
    RECT 161.31 36.765 161.52 36.835 ;
    RECT 157.53 36.045 157.74 36.115 ;
    RECT 157.53 36.405 157.74 36.475 ;
    RECT 157.53 36.765 157.74 36.835 ;
    RECT 157.99 36.045 158.2 36.115 ;
    RECT 157.99 36.405 158.2 36.475 ;
    RECT 157.99 36.765 158.2 36.835 ;
    RECT 154.21 36.045 154.42 36.115 ;
    RECT 154.21 36.405 154.42 36.475 ;
    RECT 154.21 36.765 154.42 36.835 ;
    RECT 154.67 36.045 154.88 36.115 ;
    RECT 154.67 36.405 154.88 36.475 ;
    RECT 154.67 36.765 154.88 36.835 ;
    RECT 150.89 36.045 151.1 36.115 ;
    RECT 150.89 36.405 151.1 36.475 ;
    RECT 150.89 36.765 151.1 36.835 ;
    RECT 151.35 36.045 151.56 36.115 ;
    RECT 151.35 36.405 151.56 36.475 ;
    RECT 151.35 36.765 151.56 36.835 ;
    RECT 147.57 36.045 147.78 36.115 ;
    RECT 147.57 36.405 147.78 36.475 ;
    RECT 147.57 36.765 147.78 36.835 ;
    RECT 148.03 36.045 148.24 36.115 ;
    RECT 148.03 36.405 148.24 36.475 ;
    RECT 148.03 36.765 148.24 36.835 ;
    RECT 144.25 36.045 144.46 36.115 ;
    RECT 144.25 36.405 144.46 36.475 ;
    RECT 144.25 36.765 144.46 36.835 ;
    RECT 144.71 36.045 144.92 36.115 ;
    RECT 144.71 36.405 144.92 36.475 ;
    RECT 144.71 36.765 144.92 36.835 ;
    RECT 140.93 36.045 141.14 36.115 ;
    RECT 140.93 36.405 141.14 36.475 ;
    RECT 140.93 36.765 141.14 36.835 ;
    RECT 141.39 36.045 141.6 36.115 ;
    RECT 141.39 36.405 141.6 36.475 ;
    RECT 141.39 36.765 141.6 36.835 ;
    RECT 137.61 36.045 137.82 36.115 ;
    RECT 137.61 36.405 137.82 36.475 ;
    RECT 137.61 36.765 137.82 36.835 ;
    RECT 138.07 36.045 138.28 36.115 ;
    RECT 138.07 36.405 138.28 36.475 ;
    RECT 138.07 36.765 138.28 36.835 ;
    RECT 134.29 36.045 134.5 36.115 ;
    RECT 134.29 36.405 134.5 36.475 ;
    RECT 134.29 36.765 134.5 36.835 ;
    RECT 134.75 36.045 134.96 36.115 ;
    RECT 134.75 36.405 134.96 36.475 ;
    RECT 134.75 36.765 134.96 36.835 ;
    RECT 64.57 36.045 64.78 36.115 ;
    RECT 64.57 36.405 64.78 36.475 ;
    RECT 64.57 36.765 64.78 36.835 ;
    RECT 65.03 36.045 65.24 36.115 ;
    RECT 65.03 36.405 65.24 36.475 ;
    RECT 65.03 36.765 65.24 36.835 ;
    RECT 61.25 33.165 61.46 33.235 ;
    RECT 61.25 33.525 61.46 33.595 ;
    RECT 61.25 33.885 61.46 33.955 ;
    RECT 61.71 33.165 61.92 33.235 ;
    RECT 61.71 33.525 61.92 33.595 ;
    RECT 61.71 33.885 61.92 33.955 ;
    RECT 57.93 33.165 58.14 33.235 ;
    RECT 57.93 33.525 58.14 33.595 ;
    RECT 57.93 33.885 58.14 33.955 ;
    RECT 58.39 33.165 58.6 33.235 ;
    RECT 58.39 33.525 58.6 33.595 ;
    RECT 58.39 33.885 58.6 33.955 ;
    RECT 54.61 33.165 54.82 33.235 ;
    RECT 54.61 33.525 54.82 33.595 ;
    RECT 54.61 33.885 54.82 33.955 ;
    RECT 55.07 33.165 55.28 33.235 ;
    RECT 55.07 33.525 55.28 33.595 ;
    RECT 55.07 33.885 55.28 33.955 ;
    RECT 51.29 33.165 51.5 33.235 ;
    RECT 51.29 33.525 51.5 33.595 ;
    RECT 51.29 33.885 51.5 33.955 ;
    RECT 51.75 33.165 51.96 33.235 ;
    RECT 51.75 33.525 51.96 33.595 ;
    RECT 51.75 33.885 51.96 33.955 ;
    RECT 47.97 33.165 48.18 33.235 ;
    RECT 47.97 33.525 48.18 33.595 ;
    RECT 47.97 33.885 48.18 33.955 ;
    RECT 48.43 33.165 48.64 33.235 ;
    RECT 48.43 33.525 48.64 33.595 ;
    RECT 48.43 33.885 48.64 33.955 ;
    RECT 44.65 33.165 44.86 33.235 ;
    RECT 44.65 33.525 44.86 33.595 ;
    RECT 44.65 33.885 44.86 33.955 ;
    RECT 45.11 33.165 45.32 33.235 ;
    RECT 45.11 33.525 45.32 33.595 ;
    RECT 45.11 33.885 45.32 33.955 ;
    RECT 41.33 33.165 41.54 33.235 ;
    RECT 41.33 33.525 41.54 33.595 ;
    RECT 41.33 33.885 41.54 33.955 ;
    RECT 41.79 33.165 42.0 33.235 ;
    RECT 41.79 33.525 42.0 33.595 ;
    RECT 41.79 33.885 42.0 33.955 ;
    RECT 38.01 33.165 38.22 33.235 ;
    RECT 38.01 33.525 38.22 33.595 ;
    RECT 38.01 33.885 38.22 33.955 ;
    RECT 38.47 33.165 38.68 33.235 ;
    RECT 38.47 33.525 38.68 33.595 ;
    RECT 38.47 33.885 38.68 33.955 ;
    RECT 34.69 33.165 34.9 33.235 ;
    RECT 34.69 33.525 34.9 33.595 ;
    RECT 34.69 33.885 34.9 33.955 ;
    RECT 35.15 33.165 35.36 33.235 ;
    RECT 35.15 33.525 35.36 33.595 ;
    RECT 35.15 33.885 35.36 33.955 ;
    RECT 173.945 33.525 174.015 33.595 ;
    RECT 130.97 33.165 131.18 33.235 ;
    RECT 130.97 33.525 131.18 33.595 ;
    RECT 130.97 33.885 131.18 33.955 ;
    RECT 131.43 33.165 131.64 33.235 ;
    RECT 131.43 33.525 131.64 33.595 ;
    RECT 131.43 33.885 131.64 33.955 ;
    RECT 127.65 33.165 127.86 33.235 ;
    RECT 127.65 33.525 127.86 33.595 ;
    RECT 127.65 33.885 127.86 33.955 ;
    RECT 128.11 33.165 128.32 33.235 ;
    RECT 128.11 33.525 128.32 33.595 ;
    RECT 128.11 33.885 128.32 33.955 ;
    RECT 124.33 33.165 124.54 33.235 ;
    RECT 124.33 33.525 124.54 33.595 ;
    RECT 124.33 33.885 124.54 33.955 ;
    RECT 124.79 33.165 125.0 33.235 ;
    RECT 124.79 33.525 125.0 33.595 ;
    RECT 124.79 33.885 125.0 33.955 ;
    RECT 121.01 33.165 121.22 33.235 ;
    RECT 121.01 33.525 121.22 33.595 ;
    RECT 121.01 33.885 121.22 33.955 ;
    RECT 121.47 33.165 121.68 33.235 ;
    RECT 121.47 33.525 121.68 33.595 ;
    RECT 121.47 33.885 121.68 33.955 ;
    RECT 117.69 33.165 117.9 33.235 ;
    RECT 117.69 33.525 117.9 33.595 ;
    RECT 117.69 33.885 117.9 33.955 ;
    RECT 118.15 33.165 118.36 33.235 ;
    RECT 118.15 33.525 118.36 33.595 ;
    RECT 118.15 33.885 118.36 33.955 ;
    RECT 114.37 33.165 114.58 33.235 ;
    RECT 114.37 33.525 114.58 33.595 ;
    RECT 114.37 33.885 114.58 33.955 ;
    RECT 114.83 33.165 115.04 33.235 ;
    RECT 114.83 33.525 115.04 33.595 ;
    RECT 114.83 33.885 115.04 33.955 ;
    RECT 111.05 33.165 111.26 33.235 ;
    RECT 111.05 33.525 111.26 33.595 ;
    RECT 111.05 33.885 111.26 33.955 ;
    RECT 111.51 33.165 111.72 33.235 ;
    RECT 111.51 33.525 111.72 33.595 ;
    RECT 111.51 33.885 111.72 33.955 ;
    RECT 107.73 33.165 107.94 33.235 ;
    RECT 107.73 33.525 107.94 33.595 ;
    RECT 107.73 33.885 107.94 33.955 ;
    RECT 108.19 33.165 108.4 33.235 ;
    RECT 108.19 33.525 108.4 33.595 ;
    RECT 108.19 33.885 108.4 33.955 ;
    RECT 104.41 33.165 104.62 33.235 ;
    RECT 104.41 33.525 104.62 33.595 ;
    RECT 104.41 33.885 104.62 33.955 ;
    RECT 104.87 33.165 105.08 33.235 ;
    RECT 104.87 33.525 105.08 33.595 ;
    RECT 104.87 33.885 105.08 33.955 ;
    RECT 101.09 33.165 101.3 33.235 ;
    RECT 101.09 33.525 101.3 33.595 ;
    RECT 101.09 33.885 101.3 33.955 ;
    RECT 101.55 33.165 101.76 33.235 ;
    RECT 101.55 33.525 101.76 33.595 ;
    RECT 101.55 33.885 101.76 33.955 ;
    RECT 0.4 33.525 0.47 33.595 ;
    RECT 170.81 33.165 171.02 33.235 ;
    RECT 170.81 33.525 171.02 33.595 ;
    RECT 170.81 33.885 171.02 33.955 ;
    RECT 171.27 33.165 171.48 33.235 ;
    RECT 171.27 33.525 171.48 33.595 ;
    RECT 171.27 33.885 171.48 33.955 ;
    RECT 167.49 33.165 167.7 33.235 ;
    RECT 167.49 33.525 167.7 33.595 ;
    RECT 167.49 33.885 167.7 33.955 ;
    RECT 167.95 33.165 168.16 33.235 ;
    RECT 167.95 33.525 168.16 33.595 ;
    RECT 167.95 33.885 168.16 33.955 ;
    RECT 97.77 33.165 97.98 33.235 ;
    RECT 97.77 33.525 97.98 33.595 ;
    RECT 97.77 33.885 97.98 33.955 ;
    RECT 98.23 33.165 98.44 33.235 ;
    RECT 98.23 33.525 98.44 33.595 ;
    RECT 98.23 33.885 98.44 33.955 ;
    RECT 94.45 33.165 94.66 33.235 ;
    RECT 94.45 33.525 94.66 33.595 ;
    RECT 94.45 33.885 94.66 33.955 ;
    RECT 94.91 33.165 95.12 33.235 ;
    RECT 94.91 33.525 95.12 33.595 ;
    RECT 94.91 33.885 95.12 33.955 ;
    RECT 91.13 33.165 91.34 33.235 ;
    RECT 91.13 33.525 91.34 33.595 ;
    RECT 91.13 33.885 91.34 33.955 ;
    RECT 91.59 33.165 91.8 33.235 ;
    RECT 91.59 33.525 91.8 33.595 ;
    RECT 91.59 33.885 91.8 33.955 ;
    RECT 87.81 33.165 88.02 33.235 ;
    RECT 87.81 33.525 88.02 33.595 ;
    RECT 87.81 33.885 88.02 33.955 ;
    RECT 88.27 33.165 88.48 33.235 ;
    RECT 88.27 33.525 88.48 33.595 ;
    RECT 88.27 33.885 88.48 33.955 ;
    RECT 84.49 33.165 84.7 33.235 ;
    RECT 84.49 33.525 84.7 33.595 ;
    RECT 84.49 33.885 84.7 33.955 ;
    RECT 84.95 33.165 85.16 33.235 ;
    RECT 84.95 33.525 85.16 33.595 ;
    RECT 84.95 33.885 85.16 33.955 ;
    RECT 81.17 33.165 81.38 33.235 ;
    RECT 81.17 33.525 81.38 33.595 ;
    RECT 81.17 33.885 81.38 33.955 ;
    RECT 81.63 33.165 81.84 33.235 ;
    RECT 81.63 33.525 81.84 33.595 ;
    RECT 81.63 33.885 81.84 33.955 ;
    RECT 77.85 33.165 78.06 33.235 ;
    RECT 77.85 33.525 78.06 33.595 ;
    RECT 77.85 33.885 78.06 33.955 ;
    RECT 78.31 33.165 78.52 33.235 ;
    RECT 78.31 33.525 78.52 33.595 ;
    RECT 78.31 33.885 78.52 33.955 ;
    RECT 74.53 33.165 74.74 33.235 ;
    RECT 74.53 33.525 74.74 33.595 ;
    RECT 74.53 33.885 74.74 33.955 ;
    RECT 74.99 33.165 75.2 33.235 ;
    RECT 74.99 33.525 75.2 33.595 ;
    RECT 74.99 33.885 75.2 33.955 ;
    RECT 71.21 33.165 71.42 33.235 ;
    RECT 71.21 33.525 71.42 33.595 ;
    RECT 71.21 33.885 71.42 33.955 ;
    RECT 71.67 33.165 71.88 33.235 ;
    RECT 71.67 33.525 71.88 33.595 ;
    RECT 71.67 33.885 71.88 33.955 ;
    RECT 31.37 33.165 31.58 33.235 ;
    RECT 31.37 33.525 31.58 33.595 ;
    RECT 31.37 33.885 31.58 33.955 ;
    RECT 31.83 33.165 32.04 33.235 ;
    RECT 31.83 33.525 32.04 33.595 ;
    RECT 31.83 33.885 32.04 33.955 ;
    RECT 67.89 33.165 68.1 33.235 ;
    RECT 67.89 33.525 68.1 33.595 ;
    RECT 67.89 33.885 68.1 33.955 ;
    RECT 68.35 33.165 68.56 33.235 ;
    RECT 68.35 33.525 68.56 33.595 ;
    RECT 68.35 33.885 68.56 33.955 ;
    RECT 28.05 33.165 28.26 33.235 ;
    RECT 28.05 33.525 28.26 33.595 ;
    RECT 28.05 33.885 28.26 33.955 ;
    RECT 28.51 33.165 28.72 33.235 ;
    RECT 28.51 33.525 28.72 33.595 ;
    RECT 28.51 33.885 28.72 33.955 ;
    RECT 24.73 33.165 24.94 33.235 ;
    RECT 24.73 33.525 24.94 33.595 ;
    RECT 24.73 33.885 24.94 33.955 ;
    RECT 25.19 33.165 25.4 33.235 ;
    RECT 25.19 33.525 25.4 33.595 ;
    RECT 25.19 33.885 25.4 33.955 ;
    RECT 21.41 33.165 21.62 33.235 ;
    RECT 21.41 33.525 21.62 33.595 ;
    RECT 21.41 33.885 21.62 33.955 ;
    RECT 21.87 33.165 22.08 33.235 ;
    RECT 21.87 33.525 22.08 33.595 ;
    RECT 21.87 33.885 22.08 33.955 ;
    RECT 18.09 33.165 18.3 33.235 ;
    RECT 18.09 33.525 18.3 33.595 ;
    RECT 18.09 33.885 18.3 33.955 ;
    RECT 18.55 33.165 18.76 33.235 ;
    RECT 18.55 33.525 18.76 33.595 ;
    RECT 18.55 33.885 18.76 33.955 ;
    RECT 14.77 33.165 14.98 33.235 ;
    RECT 14.77 33.525 14.98 33.595 ;
    RECT 14.77 33.885 14.98 33.955 ;
    RECT 15.23 33.165 15.44 33.235 ;
    RECT 15.23 33.525 15.44 33.595 ;
    RECT 15.23 33.885 15.44 33.955 ;
    RECT 11.45 33.165 11.66 33.235 ;
    RECT 11.45 33.525 11.66 33.595 ;
    RECT 11.45 33.885 11.66 33.955 ;
    RECT 11.91 33.165 12.12 33.235 ;
    RECT 11.91 33.525 12.12 33.595 ;
    RECT 11.91 33.885 12.12 33.955 ;
    RECT 8.13 33.165 8.34 33.235 ;
    RECT 8.13 33.525 8.34 33.595 ;
    RECT 8.13 33.885 8.34 33.955 ;
    RECT 8.59 33.165 8.8 33.235 ;
    RECT 8.59 33.525 8.8 33.595 ;
    RECT 8.59 33.885 8.8 33.955 ;
    RECT 4.81 33.165 5.02 33.235 ;
    RECT 4.81 33.525 5.02 33.595 ;
    RECT 4.81 33.885 5.02 33.955 ;
    RECT 5.27 33.165 5.48 33.235 ;
    RECT 5.27 33.525 5.48 33.595 ;
    RECT 5.27 33.885 5.48 33.955 ;
    RECT 164.17 33.165 164.38 33.235 ;
    RECT 164.17 33.525 164.38 33.595 ;
    RECT 164.17 33.885 164.38 33.955 ;
    RECT 164.63 33.165 164.84 33.235 ;
    RECT 164.63 33.525 164.84 33.595 ;
    RECT 164.63 33.885 164.84 33.955 ;
    RECT 1.49 33.165 1.7 33.235 ;
    RECT 1.49 33.525 1.7 33.595 ;
    RECT 1.49 33.885 1.7 33.955 ;
    RECT 1.95 33.165 2.16 33.235 ;
    RECT 1.95 33.525 2.16 33.595 ;
    RECT 1.95 33.885 2.16 33.955 ;
    RECT 160.85 33.165 161.06 33.235 ;
    RECT 160.85 33.525 161.06 33.595 ;
    RECT 160.85 33.885 161.06 33.955 ;
    RECT 161.31 33.165 161.52 33.235 ;
    RECT 161.31 33.525 161.52 33.595 ;
    RECT 161.31 33.885 161.52 33.955 ;
    RECT 157.53 33.165 157.74 33.235 ;
    RECT 157.53 33.525 157.74 33.595 ;
    RECT 157.53 33.885 157.74 33.955 ;
    RECT 157.99 33.165 158.2 33.235 ;
    RECT 157.99 33.525 158.2 33.595 ;
    RECT 157.99 33.885 158.2 33.955 ;
    RECT 154.21 33.165 154.42 33.235 ;
    RECT 154.21 33.525 154.42 33.595 ;
    RECT 154.21 33.885 154.42 33.955 ;
    RECT 154.67 33.165 154.88 33.235 ;
    RECT 154.67 33.525 154.88 33.595 ;
    RECT 154.67 33.885 154.88 33.955 ;
    RECT 150.89 33.165 151.1 33.235 ;
    RECT 150.89 33.525 151.1 33.595 ;
    RECT 150.89 33.885 151.1 33.955 ;
    RECT 151.35 33.165 151.56 33.235 ;
    RECT 151.35 33.525 151.56 33.595 ;
    RECT 151.35 33.885 151.56 33.955 ;
    RECT 147.57 33.165 147.78 33.235 ;
    RECT 147.57 33.525 147.78 33.595 ;
    RECT 147.57 33.885 147.78 33.955 ;
    RECT 148.03 33.165 148.24 33.235 ;
    RECT 148.03 33.525 148.24 33.595 ;
    RECT 148.03 33.885 148.24 33.955 ;
    RECT 144.25 33.165 144.46 33.235 ;
    RECT 144.25 33.525 144.46 33.595 ;
    RECT 144.25 33.885 144.46 33.955 ;
    RECT 144.71 33.165 144.92 33.235 ;
    RECT 144.71 33.525 144.92 33.595 ;
    RECT 144.71 33.885 144.92 33.955 ;
    RECT 140.93 33.165 141.14 33.235 ;
    RECT 140.93 33.525 141.14 33.595 ;
    RECT 140.93 33.885 141.14 33.955 ;
    RECT 141.39 33.165 141.6 33.235 ;
    RECT 141.39 33.525 141.6 33.595 ;
    RECT 141.39 33.885 141.6 33.955 ;
    RECT 137.61 33.165 137.82 33.235 ;
    RECT 137.61 33.525 137.82 33.595 ;
    RECT 137.61 33.885 137.82 33.955 ;
    RECT 138.07 33.165 138.28 33.235 ;
    RECT 138.07 33.525 138.28 33.595 ;
    RECT 138.07 33.885 138.28 33.955 ;
    RECT 134.29 33.165 134.5 33.235 ;
    RECT 134.29 33.525 134.5 33.595 ;
    RECT 134.29 33.885 134.5 33.955 ;
    RECT 134.75 33.165 134.96 33.235 ;
    RECT 134.75 33.525 134.96 33.595 ;
    RECT 134.75 33.885 134.96 33.955 ;
    RECT 64.57 33.165 64.78 33.235 ;
    RECT 64.57 33.525 64.78 33.595 ;
    RECT 64.57 33.885 64.78 33.955 ;
    RECT 65.03 33.165 65.24 33.235 ;
    RECT 65.03 33.525 65.24 33.595 ;
    RECT 65.03 33.885 65.24 33.955 ;
    RECT 61.25 32.445 61.46 32.515 ;
    RECT 61.25 32.805 61.46 32.875 ;
    RECT 61.25 33.165 61.46 33.235 ;
    RECT 61.71 32.445 61.92 32.515 ;
    RECT 61.71 32.805 61.92 32.875 ;
    RECT 61.71 33.165 61.92 33.235 ;
    RECT 57.93 32.445 58.14 32.515 ;
    RECT 57.93 32.805 58.14 32.875 ;
    RECT 57.93 33.165 58.14 33.235 ;
    RECT 58.39 32.445 58.6 32.515 ;
    RECT 58.39 32.805 58.6 32.875 ;
    RECT 58.39 33.165 58.6 33.235 ;
    RECT 54.61 32.445 54.82 32.515 ;
    RECT 54.61 32.805 54.82 32.875 ;
    RECT 54.61 33.165 54.82 33.235 ;
    RECT 55.07 32.445 55.28 32.515 ;
    RECT 55.07 32.805 55.28 32.875 ;
    RECT 55.07 33.165 55.28 33.235 ;
    RECT 51.29 32.445 51.5 32.515 ;
    RECT 51.29 32.805 51.5 32.875 ;
    RECT 51.29 33.165 51.5 33.235 ;
    RECT 51.75 32.445 51.96 32.515 ;
    RECT 51.75 32.805 51.96 32.875 ;
    RECT 51.75 33.165 51.96 33.235 ;
    RECT 47.97 32.445 48.18 32.515 ;
    RECT 47.97 32.805 48.18 32.875 ;
    RECT 47.97 33.165 48.18 33.235 ;
    RECT 48.43 32.445 48.64 32.515 ;
    RECT 48.43 32.805 48.64 32.875 ;
    RECT 48.43 33.165 48.64 33.235 ;
    RECT 44.65 32.445 44.86 32.515 ;
    RECT 44.65 32.805 44.86 32.875 ;
    RECT 44.65 33.165 44.86 33.235 ;
    RECT 45.11 32.445 45.32 32.515 ;
    RECT 45.11 32.805 45.32 32.875 ;
    RECT 45.11 33.165 45.32 33.235 ;
    RECT 41.33 32.445 41.54 32.515 ;
    RECT 41.33 32.805 41.54 32.875 ;
    RECT 41.33 33.165 41.54 33.235 ;
    RECT 41.79 32.445 42.0 32.515 ;
    RECT 41.79 32.805 42.0 32.875 ;
    RECT 41.79 33.165 42.0 33.235 ;
    RECT 38.01 32.445 38.22 32.515 ;
    RECT 38.01 32.805 38.22 32.875 ;
    RECT 38.01 33.165 38.22 33.235 ;
    RECT 38.47 32.445 38.68 32.515 ;
    RECT 38.47 32.805 38.68 32.875 ;
    RECT 38.47 33.165 38.68 33.235 ;
    RECT 34.69 32.445 34.9 32.515 ;
    RECT 34.69 32.805 34.9 32.875 ;
    RECT 34.69 33.165 34.9 33.235 ;
    RECT 35.15 32.445 35.36 32.515 ;
    RECT 35.15 32.805 35.36 32.875 ;
    RECT 35.15 33.165 35.36 33.235 ;
    RECT 173.945 32.805 174.015 32.875 ;
    RECT 130.97 32.445 131.18 32.515 ;
    RECT 130.97 32.805 131.18 32.875 ;
    RECT 130.97 33.165 131.18 33.235 ;
    RECT 131.43 32.445 131.64 32.515 ;
    RECT 131.43 32.805 131.64 32.875 ;
    RECT 131.43 33.165 131.64 33.235 ;
    RECT 127.65 32.445 127.86 32.515 ;
    RECT 127.65 32.805 127.86 32.875 ;
    RECT 127.65 33.165 127.86 33.235 ;
    RECT 128.11 32.445 128.32 32.515 ;
    RECT 128.11 32.805 128.32 32.875 ;
    RECT 128.11 33.165 128.32 33.235 ;
    RECT 124.33 32.445 124.54 32.515 ;
    RECT 124.33 32.805 124.54 32.875 ;
    RECT 124.33 33.165 124.54 33.235 ;
    RECT 124.79 32.445 125.0 32.515 ;
    RECT 124.79 32.805 125.0 32.875 ;
    RECT 124.79 33.165 125.0 33.235 ;
    RECT 121.01 32.445 121.22 32.515 ;
    RECT 121.01 32.805 121.22 32.875 ;
    RECT 121.01 33.165 121.22 33.235 ;
    RECT 121.47 32.445 121.68 32.515 ;
    RECT 121.47 32.805 121.68 32.875 ;
    RECT 121.47 33.165 121.68 33.235 ;
    RECT 117.69 32.445 117.9 32.515 ;
    RECT 117.69 32.805 117.9 32.875 ;
    RECT 117.69 33.165 117.9 33.235 ;
    RECT 118.15 32.445 118.36 32.515 ;
    RECT 118.15 32.805 118.36 32.875 ;
    RECT 118.15 33.165 118.36 33.235 ;
    RECT 114.37 32.445 114.58 32.515 ;
    RECT 114.37 32.805 114.58 32.875 ;
    RECT 114.37 33.165 114.58 33.235 ;
    RECT 114.83 32.445 115.04 32.515 ;
    RECT 114.83 32.805 115.04 32.875 ;
    RECT 114.83 33.165 115.04 33.235 ;
    RECT 111.05 32.445 111.26 32.515 ;
    RECT 111.05 32.805 111.26 32.875 ;
    RECT 111.05 33.165 111.26 33.235 ;
    RECT 111.51 32.445 111.72 32.515 ;
    RECT 111.51 32.805 111.72 32.875 ;
    RECT 111.51 33.165 111.72 33.235 ;
    RECT 107.73 32.445 107.94 32.515 ;
    RECT 107.73 32.805 107.94 32.875 ;
    RECT 107.73 33.165 107.94 33.235 ;
    RECT 108.19 32.445 108.4 32.515 ;
    RECT 108.19 32.805 108.4 32.875 ;
    RECT 108.19 33.165 108.4 33.235 ;
    RECT 104.41 32.445 104.62 32.515 ;
    RECT 104.41 32.805 104.62 32.875 ;
    RECT 104.41 33.165 104.62 33.235 ;
    RECT 104.87 32.445 105.08 32.515 ;
    RECT 104.87 32.805 105.08 32.875 ;
    RECT 104.87 33.165 105.08 33.235 ;
    RECT 101.09 32.445 101.3 32.515 ;
    RECT 101.09 32.805 101.3 32.875 ;
    RECT 101.09 33.165 101.3 33.235 ;
    RECT 101.55 32.445 101.76 32.515 ;
    RECT 101.55 32.805 101.76 32.875 ;
    RECT 101.55 33.165 101.76 33.235 ;
    RECT 0.4 32.805 0.47 32.875 ;
    RECT 170.81 32.445 171.02 32.515 ;
    RECT 170.81 32.805 171.02 32.875 ;
    RECT 170.81 33.165 171.02 33.235 ;
    RECT 171.27 32.445 171.48 32.515 ;
    RECT 171.27 32.805 171.48 32.875 ;
    RECT 171.27 33.165 171.48 33.235 ;
    RECT 167.49 32.445 167.7 32.515 ;
    RECT 167.49 32.805 167.7 32.875 ;
    RECT 167.49 33.165 167.7 33.235 ;
    RECT 167.95 32.445 168.16 32.515 ;
    RECT 167.95 32.805 168.16 32.875 ;
    RECT 167.95 33.165 168.16 33.235 ;
    RECT 97.77 32.445 97.98 32.515 ;
    RECT 97.77 32.805 97.98 32.875 ;
    RECT 97.77 33.165 97.98 33.235 ;
    RECT 98.23 32.445 98.44 32.515 ;
    RECT 98.23 32.805 98.44 32.875 ;
    RECT 98.23 33.165 98.44 33.235 ;
    RECT 94.45 32.445 94.66 32.515 ;
    RECT 94.45 32.805 94.66 32.875 ;
    RECT 94.45 33.165 94.66 33.235 ;
    RECT 94.91 32.445 95.12 32.515 ;
    RECT 94.91 32.805 95.12 32.875 ;
    RECT 94.91 33.165 95.12 33.235 ;
    RECT 91.13 32.445 91.34 32.515 ;
    RECT 91.13 32.805 91.34 32.875 ;
    RECT 91.13 33.165 91.34 33.235 ;
    RECT 91.59 32.445 91.8 32.515 ;
    RECT 91.59 32.805 91.8 32.875 ;
    RECT 91.59 33.165 91.8 33.235 ;
    RECT 87.81 32.445 88.02 32.515 ;
    RECT 87.81 32.805 88.02 32.875 ;
    RECT 87.81 33.165 88.02 33.235 ;
    RECT 88.27 32.445 88.48 32.515 ;
    RECT 88.27 32.805 88.48 32.875 ;
    RECT 88.27 33.165 88.48 33.235 ;
    RECT 84.49 32.445 84.7 32.515 ;
    RECT 84.49 32.805 84.7 32.875 ;
    RECT 84.49 33.165 84.7 33.235 ;
    RECT 84.95 32.445 85.16 32.515 ;
    RECT 84.95 32.805 85.16 32.875 ;
    RECT 84.95 33.165 85.16 33.235 ;
    RECT 81.17 32.445 81.38 32.515 ;
    RECT 81.17 32.805 81.38 32.875 ;
    RECT 81.17 33.165 81.38 33.235 ;
    RECT 81.63 32.445 81.84 32.515 ;
    RECT 81.63 32.805 81.84 32.875 ;
    RECT 81.63 33.165 81.84 33.235 ;
    RECT 77.85 32.445 78.06 32.515 ;
    RECT 77.85 32.805 78.06 32.875 ;
    RECT 77.85 33.165 78.06 33.235 ;
    RECT 78.31 32.445 78.52 32.515 ;
    RECT 78.31 32.805 78.52 32.875 ;
    RECT 78.31 33.165 78.52 33.235 ;
    RECT 74.53 32.445 74.74 32.515 ;
    RECT 74.53 32.805 74.74 32.875 ;
    RECT 74.53 33.165 74.74 33.235 ;
    RECT 74.99 32.445 75.2 32.515 ;
    RECT 74.99 32.805 75.2 32.875 ;
    RECT 74.99 33.165 75.2 33.235 ;
    RECT 71.21 32.445 71.42 32.515 ;
    RECT 71.21 32.805 71.42 32.875 ;
    RECT 71.21 33.165 71.42 33.235 ;
    RECT 71.67 32.445 71.88 32.515 ;
    RECT 71.67 32.805 71.88 32.875 ;
    RECT 71.67 33.165 71.88 33.235 ;
    RECT 31.37 32.445 31.58 32.515 ;
    RECT 31.37 32.805 31.58 32.875 ;
    RECT 31.37 33.165 31.58 33.235 ;
    RECT 31.83 32.445 32.04 32.515 ;
    RECT 31.83 32.805 32.04 32.875 ;
    RECT 31.83 33.165 32.04 33.235 ;
    RECT 67.89 32.445 68.1 32.515 ;
    RECT 67.89 32.805 68.1 32.875 ;
    RECT 67.89 33.165 68.1 33.235 ;
    RECT 68.35 32.445 68.56 32.515 ;
    RECT 68.35 32.805 68.56 32.875 ;
    RECT 68.35 33.165 68.56 33.235 ;
    RECT 28.05 32.445 28.26 32.515 ;
    RECT 28.05 32.805 28.26 32.875 ;
    RECT 28.05 33.165 28.26 33.235 ;
    RECT 28.51 32.445 28.72 32.515 ;
    RECT 28.51 32.805 28.72 32.875 ;
    RECT 28.51 33.165 28.72 33.235 ;
    RECT 24.73 32.445 24.94 32.515 ;
    RECT 24.73 32.805 24.94 32.875 ;
    RECT 24.73 33.165 24.94 33.235 ;
    RECT 25.19 32.445 25.4 32.515 ;
    RECT 25.19 32.805 25.4 32.875 ;
    RECT 25.19 33.165 25.4 33.235 ;
    RECT 21.41 32.445 21.62 32.515 ;
    RECT 21.41 32.805 21.62 32.875 ;
    RECT 21.41 33.165 21.62 33.235 ;
    RECT 21.87 32.445 22.08 32.515 ;
    RECT 21.87 32.805 22.08 32.875 ;
    RECT 21.87 33.165 22.08 33.235 ;
    RECT 18.09 32.445 18.3 32.515 ;
    RECT 18.09 32.805 18.3 32.875 ;
    RECT 18.09 33.165 18.3 33.235 ;
    RECT 18.55 32.445 18.76 32.515 ;
    RECT 18.55 32.805 18.76 32.875 ;
    RECT 18.55 33.165 18.76 33.235 ;
    RECT 14.77 32.445 14.98 32.515 ;
    RECT 14.77 32.805 14.98 32.875 ;
    RECT 14.77 33.165 14.98 33.235 ;
    RECT 15.23 32.445 15.44 32.515 ;
    RECT 15.23 32.805 15.44 32.875 ;
    RECT 15.23 33.165 15.44 33.235 ;
    RECT 11.45 32.445 11.66 32.515 ;
    RECT 11.45 32.805 11.66 32.875 ;
    RECT 11.45 33.165 11.66 33.235 ;
    RECT 11.91 32.445 12.12 32.515 ;
    RECT 11.91 32.805 12.12 32.875 ;
    RECT 11.91 33.165 12.12 33.235 ;
    RECT 8.13 32.445 8.34 32.515 ;
    RECT 8.13 32.805 8.34 32.875 ;
    RECT 8.13 33.165 8.34 33.235 ;
    RECT 8.59 32.445 8.8 32.515 ;
    RECT 8.59 32.805 8.8 32.875 ;
    RECT 8.59 33.165 8.8 33.235 ;
    RECT 4.81 32.445 5.02 32.515 ;
    RECT 4.81 32.805 5.02 32.875 ;
    RECT 4.81 33.165 5.02 33.235 ;
    RECT 5.27 32.445 5.48 32.515 ;
    RECT 5.27 32.805 5.48 32.875 ;
    RECT 5.27 33.165 5.48 33.235 ;
    RECT 164.17 32.445 164.38 32.515 ;
    RECT 164.17 32.805 164.38 32.875 ;
    RECT 164.17 33.165 164.38 33.235 ;
    RECT 164.63 32.445 164.84 32.515 ;
    RECT 164.63 32.805 164.84 32.875 ;
    RECT 164.63 33.165 164.84 33.235 ;
    RECT 1.49 32.445 1.7 32.515 ;
    RECT 1.49 32.805 1.7 32.875 ;
    RECT 1.49 33.165 1.7 33.235 ;
    RECT 1.95 32.445 2.16 32.515 ;
    RECT 1.95 32.805 2.16 32.875 ;
    RECT 1.95 33.165 2.16 33.235 ;
    RECT 160.85 32.445 161.06 32.515 ;
    RECT 160.85 32.805 161.06 32.875 ;
    RECT 160.85 33.165 161.06 33.235 ;
    RECT 161.31 32.445 161.52 32.515 ;
    RECT 161.31 32.805 161.52 32.875 ;
    RECT 161.31 33.165 161.52 33.235 ;
    RECT 157.53 32.445 157.74 32.515 ;
    RECT 157.53 32.805 157.74 32.875 ;
    RECT 157.53 33.165 157.74 33.235 ;
    RECT 157.99 32.445 158.2 32.515 ;
    RECT 157.99 32.805 158.2 32.875 ;
    RECT 157.99 33.165 158.2 33.235 ;
    RECT 154.21 32.445 154.42 32.515 ;
    RECT 154.21 32.805 154.42 32.875 ;
    RECT 154.21 33.165 154.42 33.235 ;
    RECT 154.67 32.445 154.88 32.515 ;
    RECT 154.67 32.805 154.88 32.875 ;
    RECT 154.67 33.165 154.88 33.235 ;
    RECT 150.89 32.445 151.1 32.515 ;
    RECT 150.89 32.805 151.1 32.875 ;
    RECT 150.89 33.165 151.1 33.235 ;
    RECT 151.35 32.445 151.56 32.515 ;
    RECT 151.35 32.805 151.56 32.875 ;
    RECT 151.35 33.165 151.56 33.235 ;
    RECT 147.57 32.445 147.78 32.515 ;
    RECT 147.57 32.805 147.78 32.875 ;
    RECT 147.57 33.165 147.78 33.235 ;
    RECT 148.03 32.445 148.24 32.515 ;
    RECT 148.03 32.805 148.24 32.875 ;
    RECT 148.03 33.165 148.24 33.235 ;
    RECT 144.25 32.445 144.46 32.515 ;
    RECT 144.25 32.805 144.46 32.875 ;
    RECT 144.25 33.165 144.46 33.235 ;
    RECT 144.71 32.445 144.92 32.515 ;
    RECT 144.71 32.805 144.92 32.875 ;
    RECT 144.71 33.165 144.92 33.235 ;
    RECT 140.93 32.445 141.14 32.515 ;
    RECT 140.93 32.805 141.14 32.875 ;
    RECT 140.93 33.165 141.14 33.235 ;
    RECT 141.39 32.445 141.6 32.515 ;
    RECT 141.39 32.805 141.6 32.875 ;
    RECT 141.39 33.165 141.6 33.235 ;
    RECT 137.61 32.445 137.82 32.515 ;
    RECT 137.61 32.805 137.82 32.875 ;
    RECT 137.61 33.165 137.82 33.235 ;
    RECT 138.07 32.445 138.28 32.515 ;
    RECT 138.07 32.805 138.28 32.875 ;
    RECT 138.07 33.165 138.28 33.235 ;
    RECT 134.29 32.445 134.5 32.515 ;
    RECT 134.29 32.805 134.5 32.875 ;
    RECT 134.29 33.165 134.5 33.235 ;
    RECT 134.75 32.445 134.96 32.515 ;
    RECT 134.75 32.805 134.96 32.875 ;
    RECT 134.75 33.165 134.96 33.235 ;
    RECT 64.57 32.445 64.78 32.515 ;
    RECT 64.57 32.805 64.78 32.875 ;
    RECT 64.57 33.165 64.78 33.235 ;
    RECT 65.03 32.445 65.24 32.515 ;
    RECT 65.03 32.805 65.24 32.875 ;
    RECT 65.03 33.165 65.24 33.235 ;
    RECT 61.25 31.725 61.46 31.795 ;
    RECT 61.25 32.085 61.46 32.155 ;
    RECT 61.25 32.445 61.46 32.515 ;
    RECT 61.71 31.725 61.92 31.795 ;
    RECT 61.71 32.085 61.92 32.155 ;
    RECT 61.71 32.445 61.92 32.515 ;
    RECT 57.93 31.725 58.14 31.795 ;
    RECT 57.93 32.085 58.14 32.155 ;
    RECT 57.93 32.445 58.14 32.515 ;
    RECT 58.39 31.725 58.6 31.795 ;
    RECT 58.39 32.085 58.6 32.155 ;
    RECT 58.39 32.445 58.6 32.515 ;
    RECT 54.61 31.725 54.82 31.795 ;
    RECT 54.61 32.085 54.82 32.155 ;
    RECT 54.61 32.445 54.82 32.515 ;
    RECT 55.07 31.725 55.28 31.795 ;
    RECT 55.07 32.085 55.28 32.155 ;
    RECT 55.07 32.445 55.28 32.515 ;
    RECT 51.29 31.725 51.5 31.795 ;
    RECT 51.29 32.085 51.5 32.155 ;
    RECT 51.29 32.445 51.5 32.515 ;
    RECT 51.75 31.725 51.96 31.795 ;
    RECT 51.75 32.085 51.96 32.155 ;
    RECT 51.75 32.445 51.96 32.515 ;
    RECT 47.97 31.725 48.18 31.795 ;
    RECT 47.97 32.085 48.18 32.155 ;
    RECT 47.97 32.445 48.18 32.515 ;
    RECT 48.43 31.725 48.64 31.795 ;
    RECT 48.43 32.085 48.64 32.155 ;
    RECT 48.43 32.445 48.64 32.515 ;
    RECT 44.65 31.725 44.86 31.795 ;
    RECT 44.65 32.085 44.86 32.155 ;
    RECT 44.65 32.445 44.86 32.515 ;
    RECT 45.11 31.725 45.32 31.795 ;
    RECT 45.11 32.085 45.32 32.155 ;
    RECT 45.11 32.445 45.32 32.515 ;
    RECT 41.33 31.725 41.54 31.795 ;
    RECT 41.33 32.085 41.54 32.155 ;
    RECT 41.33 32.445 41.54 32.515 ;
    RECT 41.79 31.725 42.0 31.795 ;
    RECT 41.79 32.085 42.0 32.155 ;
    RECT 41.79 32.445 42.0 32.515 ;
    RECT 38.01 31.725 38.22 31.795 ;
    RECT 38.01 32.085 38.22 32.155 ;
    RECT 38.01 32.445 38.22 32.515 ;
    RECT 38.47 31.725 38.68 31.795 ;
    RECT 38.47 32.085 38.68 32.155 ;
    RECT 38.47 32.445 38.68 32.515 ;
    RECT 34.69 31.725 34.9 31.795 ;
    RECT 34.69 32.085 34.9 32.155 ;
    RECT 34.69 32.445 34.9 32.515 ;
    RECT 35.15 31.725 35.36 31.795 ;
    RECT 35.15 32.085 35.36 32.155 ;
    RECT 35.15 32.445 35.36 32.515 ;
    RECT 173.945 32.085 174.015 32.155 ;
    RECT 130.97 31.725 131.18 31.795 ;
    RECT 130.97 32.085 131.18 32.155 ;
    RECT 130.97 32.445 131.18 32.515 ;
    RECT 131.43 31.725 131.64 31.795 ;
    RECT 131.43 32.085 131.64 32.155 ;
    RECT 131.43 32.445 131.64 32.515 ;
    RECT 127.65 31.725 127.86 31.795 ;
    RECT 127.65 32.085 127.86 32.155 ;
    RECT 127.65 32.445 127.86 32.515 ;
    RECT 128.11 31.725 128.32 31.795 ;
    RECT 128.11 32.085 128.32 32.155 ;
    RECT 128.11 32.445 128.32 32.515 ;
    RECT 124.33 31.725 124.54 31.795 ;
    RECT 124.33 32.085 124.54 32.155 ;
    RECT 124.33 32.445 124.54 32.515 ;
    RECT 124.79 31.725 125.0 31.795 ;
    RECT 124.79 32.085 125.0 32.155 ;
    RECT 124.79 32.445 125.0 32.515 ;
    RECT 121.01 31.725 121.22 31.795 ;
    RECT 121.01 32.085 121.22 32.155 ;
    RECT 121.01 32.445 121.22 32.515 ;
    RECT 121.47 31.725 121.68 31.795 ;
    RECT 121.47 32.085 121.68 32.155 ;
    RECT 121.47 32.445 121.68 32.515 ;
    RECT 117.69 31.725 117.9 31.795 ;
    RECT 117.69 32.085 117.9 32.155 ;
    RECT 117.69 32.445 117.9 32.515 ;
    RECT 118.15 31.725 118.36 31.795 ;
    RECT 118.15 32.085 118.36 32.155 ;
    RECT 118.15 32.445 118.36 32.515 ;
    RECT 114.37 31.725 114.58 31.795 ;
    RECT 114.37 32.085 114.58 32.155 ;
    RECT 114.37 32.445 114.58 32.515 ;
    RECT 114.83 31.725 115.04 31.795 ;
    RECT 114.83 32.085 115.04 32.155 ;
    RECT 114.83 32.445 115.04 32.515 ;
    RECT 111.05 31.725 111.26 31.795 ;
    RECT 111.05 32.085 111.26 32.155 ;
    RECT 111.05 32.445 111.26 32.515 ;
    RECT 111.51 31.725 111.72 31.795 ;
    RECT 111.51 32.085 111.72 32.155 ;
    RECT 111.51 32.445 111.72 32.515 ;
    RECT 107.73 31.725 107.94 31.795 ;
    RECT 107.73 32.085 107.94 32.155 ;
    RECT 107.73 32.445 107.94 32.515 ;
    RECT 108.19 31.725 108.4 31.795 ;
    RECT 108.19 32.085 108.4 32.155 ;
    RECT 108.19 32.445 108.4 32.515 ;
    RECT 104.41 31.725 104.62 31.795 ;
    RECT 104.41 32.085 104.62 32.155 ;
    RECT 104.41 32.445 104.62 32.515 ;
    RECT 104.87 31.725 105.08 31.795 ;
    RECT 104.87 32.085 105.08 32.155 ;
    RECT 104.87 32.445 105.08 32.515 ;
    RECT 101.09 31.725 101.3 31.795 ;
    RECT 101.09 32.085 101.3 32.155 ;
    RECT 101.09 32.445 101.3 32.515 ;
    RECT 101.55 31.725 101.76 31.795 ;
    RECT 101.55 32.085 101.76 32.155 ;
    RECT 101.55 32.445 101.76 32.515 ;
    RECT 0.4 32.085 0.47 32.155 ;
    RECT 170.81 31.725 171.02 31.795 ;
    RECT 170.81 32.085 171.02 32.155 ;
    RECT 170.81 32.445 171.02 32.515 ;
    RECT 171.27 31.725 171.48 31.795 ;
    RECT 171.27 32.085 171.48 32.155 ;
    RECT 171.27 32.445 171.48 32.515 ;
    RECT 167.49 31.725 167.7 31.795 ;
    RECT 167.49 32.085 167.7 32.155 ;
    RECT 167.49 32.445 167.7 32.515 ;
    RECT 167.95 31.725 168.16 31.795 ;
    RECT 167.95 32.085 168.16 32.155 ;
    RECT 167.95 32.445 168.16 32.515 ;
    RECT 97.77 31.725 97.98 31.795 ;
    RECT 97.77 32.085 97.98 32.155 ;
    RECT 97.77 32.445 97.98 32.515 ;
    RECT 98.23 31.725 98.44 31.795 ;
    RECT 98.23 32.085 98.44 32.155 ;
    RECT 98.23 32.445 98.44 32.515 ;
    RECT 94.45 31.725 94.66 31.795 ;
    RECT 94.45 32.085 94.66 32.155 ;
    RECT 94.45 32.445 94.66 32.515 ;
    RECT 94.91 31.725 95.12 31.795 ;
    RECT 94.91 32.085 95.12 32.155 ;
    RECT 94.91 32.445 95.12 32.515 ;
    RECT 91.13 31.725 91.34 31.795 ;
    RECT 91.13 32.085 91.34 32.155 ;
    RECT 91.13 32.445 91.34 32.515 ;
    RECT 91.59 31.725 91.8 31.795 ;
    RECT 91.59 32.085 91.8 32.155 ;
    RECT 91.59 32.445 91.8 32.515 ;
    RECT 87.81 31.725 88.02 31.795 ;
    RECT 87.81 32.085 88.02 32.155 ;
    RECT 87.81 32.445 88.02 32.515 ;
    RECT 88.27 31.725 88.48 31.795 ;
    RECT 88.27 32.085 88.48 32.155 ;
    RECT 88.27 32.445 88.48 32.515 ;
    RECT 84.49 31.725 84.7 31.795 ;
    RECT 84.49 32.085 84.7 32.155 ;
    RECT 84.49 32.445 84.7 32.515 ;
    RECT 84.95 31.725 85.16 31.795 ;
    RECT 84.95 32.085 85.16 32.155 ;
    RECT 84.95 32.445 85.16 32.515 ;
    RECT 81.17 31.725 81.38 31.795 ;
    RECT 81.17 32.085 81.38 32.155 ;
    RECT 81.17 32.445 81.38 32.515 ;
    RECT 81.63 31.725 81.84 31.795 ;
    RECT 81.63 32.085 81.84 32.155 ;
    RECT 81.63 32.445 81.84 32.515 ;
    RECT 77.85 31.725 78.06 31.795 ;
    RECT 77.85 32.085 78.06 32.155 ;
    RECT 77.85 32.445 78.06 32.515 ;
    RECT 78.31 31.725 78.52 31.795 ;
    RECT 78.31 32.085 78.52 32.155 ;
    RECT 78.31 32.445 78.52 32.515 ;
    RECT 74.53 31.725 74.74 31.795 ;
    RECT 74.53 32.085 74.74 32.155 ;
    RECT 74.53 32.445 74.74 32.515 ;
    RECT 74.99 31.725 75.2 31.795 ;
    RECT 74.99 32.085 75.2 32.155 ;
    RECT 74.99 32.445 75.2 32.515 ;
    RECT 71.21 31.725 71.42 31.795 ;
    RECT 71.21 32.085 71.42 32.155 ;
    RECT 71.21 32.445 71.42 32.515 ;
    RECT 71.67 31.725 71.88 31.795 ;
    RECT 71.67 32.085 71.88 32.155 ;
    RECT 71.67 32.445 71.88 32.515 ;
    RECT 31.37 31.725 31.58 31.795 ;
    RECT 31.37 32.085 31.58 32.155 ;
    RECT 31.37 32.445 31.58 32.515 ;
    RECT 31.83 31.725 32.04 31.795 ;
    RECT 31.83 32.085 32.04 32.155 ;
    RECT 31.83 32.445 32.04 32.515 ;
    RECT 67.89 31.725 68.1 31.795 ;
    RECT 67.89 32.085 68.1 32.155 ;
    RECT 67.89 32.445 68.1 32.515 ;
    RECT 68.35 31.725 68.56 31.795 ;
    RECT 68.35 32.085 68.56 32.155 ;
    RECT 68.35 32.445 68.56 32.515 ;
    RECT 28.05 31.725 28.26 31.795 ;
    RECT 28.05 32.085 28.26 32.155 ;
    RECT 28.05 32.445 28.26 32.515 ;
    RECT 28.51 31.725 28.72 31.795 ;
    RECT 28.51 32.085 28.72 32.155 ;
    RECT 28.51 32.445 28.72 32.515 ;
    RECT 24.73 31.725 24.94 31.795 ;
    RECT 24.73 32.085 24.94 32.155 ;
    RECT 24.73 32.445 24.94 32.515 ;
    RECT 25.19 31.725 25.4 31.795 ;
    RECT 25.19 32.085 25.4 32.155 ;
    RECT 25.19 32.445 25.4 32.515 ;
    RECT 21.41 31.725 21.62 31.795 ;
    RECT 21.41 32.085 21.62 32.155 ;
    RECT 21.41 32.445 21.62 32.515 ;
    RECT 21.87 31.725 22.08 31.795 ;
    RECT 21.87 32.085 22.08 32.155 ;
    RECT 21.87 32.445 22.08 32.515 ;
    RECT 18.09 31.725 18.3 31.795 ;
    RECT 18.09 32.085 18.3 32.155 ;
    RECT 18.09 32.445 18.3 32.515 ;
    RECT 18.55 31.725 18.76 31.795 ;
    RECT 18.55 32.085 18.76 32.155 ;
    RECT 18.55 32.445 18.76 32.515 ;
    RECT 14.77 31.725 14.98 31.795 ;
    RECT 14.77 32.085 14.98 32.155 ;
    RECT 14.77 32.445 14.98 32.515 ;
    RECT 15.23 31.725 15.44 31.795 ;
    RECT 15.23 32.085 15.44 32.155 ;
    RECT 15.23 32.445 15.44 32.515 ;
    RECT 11.45 31.725 11.66 31.795 ;
    RECT 11.45 32.085 11.66 32.155 ;
    RECT 11.45 32.445 11.66 32.515 ;
    RECT 11.91 31.725 12.12 31.795 ;
    RECT 11.91 32.085 12.12 32.155 ;
    RECT 11.91 32.445 12.12 32.515 ;
    RECT 8.13 31.725 8.34 31.795 ;
    RECT 8.13 32.085 8.34 32.155 ;
    RECT 8.13 32.445 8.34 32.515 ;
    RECT 8.59 31.725 8.8 31.795 ;
    RECT 8.59 32.085 8.8 32.155 ;
    RECT 8.59 32.445 8.8 32.515 ;
    RECT 4.81 31.725 5.02 31.795 ;
    RECT 4.81 32.085 5.02 32.155 ;
    RECT 4.81 32.445 5.02 32.515 ;
    RECT 5.27 31.725 5.48 31.795 ;
    RECT 5.27 32.085 5.48 32.155 ;
    RECT 5.27 32.445 5.48 32.515 ;
    RECT 164.17 31.725 164.38 31.795 ;
    RECT 164.17 32.085 164.38 32.155 ;
    RECT 164.17 32.445 164.38 32.515 ;
    RECT 164.63 31.725 164.84 31.795 ;
    RECT 164.63 32.085 164.84 32.155 ;
    RECT 164.63 32.445 164.84 32.515 ;
    RECT 1.49 31.725 1.7 31.795 ;
    RECT 1.49 32.085 1.7 32.155 ;
    RECT 1.49 32.445 1.7 32.515 ;
    RECT 1.95 31.725 2.16 31.795 ;
    RECT 1.95 32.085 2.16 32.155 ;
    RECT 1.95 32.445 2.16 32.515 ;
    RECT 160.85 31.725 161.06 31.795 ;
    RECT 160.85 32.085 161.06 32.155 ;
    RECT 160.85 32.445 161.06 32.515 ;
    RECT 161.31 31.725 161.52 31.795 ;
    RECT 161.31 32.085 161.52 32.155 ;
    RECT 161.31 32.445 161.52 32.515 ;
    RECT 157.53 31.725 157.74 31.795 ;
    RECT 157.53 32.085 157.74 32.155 ;
    RECT 157.53 32.445 157.74 32.515 ;
    RECT 157.99 31.725 158.2 31.795 ;
    RECT 157.99 32.085 158.2 32.155 ;
    RECT 157.99 32.445 158.2 32.515 ;
    RECT 154.21 31.725 154.42 31.795 ;
    RECT 154.21 32.085 154.42 32.155 ;
    RECT 154.21 32.445 154.42 32.515 ;
    RECT 154.67 31.725 154.88 31.795 ;
    RECT 154.67 32.085 154.88 32.155 ;
    RECT 154.67 32.445 154.88 32.515 ;
    RECT 150.89 31.725 151.1 31.795 ;
    RECT 150.89 32.085 151.1 32.155 ;
    RECT 150.89 32.445 151.1 32.515 ;
    RECT 151.35 31.725 151.56 31.795 ;
    RECT 151.35 32.085 151.56 32.155 ;
    RECT 151.35 32.445 151.56 32.515 ;
    RECT 147.57 31.725 147.78 31.795 ;
    RECT 147.57 32.085 147.78 32.155 ;
    RECT 147.57 32.445 147.78 32.515 ;
    RECT 148.03 31.725 148.24 31.795 ;
    RECT 148.03 32.085 148.24 32.155 ;
    RECT 148.03 32.445 148.24 32.515 ;
    RECT 144.25 31.725 144.46 31.795 ;
    RECT 144.25 32.085 144.46 32.155 ;
    RECT 144.25 32.445 144.46 32.515 ;
    RECT 144.71 31.725 144.92 31.795 ;
    RECT 144.71 32.085 144.92 32.155 ;
    RECT 144.71 32.445 144.92 32.515 ;
    RECT 140.93 31.725 141.14 31.795 ;
    RECT 140.93 32.085 141.14 32.155 ;
    RECT 140.93 32.445 141.14 32.515 ;
    RECT 141.39 31.725 141.6 31.795 ;
    RECT 141.39 32.085 141.6 32.155 ;
    RECT 141.39 32.445 141.6 32.515 ;
    RECT 137.61 31.725 137.82 31.795 ;
    RECT 137.61 32.085 137.82 32.155 ;
    RECT 137.61 32.445 137.82 32.515 ;
    RECT 138.07 31.725 138.28 31.795 ;
    RECT 138.07 32.085 138.28 32.155 ;
    RECT 138.07 32.445 138.28 32.515 ;
    RECT 134.29 31.725 134.5 31.795 ;
    RECT 134.29 32.085 134.5 32.155 ;
    RECT 134.29 32.445 134.5 32.515 ;
    RECT 134.75 31.725 134.96 31.795 ;
    RECT 134.75 32.085 134.96 32.155 ;
    RECT 134.75 32.445 134.96 32.515 ;
    RECT 64.57 31.725 64.78 31.795 ;
    RECT 64.57 32.085 64.78 32.155 ;
    RECT 64.57 32.445 64.78 32.515 ;
    RECT 65.03 31.725 65.24 31.795 ;
    RECT 65.03 32.085 65.24 32.155 ;
    RECT 65.03 32.445 65.24 32.515 ;
    RECT 61.25 31.005 61.46 31.075 ;
    RECT 61.25 31.365 61.46 31.435 ;
    RECT 61.25 31.725 61.46 31.795 ;
    RECT 61.71 31.005 61.92 31.075 ;
    RECT 61.71 31.365 61.92 31.435 ;
    RECT 61.71 31.725 61.92 31.795 ;
    RECT 57.93 31.005 58.14 31.075 ;
    RECT 57.93 31.365 58.14 31.435 ;
    RECT 57.93 31.725 58.14 31.795 ;
    RECT 58.39 31.005 58.6 31.075 ;
    RECT 58.39 31.365 58.6 31.435 ;
    RECT 58.39 31.725 58.6 31.795 ;
    RECT 54.61 31.005 54.82 31.075 ;
    RECT 54.61 31.365 54.82 31.435 ;
    RECT 54.61 31.725 54.82 31.795 ;
    RECT 55.07 31.005 55.28 31.075 ;
    RECT 55.07 31.365 55.28 31.435 ;
    RECT 55.07 31.725 55.28 31.795 ;
    RECT 51.29 31.005 51.5 31.075 ;
    RECT 51.29 31.365 51.5 31.435 ;
    RECT 51.29 31.725 51.5 31.795 ;
    RECT 51.75 31.005 51.96 31.075 ;
    RECT 51.75 31.365 51.96 31.435 ;
    RECT 51.75 31.725 51.96 31.795 ;
    RECT 47.97 31.005 48.18 31.075 ;
    RECT 47.97 31.365 48.18 31.435 ;
    RECT 47.97 31.725 48.18 31.795 ;
    RECT 48.43 31.005 48.64 31.075 ;
    RECT 48.43 31.365 48.64 31.435 ;
    RECT 48.43 31.725 48.64 31.795 ;
    RECT 44.65 31.005 44.86 31.075 ;
    RECT 44.65 31.365 44.86 31.435 ;
    RECT 44.65 31.725 44.86 31.795 ;
    RECT 45.11 31.005 45.32 31.075 ;
    RECT 45.11 31.365 45.32 31.435 ;
    RECT 45.11 31.725 45.32 31.795 ;
    RECT 41.33 31.005 41.54 31.075 ;
    RECT 41.33 31.365 41.54 31.435 ;
    RECT 41.33 31.725 41.54 31.795 ;
    RECT 41.79 31.005 42.0 31.075 ;
    RECT 41.79 31.365 42.0 31.435 ;
    RECT 41.79 31.725 42.0 31.795 ;
    RECT 38.01 31.005 38.22 31.075 ;
    RECT 38.01 31.365 38.22 31.435 ;
    RECT 38.01 31.725 38.22 31.795 ;
    RECT 38.47 31.005 38.68 31.075 ;
    RECT 38.47 31.365 38.68 31.435 ;
    RECT 38.47 31.725 38.68 31.795 ;
    RECT 34.69 31.005 34.9 31.075 ;
    RECT 34.69 31.365 34.9 31.435 ;
    RECT 34.69 31.725 34.9 31.795 ;
    RECT 35.15 31.005 35.36 31.075 ;
    RECT 35.15 31.365 35.36 31.435 ;
    RECT 35.15 31.725 35.36 31.795 ;
    RECT 173.945 31.365 174.015 31.435 ;
    RECT 130.97 31.005 131.18 31.075 ;
    RECT 130.97 31.365 131.18 31.435 ;
    RECT 130.97 31.725 131.18 31.795 ;
    RECT 131.43 31.005 131.64 31.075 ;
    RECT 131.43 31.365 131.64 31.435 ;
    RECT 131.43 31.725 131.64 31.795 ;
    RECT 127.65 31.005 127.86 31.075 ;
    RECT 127.65 31.365 127.86 31.435 ;
    RECT 127.65 31.725 127.86 31.795 ;
    RECT 128.11 31.005 128.32 31.075 ;
    RECT 128.11 31.365 128.32 31.435 ;
    RECT 128.11 31.725 128.32 31.795 ;
    RECT 124.33 31.005 124.54 31.075 ;
    RECT 124.33 31.365 124.54 31.435 ;
    RECT 124.33 31.725 124.54 31.795 ;
    RECT 124.79 31.005 125.0 31.075 ;
    RECT 124.79 31.365 125.0 31.435 ;
    RECT 124.79 31.725 125.0 31.795 ;
    RECT 121.01 31.005 121.22 31.075 ;
    RECT 121.01 31.365 121.22 31.435 ;
    RECT 121.01 31.725 121.22 31.795 ;
    RECT 121.47 31.005 121.68 31.075 ;
    RECT 121.47 31.365 121.68 31.435 ;
    RECT 121.47 31.725 121.68 31.795 ;
    RECT 117.69 31.005 117.9 31.075 ;
    RECT 117.69 31.365 117.9 31.435 ;
    RECT 117.69 31.725 117.9 31.795 ;
    RECT 118.15 31.005 118.36 31.075 ;
    RECT 118.15 31.365 118.36 31.435 ;
    RECT 118.15 31.725 118.36 31.795 ;
    RECT 114.37 31.005 114.58 31.075 ;
    RECT 114.37 31.365 114.58 31.435 ;
    RECT 114.37 31.725 114.58 31.795 ;
    RECT 114.83 31.005 115.04 31.075 ;
    RECT 114.83 31.365 115.04 31.435 ;
    RECT 114.83 31.725 115.04 31.795 ;
    RECT 111.05 31.005 111.26 31.075 ;
    RECT 111.05 31.365 111.26 31.435 ;
    RECT 111.05 31.725 111.26 31.795 ;
    RECT 111.51 31.005 111.72 31.075 ;
    RECT 111.51 31.365 111.72 31.435 ;
    RECT 111.51 31.725 111.72 31.795 ;
    RECT 107.73 31.005 107.94 31.075 ;
    RECT 107.73 31.365 107.94 31.435 ;
    RECT 107.73 31.725 107.94 31.795 ;
    RECT 108.19 31.005 108.4 31.075 ;
    RECT 108.19 31.365 108.4 31.435 ;
    RECT 108.19 31.725 108.4 31.795 ;
    RECT 104.41 31.005 104.62 31.075 ;
    RECT 104.41 31.365 104.62 31.435 ;
    RECT 104.41 31.725 104.62 31.795 ;
    RECT 104.87 31.005 105.08 31.075 ;
    RECT 104.87 31.365 105.08 31.435 ;
    RECT 104.87 31.725 105.08 31.795 ;
    RECT 101.09 31.005 101.3 31.075 ;
    RECT 101.09 31.365 101.3 31.435 ;
    RECT 101.09 31.725 101.3 31.795 ;
    RECT 101.55 31.005 101.76 31.075 ;
    RECT 101.55 31.365 101.76 31.435 ;
    RECT 101.55 31.725 101.76 31.795 ;
    RECT 0.4 31.365 0.47 31.435 ;
    RECT 170.81 31.005 171.02 31.075 ;
    RECT 170.81 31.365 171.02 31.435 ;
    RECT 170.81 31.725 171.02 31.795 ;
    RECT 171.27 31.005 171.48 31.075 ;
    RECT 171.27 31.365 171.48 31.435 ;
    RECT 171.27 31.725 171.48 31.795 ;
    RECT 167.49 31.005 167.7 31.075 ;
    RECT 167.49 31.365 167.7 31.435 ;
    RECT 167.49 31.725 167.7 31.795 ;
    RECT 167.95 31.005 168.16 31.075 ;
    RECT 167.95 31.365 168.16 31.435 ;
    RECT 167.95 31.725 168.16 31.795 ;
    RECT 97.77 31.005 97.98 31.075 ;
    RECT 97.77 31.365 97.98 31.435 ;
    RECT 97.77 31.725 97.98 31.795 ;
    RECT 98.23 31.005 98.44 31.075 ;
    RECT 98.23 31.365 98.44 31.435 ;
    RECT 98.23 31.725 98.44 31.795 ;
    RECT 94.45 31.005 94.66 31.075 ;
    RECT 94.45 31.365 94.66 31.435 ;
    RECT 94.45 31.725 94.66 31.795 ;
    RECT 94.91 31.005 95.12 31.075 ;
    RECT 94.91 31.365 95.12 31.435 ;
    RECT 94.91 31.725 95.12 31.795 ;
    RECT 91.13 31.005 91.34 31.075 ;
    RECT 91.13 31.365 91.34 31.435 ;
    RECT 91.13 31.725 91.34 31.795 ;
    RECT 91.59 31.005 91.8 31.075 ;
    RECT 91.59 31.365 91.8 31.435 ;
    RECT 91.59 31.725 91.8 31.795 ;
    RECT 87.81 31.005 88.02 31.075 ;
    RECT 87.81 31.365 88.02 31.435 ;
    RECT 87.81 31.725 88.02 31.795 ;
    RECT 88.27 31.005 88.48 31.075 ;
    RECT 88.27 31.365 88.48 31.435 ;
    RECT 88.27 31.725 88.48 31.795 ;
    RECT 84.49 31.005 84.7 31.075 ;
    RECT 84.49 31.365 84.7 31.435 ;
    RECT 84.49 31.725 84.7 31.795 ;
    RECT 84.95 31.005 85.16 31.075 ;
    RECT 84.95 31.365 85.16 31.435 ;
    RECT 84.95 31.725 85.16 31.795 ;
    RECT 81.17 31.005 81.38 31.075 ;
    RECT 81.17 31.365 81.38 31.435 ;
    RECT 81.17 31.725 81.38 31.795 ;
    RECT 81.63 31.005 81.84 31.075 ;
    RECT 81.63 31.365 81.84 31.435 ;
    RECT 81.63 31.725 81.84 31.795 ;
    RECT 77.85 31.005 78.06 31.075 ;
    RECT 77.85 31.365 78.06 31.435 ;
    RECT 77.85 31.725 78.06 31.795 ;
    RECT 78.31 31.005 78.52 31.075 ;
    RECT 78.31 31.365 78.52 31.435 ;
    RECT 78.31 31.725 78.52 31.795 ;
    RECT 74.53 31.005 74.74 31.075 ;
    RECT 74.53 31.365 74.74 31.435 ;
    RECT 74.53 31.725 74.74 31.795 ;
    RECT 74.99 31.005 75.2 31.075 ;
    RECT 74.99 31.365 75.2 31.435 ;
    RECT 74.99 31.725 75.2 31.795 ;
    RECT 71.21 31.005 71.42 31.075 ;
    RECT 71.21 31.365 71.42 31.435 ;
    RECT 71.21 31.725 71.42 31.795 ;
    RECT 71.67 31.005 71.88 31.075 ;
    RECT 71.67 31.365 71.88 31.435 ;
    RECT 71.67 31.725 71.88 31.795 ;
    RECT 31.37 31.005 31.58 31.075 ;
    RECT 31.37 31.365 31.58 31.435 ;
    RECT 31.37 31.725 31.58 31.795 ;
    RECT 31.83 31.005 32.04 31.075 ;
    RECT 31.83 31.365 32.04 31.435 ;
    RECT 31.83 31.725 32.04 31.795 ;
    RECT 67.89 31.005 68.1 31.075 ;
    RECT 67.89 31.365 68.1 31.435 ;
    RECT 67.89 31.725 68.1 31.795 ;
    RECT 68.35 31.005 68.56 31.075 ;
    RECT 68.35 31.365 68.56 31.435 ;
    RECT 68.35 31.725 68.56 31.795 ;
    RECT 28.05 31.005 28.26 31.075 ;
    RECT 28.05 31.365 28.26 31.435 ;
    RECT 28.05 31.725 28.26 31.795 ;
    RECT 28.51 31.005 28.72 31.075 ;
    RECT 28.51 31.365 28.72 31.435 ;
    RECT 28.51 31.725 28.72 31.795 ;
    RECT 24.73 31.005 24.94 31.075 ;
    RECT 24.73 31.365 24.94 31.435 ;
    RECT 24.73 31.725 24.94 31.795 ;
    RECT 25.19 31.005 25.4 31.075 ;
    RECT 25.19 31.365 25.4 31.435 ;
    RECT 25.19 31.725 25.4 31.795 ;
    RECT 21.41 31.005 21.62 31.075 ;
    RECT 21.41 31.365 21.62 31.435 ;
    RECT 21.41 31.725 21.62 31.795 ;
    RECT 21.87 31.005 22.08 31.075 ;
    RECT 21.87 31.365 22.08 31.435 ;
    RECT 21.87 31.725 22.08 31.795 ;
    RECT 18.09 31.005 18.3 31.075 ;
    RECT 18.09 31.365 18.3 31.435 ;
    RECT 18.09 31.725 18.3 31.795 ;
    RECT 18.55 31.005 18.76 31.075 ;
    RECT 18.55 31.365 18.76 31.435 ;
    RECT 18.55 31.725 18.76 31.795 ;
    RECT 14.77 31.005 14.98 31.075 ;
    RECT 14.77 31.365 14.98 31.435 ;
    RECT 14.77 31.725 14.98 31.795 ;
    RECT 15.23 31.005 15.44 31.075 ;
    RECT 15.23 31.365 15.44 31.435 ;
    RECT 15.23 31.725 15.44 31.795 ;
    RECT 11.45 31.005 11.66 31.075 ;
    RECT 11.45 31.365 11.66 31.435 ;
    RECT 11.45 31.725 11.66 31.795 ;
    RECT 11.91 31.005 12.12 31.075 ;
    RECT 11.91 31.365 12.12 31.435 ;
    RECT 11.91 31.725 12.12 31.795 ;
    RECT 8.13 31.005 8.34 31.075 ;
    RECT 8.13 31.365 8.34 31.435 ;
    RECT 8.13 31.725 8.34 31.795 ;
    RECT 8.59 31.005 8.8 31.075 ;
    RECT 8.59 31.365 8.8 31.435 ;
    RECT 8.59 31.725 8.8 31.795 ;
    RECT 4.81 31.005 5.02 31.075 ;
    RECT 4.81 31.365 5.02 31.435 ;
    RECT 4.81 31.725 5.02 31.795 ;
    RECT 5.27 31.005 5.48 31.075 ;
    RECT 5.27 31.365 5.48 31.435 ;
    RECT 5.27 31.725 5.48 31.795 ;
    RECT 164.17 31.005 164.38 31.075 ;
    RECT 164.17 31.365 164.38 31.435 ;
    RECT 164.17 31.725 164.38 31.795 ;
    RECT 164.63 31.005 164.84 31.075 ;
    RECT 164.63 31.365 164.84 31.435 ;
    RECT 164.63 31.725 164.84 31.795 ;
    RECT 1.49 31.005 1.7 31.075 ;
    RECT 1.49 31.365 1.7 31.435 ;
    RECT 1.49 31.725 1.7 31.795 ;
    RECT 1.95 31.005 2.16 31.075 ;
    RECT 1.95 31.365 2.16 31.435 ;
    RECT 1.95 31.725 2.16 31.795 ;
    RECT 160.85 31.005 161.06 31.075 ;
    RECT 160.85 31.365 161.06 31.435 ;
    RECT 160.85 31.725 161.06 31.795 ;
    RECT 161.31 31.005 161.52 31.075 ;
    RECT 161.31 31.365 161.52 31.435 ;
    RECT 161.31 31.725 161.52 31.795 ;
    RECT 157.53 31.005 157.74 31.075 ;
    RECT 157.53 31.365 157.74 31.435 ;
    RECT 157.53 31.725 157.74 31.795 ;
    RECT 157.99 31.005 158.2 31.075 ;
    RECT 157.99 31.365 158.2 31.435 ;
    RECT 157.99 31.725 158.2 31.795 ;
    RECT 154.21 31.005 154.42 31.075 ;
    RECT 154.21 31.365 154.42 31.435 ;
    RECT 154.21 31.725 154.42 31.795 ;
    RECT 154.67 31.005 154.88 31.075 ;
    RECT 154.67 31.365 154.88 31.435 ;
    RECT 154.67 31.725 154.88 31.795 ;
    RECT 150.89 31.005 151.1 31.075 ;
    RECT 150.89 31.365 151.1 31.435 ;
    RECT 150.89 31.725 151.1 31.795 ;
    RECT 151.35 31.005 151.56 31.075 ;
    RECT 151.35 31.365 151.56 31.435 ;
    RECT 151.35 31.725 151.56 31.795 ;
    RECT 147.57 31.005 147.78 31.075 ;
    RECT 147.57 31.365 147.78 31.435 ;
    RECT 147.57 31.725 147.78 31.795 ;
    RECT 148.03 31.005 148.24 31.075 ;
    RECT 148.03 31.365 148.24 31.435 ;
    RECT 148.03 31.725 148.24 31.795 ;
    RECT 144.25 31.005 144.46 31.075 ;
    RECT 144.25 31.365 144.46 31.435 ;
    RECT 144.25 31.725 144.46 31.795 ;
    RECT 144.71 31.005 144.92 31.075 ;
    RECT 144.71 31.365 144.92 31.435 ;
    RECT 144.71 31.725 144.92 31.795 ;
    RECT 140.93 31.005 141.14 31.075 ;
    RECT 140.93 31.365 141.14 31.435 ;
    RECT 140.93 31.725 141.14 31.795 ;
    RECT 141.39 31.005 141.6 31.075 ;
    RECT 141.39 31.365 141.6 31.435 ;
    RECT 141.39 31.725 141.6 31.795 ;
    RECT 137.61 31.005 137.82 31.075 ;
    RECT 137.61 31.365 137.82 31.435 ;
    RECT 137.61 31.725 137.82 31.795 ;
    RECT 138.07 31.005 138.28 31.075 ;
    RECT 138.07 31.365 138.28 31.435 ;
    RECT 138.07 31.725 138.28 31.795 ;
    RECT 134.29 31.005 134.5 31.075 ;
    RECT 134.29 31.365 134.5 31.435 ;
    RECT 134.29 31.725 134.5 31.795 ;
    RECT 134.75 31.005 134.96 31.075 ;
    RECT 134.75 31.365 134.96 31.435 ;
    RECT 134.75 31.725 134.96 31.795 ;
    RECT 64.57 31.005 64.78 31.075 ;
    RECT 64.57 31.365 64.78 31.435 ;
    RECT 64.57 31.725 64.78 31.795 ;
    RECT 65.03 31.005 65.24 31.075 ;
    RECT 65.03 31.365 65.24 31.435 ;
    RECT 65.03 31.725 65.24 31.795 ;
    RECT 61.25 30.285 61.46 30.355 ;
    RECT 61.25 30.645 61.46 30.715 ;
    RECT 61.25 31.005 61.46 31.075 ;
    RECT 61.71 30.285 61.92 30.355 ;
    RECT 61.71 30.645 61.92 30.715 ;
    RECT 61.71 31.005 61.92 31.075 ;
    RECT 57.93 30.285 58.14 30.355 ;
    RECT 57.93 30.645 58.14 30.715 ;
    RECT 57.93 31.005 58.14 31.075 ;
    RECT 58.39 30.285 58.6 30.355 ;
    RECT 58.39 30.645 58.6 30.715 ;
    RECT 58.39 31.005 58.6 31.075 ;
    RECT 54.61 30.285 54.82 30.355 ;
    RECT 54.61 30.645 54.82 30.715 ;
    RECT 54.61 31.005 54.82 31.075 ;
    RECT 55.07 30.285 55.28 30.355 ;
    RECT 55.07 30.645 55.28 30.715 ;
    RECT 55.07 31.005 55.28 31.075 ;
    RECT 51.29 30.285 51.5 30.355 ;
    RECT 51.29 30.645 51.5 30.715 ;
    RECT 51.29 31.005 51.5 31.075 ;
    RECT 51.75 30.285 51.96 30.355 ;
    RECT 51.75 30.645 51.96 30.715 ;
    RECT 51.75 31.005 51.96 31.075 ;
    RECT 47.97 30.285 48.18 30.355 ;
    RECT 47.97 30.645 48.18 30.715 ;
    RECT 47.97 31.005 48.18 31.075 ;
    RECT 48.43 30.285 48.64 30.355 ;
    RECT 48.43 30.645 48.64 30.715 ;
    RECT 48.43 31.005 48.64 31.075 ;
    RECT 44.65 30.285 44.86 30.355 ;
    RECT 44.65 30.645 44.86 30.715 ;
    RECT 44.65 31.005 44.86 31.075 ;
    RECT 45.11 30.285 45.32 30.355 ;
    RECT 45.11 30.645 45.32 30.715 ;
    RECT 45.11 31.005 45.32 31.075 ;
    RECT 41.33 30.285 41.54 30.355 ;
    RECT 41.33 30.645 41.54 30.715 ;
    RECT 41.33 31.005 41.54 31.075 ;
    RECT 41.79 30.285 42.0 30.355 ;
    RECT 41.79 30.645 42.0 30.715 ;
    RECT 41.79 31.005 42.0 31.075 ;
    RECT 38.01 30.285 38.22 30.355 ;
    RECT 38.01 30.645 38.22 30.715 ;
    RECT 38.01 31.005 38.22 31.075 ;
    RECT 38.47 30.285 38.68 30.355 ;
    RECT 38.47 30.645 38.68 30.715 ;
    RECT 38.47 31.005 38.68 31.075 ;
    RECT 34.69 30.285 34.9 30.355 ;
    RECT 34.69 30.645 34.9 30.715 ;
    RECT 34.69 31.005 34.9 31.075 ;
    RECT 35.15 30.285 35.36 30.355 ;
    RECT 35.15 30.645 35.36 30.715 ;
    RECT 35.15 31.005 35.36 31.075 ;
    RECT 173.945 30.645 174.015 30.715 ;
    RECT 130.97 30.285 131.18 30.355 ;
    RECT 130.97 30.645 131.18 30.715 ;
    RECT 130.97 31.005 131.18 31.075 ;
    RECT 131.43 30.285 131.64 30.355 ;
    RECT 131.43 30.645 131.64 30.715 ;
    RECT 131.43 31.005 131.64 31.075 ;
    RECT 127.65 30.285 127.86 30.355 ;
    RECT 127.65 30.645 127.86 30.715 ;
    RECT 127.65 31.005 127.86 31.075 ;
    RECT 128.11 30.285 128.32 30.355 ;
    RECT 128.11 30.645 128.32 30.715 ;
    RECT 128.11 31.005 128.32 31.075 ;
    RECT 124.33 30.285 124.54 30.355 ;
    RECT 124.33 30.645 124.54 30.715 ;
    RECT 124.33 31.005 124.54 31.075 ;
    RECT 124.79 30.285 125.0 30.355 ;
    RECT 124.79 30.645 125.0 30.715 ;
    RECT 124.79 31.005 125.0 31.075 ;
    RECT 121.01 30.285 121.22 30.355 ;
    RECT 121.01 30.645 121.22 30.715 ;
    RECT 121.01 31.005 121.22 31.075 ;
    RECT 121.47 30.285 121.68 30.355 ;
    RECT 121.47 30.645 121.68 30.715 ;
    RECT 121.47 31.005 121.68 31.075 ;
    RECT 117.69 30.285 117.9 30.355 ;
    RECT 117.69 30.645 117.9 30.715 ;
    RECT 117.69 31.005 117.9 31.075 ;
    RECT 118.15 30.285 118.36 30.355 ;
    RECT 118.15 30.645 118.36 30.715 ;
    RECT 118.15 31.005 118.36 31.075 ;
    RECT 114.37 30.285 114.58 30.355 ;
    RECT 114.37 30.645 114.58 30.715 ;
    RECT 114.37 31.005 114.58 31.075 ;
    RECT 114.83 30.285 115.04 30.355 ;
    RECT 114.83 30.645 115.04 30.715 ;
    RECT 114.83 31.005 115.04 31.075 ;
    RECT 111.05 30.285 111.26 30.355 ;
    RECT 111.05 30.645 111.26 30.715 ;
    RECT 111.05 31.005 111.26 31.075 ;
    RECT 111.51 30.285 111.72 30.355 ;
    RECT 111.51 30.645 111.72 30.715 ;
    RECT 111.51 31.005 111.72 31.075 ;
    RECT 107.73 30.285 107.94 30.355 ;
    RECT 107.73 30.645 107.94 30.715 ;
    RECT 107.73 31.005 107.94 31.075 ;
    RECT 108.19 30.285 108.4 30.355 ;
    RECT 108.19 30.645 108.4 30.715 ;
    RECT 108.19 31.005 108.4 31.075 ;
    RECT 104.41 30.285 104.62 30.355 ;
    RECT 104.41 30.645 104.62 30.715 ;
    RECT 104.41 31.005 104.62 31.075 ;
    RECT 104.87 30.285 105.08 30.355 ;
    RECT 104.87 30.645 105.08 30.715 ;
    RECT 104.87 31.005 105.08 31.075 ;
    RECT 101.09 30.285 101.3 30.355 ;
    RECT 101.09 30.645 101.3 30.715 ;
    RECT 101.09 31.005 101.3 31.075 ;
    RECT 101.55 30.285 101.76 30.355 ;
    RECT 101.55 30.645 101.76 30.715 ;
    RECT 101.55 31.005 101.76 31.075 ;
    RECT 0.4 30.645 0.47 30.715 ;
    RECT 170.81 30.285 171.02 30.355 ;
    RECT 170.81 30.645 171.02 30.715 ;
    RECT 170.81 31.005 171.02 31.075 ;
    RECT 171.27 30.285 171.48 30.355 ;
    RECT 171.27 30.645 171.48 30.715 ;
    RECT 171.27 31.005 171.48 31.075 ;
    RECT 167.49 30.285 167.7 30.355 ;
    RECT 167.49 30.645 167.7 30.715 ;
    RECT 167.49 31.005 167.7 31.075 ;
    RECT 167.95 30.285 168.16 30.355 ;
    RECT 167.95 30.645 168.16 30.715 ;
    RECT 167.95 31.005 168.16 31.075 ;
    RECT 97.77 30.285 97.98 30.355 ;
    RECT 97.77 30.645 97.98 30.715 ;
    RECT 97.77 31.005 97.98 31.075 ;
    RECT 98.23 30.285 98.44 30.355 ;
    RECT 98.23 30.645 98.44 30.715 ;
    RECT 98.23 31.005 98.44 31.075 ;
    RECT 94.45 30.285 94.66 30.355 ;
    RECT 94.45 30.645 94.66 30.715 ;
    RECT 94.45 31.005 94.66 31.075 ;
    RECT 94.91 30.285 95.12 30.355 ;
    RECT 94.91 30.645 95.12 30.715 ;
    RECT 94.91 31.005 95.12 31.075 ;
    RECT 91.13 30.285 91.34 30.355 ;
    RECT 91.13 30.645 91.34 30.715 ;
    RECT 91.13 31.005 91.34 31.075 ;
    RECT 91.59 30.285 91.8 30.355 ;
    RECT 91.59 30.645 91.8 30.715 ;
    RECT 91.59 31.005 91.8 31.075 ;
    RECT 87.81 30.285 88.02 30.355 ;
    RECT 87.81 30.645 88.02 30.715 ;
    RECT 87.81 31.005 88.02 31.075 ;
    RECT 88.27 30.285 88.48 30.355 ;
    RECT 88.27 30.645 88.48 30.715 ;
    RECT 88.27 31.005 88.48 31.075 ;
    RECT 84.49 30.285 84.7 30.355 ;
    RECT 84.49 30.645 84.7 30.715 ;
    RECT 84.49 31.005 84.7 31.075 ;
    RECT 84.95 30.285 85.16 30.355 ;
    RECT 84.95 30.645 85.16 30.715 ;
    RECT 84.95 31.005 85.16 31.075 ;
    RECT 81.17 30.285 81.38 30.355 ;
    RECT 81.17 30.645 81.38 30.715 ;
    RECT 81.17 31.005 81.38 31.075 ;
    RECT 81.63 30.285 81.84 30.355 ;
    RECT 81.63 30.645 81.84 30.715 ;
    RECT 81.63 31.005 81.84 31.075 ;
    RECT 77.85 30.285 78.06 30.355 ;
    RECT 77.85 30.645 78.06 30.715 ;
    RECT 77.85 31.005 78.06 31.075 ;
    RECT 78.31 30.285 78.52 30.355 ;
    RECT 78.31 30.645 78.52 30.715 ;
    RECT 78.31 31.005 78.52 31.075 ;
    RECT 74.53 30.285 74.74 30.355 ;
    RECT 74.53 30.645 74.74 30.715 ;
    RECT 74.53 31.005 74.74 31.075 ;
    RECT 74.99 30.285 75.2 30.355 ;
    RECT 74.99 30.645 75.2 30.715 ;
    RECT 74.99 31.005 75.2 31.075 ;
    RECT 71.21 30.285 71.42 30.355 ;
    RECT 71.21 30.645 71.42 30.715 ;
    RECT 71.21 31.005 71.42 31.075 ;
    RECT 71.67 30.285 71.88 30.355 ;
    RECT 71.67 30.645 71.88 30.715 ;
    RECT 71.67 31.005 71.88 31.075 ;
    RECT 31.37 30.285 31.58 30.355 ;
    RECT 31.37 30.645 31.58 30.715 ;
    RECT 31.37 31.005 31.58 31.075 ;
    RECT 31.83 30.285 32.04 30.355 ;
    RECT 31.83 30.645 32.04 30.715 ;
    RECT 31.83 31.005 32.04 31.075 ;
    RECT 67.89 30.285 68.1 30.355 ;
    RECT 67.89 30.645 68.1 30.715 ;
    RECT 67.89 31.005 68.1 31.075 ;
    RECT 68.35 30.285 68.56 30.355 ;
    RECT 68.35 30.645 68.56 30.715 ;
    RECT 68.35 31.005 68.56 31.075 ;
    RECT 28.05 30.285 28.26 30.355 ;
    RECT 28.05 30.645 28.26 30.715 ;
    RECT 28.05 31.005 28.26 31.075 ;
    RECT 28.51 30.285 28.72 30.355 ;
    RECT 28.51 30.645 28.72 30.715 ;
    RECT 28.51 31.005 28.72 31.075 ;
    RECT 24.73 30.285 24.94 30.355 ;
    RECT 24.73 30.645 24.94 30.715 ;
    RECT 24.73 31.005 24.94 31.075 ;
    RECT 25.19 30.285 25.4 30.355 ;
    RECT 25.19 30.645 25.4 30.715 ;
    RECT 25.19 31.005 25.4 31.075 ;
    RECT 21.41 30.285 21.62 30.355 ;
    RECT 21.41 30.645 21.62 30.715 ;
    RECT 21.41 31.005 21.62 31.075 ;
    RECT 21.87 30.285 22.08 30.355 ;
    RECT 21.87 30.645 22.08 30.715 ;
    RECT 21.87 31.005 22.08 31.075 ;
    RECT 18.09 30.285 18.3 30.355 ;
    RECT 18.09 30.645 18.3 30.715 ;
    RECT 18.09 31.005 18.3 31.075 ;
    RECT 18.55 30.285 18.76 30.355 ;
    RECT 18.55 30.645 18.76 30.715 ;
    RECT 18.55 31.005 18.76 31.075 ;
    RECT 14.77 30.285 14.98 30.355 ;
    RECT 14.77 30.645 14.98 30.715 ;
    RECT 14.77 31.005 14.98 31.075 ;
    RECT 15.23 30.285 15.44 30.355 ;
    RECT 15.23 30.645 15.44 30.715 ;
    RECT 15.23 31.005 15.44 31.075 ;
    RECT 11.45 30.285 11.66 30.355 ;
    RECT 11.45 30.645 11.66 30.715 ;
    RECT 11.45 31.005 11.66 31.075 ;
    RECT 11.91 30.285 12.12 30.355 ;
    RECT 11.91 30.645 12.12 30.715 ;
    RECT 11.91 31.005 12.12 31.075 ;
    RECT 8.13 30.285 8.34 30.355 ;
    RECT 8.13 30.645 8.34 30.715 ;
    RECT 8.13 31.005 8.34 31.075 ;
    RECT 8.59 30.285 8.8 30.355 ;
    RECT 8.59 30.645 8.8 30.715 ;
    RECT 8.59 31.005 8.8 31.075 ;
    RECT 4.81 30.285 5.02 30.355 ;
    RECT 4.81 30.645 5.02 30.715 ;
    RECT 4.81 31.005 5.02 31.075 ;
    RECT 5.27 30.285 5.48 30.355 ;
    RECT 5.27 30.645 5.48 30.715 ;
    RECT 5.27 31.005 5.48 31.075 ;
    RECT 164.17 30.285 164.38 30.355 ;
    RECT 164.17 30.645 164.38 30.715 ;
    RECT 164.17 31.005 164.38 31.075 ;
    RECT 164.63 30.285 164.84 30.355 ;
    RECT 164.63 30.645 164.84 30.715 ;
    RECT 164.63 31.005 164.84 31.075 ;
    RECT 1.49 30.285 1.7 30.355 ;
    RECT 1.49 30.645 1.7 30.715 ;
    RECT 1.49 31.005 1.7 31.075 ;
    RECT 1.95 30.285 2.16 30.355 ;
    RECT 1.95 30.645 2.16 30.715 ;
    RECT 1.95 31.005 2.16 31.075 ;
    RECT 160.85 30.285 161.06 30.355 ;
    RECT 160.85 30.645 161.06 30.715 ;
    RECT 160.85 31.005 161.06 31.075 ;
    RECT 161.31 30.285 161.52 30.355 ;
    RECT 161.31 30.645 161.52 30.715 ;
    RECT 161.31 31.005 161.52 31.075 ;
    RECT 157.53 30.285 157.74 30.355 ;
    RECT 157.53 30.645 157.74 30.715 ;
    RECT 157.53 31.005 157.74 31.075 ;
    RECT 157.99 30.285 158.2 30.355 ;
    RECT 157.99 30.645 158.2 30.715 ;
    RECT 157.99 31.005 158.2 31.075 ;
    RECT 154.21 30.285 154.42 30.355 ;
    RECT 154.21 30.645 154.42 30.715 ;
    RECT 154.21 31.005 154.42 31.075 ;
    RECT 154.67 30.285 154.88 30.355 ;
    RECT 154.67 30.645 154.88 30.715 ;
    RECT 154.67 31.005 154.88 31.075 ;
    RECT 150.89 30.285 151.1 30.355 ;
    RECT 150.89 30.645 151.1 30.715 ;
    RECT 150.89 31.005 151.1 31.075 ;
    RECT 151.35 30.285 151.56 30.355 ;
    RECT 151.35 30.645 151.56 30.715 ;
    RECT 151.35 31.005 151.56 31.075 ;
    RECT 147.57 30.285 147.78 30.355 ;
    RECT 147.57 30.645 147.78 30.715 ;
    RECT 147.57 31.005 147.78 31.075 ;
    RECT 148.03 30.285 148.24 30.355 ;
    RECT 148.03 30.645 148.24 30.715 ;
    RECT 148.03 31.005 148.24 31.075 ;
    RECT 144.25 30.285 144.46 30.355 ;
    RECT 144.25 30.645 144.46 30.715 ;
    RECT 144.25 31.005 144.46 31.075 ;
    RECT 144.71 30.285 144.92 30.355 ;
    RECT 144.71 30.645 144.92 30.715 ;
    RECT 144.71 31.005 144.92 31.075 ;
    RECT 140.93 30.285 141.14 30.355 ;
    RECT 140.93 30.645 141.14 30.715 ;
    RECT 140.93 31.005 141.14 31.075 ;
    RECT 141.39 30.285 141.6 30.355 ;
    RECT 141.39 30.645 141.6 30.715 ;
    RECT 141.39 31.005 141.6 31.075 ;
    RECT 137.61 30.285 137.82 30.355 ;
    RECT 137.61 30.645 137.82 30.715 ;
    RECT 137.61 31.005 137.82 31.075 ;
    RECT 138.07 30.285 138.28 30.355 ;
    RECT 138.07 30.645 138.28 30.715 ;
    RECT 138.07 31.005 138.28 31.075 ;
    RECT 134.29 30.285 134.5 30.355 ;
    RECT 134.29 30.645 134.5 30.715 ;
    RECT 134.29 31.005 134.5 31.075 ;
    RECT 134.75 30.285 134.96 30.355 ;
    RECT 134.75 30.645 134.96 30.715 ;
    RECT 134.75 31.005 134.96 31.075 ;
    RECT 64.57 30.285 64.78 30.355 ;
    RECT 64.57 30.645 64.78 30.715 ;
    RECT 64.57 31.005 64.78 31.075 ;
    RECT 65.03 30.285 65.24 30.355 ;
    RECT 65.03 30.645 65.24 30.715 ;
    RECT 65.03 31.005 65.24 31.075 ;
    RECT 61.25 29.565 61.46 29.635 ;
    RECT 61.25 29.925 61.46 29.995 ;
    RECT 61.25 30.285 61.46 30.355 ;
    RECT 61.71 29.565 61.92 29.635 ;
    RECT 61.71 29.925 61.92 29.995 ;
    RECT 61.71 30.285 61.92 30.355 ;
    RECT 57.93 29.565 58.14 29.635 ;
    RECT 57.93 29.925 58.14 29.995 ;
    RECT 57.93 30.285 58.14 30.355 ;
    RECT 58.39 29.565 58.6 29.635 ;
    RECT 58.39 29.925 58.6 29.995 ;
    RECT 58.39 30.285 58.6 30.355 ;
    RECT 54.61 29.565 54.82 29.635 ;
    RECT 54.61 29.925 54.82 29.995 ;
    RECT 54.61 30.285 54.82 30.355 ;
    RECT 55.07 29.565 55.28 29.635 ;
    RECT 55.07 29.925 55.28 29.995 ;
    RECT 55.07 30.285 55.28 30.355 ;
    RECT 51.29 29.565 51.5 29.635 ;
    RECT 51.29 29.925 51.5 29.995 ;
    RECT 51.29 30.285 51.5 30.355 ;
    RECT 51.75 29.565 51.96 29.635 ;
    RECT 51.75 29.925 51.96 29.995 ;
    RECT 51.75 30.285 51.96 30.355 ;
    RECT 47.97 29.565 48.18 29.635 ;
    RECT 47.97 29.925 48.18 29.995 ;
    RECT 47.97 30.285 48.18 30.355 ;
    RECT 48.43 29.565 48.64 29.635 ;
    RECT 48.43 29.925 48.64 29.995 ;
    RECT 48.43 30.285 48.64 30.355 ;
    RECT 44.65 29.565 44.86 29.635 ;
    RECT 44.65 29.925 44.86 29.995 ;
    RECT 44.65 30.285 44.86 30.355 ;
    RECT 45.11 29.565 45.32 29.635 ;
    RECT 45.11 29.925 45.32 29.995 ;
    RECT 45.11 30.285 45.32 30.355 ;
    RECT 41.33 29.565 41.54 29.635 ;
    RECT 41.33 29.925 41.54 29.995 ;
    RECT 41.33 30.285 41.54 30.355 ;
    RECT 41.79 29.565 42.0 29.635 ;
    RECT 41.79 29.925 42.0 29.995 ;
    RECT 41.79 30.285 42.0 30.355 ;
    RECT 38.01 29.565 38.22 29.635 ;
    RECT 38.01 29.925 38.22 29.995 ;
    RECT 38.01 30.285 38.22 30.355 ;
    RECT 38.47 29.565 38.68 29.635 ;
    RECT 38.47 29.925 38.68 29.995 ;
    RECT 38.47 30.285 38.68 30.355 ;
    RECT 34.69 29.565 34.9 29.635 ;
    RECT 34.69 29.925 34.9 29.995 ;
    RECT 34.69 30.285 34.9 30.355 ;
    RECT 35.15 29.565 35.36 29.635 ;
    RECT 35.15 29.925 35.36 29.995 ;
    RECT 35.15 30.285 35.36 30.355 ;
    RECT 173.945 29.925 174.015 29.995 ;
    RECT 130.97 29.565 131.18 29.635 ;
    RECT 130.97 29.925 131.18 29.995 ;
    RECT 130.97 30.285 131.18 30.355 ;
    RECT 131.43 29.565 131.64 29.635 ;
    RECT 131.43 29.925 131.64 29.995 ;
    RECT 131.43 30.285 131.64 30.355 ;
    RECT 127.65 29.565 127.86 29.635 ;
    RECT 127.65 29.925 127.86 29.995 ;
    RECT 127.65 30.285 127.86 30.355 ;
    RECT 128.11 29.565 128.32 29.635 ;
    RECT 128.11 29.925 128.32 29.995 ;
    RECT 128.11 30.285 128.32 30.355 ;
    RECT 124.33 29.565 124.54 29.635 ;
    RECT 124.33 29.925 124.54 29.995 ;
    RECT 124.33 30.285 124.54 30.355 ;
    RECT 124.79 29.565 125.0 29.635 ;
    RECT 124.79 29.925 125.0 29.995 ;
    RECT 124.79 30.285 125.0 30.355 ;
    RECT 121.01 29.565 121.22 29.635 ;
    RECT 121.01 29.925 121.22 29.995 ;
    RECT 121.01 30.285 121.22 30.355 ;
    RECT 121.47 29.565 121.68 29.635 ;
    RECT 121.47 29.925 121.68 29.995 ;
    RECT 121.47 30.285 121.68 30.355 ;
    RECT 117.69 29.565 117.9 29.635 ;
    RECT 117.69 29.925 117.9 29.995 ;
    RECT 117.69 30.285 117.9 30.355 ;
    RECT 118.15 29.565 118.36 29.635 ;
    RECT 118.15 29.925 118.36 29.995 ;
    RECT 118.15 30.285 118.36 30.355 ;
    RECT 114.37 29.565 114.58 29.635 ;
    RECT 114.37 29.925 114.58 29.995 ;
    RECT 114.37 30.285 114.58 30.355 ;
    RECT 114.83 29.565 115.04 29.635 ;
    RECT 114.83 29.925 115.04 29.995 ;
    RECT 114.83 30.285 115.04 30.355 ;
    RECT 111.05 29.565 111.26 29.635 ;
    RECT 111.05 29.925 111.26 29.995 ;
    RECT 111.05 30.285 111.26 30.355 ;
    RECT 111.51 29.565 111.72 29.635 ;
    RECT 111.51 29.925 111.72 29.995 ;
    RECT 111.51 30.285 111.72 30.355 ;
    RECT 107.73 29.565 107.94 29.635 ;
    RECT 107.73 29.925 107.94 29.995 ;
    RECT 107.73 30.285 107.94 30.355 ;
    RECT 108.19 29.565 108.4 29.635 ;
    RECT 108.19 29.925 108.4 29.995 ;
    RECT 108.19 30.285 108.4 30.355 ;
    RECT 104.41 29.565 104.62 29.635 ;
    RECT 104.41 29.925 104.62 29.995 ;
    RECT 104.41 30.285 104.62 30.355 ;
    RECT 104.87 29.565 105.08 29.635 ;
    RECT 104.87 29.925 105.08 29.995 ;
    RECT 104.87 30.285 105.08 30.355 ;
    RECT 101.09 29.565 101.3 29.635 ;
    RECT 101.09 29.925 101.3 29.995 ;
    RECT 101.09 30.285 101.3 30.355 ;
    RECT 101.55 29.565 101.76 29.635 ;
    RECT 101.55 29.925 101.76 29.995 ;
    RECT 101.55 30.285 101.76 30.355 ;
    RECT 0.4 29.925 0.47 29.995 ;
    RECT 170.81 29.565 171.02 29.635 ;
    RECT 170.81 29.925 171.02 29.995 ;
    RECT 170.81 30.285 171.02 30.355 ;
    RECT 171.27 29.565 171.48 29.635 ;
    RECT 171.27 29.925 171.48 29.995 ;
    RECT 171.27 30.285 171.48 30.355 ;
    RECT 167.49 29.565 167.7 29.635 ;
    RECT 167.49 29.925 167.7 29.995 ;
    RECT 167.49 30.285 167.7 30.355 ;
    RECT 167.95 29.565 168.16 29.635 ;
    RECT 167.95 29.925 168.16 29.995 ;
    RECT 167.95 30.285 168.16 30.355 ;
    RECT 97.77 29.565 97.98 29.635 ;
    RECT 97.77 29.925 97.98 29.995 ;
    RECT 97.77 30.285 97.98 30.355 ;
    RECT 98.23 29.565 98.44 29.635 ;
    RECT 98.23 29.925 98.44 29.995 ;
    RECT 98.23 30.285 98.44 30.355 ;
    RECT 94.45 29.565 94.66 29.635 ;
    RECT 94.45 29.925 94.66 29.995 ;
    RECT 94.45 30.285 94.66 30.355 ;
    RECT 94.91 29.565 95.12 29.635 ;
    RECT 94.91 29.925 95.12 29.995 ;
    RECT 94.91 30.285 95.12 30.355 ;
    RECT 91.13 29.565 91.34 29.635 ;
    RECT 91.13 29.925 91.34 29.995 ;
    RECT 91.13 30.285 91.34 30.355 ;
    RECT 91.59 29.565 91.8 29.635 ;
    RECT 91.59 29.925 91.8 29.995 ;
    RECT 91.59 30.285 91.8 30.355 ;
    RECT 87.81 29.565 88.02 29.635 ;
    RECT 87.81 29.925 88.02 29.995 ;
    RECT 87.81 30.285 88.02 30.355 ;
    RECT 88.27 29.565 88.48 29.635 ;
    RECT 88.27 29.925 88.48 29.995 ;
    RECT 88.27 30.285 88.48 30.355 ;
    RECT 84.49 29.565 84.7 29.635 ;
    RECT 84.49 29.925 84.7 29.995 ;
    RECT 84.49 30.285 84.7 30.355 ;
    RECT 84.95 29.565 85.16 29.635 ;
    RECT 84.95 29.925 85.16 29.995 ;
    RECT 84.95 30.285 85.16 30.355 ;
    RECT 81.17 29.565 81.38 29.635 ;
    RECT 81.17 29.925 81.38 29.995 ;
    RECT 81.17 30.285 81.38 30.355 ;
    RECT 81.63 29.565 81.84 29.635 ;
    RECT 81.63 29.925 81.84 29.995 ;
    RECT 81.63 30.285 81.84 30.355 ;
    RECT 77.85 29.565 78.06 29.635 ;
    RECT 77.85 29.925 78.06 29.995 ;
    RECT 77.85 30.285 78.06 30.355 ;
    RECT 78.31 29.565 78.52 29.635 ;
    RECT 78.31 29.925 78.52 29.995 ;
    RECT 78.31 30.285 78.52 30.355 ;
    RECT 74.53 29.565 74.74 29.635 ;
    RECT 74.53 29.925 74.74 29.995 ;
    RECT 74.53 30.285 74.74 30.355 ;
    RECT 74.99 29.565 75.2 29.635 ;
    RECT 74.99 29.925 75.2 29.995 ;
    RECT 74.99 30.285 75.2 30.355 ;
    RECT 71.21 29.565 71.42 29.635 ;
    RECT 71.21 29.925 71.42 29.995 ;
    RECT 71.21 30.285 71.42 30.355 ;
    RECT 71.67 29.565 71.88 29.635 ;
    RECT 71.67 29.925 71.88 29.995 ;
    RECT 71.67 30.285 71.88 30.355 ;
    RECT 31.37 29.565 31.58 29.635 ;
    RECT 31.37 29.925 31.58 29.995 ;
    RECT 31.37 30.285 31.58 30.355 ;
    RECT 31.83 29.565 32.04 29.635 ;
    RECT 31.83 29.925 32.04 29.995 ;
    RECT 31.83 30.285 32.04 30.355 ;
    RECT 67.89 29.565 68.1 29.635 ;
    RECT 67.89 29.925 68.1 29.995 ;
    RECT 67.89 30.285 68.1 30.355 ;
    RECT 68.35 29.565 68.56 29.635 ;
    RECT 68.35 29.925 68.56 29.995 ;
    RECT 68.35 30.285 68.56 30.355 ;
    RECT 28.05 29.565 28.26 29.635 ;
    RECT 28.05 29.925 28.26 29.995 ;
    RECT 28.05 30.285 28.26 30.355 ;
    RECT 28.51 29.565 28.72 29.635 ;
    RECT 28.51 29.925 28.72 29.995 ;
    RECT 28.51 30.285 28.72 30.355 ;
    RECT 24.73 29.565 24.94 29.635 ;
    RECT 24.73 29.925 24.94 29.995 ;
    RECT 24.73 30.285 24.94 30.355 ;
    RECT 25.19 29.565 25.4 29.635 ;
    RECT 25.19 29.925 25.4 29.995 ;
    RECT 25.19 30.285 25.4 30.355 ;
    RECT 21.41 29.565 21.62 29.635 ;
    RECT 21.41 29.925 21.62 29.995 ;
    RECT 21.41 30.285 21.62 30.355 ;
    RECT 21.87 29.565 22.08 29.635 ;
    RECT 21.87 29.925 22.08 29.995 ;
    RECT 21.87 30.285 22.08 30.355 ;
    RECT 18.09 29.565 18.3 29.635 ;
    RECT 18.09 29.925 18.3 29.995 ;
    RECT 18.09 30.285 18.3 30.355 ;
    RECT 18.55 29.565 18.76 29.635 ;
    RECT 18.55 29.925 18.76 29.995 ;
    RECT 18.55 30.285 18.76 30.355 ;
    RECT 14.77 29.565 14.98 29.635 ;
    RECT 14.77 29.925 14.98 29.995 ;
    RECT 14.77 30.285 14.98 30.355 ;
    RECT 15.23 29.565 15.44 29.635 ;
    RECT 15.23 29.925 15.44 29.995 ;
    RECT 15.23 30.285 15.44 30.355 ;
    RECT 11.45 29.565 11.66 29.635 ;
    RECT 11.45 29.925 11.66 29.995 ;
    RECT 11.45 30.285 11.66 30.355 ;
    RECT 11.91 29.565 12.12 29.635 ;
    RECT 11.91 29.925 12.12 29.995 ;
    RECT 11.91 30.285 12.12 30.355 ;
    RECT 8.13 29.565 8.34 29.635 ;
    RECT 8.13 29.925 8.34 29.995 ;
    RECT 8.13 30.285 8.34 30.355 ;
    RECT 8.59 29.565 8.8 29.635 ;
    RECT 8.59 29.925 8.8 29.995 ;
    RECT 8.59 30.285 8.8 30.355 ;
    RECT 4.81 29.565 5.02 29.635 ;
    RECT 4.81 29.925 5.02 29.995 ;
    RECT 4.81 30.285 5.02 30.355 ;
    RECT 5.27 29.565 5.48 29.635 ;
    RECT 5.27 29.925 5.48 29.995 ;
    RECT 5.27 30.285 5.48 30.355 ;
    RECT 164.17 29.565 164.38 29.635 ;
    RECT 164.17 29.925 164.38 29.995 ;
    RECT 164.17 30.285 164.38 30.355 ;
    RECT 164.63 29.565 164.84 29.635 ;
    RECT 164.63 29.925 164.84 29.995 ;
    RECT 164.63 30.285 164.84 30.355 ;
    RECT 1.49 29.565 1.7 29.635 ;
    RECT 1.49 29.925 1.7 29.995 ;
    RECT 1.49 30.285 1.7 30.355 ;
    RECT 1.95 29.565 2.16 29.635 ;
    RECT 1.95 29.925 2.16 29.995 ;
    RECT 1.95 30.285 2.16 30.355 ;
    RECT 160.85 29.565 161.06 29.635 ;
    RECT 160.85 29.925 161.06 29.995 ;
    RECT 160.85 30.285 161.06 30.355 ;
    RECT 161.31 29.565 161.52 29.635 ;
    RECT 161.31 29.925 161.52 29.995 ;
    RECT 161.31 30.285 161.52 30.355 ;
    RECT 157.53 29.565 157.74 29.635 ;
    RECT 157.53 29.925 157.74 29.995 ;
    RECT 157.53 30.285 157.74 30.355 ;
    RECT 157.99 29.565 158.2 29.635 ;
    RECT 157.99 29.925 158.2 29.995 ;
    RECT 157.99 30.285 158.2 30.355 ;
    RECT 154.21 29.565 154.42 29.635 ;
    RECT 154.21 29.925 154.42 29.995 ;
    RECT 154.21 30.285 154.42 30.355 ;
    RECT 154.67 29.565 154.88 29.635 ;
    RECT 154.67 29.925 154.88 29.995 ;
    RECT 154.67 30.285 154.88 30.355 ;
    RECT 150.89 29.565 151.1 29.635 ;
    RECT 150.89 29.925 151.1 29.995 ;
    RECT 150.89 30.285 151.1 30.355 ;
    RECT 151.35 29.565 151.56 29.635 ;
    RECT 151.35 29.925 151.56 29.995 ;
    RECT 151.35 30.285 151.56 30.355 ;
    RECT 147.57 29.565 147.78 29.635 ;
    RECT 147.57 29.925 147.78 29.995 ;
    RECT 147.57 30.285 147.78 30.355 ;
    RECT 148.03 29.565 148.24 29.635 ;
    RECT 148.03 29.925 148.24 29.995 ;
    RECT 148.03 30.285 148.24 30.355 ;
    RECT 144.25 29.565 144.46 29.635 ;
    RECT 144.25 29.925 144.46 29.995 ;
    RECT 144.25 30.285 144.46 30.355 ;
    RECT 144.71 29.565 144.92 29.635 ;
    RECT 144.71 29.925 144.92 29.995 ;
    RECT 144.71 30.285 144.92 30.355 ;
    RECT 140.93 29.565 141.14 29.635 ;
    RECT 140.93 29.925 141.14 29.995 ;
    RECT 140.93 30.285 141.14 30.355 ;
    RECT 141.39 29.565 141.6 29.635 ;
    RECT 141.39 29.925 141.6 29.995 ;
    RECT 141.39 30.285 141.6 30.355 ;
    RECT 137.61 29.565 137.82 29.635 ;
    RECT 137.61 29.925 137.82 29.995 ;
    RECT 137.61 30.285 137.82 30.355 ;
    RECT 138.07 29.565 138.28 29.635 ;
    RECT 138.07 29.925 138.28 29.995 ;
    RECT 138.07 30.285 138.28 30.355 ;
    RECT 134.29 29.565 134.5 29.635 ;
    RECT 134.29 29.925 134.5 29.995 ;
    RECT 134.29 30.285 134.5 30.355 ;
    RECT 134.75 29.565 134.96 29.635 ;
    RECT 134.75 29.925 134.96 29.995 ;
    RECT 134.75 30.285 134.96 30.355 ;
    RECT 64.57 29.565 64.78 29.635 ;
    RECT 64.57 29.925 64.78 29.995 ;
    RECT 64.57 30.285 64.78 30.355 ;
    RECT 65.03 29.565 65.24 29.635 ;
    RECT 65.03 29.925 65.24 29.995 ;
    RECT 65.03 30.285 65.24 30.355 ;
    RECT 61.25 28.845 61.46 28.915 ;
    RECT 61.25 29.205 61.46 29.275 ;
    RECT 61.25 29.565 61.46 29.635 ;
    RECT 61.71 28.845 61.92 28.915 ;
    RECT 61.71 29.205 61.92 29.275 ;
    RECT 61.71 29.565 61.92 29.635 ;
    RECT 57.93 28.845 58.14 28.915 ;
    RECT 57.93 29.205 58.14 29.275 ;
    RECT 57.93 29.565 58.14 29.635 ;
    RECT 58.39 28.845 58.6 28.915 ;
    RECT 58.39 29.205 58.6 29.275 ;
    RECT 58.39 29.565 58.6 29.635 ;
    RECT 54.61 28.845 54.82 28.915 ;
    RECT 54.61 29.205 54.82 29.275 ;
    RECT 54.61 29.565 54.82 29.635 ;
    RECT 55.07 28.845 55.28 28.915 ;
    RECT 55.07 29.205 55.28 29.275 ;
    RECT 55.07 29.565 55.28 29.635 ;
    RECT 51.29 28.845 51.5 28.915 ;
    RECT 51.29 29.205 51.5 29.275 ;
    RECT 51.29 29.565 51.5 29.635 ;
    RECT 51.75 28.845 51.96 28.915 ;
    RECT 51.75 29.205 51.96 29.275 ;
    RECT 51.75 29.565 51.96 29.635 ;
    RECT 47.97 28.845 48.18 28.915 ;
    RECT 47.97 29.205 48.18 29.275 ;
    RECT 47.97 29.565 48.18 29.635 ;
    RECT 48.43 28.845 48.64 28.915 ;
    RECT 48.43 29.205 48.64 29.275 ;
    RECT 48.43 29.565 48.64 29.635 ;
    RECT 44.65 28.845 44.86 28.915 ;
    RECT 44.65 29.205 44.86 29.275 ;
    RECT 44.65 29.565 44.86 29.635 ;
    RECT 45.11 28.845 45.32 28.915 ;
    RECT 45.11 29.205 45.32 29.275 ;
    RECT 45.11 29.565 45.32 29.635 ;
    RECT 41.33 28.845 41.54 28.915 ;
    RECT 41.33 29.205 41.54 29.275 ;
    RECT 41.33 29.565 41.54 29.635 ;
    RECT 41.79 28.845 42.0 28.915 ;
    RECT 41.79 29.205 42.0 29.275 ;
    RECT 41.79 29.565 42.0 29.635 ;
    RECT 38.01 28.845 38.22 28.915 ;
    RECT 38.01 29.205 38.22 29.275 ;
    RECT 38.01 29.565 38.22 29.635 ;
    RECT 38.47 28.845 38.68 28.915 ;
    RECT 38.47 29.205 38.68 29.275 ;
    RECT 38.47 29.565 38.68 29.635 ;
    RECT 34.69 28.845 34.9 28.915 ;
    RECT 34.69 29.205 34.9 29.275 ;
    RECT 34.69 29.565 34.9 29.635 ;
    RECT 35.15 28.845 35.36 28.915 ;
    RECT 35.15 29.205 35.36 29.275 ;
    RECT 35.15 29.565 35.36 29.635 ;
    RECT 173.945 29.205 174.015 29.275 ;
    RECT 130.97 28.845 131.18 28.915 ;
    RECT 130.97 29.205 131.18 29.275 ;
    RECT 130.97 29.565 131.18 29.635 ;
    RECT 131.43 28.845 131.64 28.915 ;
    RECT 131.43 29.205 131.64 29.275 ;
    RECT 131.43 29.565 131.64 29.635 ;
    RECT 127.65 28.845 127.86 28.915 ;
    RECT 127.65 29.205 127.86 29.275 ;
    RECT 127.65 29.565 127.86 29.635 ;
    RECT 128.11 28.845 128.32 28.915 ;
    RECT 128.11 29.205 128.32 29.275 ;
    RECT 128.11 29.565 128.32 29.635 ;
    RECT 124.33 28.845 124.54 28.915 ;
    RECT 124.33 29.205 124.54 29.275 ;
    RECT 124.33 29.565 124.54 29.635 ;
    RECT 124.79 28.845 125.0 28.915 ;
    RECT 124.79 29.205 125.0 29.275 ;
    RECT 124.79 29.565 125.0 29.635 ;
    RECT 121.01 28.845 121.22 28.915 ;
    RECT 121.01 29.205 121.22 29.275 ;
    RECT 121.01 29.565 121.22 29.635 ;
    RECT 121.47 28.845 121.68 28.915 ;
    RECT 121.47 29.205 121.68 29.275 ;
    RECT 121.47 29.565 121.68 29.635 ;
    RECT 117.69 28.845 117.9 28.915 ;
    RECT 117.69 29.205 117.9 29.275 ;
    RECT 117.69 29.565 117.9 29.635 ;
    RECT 118.15 28.845 118.36 28.915 ;
    RECT 118.15 29.205 118.36 29.275 ;
    RECT 118.15 29.565 118.36 29.635 ;
    RECT 114.37 28.845 114.58 28.915 ;
    RECT 114.37 29.205 114.58 29.275 ;
    RECT 114.37 29.565 114.58 29.635 ;
    RECT 114.83 28.845 115.04 28.915 ;
    RECT 114.83 29.205 115.04 29.275 ;
    RECT 114.83 29.565 115.04 29.635 ;
    RECT 111.05 28.845 111.26 28.915 ;
    RECT 111.05 29.205 111.26 29.275 ;
    RECT 111.05 29.565 111.26 29.635 ;
    RECT 111.51 28.845 111.72 28.915 ;
    RECT 111.51 29.205 111.72 29.275 ;
    RECT 111.51 29.565 111.72 29.635 ;
    RECT 107.73 28.845 107.94 28.915 ;
    RECT 107.73 29.205 107.94 29.275 ;
    RECT 107.73 29.565 107.94 29.635 ;
    RECT 108.19 28.845 108.4 28.915 ;
    RECT 108.19 29.205 108.4 29.275 ;
    RECT 108.19 29.565 108.4 29.635 ;
    RECT 104.41 28.845 104.62 28.915 ;
    RECT 104.41 29.205 104.62 29.275 ;
    RECT 104.41 29.565 104.62 29.635 ;
    RECT 104.87 28.845 105.08 28.915 ;
    RECT 104.87 29.205 105.08 29.275 ;
    RECT 104.87 29.565 105.08 29.635 ;
    RECT 101.09 28.845 101.3 28.915 ;
    RECT 101.09 29.205 101.3 29.275 ;
    RECT 101.09 29.565 101.3 29.635 ;
    RECT 101.55 28.845 101.76 28.915 ;
    RECT 101.55 29.205 101.76 29.275 ;
    RECT 101.55 29.565 101.76 29.635 ;
    RECT 0.4 29.205 0.47 29.275 ;
    RECT 170.81 28.845 171.02 28.915 ;
    RECT 170.81 29.205 171.02 29.275 ;
    RECT 170.81 29.565 171.02 29.635 ;
    RECT 171.27 28.845 171.48 28.915 ;
    RECT 171.27 29.205 171.48 29.275 ;
    RECT 171.27 29.565 171.48 29.635 ;
    RECT 167.49 28.845 167.7 28.915 ;
    RECT 167.49 29.205 167.7 29.275 ;
    RECT 167.49 29.565 167.7 29.635 ;
    RECT 167.95 28.845 168.16 28.915 ;
    RECT 167.95 29.205 168.16 29.275 ;
    RECT 167.95 29.565 168.16 29.635 ;
    RECT 97.77 28.845 97.98 28.915 ;
    RECT 97.77 29.205 97.98 29.275 ;
    RECT 97.77 29.565 97.98 29.635 ;
    RECT 98.23 28.845 98.44 28.915 ;
    RECT 98.23 29.205 98.44 29.275 ;
    RECT 98.23 29.565 98.44 29.635 ;
    RECT 94.45 28.845 94.66 28.915 ;
    RECT 94.45 29.205 94.66 29.275 ;
    RECT 94.45 29.565 94.66 29.635 ;
    RECT 94.91 28.845 95.12 28.915 ;
    RECT 94.91 29.205 95.12 29.275 ;
    RECT 94.91 29.565 95.12 29.635 ;
    RECT 91.13 28.845 91.34 28.915 ;
    RECT 91.13 29.205 91.34 29.275 ;
    RECT 91.13 29.565 91.34 29.635 ;
    RECT 91.59 28.845 91.8 28.915 ;
    RECT 91.59 29.205 91.8 29.275 ;
    RECT 91.59 29.565 91.8 29.635 ;
    RECT 87.81 28.845 88.02 28.915 ;
    RECT 87.81 29.205 88.02 29.275 ;
    RECT 87.81 29.565 88.02 29.635 ;
    RECT 88.27 28.845 88.48 28.915 ;
    RECT 88.27 29.205 88.48 29.275 ;
    RECT 88.27 29.565 88.48 29.635 ;
    RECT 84.49 28.845 84.7 28.915 ;
    RECT 84.49 29.205 84.7 29.275 ;
    RECT 84.49 29.565 84.7 29.635 ;
    RECT 84.95 28.845 85.16 28.915 ;
    RECT 84.95 29.205 85.16 29.275 ;
    RECT 84.95 29.565 85.16 29.635 ;
    RECT 81.17 28.845 81.38 28.915 ;
    RECT 81.17 29.205 81.38 29.275 ;
    RECT 81.17 29.565 81.38 29.635 ;
    RECT 81.63 28.845 81.84 28.915 ;
    RECT 81.63 29.205 81.84 29.275 ;
    RECT 81.63 29.565 81.84 29.635 ;
    RECT 77.85 28.845 78.06 28.915 ;
    RECT 77.85 29.205 78.06 29.275 ;
    RECT 77.85 29.565 78.06 29.635 ;
    RECT 78.31 28.845 78.52 28.915 ;
    RECT 78.31 29.205 78.52 29.275 ;
    RECT 78.31 29.565 78.52 29.635 ;
    RECT 74.53 28.845 74.74 28.915 ;
    RECT 74.53 29.205 74.74 29.275 ;
    RECT 74.53 29.565 74.74 29.635 ;
    RECT 74.99 28.845 75.2 28.915 ;
    RECT 74.99 29.205 75.2 29.275 ;
    RECT 74.99 29.565 75.2 29.635 ;
    RECT 71.21 28.845 71.42 28.915 ;
    RECT 71.21 29.205 71.42 29.275 ;
    RECT 71.21 29.565 71.42 29.635 ;
    RECT 71.67 28.845 71.88 28.915 ;
    RECT 71.67 29.205 71.88 29.275 ;
    RECT 71.67 29.565 71.88 29.635 ;
    RECT 31.37 28.845 31.58 28.915 ;
    RECT 31.37 29.205 31.58 29.275 ;
    RECT 31.37 29.565 31.58 29.635 ;
    RECT 31.83 28.845 32.04 28.915 ;
    RECT 31.83 29.205 32.04 29.275 ;
    RECT 31.83 29.565 32.04 29.635 ;
    RECT 67.89 28.845 68.1 28.915 ;
    RECT 67.89 29.205 68.1 29.275 ;
    RECT 67.89 29.565 68.1 29.635 ;
    RECT 68.35 28.845 68.56 28.915 ;
    RECT 68.35 29.205 68.56 29.275 ;
    RECT 68.35 29.565 68.56 29.635 ;
    RECT 28.05 28.845 28.26 28.915 ;
    RECT 28.05 29.205 28.26 29.275 ;
    RECT 28.05 29.565 28.26 29.635 ;
    RECT 28.51 28.845 28.72 28.915 ;
    RECT 28.51 29.205 28.72 29.275 ;
    RECT 28.51 29.565 28.72 29.635 ;
    RECT 24.73 28.845 24.94 28.915 ;
    RECT 24.73 29.205 24.94 29.275 ;
    RECT 24.73 29.565 24.94 29.635 ;
    RECT 25.19 28.845 25.4 28.915 ;
    RECT 25.19 29.205 25.4 29.275 ;
    RECT 25.19 29.565 25.4 29.635 ;
    RECT 21.41 28.845 21.62 28.915 ;
    RECT 21.41 29.205 21.62 29.275 ;
    RECT 21.41 29.565 21.62 29.635 ;
    RECT 21.87 28.845 22.08 28.915 ;
    RECT 21.87 29.205 22.08 29.275 ;
    RECT 21.87 29.565 22.08 29.635 ;
    RECT 18.09 28.845 18.3 28.915 ;
    RECT 18.09 29.205 18.3 29.275 ;
    RECT 18.09 29.565 18.3 29.635 ;
    RECT 18.55 28.845 18.76 28.915 ;
    RECT 18.55 29.205 18.76 29.275 ;
    RECT 18.55 29.565 18.76 29.635 ;
    RECT 14.77 28.845 14.98 28.915 ;
    RECT 14.77 29.205 14.98 29.275 ;
    RECT 14.77 29.565 14.98 29.635 ;
    RECT 15.23 28.845 15.44 28.915 ;
    RECT 15.23 29.205 15.44 29.275 ;
    RECT 15.23 29.565 15.44 29.635 ;
    RECT 11.45 28.845 11.66 28.915 ;
    RECT 11.45 29.205 11.66 29.275 ;
    RECT 11.45 29.565 11.66 29.635 ;
    RECT 11.91 28.845 12.12 28.915 ;
    RECT 11.91 29.205 12.12 29.275 ;
    RECT 11.91 29.565 12.12 29.635 ;
    RECT 8.13 28.845 8.34 28.915 ;
    RECT 8.13 29.205 8.34 29.275 ;
    RECT 8.13 29.565 8.34 29.635 ;
    RECT 8.59 28.845 8.8 28.915 ;
    RECT 8.59 29.205 8.8 29.275 ;
    RECT 8.59 29.565 8.8 29.635 ;
    RECT 4.81 28.845 5.02 28.915 ;
    RECT 4.81 29.205 5.02 29.275 ;
    RECT 4.81 29.565 5.02 29.635 ;
    RECT 5.27 28.845 5.48 28.915 ;
    RECT 5.27 29.205 5.48 29.275 ;
    RECT 5.27 29.565 5.48 29.635 ;
    RECT 164.17 28.845 164.38 28.915 ;
    RECT 164.17 29.205 164.38 29.275 ;
    RECT 164.17 29.565 164.38 29.635 ;
    RECT 164.63 28.845 164.84 28.915 ;
    RECT 164.63 29.205 164.84 29.275 ;
    RECT 164.63 29.565 164.84 29.635 ;
    RECT 1.49 28.845 1.7 28.915 ;
    RECT 1.49 29.205 1.7 29.275 ;
    RECT 1.49 29.565 1.7 29.635 ;
    RECT 1.95 28.845 2.16 28.915 ;
    RECT 1.95 29.205 2.16 29.275 ;
    RECT 1.95 29.565 2.16 29.635 ;
    RECT 160.85 28.845 161.06 28.915 ;
    RECT 160.85 29.205 161.06 29.275 ;
    RECT 160.85 29.565 161.06 29.635 ;
    RECT 161.31 28.845 161.52 28.915 ;
    RECT 161.31 29.205 161.52 29.275 ;
    RECT 161.31 29.565 161.52 29.635 ;
    RECT 157.53 28.845 157.74 28.915 ;
    RECT 157.53 29.205 157.74 29.275 ;
    RECT 157.53 29.565 157.74 29.635 ;
    RECT 157.99 28.845 158.2 28.915 ;
    RECT 157.99 29.205 158.2 29.275 ;
    RECT 157.99 29.565 158.2 29.635 ;
    RECT 154.21 28.845 154.42 28.915 ;
    RECT 154.21 29.205 154.42 29.275 ;
    RECT 154.21 29.565 154.42 29.635 ;
    RECT 154.67 28.845 154.88 28.915 ;
    RECT 154.67 29.205 154.88 29.275 ;
    RECT 154.67 29.565 154.88 29.635 ;
    RECT 150.89 28.845 151.1 28.915 ;
    RECT 150.89 29.205 151.1 29.275 ;
    RECT 150.89 29.565 151.1 29.635 ;
    RECT 151.35 28.845 151.56 28.915 ;
    RECT 151.35 29.205 151.56 29.275 ;
    RECT 151.35 29.565 151.56 29.635 ;
    RECT 147.57 28.845 147.78 28.915 ;
    RECT 147.57 29.205 147.78 29.275 ;
    RECT 147.57 29.565 147.78 29.635 ;
    RECT 148.03 28.845 148.24 28.915 ;
    RECT 148.03 29.205 148.24 29.275 ;
    RECT 148.03 29.565 148.24 29.635 ;
    RECT 144.25 28.845 144.46 28.915 ;
    RECT 144.25 29.205 144.46 29.275 ;
    RECT 144.25 29.565 144.46 29.635 ;
    RECT 144.71 28.845 144.92 28.915 ;
    RECT 144.71 29.205 144.92 29.275 ;
    RECT 144.71 29.565 144.92 29.635 ;
    RECT 140.93 28.845 141.14 28.915 ;
    RECT 140.93 29.205 141.14 29.275 ;
    RECT 140.93 29.565 141.14 29.635 ;
    RECT 141.39 28.845 141.6 28.915 ;
    RECT 141.39 29.205 141.6 29.275 ;
    RECT 141.39 29.565 141.6 29.635 ;
    RECT 137.61 28.845 137.82 28.915 ;
    RECT 137.61 29.205 137.82 29.275 ;
    RECT 137.61 29.565 137.82 29.635 ;
    RECT 138.07 28.845 138.28 28.915 ;
    RECT 138.07 29.205 138.28 29.275 ;
    RECT 138.07 29.565 138.28 29.635 ;
    RECT 134.29 28.845 134.5 28.915 ;
    RECT 134.29 29.205 134.5 29.275 ;
    RECT 134.29 29.565 134.5 29.635 ;
    RECT 134.75 28.845 134.96 28.915 ;
    RECT 134.75 29.205 134.96 29.275 ;
    RECT 134.75 29.565 134.96 29.635 ;
    RECT 64.57 28.845 64.78 28.915 ;
    RECT 64.57 29.205 64.78 29.275 ;
    RECT 64.57 29.565 64.78 29.635 ;
    RECT 65.03 28.845 65.24 28.915 ;
    RECT 65.03 29.205 65.24 29.275 ;
    RECT 65.03 29.565 65.24 29.635 ;
    RECT 61.25 28.125 61.46 28.195 ;
    RECT 61.25 28.485 61.46 28.555 ;
    RECT 61.25 28.845 61.46 28.915 ;
    RECT 61.71 28.125 61.92 28.195 ;
    RECT 61.71 28.485 61.92 28.555 ;
    RECT 61.71 28.845 61.92 28.915 ;
    RECT 57.93 28.125 58.14 28.195 ;
    RECT 57.93 28.485 58.14 28.555 ;
    RECT 57.93 28.845 58.14 28.915 ;
    RECT 58.39 28.125 58.6 28.195 ;
    RECT 58.39 28.485 58.6 28.555 ;
    RECT 58.39 28.845 58.6 28.915 ;
    RECT 54.61 28.125 54.82 28.195 ;
    RECT 54.61 28.485 54.82 28.555 ;
    RECT 54.61 28.845 54.82 28.915 ;
    RECT 55.07 28.125 55.28 28.195 ;
    RECT 55.07 28.485 55.28 28.555 ;
    RECT 55.07 28.845 55.28 28.915 ;
    RECT 51.29 28.125 51.5 28.195 ;
    RECT 51.29 28.485 51.5 28.555 ;
    RECT 51.29 28.845 51.5 28.915 ;
    RECT 51.75 28.125 51.96 28.195 ;
    RECT 51.75 28.485 51.96 28.555 ;
    RECT 51.75 28.845 51.96 28.915 ;
    RECT 47.97 28.125 48.18 28.195 ;
    RECT 47.97 28.485 48.18 28.555 ;
    RECT 47.97 28.845 48.18 28.915 ;
    RECT 48.43 28.125 48.64 28.195 ;
    RECT 48.43 28.485 48.64 28.555 ;
    RECT 48.43 28.845 48.64 28.915 ;
    RECT 44.65 28.125 44.86 28.195 ;
    RECT 44.65 28.485 44.86 28.555 ;
    RECT 44.65 28.845 44.86 28.915 ;
    RECT 45.11 28.125 45.32 28.195 ;
    RECT 45.11 28.485 45.32 28.555 ;
    RECT 45.11 28.845 45.32 28.915 ;
    RECT 41.33 28.125 41.54 28.195 ;
    RECT 41.33 28.485 41.54 28.555 ;
    RECT 41.33 28.845 41.54 28.915 ;
    RECT 41.79 28.125 42.0 28.195 ;
    RECT 41.79 28.485 42.0 28.555 ;
    RECT 41.79 28.845 42.0 28.915 ;
    RECT 38.01 28.125 38.22 28.195 ;
    RECT 38.01 28.485 38.22 28.555 ;
    RECT 38.01 28.845 38.22 28.915 ;
    RECT 38.47 28.125 38.68 28.195 ;
    RECT 38.47 28.485 38.68 28.555 ;
    RECT 38.47 28.845 38.68 28.915 ;
    RECT 34.69 28.125 34.9 28.195 ;
    RECT 34.69 28.485 34.9 28.555 ;
    RECT 34.69 28.845 34.9 28.915 ;
    RECT 35.15 28.125 35.36 28.195 ;
    RECT 35.15 28.485 35.36 28.555 ;
    RECT 35.15 28.845 35.36 28.915 ;
    RECT 173.945 28.485 174.015 28.555 ;
    RECT 130.97 28.125 131.18 28.195 ;
    RECT 130.97 28.485 131.18 28.555 ;
    RECT 130.97 28.845 131.18 28.915 ;
    RECT 131.43 28.125 131.64 28.195 ;
    RECT 131.43 28.485 131.64 28.555 ;
    RECT 131.43 28.845 131.64 28.915 ;
    RECT 127.65 28.125 127.86 28.195 ;
    RECT 127.65 28.485 127.86 28.555 ;
    RECT 127.65 28.845 127.86 28.915 ;
    RECT 128.11 28.125 128.32 28.195 ;
    RECT 128.11 28.485 128.32 28.555 ;
    RECT 128.11 28.845 128.32 28.915 ;
    RECT 124.33 28.125 124.54 28.195 ;
    RECT 124.33 28.485 124.54 28.555 ;
    RECT 124.33 28.845 124.54 28.915 ;
    RECT 124.79 28.125 125.0 28.195 ;
    RECT 124.79 28.485 125.0 28.555 ;
    RECT 124.79 28.845 125.0 28.915 ;
    RECT 121.01 28.125 121.22 28.195 ;
    RECT 121.01 28.485 121.22 28.555 ;
    RECT 121.01 28.845 121.22 28.915 ;
    RECT 121.47 28.125 121.68 28.195 ;
    RECT 121.47 28.485 121.68 28.555 ;
    RECT 121.47 28.845 121.68 28.915 ;
    RECT 117.69 28.125 117.9 28.195 ;
    RECT 117.69 28.485 117.9 28.555 ;
    RECT 117.69 28.845 117.9 28.915 ;
    RECT 118.15 28.125 118.36 28.195 ;
    RECT 118.15 28.485 118.36 28.555 ;
    RECT 118.15 28.845 118.36 28.915 ;
    RECT 114.37 28.125 114.58 28.195 ;
    RECT 114.37 28.485 114.58 28.555 ;
    RECT 114.37 28.845 114.58 28.915 ;
    RECT 114.83 28.125 115.04 28.195 ;
    RECT 114.83 28.485 115.04 28.555 ;
    RECT 114.83 28.845 115.04 28.915 ;
    RECT 111.05 28.125 111.26 28.195 ;
    RECT 111.05 28.485 111.26 28.555 ;
    RECT 111.05 28.845 111.26 28.915 ;
    RECT 111.51 28.125 111.72 28.195 ;
    RECT 111.51 28.485 111.72 28.555 ;
    RECT 111.51 28.845 111.72 28.915 ;
    RECT 107.73 28.125 107.94 28.195 ;
    RECT 107.73 28.485 107.94 28.555 ;
    RECT 107.73 28.845 107.94 28.915 ;
    RECT 108.19 28.125 108.4 28.195 ;
    RECT 108.19 28.485 108.4 28.555 ;
    RECT 108.19 28.845 108.4 28.915 ;
    RECT 104.41 28.125 104.62 28.195 ;
    RECT 104.41 28.485 104.62 28.555 ;
    RECT 104.41 28.845 104.62 28.915 ;
    RECT 104.87 28.125 105.08 28.195 ;
    RECT 104.87 28.485 105.08 28.555 ;
    RECT 104.87 28.845 105.08 28.915 ;
    RECT 101.09 28.125 101.3 28.195 ;
    RECT 101.09 28.485 101.3 28.555 ;
    RECT 101.09 28.845 101.3 28.915 ;
    RECT 101.55 28.125 101.76 28.195 ;
    RECT 101.55 28.485 101.76 28.555 ;
    RECT 101.55 28.845 101.76 28.915 ;
    RECT 0.4 28.485 0.47 28.555 ;
    RECT 170.81 28.125 171.02 28.195 ;
    RECT 170.81 28.485 171.02 28.555 ;
    RECT 170.81 28.845 171.02 28.915 ;
    RECT 171.27 28.125 171.48 28.195 ;
    RECT 171.27 28.485 171.48 28.555 ;
    RECT 171.27 28.845 171.48 28.915 ;
    RECT 167.49 28.125 167.7 28.195 ;
    RECT 167.49 28.485 167.7 28.555 ;
    RECT 167.49 28.845 167.7 28.915 ;
    RECT 167.95 28.125 168.16 28.195 ;
    RECT 167.95 28.485 168.16 28.555 ;
    RECT 167.95 28.845 168.16 28.915 ;
    RECT 97.77 28.125 97.98 28.195 ;
    RECT 97.77 28.485 97.98 28.555 ;
    RECT 97.77 28.845 97.98 28.915 ;
    RECT 98.23 28.125 98.44 28.195 ;
    RECT 98.23 28.485 98.44 28.555 ;
    RECT 98.23 28.845 98.44 28.915 ;
    RECT 94.45 28.125 94.66 28.195 ;
    RECT 94.45 28.485 94.66 28.555 ;
    RECT 94.45 28.845 94.66 28.915 ;
    RECT 94.91 28.125 95.12 28.195 ;
    RECT 94.91 28.485 95.12 28.555 ;
    RECT 94.91 28.845 95.12 28.915 ;
    RECT 91.13 28.125 91.34 28.195 ;
    RECT 91.13 28.485 91.34 28.555 ;
    RECT 91.13 28.845 91.34 28.915 ;
    RECT 91.59 28.125 91.8 28.195 ;
    RECT 91.59 28.485 91.8 28.555 ;
    RECT 91.59 28.845 91.8 28.915 ;
    RECT 87.81 28.125 88.02 28.195 ;
    RECT 87.81 28.485 88.02 28.555 ;
    RECT 87.81 28.845 88.02 28.915 ;
    RECT 88.27 28.125 88.48 28.195 ;
    RECT 88.27 28.485 88.48 28.555 ;
    RECT 88.27 28.845 88.48 28.915 ;
    RECT 84.49 28.125 84.7 28.195 ;
    RECT 84.49 28.485 84.7 28.555 ;
    RECT 84.49 28.845 84.7 28.915 ;
    RECT 84.95 28.125 85.16 28.195 ;
    RECT 84.95 28.485 85.16 28.555 ;
    RECT 84.95 28.845 85.16 28.915 ;
    RECT 81.17 28.125 81.38 28.195 ;
    RECT 81.17 28.485 81.38 28.555 ;
    RECT 81.17 28.845 81.38 28.915 ;
    RECT 81.63 28.125 81.84 28.195 ;
    RECT 81.63 28.485 81.84 28.555 ;
    RECT 81.63 28.845 81.84 28.915 ;
    RECT 77.85 28.125 78.06 28.195 ;
    RECT 77.85 28.485 78.06 28.555 ;
    RECT 77.85 28.845 78.06 28.915 ;
    RECT 78.31 28.125 78.52 28.195 ;
    RECT 78.31 28.485 78.52 28.555 ;
    RECT 78.31 28.845 78.52 28.915 ;
    RECT 74.53 28.125 74.74 28.195 ;
    RECT 74.53 28.485 74.74 28.555 ;
    RECT 74.53 28.845 74.74 28.915 ;
    RECT 74.99 28.125 75.2 28.195 ;
    RECT 74.99 28.485 75.2 28.555 ;
    RECT 74.99 28.845 75.2 28.915 ;
    RECT 71.21 28.125 71.42 28.195 ;
    RECT 71.21 28.485 71.42 28.555 ;
    RECT 71.21 28.845 71.42 28.915 ;
    RECT 71.67 28.125 71.88 28.195 ;
    RECT 71.67 28.485 71.88 28.555 ;
    RECT 71.67 28.845 71.88 28.915 ;
    RECT 31.37 28.125 31.58 28.195 ;
    RECT 31.37 28.485 31.58 28.555 ;
    RECT 31.37 28.845 31.58 28.915 ;
    RECT 31.83 28.125 32.04 28.195 ;
    RECT 31.83 28.485 32.04 28.555 ;
    RECT 31.83 28.845 32.04 28.915 ;
    RECT 67.89 28.125 68.1 28.195 ;
    RECT 67.89 28.485 68.1 28.555 ;
    RECT 67.89 28.845 68.1 28.915 ;
    RECT 68.35 28.125 68.56 28.195 ;
    RECT 68.35 28.485 68.56 28.555 ;
    RECT 68.35 28.845 68.56 28.915 ;
    RECT 28.05 28.125 28.26 28.195 ;
    RECT 28.05 28.485 28.26 28.555 ;
    RECT 28.05 28.845 28.26 28.915 ;
    RECT 28.51 28.125 28.72 28.195 ;
    RECT 28.51 28.485 28.72 28.555 ;
    RECT 28.51 28.845 28.72 28.915 ;
    RECT 24.73 28.125 24.94 28.195 ;
    RECT 24.73 28.485 24.94 28.555 ;
    RECT 24.73 28.845 24.94 28.915 ;
    RECT 25.19 28.125 25.4 28.195 ;
    RECT 25.19 28.485 25.4 28.555 ;
    RECT 25.19 28.845 25.4 28.915 ;
    RECT 21.41 28.125 21.62 28.195 ;
    RECT 21.41 28.485 21.62 28.555 ;
    RECT 21.41 28.845 21.62 28.915 ;
    RECT 21.87 28.125 22.08 28.195 ;
    RECT 21.87 28.485 22.08 28.555 ;
    RECT 21.87 28.845 22.08 28.915 ;
    RECT 18.09 28.125 18.3 28.195 ;
    RECT 18.09 28.485 18.3 28.555 ;
    RECT 18.09 28.845 18.3 28.915 ;
    RECT 18.55 28.125 18.76 28.195 ;
    RECT 18.55 28.485 18.76 28.555 ;
    RECT 18.55 28.845 18.76 28.915 ;
    RECT 14.77 28.125 14.98 28.195 ;
    RECT 14.77 28.485 14.98 28.555 ;
    RECT 14.77 28.845 14.98 28.915 ;
    RECT 15.23 28.125 15.44 28.195 ;
    RECT 15.23 28.485 15.44 28.555 ;
    RECT 15.23 28.845 15.44 28.915 ;
    RECT 11.45 28.125 11.66 28.195 ;
    RECT 11.45 28.485 11.66 28.555 ;
    RECT 11.45 28.845 11.66 28.915 ;
    RECT 11.91 28.125 12.12 28.195 ;
    RECT 11.91 28.485 12.12 28.555 ;
    RECT 11.91 28.845 12.12 28.915 ;
    RECT 8.13 28.125 8.34 28.195 ;
    RECT 8.13 28.485 8.34 28.555 ;
    RECT 8.13 28.845 8.34 28.915 ;
    RECT 8.59 28.125 8.8 28.195 ;
    RECT 8.59 28.485 8.8 28.555 ;
    RECT 8.59 28.845 8.8 28.915 ;
    RECT 4.81 28.125 5.02 28.195 ;
    RECT 4.81 28.485 5.02 28.555 ;
    RECT 4.81 28.845 5.02 28.915 ;
    RECT 5.27 28.125 5.48 28.195 ;
    RECT 5.27 28.485 5.48 28.555 ;
    RECT 5.27 28.845 5.48 28.915 ;
    RECT 164.17 28.125 164.38 28.195 ;
    RECT 164.17 28.485 164.38 28.555 ;
    RECT 164.17 28.845 164.38 28.915 ;
    RECT 164.63 28.125 164.84 28.195 ;
    RECT 164.63 28.485 164.84 28.555 ;
    RECT 164.63 28.845 164.84 28.915 ;
    RECT 1.49 28.125 1.7 28.195 ;
    RECT 1.49 28.485 1.7 28.555 ;
    RECT 1.49 28.845 1.7 28.915 ;
    RECT 1.95 28.125 2.16 28.195 ;
    RECT 1.95 28.485 2.16 28.555 ;
    RECT 1.95 28.845 2.16 28.915 ;
    RECT 160.85 28.125 161.06 28.195 ;
    RECT 160.85 28.485 161.06 28.555 ;
    RECT 160.85 28.845 161.06 28.915 ;
    RECT 161.31 28.125 161.52 28.195 ;
    RECT 161.31 28.485 161.52 28.555 ;
    RECT 161.31 28.845 161.52 28.915 ;
    RECT 157.53 28.125 157.74 28.195 ;
    RECT 157.53 28.485 157.74 28.555 ;
    RECT 157.53 28.845 157.74 28.915 ;
    RECT 157.99 28.125 158.2 28.195 ;
    RECT 157.99 28.485 158.2 28.555 ;
    RECT 157.99 28.845 158.2 28.915 ;
    RECT 154.21 28.125 154.42 28.195 ;
    RECT 154.21 28.485 154.42 28.555 ;
    RECT 154.21 28.845 154.42 28.915 ;
    RECT 154.67 28.125 154.88 28.195 ;
    RECT 154.67 28.485 154.88 28.555 ;
    RECT 154.67 28.845 154.88 28.915 ;
    RECT 150.89 28.125 151.1 28.195 ;
    RECT 150.89 28.485 151.1 28.555 ;
    RECT 150.89 28.845 151.1 28.915 ;
    RECT 151.35 28.125 151.56 28.195 ;
    RECT 151.35 28.485 151.56 28.555 ;
    RECT 151.35 28.845 151.56 28.915 ;
    RECT 147.57 28.125 147.78 28.195 ;
    RECT 147.57 28.485 147.78 28.555 ;
    RECT 147.57 28.845 147.78 28.915 ;
    RECT 148.03 28.125 148.24 28.195 ;
    RECT 148.03 28.485 148.24 28.555 ;
    RECT 148.03 28.845 148.24 28.915 ;
    RECT 144.25 28.125 144.46 28.195 ;
    RECT 144.25 28.485 144.46 28.555 ;
    RECT 144.25 28.845 144.46 28.915 ;
    RECT 144.71 28.125 144.92 28.195 ;
    RECT 144.71 28.485 144.92 28.555 ;
    RECT 144.71 28.845 144.92 28.915 ;
    RECT 140.93 28.125 141.14 28.195 ;
    RECT 140.93 28.485 141.14 28.555 ;
    RECT 140.93 28.845 141.14 28.915 ;
    RECT 141.39 28.125 141.6 28.195 ;
    RECT 141.39 28.485 141.6 28.555 ;
    RECT 141.39 28.845 141.6 28.915 ;
    RECT 137.61 28.125 137.82 28.195 ;
    RECT 137.61 28.485 137.82 28.555 ;
    RECT 137.61 28.845 137.82 28.915 ;
    RECT 138.07 28.125 138.28 28.195 ;
    RECT 138.07 28.485 138.28 28.555 ;
    RECT 138.07 28.845 138.28 28.915 ;
    RECT 134.29 28.125 134.5 28.195 ;
    RECT 134.29 28.485 134.5 28.555 ;
    RECT 134.29 28.845 134.5 28.915 ;
    RECT 134.75 28.125 134.96 28.195 ;
    RECT 134.75 28.485 134.96 28.555 ;
    RECT 134.75 28.845 134.96 28.915 ;
    RECT 64.57 28.125 64.78 28.195 ;
    RECT 64.57 28.485 64.78 28.555 ;
    RECT 64.57 28.845 64.78 28.915 ;
    RECT 65.03 28.125 65.24 28.195 ;
    RECT 65.03 28.485 65.24 28.555 ;
    RECT 65.03 28.845 65.24 28.915 ;
    RECT 61.25 27.405 61.46 27.475 ;
    RECT 61.25 27.765 61.46 27.835 ;
    RECT 61.25 28.125 61.46 28.195 ;
    RECT 61.71 27.405 61.92 27.475 ;
    RECT 61.71 27.765 61.92 27.835 ;
    RECT 61.71 28.125 61.92 28.195 ;
    RECT 57.93 27.405 58.14 27.475 ;
    RECT 57.93 27.765 58.14 27.835 ;
    RECT 57.93 28.125 58.14 28.195 ;
    RECT 58.39 27.405 58.6 27.475 ;
    RECT 58.39 27.765 58.6 27.835 ;
    RECT 58.39 28.125 58.6 28.195 ;
    RECT 54.61 27.405 54.82 27.475 ;
    RECT 54.61 27.765 54.82 27.835 ;
    RECT 54.61 28.125 54.82 28.195 ;
    RECT 55.07 27.405 55.28 27.475 ;
    RECT 55.07 27.765 55.28 27.835 ;
    RECT 55.07 28.125 55.28 28.195 ;
    RECT 51.29 27.405 51.5 27.475 ;
    RECT 51.29 27.765 51.5 27.835 ;
    RECT 51.29 28.125 51.5 28.195 ;
    RECT 51.75 27.405 51.96 27.475 ;
    RECT 51.75 27.765 51.96 27.835 ;
    RECT 51.75 28.125 51.96 28.195 ;
    RECT 47.97 27.405 48.18 27.475 ;
    RECT 47.97 27.765 48.18 27.835 ;
    RECT 47.97 28.125 48.18 28.195 ;
    RECT 48.43 27.405 48.64 27.475 ;
    RECT 48.43 27.765 48.64 27.835 ;
    RECT 48.43 28.125 48.64 28.195 ;
    RECT 44.65 27.405 44.86 27.475 ;
    RECT 44.65 27.765 44.86 27.835 ;
    RECT 44.65 28.125 44.86 28.195 ;
    RECT 45.11 27.405 45.32 27.475 ;
    RECT 45.11 27.765 45.32 27.835 ;
    RECT 45.11 28.125 45.32 28.195 ;
    RECT 41.33 27.405 41.54 27.475 ;
    RECT 41.33 27.765 41.54 27.835 ;
    RECT 41.33 28.125 41.54 28.195 ;
    RECT 41.79 27.405 42.0 27.475 ;
    RECT 41.79 27.765 42.0 27.835 ;
    RECT 41.79 28.125 42.0 28.195 ;
    RECT 38.01 27.405 38.22 27.475 ;
    RECT 38.01 27.765 38.22 27.835 ;
    RECT 38.01 28.125 38.22 28.195 ;
    RECT 38.47 27.405 38.68 27.475 ;
    RECT 38.47 27.765 38.68 27.835 ;
    RECT 38.47 28.125 38.68 28.195 ;
    RECT 34.69 27.405 34.9 27.475 ;
    RECT 34.69 27.765 34.9 27.835 ;
    RECT 34.69 28.125 34.9 28.195 ;
    RECT 35.15 27.405 35.36 27.475 ;
    RECT 35.15 27.765 35.36 27.835 ;
    RECT 35.15 28.125 35.36 28.195 ;
    RECT 173.945 27.765 174.015 27.835 ;
    RECT 130.97 27.405 131.18 27.475 ;
    RECT 130.97 27.765 131.18 27.835 ;
    RECT 130.97 28.125 131.18 28.195 ;
    RECT 131.43 27.405 131.64 27.475 ;
    RECT 131.43 27.765 131.64 27.835 ;
    RECT 131.43 28.125 131.64 28.195 ;
    RECT 127.65 27.405 127.86 27.475 ;
    RECT 127.65 27.765 127.86 27.835 ;
    RECT 127.65 28.125 127.86 28.195 ;
    RECT 128.11 27.405 128.32 27.475 ;
    RECT 128.11 27.765 128.32 27.835 ;
    RECT 128.11 28.125 128.32 28.195 ;
    RECT 124.33 27.405 124.54 27.475 ;
    RECT 124.33 27.765 124.54 27.835 ;
    RECT 124.33 28.125 124.54 28.195 ;
    RECT 124.79 27.405 125.0 27.475 ;
    RECT 124.79 27.765 125.0 27.835 ;
    RECT 124.79 28.125 125.0 28.195 ;
    RECT 121.01 27.405 121.22 27.475 ;
    RECT 121.01 27.765 121.22 27.835 ;
    RECT 121.01 28.125 121.22 28.195 ;
    RECT 121.47 27.405 121.68 27.475 ;
    RECT 121.47 27.765 121.68 27.835 ;
    RECT 121.47 28.125 121.68 28.195 ;
    RECT 117.69 27.405 117.9 27.475 ;
    RECT 117.69 27.765 117.9 27.835 ;
    RECT 117.69 28.125 117.9 28.195 ;
    RECT 118.15 27.405 118.36 27.475 ;
    RECT 118.15 27.765 118.36 27.835 ;
    RECT 118.15 28.125 118.36 28.195 ;
    RECT 114.37 27.405 114.58 27.475 ;
    RECT 114.37 27.765 114.58 27.835 ;
    RECT 114.37 28.125 114.58 28.195 ;
    RECT 114.83 27.405 115.04 27.475 ;
    RECT 114.83 27.765 115.04 27.835 ;
    RECT 114.83 28.125 115.04 28.195 ;
    RECT 111.05 27.405 111.26 27.475 ;
    RECT 111.05 27.765 111.26 27.835 ;
    RECT 111.05 28.125 111.26 28.195 ;
    RECT 111.51 27.405 111.72 27.475 ;
    RECT 111.51 27.765 111.72 27.835 ;
    RECT 111.51 28.125 111.72 28.195 ;
    RECT 107.73 27.405 107.94 27.475 ;
    RECT 107.73 27.765 107.94 27.835 ;
    RECT 107.73 28.125 107.94 28.195 ;
    RECT 108.19 27.405 108.4 27.475 ;
    RECT 108.19 27.765 108.4 27.835 ;
    RECT 108.19 28.125 108.4 28.195 ;
    RECT 104.41 27.405 104.62 27.475 ;
    RECT 104.41 27.765 104.62 27.835 ;
    RECT 104.41 28.125 104.62 28.195 ;
    RECT 104.87 27.405 105.08 27.475 ;
    RECT 104.87 27.765 105.08 27.835 ;
    RECT 104.87 28.125 105.08 28.195 ;
    RECT 101.09 27.405 101.3 27.475 ;
    RECT 101.09 27.765 101.3 27.835 ;
    RECT 101.09 28.125 101.3 28.195 ;
    RECT 101.55 27.405 101.76 27.475 ;
    RECT 101.55 27.765 101.76 27.835 ;
    RECT 101.55 28.125 101.76 28.195 ;
    RECT 0.4 27.765 0.47 27.835 ;
    RECT 170.81 27.405 171.02 27.475 ;
    RECT 170.81 27.765 171.02 27.835 ;
    RECT 170.81 28.125 171.02 28.195 ;
    RECT 171.27 27.405 171.48 27.475 ;
    RECT 171.27 27.765 171.48 27.835 ;
    RECT 171.27 28.125 171.48 28.195 ;
    RECT 167.49 27.405 167.7 27.475 ;
    RECT 167.49 27.765 167.7 27.835 ;
    RECT 167.49 28.125 167.7 28.195 ;
    RECT 167.95 27.405 168.16 27.475 ;
    RECT 167.95 27.765 168.16 27.835 ;
    RECT 167.95 28.125 168.16 28.195 ;
    RECT 97.77 27.405 97.98 27.475 ;
    RECT 97.77 27.765 97.98 27.835 ;
    RECT 97.77 28.125 97.98 28.195 ;
    RECT 98.23 27.405 98.44 27.475 ;
    RECT 98.23 27.765 98.44 27.835 ;
    RECT 98.23 28.125 98.44 28.195 ;
    RECT 94.45 27.405 94.66 27.475 ;
    RECT 94.45 27.765 94.66 27.835 ;
    RECT 94.45 28.125 94.66 28.195 ;
    RECT 94.91 27.405 95.12 27.475 ;
    RECT 94.91 27.765 95.12 27.835 ;
    RECT 94.91 28.125 95.12 28.195 ;
    RECT 91.13 27.405 91.34 27.475 ;
    RECT 91.13 27.765 91.34 27.835 ;
    RECT 91.13 28.125 91.34 28.195 ;
    RECT 91.59 27.405 91.8 27.475 ;
    RECT 91.59 27.765 91.8 27.835 ;
    RECT 91.59 28.125 91.8 28.195 ;
    RECT 87.81 27.405 88.02 27.475 ;
    RECT 87.81 27.765 88.02 27.835 ;
    RECT 87.81 28.125 88.02 28.195 ;
    RECT 88.27 27.405 88.48 27.475 ;
    RECT 88.27 27.765 88.48 27.835 ;
    RECT 88.27 28.125 88.48 28.195 ;
    RECT 84.49 27.405 84.7 27.475 ;
    RECT 84.49 27.765 84.7 27.835 ;
    RECT 84.49 28.125 84.7 28.195 ;
    RECT 84.95 27.405 85.16 27.475 ;
    RECT 84.95 27.765 85.16 27.835 ;
    RECT 84.95 28.125 85.16 28.195 ;
    RECT 81.17 27.405 81.38 27.475 ;
    RECT 81.17 27.765 81.38 27.835 ;
    RECT 81.17 28.125 81.38 28.195 ;
    RECT 81.63 27.405 81.84 27.475 ;
    RECT 81.63 27.765 81.84 27.835 ;
    RECT 81.63 28.125 81.84 28.195 ;
    RECT 77.85 27.405 78.06 27.475 ;
    RECT 77.85 27.765 78.06 27.835 ;
    RECT 77.85 28.125 78.06 28.195 ;
    RECT 78.31 27.405 78.52 27.475 ;
    RECT 78.31 27.765 78.52 27.835 ;
    RECT 78.31 28.125 78.52 28.195 ;
    RECT 74.53 27.405 74.74 27.475 ;
    RECT 74.53 27.765 74.74 27.835 ;
    RECT 74.53 28.125 74.74 28.195 ;
    RECT 74.99 27.405 75.2 27.475 ;
    RECT 74.99 27.765 75.2 27.835 ;
    RECT 74.99 28.125 75.2 28.195 ;
    RECT 71.21 27.405 71.42 27.475 ;
    RECT 71.21 27.765 71.42 27.835 ;
    RECT 71.21 28.125 71.42 28.195 ;
    RECT 71.67 27.405 71.88 27.475 ;
    RECT 71.67 27.765 71.88 27.835 ;
    RECT 71.67 28.125 71.88 28.195 ;
    RECT 31.37 27.405 31.58 27.475 ;
    RECT 31.37 27.765 31.58 27.835 ;
    RECT 31.37 28.125 31.58 28.195 ;
    RECT 31.83 27.405 32.04 27.475 ;
    RECT 31.83 27.765 32.04 27.835 ;
    RECT 31.83 28.125 32.04 28.195 ;
    RECT 67.89 27.405 68.1 27.475 ;
    RECT 67.89 27.765 68.1 27.835 ;
    RECT 67.89 28.125 68.1 28.195 ;
    RECT 68.35 27.405 68.56 27.475 ;
    RECT 68.35 27.765 68.56 27.835 ;
    RECT 68.35 28.125 68.56 28.195 ;
    RECT 28.05 27.405 28.26 27.475 ;
    RECT 28.05 27.765 28.26 27.835 ;
    RECT 28.05 28.125 28.26 28.195 ;
    RECT 28.51 27.405 28.72 27.475 ;
    RECT 28.51 27.765 28.72 27.835 ;
    RECT 28.51 28.125 28.72 28.195 ;
    RECT 24.73 27.405 24.94 27.475 ;
    RECT 24.73 27.765 24.94 27.835 ;
    RECT 24.73 28.125 24.94 28.195 ;
    RECT 25.19 27.405 25.4 27.475 ;
    RECT 25.19 27.765 25.4 27.835 ;
    RECT 25.19 28.125 25.4 28.195 ;
    RECT 21.41 27.405 21.62 27.475 ;
    RECT 21.41 27.765 21.62 27.835 ;
    RECT 21.41 28.125 21.62 28.195 ;
    RECT 21.87 27.405 22.08 27.475 ;
    RECT 21.87 27.765 22.08 27.835 ;
    RECT 21.87 28.125 22.08 28.195 ;
    RECT 18.09 27.405 18.3 27.475 ;
    RECT 18.09 27.765 18.3 27.835 ;
    RECT 18.09 28.125 18.3 28.195 ;
    RECT 18.55 27.405 18.76 27.475 ;
    RECT 18.55 27.765 18.76 27.835 ;
    RECT 18.55 28.125 18.76 28.195 ;
    RECT 14.77 27.405 14.98 27.475 ;
    RECT 14.77 27.765 14.98 27.835 ;
    RECT 14.77 28.125 14.98 28.195 ;
    RECT 15.23 27.405 15.44 27.475 ;
    RECT 15.23 27.765 15.44 27.835 ;
    RECT 15.23 28.125 15.44 28.195 ;
    RECT 11.45 27.405 11.66 27.475 ;
    RECT 11.45 27.765 11.66 27.835 ;
    RECT 11.45 28.125 11.66 28.195 ;
    RECT 11.91 27.405 12.12 27.475 ;
    RECT 11.91 27.765 12.12 27.835 ;
    RECT 11.91 28.125 12.12 28.195 ;
    RECT 8.13 27.405 8.34 27.475 ;
    RECT 8.13 27.765 8.34 27.835 ;
    RECT 8.13 28.125 8.34 28.195 ;
    RECT 8.59 27.405 8.8 27.475 ;
    RECT 8.59 27.765 8.8 27.835 ;
    RECT 8.59 28.125 8.8 28.195 ;
    RECT 4.81 27.405 5.02 27.475 ;
    RECT 4.81 27.765 5.02 27.835 ;
    RECT 4.81 28.125 5.02 28.195 ;
    RECT 5.27 27.405 5.48 27.475 ;
    RECT 5.27 27.765 5.48 27.835 ;
    RECT 5.27 28.125 5.48 28.195 ;
    RECT 164.17 27.405 164.38 27.475 ;
    RECT 164.17 27.765 164.38 27.835 ;
    RECT 164.17 28.125 164.38 28.195 ;
    RECT 164.63 27.405 164.84 27.475 ;
    RECT 164.63 27.765 164.84 27.835 ;
    RECT 164.63 28.125 164.84 28.195 ;
    RECT 1.49 27.405 1.7 27.475 ;
    RECT 1.49 27.765 1.7 27.835 ;
    RECT 1.49 28.125 1.7 28.195 ;
    RECT 1.95 27.405 2.16 27.475 ;
    RECT 1.95 27.765 2.16 27.835 ;
    RECT 1.95 28.125 2.16 28.195 ;
    RECT 160.85 27.405 161.06 27.475 ;
    RECT 160.85 27.765 161.06 27.835 ;
    RECT 160.85 28.125 161.06 28.195 ;
    RECT 161.31 27.405 161.52 27.475 ;
    RECT 161.31 27.765 161.52 27.835 ;
    RECT 161.31 28.125 161.52 28.195 ;
    RECT 157.53 27.405 157.74 27.475 ;
    RECT 157.53 27.765 157.74 27.835 ;
    RECT 157.53 28.125 157.74 28.195 ;
    RECT 157.99 27.405 158.2 27.475 ;
    RECT 157.99 27.765 158.2 27.835 ;
    RECT 157.99 28.125 158.2 28.195 ;
    RECT 154.21 27.405 154.42 27.475 ;
    RECT 154.21 27.765 154.42 27.835 ;
    RECT 154.21 28.125 154.42 28.195 ;
    RECT 154.67 27.405 154.88 27.475 ;
    RECT 154.67 27.765 154.88 27.835 ;
    RECT 154.67 28.125 154.88 28.195 ;
    RECT 150.89 27.405 151.1 27.475 ;
    RECT 150.89 27.765 151.1 27.835 ;
    RECT 150.89 28.125 151.1 28.195 ;
    RECT 151.35 27.405 151.56 27.475 ;
    RECT 151.35 27.765 151.56 27.835 ;
    RECT 151.35 28.125 151.56 28.195 ;
    RECT 147.57 27.405 147.78 27.475 ;
    RECT 147.57 27.765 147.78 27.835 ;
    RECT 147.57 28.125 147.78 28.195 ;
    RECT 148.03 27.405 148.24 27.475 ;
    RECT 148.03 27.765 148.24 27.835 ;
    RECT 148.03 28.125 148.24 28.195 ;
    RECT 144.25 27.405 144.46 27.475 ;
    RECT 144.25 27.765 144.46 27.835 ;
    RECT 144.25 28.125 144.46 28.195 ;
    RECT 144.71 27.405 144.92 27.475 ;
    RECT 144.71 27.765 144.92 27.835 ;
    RECT 144.71 28.125 144.92 28.195 ;
    RECT 140.93 27.405 141.14 27.475 ;
    RECT 140.93 27.765 141.14 27.835 ;
    RECT 140.93 28.125 141.14 28.195 ;
    RECT 141.39 27.405 141.6 27.475 ;
    RECT 141.39 27.765 141.6 27.835 ;
    RECT 141.39 28.125 141.6 28.195 ;
    RECT 137.61 27.405 137.82 27.475 ;
    RECT 137.61 27.765 137.82 27.835 ;
    RECT 137.61 28.125 137.82 28.195 ;
    RECT 138.07 27.405 138.28 27.475 ;
    RECT 138.07 27.765 138.28 27.835 ;
    RECT 138.07 28.125 138.28 28.195 ;
    RECT 134.29 27.405 134.5 27.475 ;
    RECT 134.29 27.765 134.5 27.835 ;
    RECT 134.29 28.125 134.5 28.195 ;
    RECT 134.75 27.405 134.96 27.475 ;
    RECT 134.75 27.765 134.96 27.835 ;
    RECT 134.75 28.125 134.96 28.195 ;
    RECT 64.57 27.405 64.78 27.475 ;
    RECT 64.57 27.765 64.78 27.835 ;
    RECT 64.57 28.125 64.78 28.195 ;
    RECT 65.03 27.405 65.24 27.475 ;
    RECT 65.03 27.765 65.24 27.835 ;
    RECT 65.03 28.125 65.24 28.195 ;
    RECT 61.25 26.685 61.46 26.755 ;
    RECT 61.25 27.045 61.46 27.115 ;
    RECT 61.25 27.405 61.46 27.475 ;
    RECT 61.71 26.685 61.92 26.755 ;
    RECT 61.71 27.045 61.92 27.115 ;
    RECT 61.71 27.405 61.92 27.475 ;
    RECT 57.93 26.685 58.14 26.755 ;
    RECT 57.93 27.045 58.14 27.115 ;
    RECT 57.93 27.405 58.14 27.475 ;
    RECT 58.39 26.685 58.6 26.755 ;
    RECT 58.39 27.045 58.6 27.115 ;
    RECT 58.39 27.405 58.6 27.475 ;
    RECT 54.61 26.685 54.82 26.755 ;
    RECT 54.61 27.045 54.82 27.115 ;
    RECT 54.61 27.405 54.82 27.475 ;
    RECT 55.07 26.685 55.28 26.755 ;
    RECT 55.07 27.045 55.28 27.115 ;
    RECT 55.07 27.405 55.28 27.475 ;
    RECT 51.29 26.685 51.5 26.755 ;
    RECT 51.29 27.045 51.5 27.115 ;
    RECT 51.29 27.405 51.5 27.475 ;
    RECT 51.75 26.685 51.96 26.755 ;
    RECT 51.75 27.045 51.96 27.115 ;
    RECT 51.75 27.405 51.96 27.475 ;
    RECT 47.97 26.685 48.18 26.755 ;
    RECT 47.97 27.045 48.18 27.115 ;
    RECT 47.97 27.405 48.18 27.475 ;
    RECT 48.43 26.685 48.64 26.755 ;
    RECT 48.43 27.045 48.64 27.115 ;
    RECT 48.43 27.405 48.64 27.475 ;
    RECT 44.65 26.685 44.86 26.755 ;
    RECT 44.65 27.045 44.86 27.115 ;
    RECT 44.65 27.405 44.86 27.475 ;
    RECT 45.11 26.685 45.32 26.755 ;
    RECT 45.11 27.045 45.32 27.115 ;
    RECT 45.11 27.405 45.32 27.475 ;
    RECT 41.33 26.685 41.54 26.755 ;
    RECT 41.33 27.045 41.54 27.115 ;
    RECT 41.33 27.405 41.54 27.475 ;
    RECT 41.79 26.685 42.0 26.755 ;
    RECT 41.79 27.045 42.0 27.115 ;
    RECT 41.79 27.405 42.0 27.475 ;
    RECT 38.01 26.685 38.22 26.755 ;
    RECT 38.01 27.045 38.22 27.115 ;
    RECT 38.01 27.405 38.22 27.475 ;
    RECT 38.47 26.685 38.68 26.755 ;
    RECT 38.47 27.045 38.68 27.115 ;
    RECT 38.47 27.405 38.68 27.475 ;
    RECT 34.69 26.685 34.9 26.755 ;
    RECT 34.69 27.045 34.9 27.115 ;
    RECT 34.69 27.405 34.9 27.475 ;
    RECT 35.15 26.685 35.36 26.755 ;
    RECT 35.15 27.045 35.36 27.115 ;
    RECT 35.15 27.405 35.36 27.475 ;
    RECT 173.945 27.045 174.015 27.115 ;
    RECT 130.97 26.685 131.18 26.755 ;
    RECT 130.97 27.045 131.18 27.115 ;
    RECT 130.97 27.405 131.18 27.475 ;
    RECT 131.43 26.685 131.64 26.755 ;
    RECT 131.43 27.045 131.64 27.115 ;
    RECT 131.43 27.405 131.64 27.475 ;
    RECT 127.65 26.685 127.86 26.755 ;
    RECT 127.65 27.045 127.86 27.115 ;
    RECT 127.65 27.405 127.86 27.475 ;
    RECT 128.11 26.685 128.32 26.755 ;
    RECT 128.11 27.045 128.32 27.115 ;
    RECT 128.11 27.405 128.32 27.475 ;
    RECT 124.33 26.685 124.54 26.755 ;
    RECT 124.33 27.045 124.54 27.115 ;
    RECT 124.33 27.405 124.54 27.475 ;
    RECT 124.79 26.685 125.0 26.755 ;
    RECT 124.79 27.045 125.0 27.115 ;
    RECT 124.79 27.405 125.0 27.475 ;
    RECT 121.01 26.685 121.22 26.755 ;
    RECT 121.01 27.045 121.22 27.115 ;
    RECT 121.01 27.405 121.22 27.475 ;
    RECT 121.47 26.685 121.68 26.755 ;
    RECT 121.47 27.045 121.68 27.115 ;
    RECT 121.47 27.405 121.68 27.475 ;
    RECT 117.69 26.685 117.9 26.755 ;
    RECT 117.69 27.045 117.9 27.115 ;
    RECT 117.69 27.405 117.9 27.475 ;
    RECT 118.15 26.685 118.36 26.755 ;
    RECT 118.15 27.045 118.36 27.115 ;
    RECT 118.15 27.405 118.36 27.475 ;
    RECT 114.37 26.685 114.58 26.755 ;
    RECT 114.37 27.045 114.58 27.115 ;
    RECT 114.37 27.405 114.58 27.475 ;
    RECT 114.83 26.685 115.04 26.755 ;
    RECT 114.83 27.045 115.04 27.115 ;
    RECT 114.83 27.405 115.04 27.475 ;
    RECT 111.05 26.685 111.26 26.755 ;
    RECT 111.05 27.045 111.26 27.115 ;
    RECT 111.05 27.405 111.26 27.475 ;
    RECT 111.51 26.685 111.72 26.755 ;
    RECT 111.51 27.045 111.72 27.115 ;
    RECT 111.51 27.405 111.72 27.475 ;
    RECT 107.73 26.685 107.94 26.755 ;
    RECT 107.73 27.045 107.94 27.115 ;
    RECT 107.73 27.405 107.94 27.475 ;
    RECT 108.19 26.685 108.4 26.755 ;
    RECT 108.19 27.045 108.4 27.115 ;
    RECT 108.19 27.405 108.4 27.475 ;
    RECT 104.41 26.685 104.62 26.755 ;
    RECT 104.41 27.045 104.62 27.115 ;
    RECT 104.41 27.405 104.62 27.475 ;
    RECT 104.87 26.685 105.08 26.755 ;
    RECT 104.87 27.045 105.08 27.115 ;
    RECT 104.87 27.405 105.08 27.475 ;
    RECT 101.09 26.685 101.3 26.755 ;
    RECT 101.09 27.045 101.3 27.115 ;
    RECT 101.09 27.405 101.3 27.475 ;
    RECT 101.55 26.685 101.76 26.755 ;
    RECT 101.55 27.045 101.76 27.115 ;
    RECT 101.55 27.405 101.76 27.475 ;
    RECT 0.4 27.045 0.47 27.115 ;
    RECT 170.81 26.685 171.02 26.755 ;
    RECT 170.81 27.045 171.02 27.115 ;
    RECT 170.81 27.405 171.02 27.475 ;
    RECT 171.27 26.685 171.48 26.755 ;
    RECT 171.27 27.045 171.48 27.115 ;
    RECT 171.27 27.405 171.48 27.475 ;
    RECT 167.49 26.685 167.7 26.755 ;
    RECT 167.49 27.045 167.7 27.115 ;
    RECT 167.49 27.405 167.7 27.475 ;
    RECT 167.95 26.685 168.16 26.755 ;
    RECT 167.95 27.045 168.16 27.115 ;
    RECT 167.95 27.405 168.16 27.475 ;
    RECT 97.77 26.685 97.98 26.755 ;
    RECT 97.77 27.045 97.98 27.115 ;
    RECT 97.77 27.405 97.98 27.475 ;
    RECT 98.23 26.685 98.44 26.755 ;
    RECT 98.23 27.045 98.44 27.115 ;
    RECT 98.23 27.405 98.44 27.475 ;
    RECT 94.45 26.685 94.66 26.755 ;
    RECT 94.45 27.045 94.66 27.115 ;
    RECT 94.45 27.405 94.66 27.475 ;
    RECT 94.91 26.685 95.12 26.755 ;
    RECT 94.91 27.045 95.12 27.115 ;
    RECT 94.91 27.405 95.12 27.475 ;
    RECT 91.13 26.685 91.34 26.755 ;
    RECT 91.13 27.045 91.34 27.115 ;
    RECT 91.13 27.405 91.34 27.475 ;
    RECT 91.59 26.685 91.8 26.755 ;
    RECT 91.59 27.045 91.8 27.115 ;
    RECT 91.59 27.405 91.8 27.475 ;
    RECT 87.81 26.685 88.02 26.755 ;
    RECT 87.81 27.045 88.02 27.115 ;
    RECT 87.81 27.405 88.02 27.475 ;
    RECT 88.27 26.685 88.48 26.755 ;
    RECT 88.27 27.045 88.48 27.115 ;
    RECT 88.27 27.405 88.48 27.475 ;
    RECT 84.49 26.685 84.7 26.755 ;
    RECT 84.49 27.045 84.7 27.115 ;
    RECT 84.49 27.405 84.7 27.475 ;
    RECT 84.95 26.685 85.16 26.755 ;
    RECT 84.95 27.045 85.16 27.115 ;
    RECT 84.95 27.405 85.16 27.475 ;
    RECT 81.17 26.685 81.38 26.755 ;
    RECT 81.17 27.045 81.38 27.115 ;
    RECT 81.17 27.405 81.38 27.475 ;
    RECT 81.63 26.685 81.84 26.755 ;
    RECT 81.63 27.045 81.84 27.115 ;
    RECT 81.63 27.405 81.84 27.475 ;
    RECT 77.85 26.685 78.06 26.755 ;
    RECT 77.85 27.045 78.06 27.115 ;
    RECT 77.85 27.405 78.06 27.475 ;
    RECT 78.31 26.685 78.52 26.755 ;
    RECT 78.31 27.045 78.52 27.115 ;
    RECT 78.31 27.405 78.52 27.475 ;
    RECT 74.53 26.685 74.74 26.755 ;
    RECT 74.53 27.045 74.74 27.115 ;
    RECT 74.53 27.405 74.74 27.475 ;
    RECT 74.99 26.685 75.2 26.755 ;
    RECT 74.99 27.045 75.2 27.115 ;
    RECT 74.99 27.405 75.2 27.475 ;
    RECT 71.21 26.685 71.42 26.755 ;
    RECT 71.21 27.045 71.42 27.115 ;
    RECT 71.21 27.405 71.42 27.475 ;
    RECT 71.67 26.685 71.88 26.755 ;
    RECT 71.67 27.045 71.88 27.115 ;
    RECT 71.67 27.405 71.88 27.475 ;
    RECT 31.37 26.685 31.58 26.755 ;
    RECT 31.37 27.045 31.58 27.115 ;
    RECT 31.37 27.405 31.58 27.475 ;
    RECT 31.83 26.685 32.04 26.755 ;
    RECT 31.83 27.045 32.04 27.115 ;
    RECT 31.83 27.405 32.04 27.475 ;
    RECT 67.89 26.685 68.1 26.755 ;
    RECT 67.89 27.045 68.1 27.115 ;
    RECT 67.89 27.405 68.1 27.475 ;
    RECT 68.35 26.685 68.56 26.755 ;
    RECT 68.35 27.045 68.56 27.115 ;
    RECT 68.35 27.405 68.56 27.475 ;
    RECT 28.05 26.685 28.26 26.755 ;
    RECT 28.05 27.045 28.26 27.115 ;
    RECT 28.05 27.405 28.26 27.475 ;
    RECT 28.51 26.685 28.72 26.755 ;
    RECT 28.51 27.045 28.72 27.115 ;
    RECT 28.51 27.405 28.72 27.475 ;
    RECT 24.73 26.685 24.94 26.755 ;
    RECT 24.73 27.045 24.94 27.115 ;
    RECT 24.73 27.405 24.94 27.475 ;
    RECT 25.19 26.685 25.4 26.755 ;
    RECT 25.19 27.045 25.4 27.115 ;
    RECT 25.19 27.405 25.4 27.475 ;
    RECT 21.41 26.685 21.62 26.755 ;
    RECT 21.41 27.045 21.62 27.115 ;
    RECT 21.41 27.405 21.62 27.475 ;
    RECT 21.87 26.685 22.08 26.755 ;
    RECT 21.87 27.045 22.08 27.115 ;
    RECT 21.87 27.405 22.08 27.475 ;
    RECT 18.09 26.685 18.3 26.755 ;
    RECT 18.09 27.045 18.3 27.115 ;
    RECT 18.09 27.405 18.3 27.475 ;
    RECT 18.55 26.685 18.76 26.755 ;
    RECT 18.55 27.045 18.76 27.115 ;
    RECT 18.55 27.405 18.76 27.475 ;
    RECT 14.77 26.685 14.98 26.755 ;
    RECT 14.77 27.045 14.98 27.115 ;
    RECT 14.77 27.405 14.98 27.475 ;
    RECT 15.23 26.685 15.44 26.755 ;
    RECT 15.23 27.045 15.44 27.115 ;
    RECT 15.23 27.405 15.44 27.475 ;
    RECT 11.45 26.685 11.66 26.755 ;
    RECT 11.45 27.045 11.66 27.115 ;
    RECT 11.45 27.405 11.66 27.475 ;
    RECT 11.91 26.685 12.12 26.755 ;
    RECT 11.91 27.045 12.12 27.115 ;
    RECT 11.91 27.405 12.12 27.475 ;
    RECT 8.13 26.685 8.34 26.755 ;
    RECT 8.13 27.045 8.34 27.115 ;
    RECT 8.13 27.405 8.34 27.475 ;
    RECT 8.59 26.685 8.8 26.755 ;
    RECT 8.59 27.045 8.8 27.115 ;
    RECT 8.59 27.405 8.8 27.475 ;
    RECT 4.81 26.685 5.02 26.755 ;
    RECT 4.81 27.045 5.02 27.115 ;
    RECT 4.81 27.405 5.02 27.475 ;
    RECT 5.27 26.685 5.48 26.755 ;
    RECT 5.27 27.045 5.48 27.115 ;
    RECT 5.27 27.405 5.48 27.475 ;
    RECT 164.17 26.685 164.38 26.755 ;
    RECT 164.17 27.045 164.38 27.115 ;
    RECT 164.17 27.405 164.38 27.475 ;
    RECT 164.63 26.685 164.84 26.755 ;
    RECT 164.63 27.045 164.84 27.115 ;
    RECT 164.63 27.405 164.84 27.475 ;
    RECT 1.49 26.685 1.7 26.755 ;
    RECT 1.49 27.045 1.7 27.115 ;
    RECT 1.49 27.405 1.7 27.475 ;
    RECT 1.95 26.685 2.16 26.755 ;
    RECT 1.95 27.045 2.16 27.115 ;
    RECT 1.95 27.405 2.16 27.475 ;
    RECT 160.85 26.685 161.06 26.755 ;
    RECT 160.85 27.045 161.06 27.115 ;
    RECT 160.85 27.405 161.06 27.475 ;
    RECT 161.31 26.685 161.52 26.755 ;
    RECT 161.31 27.045 161.52 27.115 ;
    RECT 161.31 27.405 161.52 27.475 ;
    RECT 157.53 26.685 157.74 26.755 ;
    RECT 157.53 27.045 157.74 27.115 ;
    RECT 157.53 27.405 157.74 27.475 ;
    RECT 157.99 26.685 158.2 26.755 ;
    RECT 157.99 27.045 158.2 27.115 ;
    RECT 157.99 27.405 158.2 27.475 ;
    RECT 154.21 26.685 154.42 26.755 ;
    RECT 154.21 27.045 154.42 27.115 ;
    RECT 154.21 27.405 154.42 27.475 ;
    RECT 154.67 26.685 154.88 26.755 ;
    RECT 154.67 27.045 154.88 27.115 ;
    RECT 154.67 27.405 154.88 27.475 ;
    RECT 150.89 26.685 151.1 26.755 ;
    RECT 150.89 27.045 151.1 27.115 ;
    RECT 150.89 27.405 151.1 27.475 ;
    RECT 151.35 26.685 151.56 26.755 ;
    RECT 151.35 27.045 151.56 27.115 ;
    RECT 151.35 27.405 151.56 27.475 ;
    RECT 147.57 26.685 147.78 26.755 ;
    RECT 147.57 27.045 147.78 27.115 ;
    RECT 147.57 27.405 147.78 27.475 ;
    RECT 148.03 26.685 148.24 26.755 ;
    RECT 148.03 27.045 148.24 27.115 ;
    RECT 148.03 27.405 148.24 27.475 ;
    RECT 144.25 26.685 144.46 26.755 ;
    RECT 144.25 27.045 144.46 27.115 ;
    RECT 144.25 27.405 144.46 27.475 ;
    RECT 144.71 26.685 144.92 26.755 ;
    RECT 144.71 27.045 144.92 27.115 ;
    RECT 144.71 27.405 144.92 27.475 ;
    RECT 140.93 26.685 141.14 26.755 ;
    RECT 140.93 27.045 141.14 27.115 ;
    RECT 140.93 27.405 141.14 27.475 ;
    RECT 141.39 26.685 141.6 26.755 ;
    RECT 141.39 27.045 141.6 27.115 ;
    RECT 141.39 27.405 141.6 27.475 ;
    RECT 137.61 26.685 137.82 26.755 ;
    RECT 137.61 27.045 137.82 27.115 ;
    RECT 137.61 27.405 137.82 27.475 ;
    RECT 138.07 26.685 138.28 26.755 ;
    RECT 138.07 27.045 138.28 27.115 ;
    RECT 138.07 27.405 138.28 27.475 ;
    RECT 134.29 26.685 134.5 26.755 ;
    RECT 134.29 27.045 134.5 27.115 ;
    RECT 134.29 27.405 134.5 27.475 ;
    RECT 134.75 26.685 134.96 26.755 ;
    RECT 134.75 27.045 134.96 27.115 ;
    RECT 134.75 27.405 134.96 27.475 ;
    RECT 64.57 26.685 64.78 26.755 ;
    RECT 64.57 27.045 64.78 27.115 ;
    RECT 64.57 27.405 64.78 27.475 ;
    RECT 65.03 26.685 65.24 26.755 ;
    RECT 65.03 27.045 65.24 27.115 ;
    RECT 65.03 27.405 65.24 27.475 ;
    RECT 61.25 25.965 61.46 26.035 ;
    RECT 61.25 26.325 61.46 26.395 ;
    RECT 61.25 26.685 61.46 26.755 ;
    RECT 61.71 25.965 61.92 26.035 ;
    RECT 61.71 26.325 61.92 26.395 ;
    RECT 61.71 26.685 61.92 26.755 ;
    RECT 57.93 25.965 58.14 26.035 ;
    RECT 57.93 26.325 58.14 26.395 ;
    RECT 57.93 26.685 58.14 26.755 ;
    RECT 58.39 25.965 58.6 26.035 ;
    RECT 58.39 26.325 58.6 26.395 ;
    RECT 58.39 26.685 58.6 26.755 ;
    RECT 54.61 25.965 54.82 26.035 ;
    RECT 54.61 26.325 54.82 26.395 ;
    RECT 54.61 26.685 54.82 26.755 ;
    RECT 55.07 25.965 55.28 26.035 ;
    RECT 55.07 26.325 55.28 26.395 ;
    RECT 55.07 26.685 55.28 26.755 ;
    RECT 51.29 25.965 51.5 26.035 ;
    RECT 51.29 26.325 51.5 26.395 ;
    RECT 51.29 26.685 51.5 26.755 ;
    RECT 51.75 25.965 51.96 26.035 ;
    RECT 51.75 26.325 51.96 26.395 ;
    RECT 51.75 26.685 51.96 26.755 ;
    RECT 47.97 25.965 48.18 26.035 ;
    RECT 47.97 26.325 48.18 26.395 ;
    RECT 47.97 26.685 48.18 26.755 ;
    RECT 48.43 25.965 48.64 26.035 ;
    RECT 48.43 26.325 48.64 26.395 ;
    RECT 48.43 26.685 48.64 26.755 ;
    RECT 44.65 25.965 44.86 26.035 ;
    RECT 44.65 26.325 44.86 26.395 ;
    RECT 44.65 26.685 44.86 26.755 ;
    RECT 45.11 25.965 45.32 26.035 ;
    RECT 45.11 26.325 45.32 26.395 ;
    RECT 45.11 26.685 45.32 26.755 ;
    RECT 41.33 25.965 41.54 26.035 ;
    RECT 41.33 26.325 41.54 26.395 ;
    RECT 41.33 26.685 41.54 26.755 ;
    RECT 41.79 25.965 42.0 26.035 ;
    RECT 41.79 26.325 42.0 26.395 ;
    RECT 41.79 26.685 42.0 26.755 ;
    RECT 38.01 25.965 38.22 26.035 ;
    RECT 38.01 26.325 38.22 26.395 ;
    RECT 38.01 26.685 38.22 26.755 ;
    RECT 38.47 25.965 38.68 26.035 ;
    RECT 38.47 26.325 38.68 26.395 ;
    RECT 38.47 26.685 38.68 26.755 ;
    RECT 34.69 25.965 34.9 26.035 ;
    RECT 34.69 26.325 34.9 26.395 ;
    RECT 34.69 26.685 34.9 26.755 ;
    RECT 35.15 25.965 35.36 26.035 ;
    RECT 35.15 26.325 35.36 26.395 ;
    RECT 35.15 26.685 35.36 26.755 ;
    RECT 173.945 26.325 174.015 26.395 ;
    RECT 130.97 25.965 131.18 26.035 ;
    RECT 130.97 26.325 131.18 26.395 ;
    RECT 130.97 26.685 131.18 26.755 ;
    RECT 131.43 25.965 131.64 26.035 ;
    RECT 131.43 26.325 131.64 26.395 ;
    RECT 131.43 26.685 131.64 26.755 ;
    RECT 127.65 25.965 127.86 26.035 ;
    RECT 127.65 26.325 127.86 26.395 ;
    RECT 127.65 26.685 127.86 26.755 ;
    RECT 128.11 25.965 128.32 26.035 ;
    RECT 128.11 26.325 128.32 26.395 ;
    RECT 128.11 26.685 128.32 26.755 ;
    RECT 124.33 25.965 124.54 26.035 ;
    RECT 124.33 26.325 124.54 26.395 ;
    RECT 124.33 26.685 124.54 26.755 ;
    RECT 124.79 25.965 125.0 26.035 ;
    RECT 124.79 26.325 125.0 26.395 ;
    RECT 124.79 26.685 125.0 26.755 ;
    RECT 121.01 25.965 121.22 26.035 ;
    RECT 121.01 26.325 121.22 26.395 ;
    RECT 121.01 26.685 121.22 26.755 ;
    RECT 121.47 25.965 121.68 26.035 ;
    RECT 121.47 26.325 121.68 26.395 ;
    RECT 121.47 26.685 121.68 26.755 ;
    RECT 117.69 25.965 117.9 26.035 ;
    RECT 117.69 26.325 117.9 26.395 ;
    RECT 117.69 26.685 117.9 26.755 ;
    RECT 118.15 25.965 118.36 26.035 ;
    RECT 118.15 26.325 118.36 26.395 ;
    RECT 118.15 26.685 118.36 26.755 ;
    RECT 114.37 25.965 114.58 26.035 ;
    RECT 114.37 26.325 114.58 26.395 ;
    RECT 114.37 26.685 114.58 26.755 ;
    RECT 114.83 25.965 115.04 26.035 ;
    RECT 114.83 26.325 115.04 26.395 ;
    RECT 114.83 26.685 115.04 26.755 ;
    RECT 111.05 25.965 111.26 26.035 ;
    RECT 111.05 26.325 111.26 26.395 ;
    RECT 111.05 26.685 111.26 26.755 ;
    RECT 111.51 25.965 111.72 26.035 ;
    RECT 111.51 26.325 111.72 26.395 ;
    RECT 111.51 26.685 111.72 26.755 ;
    RECT 107.73 25.965 107.94 26.035 ;
    RECT 107.73 26.325 107.94 26.395 ;
    RECT 107.73 26.685 107.94 26.755 ;
    RECT 108.19 25.965 108.4 26.035 ;
    RECT 108.19 26.325 108.4 26.395 ;
    RECT 108.19 26.685 108.4 26.755 ;
    RECT 104.41 25.965 104.62 26.035 ;
    RECT 104.41 26.325 104.62 26.395 ;
    RECT 104.41 26.685 104.62 26.755 ;
    RECT 104.87 25.965 105.08 26.035 ;
    RECT 104.87 26.325 105.08 26.395 ;
    RECT 104.87 26.685 105.08 26.755 ;
    RECT 101.09 25.965 101.3 26.035 ;
    RECT 101.09 26.325 101.3 26.395 ;
    RECT 101.09 26.685 101.3 26.755 ;
    RECT 101.55 25.965 101.76 26.035 ;
    RECT 101.55 26.325 101.76 26.395 ;
    RECT 101.55 26.685 101.76 26.755 ;
    RECT 0.4 26.325 0.47 26.395 ;
    RECT 170.81 25.965 171.02 26.035 ;
    RECT 170.81 26.325 171.02 26.395 ;
    RECT 170.81 26.685 171.02 26.755 ;
    RECT 171.27 25.965 171.48 26.035 ;
    RECT 171.27 26.325 171.48 26.395 ;
    RECT 171.27 26.685 171.48 26.755 ;
    RECT 167.49 25.965 167.7 26.035 ;
    RECT 167.49 26.325 167.7 26.395 ;
    RECT 167.49 26.685 167.7 26.755 ;
    RECT 167.95 25.965 168.16 26.035 ;
    RECT 167.95 26.325 168.16 26.395 ;
    RECT 167.95 26.685 168.16 26.755 ;
    RECT 97.77 25.965 97.98 26.035 ;
    RECT 97.77 26.325 97.98 26.395 ;
    RECT 97.77 26.685 97.98 26.755 ;
    RECT 98.23 25.965 98.44 26.035 ;
    RECT 98.23 26.325 98.44 26.395 ;
    RECT 98.23 26.685 98.44 26.755 ;
    RECT 94.45 25.965 94.66 26.035 ;
    RECT 94.45 26.325 94.66 26.395 ;
    RECT 94.45 26.685 94.66 26.755 ;
    RECT 94.91 25.965 95.12 26.035 ;
    RECT 94.91 26.325 95.12 26.395 ;
    RECT 94.91 26.685 95.12 26.755 ;
    RECT 91.13 25.965 91.34 26.035 ;
    RECT 91.13 26.325 91.34 26.395 ;
    RECT 91.13 26.685 91.34 26.755 ;
    RECT 91.59 25.965 91.8 26.035 ;
    RECT 91.59 26.325 91.8 26.395 ;
    RECT 91.59 26.685 91.8 26.755 ;
    RECT 87.81 25.965 88.02 26.035 ;
    RECT 87.81 26.325 88.02 26.395 ;
    RECT 87.81 26.685 88.02 26.755 ;
    RECT 88.27 25.965 88.48 26.035 ;
    RECT 88.27 26.325 88.48 26.395 ;
    RECT 88.27 26.685 88.48 26.755 ;
    RECT 84.49 25.965 84.7 26.035 ;
    RECT 84.49 26.325 84.7 26.395 ;
    RECT 84.49 26.685 84.7 26.755 ;
    RECT 84.95 25.965 85.16 26.035 ;
    RECT 84.95 26.325 85.16 26.395 ;
    RECT 84.95 26.685 85.16 26.755 ;
    RECT 81.17 25.965 81.38 26.035 ;
    RECT 81.17 26.325 81.38 26.395 ;
    RECT 81.17 26.685 81.38 26.755 ;
    RECT 81.63 25.965 81.84 26.035 ;
    RECT 81.63 26.325 81.84 26.395 ;
    RECT 81.63 26.685 81.84 26.755 ;
    RECT 77.85 25.965 78.06 26.035 ;
    RECT 77.85 26.325 78.06 26.395 ;
    RECT 77.85 26.685 78.06 26.755 ;
    RECT 78.31 25.965 78.52 26.035 ;
    RECT 78.31 26.325 78.52 26.395 ;
    RECT 78.31 26.685 78.52 26.755 ;
    RECT 74.53 25.965 74.74 26.035 ;
    RECT 74.53 26.325 74.74 26.395 ;
    RECT 74.53 26.685 74.74 26.755 ;
    RECT 74.99 25.965 75.2 26.035 ;
    RECT 74.99 26.325 75.2 26.395 ;
    RECT 74.99 26.685 75.2 26.755 ;
    RECT 71.21 25.965 71.42 26.035 ;
    RECT 71.21 26.325 71.42 26.395 ;
    RECT 71.21 26.685 71.42 26.755 ;
    RECT 71.67 25.965 71.88 26.035 ;
    RECT 71.67 26.325 71.88 26.395 ;
    RECT 71.67 26.685 71.88 26.755 ;
    RECT 31.37 25.965 31.58 26.035 ;
    RECT 31.37 26.325 31.58 26.395 ;
    RECT 31.37 26.685 31.58 26.755 ;
    RECT 31.83 25.965 32.04 26.035 ;
    RECT 31.83 26.325 32.04 26.395 ;
    RECT 31.83 26.685 32.04 26.755 ;
    RECT 67.89 25.965 68.1 26.035 ;
    RECT 67.89 26.325 68.1 26.395 ;
    RECT 67.89 26.685 68.1 26.755 ;
    RECT 68.35 25.965 68.56 26.035 ;
    RECT 68.35 26.325 68.56 26.395 ;
    RECT 68.35 26.685 68.56 26.755 ;
    RECT 28.05 25.965 28.26 26.035 ;
    RECT 28.05 26.325 28.26 26.395 ;
    RECT 28.05 26.685 28.26 26.755 ;
    RECT 28.51 25.965 28.72 26.035 ;
    RECT 28.51 26.325 28.72 26.395 ;
    RECT 28.51 26.685 28.72 26.755 ;
    RECT 24.73 25.965 24.94 26.035 ;
    RECT 24.73 26.325 24.94 26.395 ;
    RECT 24.73 26.685 24.94 26.755 ;
    RECT 25.19 25.965 25.4 26.035 ;
    RECT 25.19 26.325 25.4 26.395 ;
    RECT 25.19 26.685 25.4 26.755 ;
    RECT 21.41 25.965 21.62 26.035 ;
    RECT 21.41 26.325 21.62 26.395 ;
    RECT 21.41 26.685 21.62 26.755 ;
    RECT 21.87 25.965 22.08 26.035 ;
    RECT 21.87 26.325 22.08 26.395 ;
    RECT 21.87 26.685 22.08 26.755 ;
    RECT 18.09 25.965 18.3 26.035 ;
    RECT 18.09 26.325 18.3 26.395 ;
    RECT 18.09 26.685 18.3 26.755 ;
    RECT 18.55 25.965 18.76 26.035 ;
    RECT 18.55 26.325 18.76 26.395 ;
    RECT 18.55 26.685 18.76 26.755 ;
    RECT 14.77 25.965 14.98 26.035 ;
    RECT 14.77 26.325 14.98 26.395 ;
    RECT 14.77 26.685 14.98 26.755 ;
    RECT 15.23 25.965 15.44 26.035 ;
    RECT 15.23 26.325 15.44 26.395 ;
    RECT 15.23 26.685 15.44 26.755 ;
    RECT 11.45 25.965 11.66 26.035 ;
    RECT 11.45 26.325 11.66 26.395 ;
    RECT 11.45 26.685 11.66 26.755 ;
    RECT 11.91 25.965 12.12 26.035 ;
    RECT 11.91 26.325 12.12 26.395 ;
    RECT 11.91 26.685 12.12 26.755 ;
    RECT 8.13 25.965 8.34 26.035 ;
    RECT 8.13 26.325 8.34 26.395 ;
    RECT 8.13 26.685 8.34 26.755 ;
    RECT 8.59 25.965 8.8 26.035 ;
    RECT 8.59 26.325 8.8 26.395 ;
    RECT 8.59 26.685 8.8 26.755 ;
    RECT 4.81 25.965 5.02 26.035 ;
    RECT 4.81 26.325 5.02 26.395 ;
    RECT 4.81 26.685 5.02 26.755 ;
    RECT 5.27 25.965 5.48 26.035 ;
    RECT 5.27 26.325 5.48 26.395 ;
    RECT 5.27 26.685 5.48 26.755 ;
    RECT 164.17 25.965 164.38 26.035 ;
    RECT 164.17 26.325 164.38 26.395 ;
    RECT 164.17 26.685 164.38 26.755 ;
    RECT 164.63 25.965 164.84 26.035 ;
    RECT 164.63 26.325 164.84 26.395 ;
    RECT 164.63 26.685 164.84 26.755 ;
    RECT 1.49 25.965 1.7 26.035 ;
    RECT 1.49 26.325 1.7 26.395 ;
    RECT 1.49 26.685 1.7 26.755 ;
    RECT 1.95 25.965 2.16 26.035 ;
    RECT 1.95 26.325 2.16 26.395 ;
    RECT 1.95 26.685 2.16 26.755 ;
    RECT 160.85 25.965 161.06 26.035 ;
    RECT 160.85 26.325 161.06 26.395 ;
    RECT 160.85 26.685 161.06 26.755 ;
    RECT 161.31 25.965 161.52 26.035 ;
    RECT 161.31 26.325 161.52 26.395 ;
    RECT 161.31 26.685 161.52 26.755 ;
    RECT 157.53 25.965 157.74 26.035 ;
    RECT 157.53 26.325 157.74 26.395 ;
    RECT 157.53 26.685 157.74 26.755 ;
    RECT 157.99 25.965 158.2 26.035 ;
    RECT 157.99 26.325 158.2 26.395 ;
    RECT 157.99 26.685 158.2 26.755 ;
    RECT 154.21 25.965 154.42 26.035 ;
    RECT 154.21 26.325 154.42 26.395 ;
    RECT 154.21 26.685 154.42 26.755 ;
    RECT 154.67 25.965 154.88 26.035 ;
    RECT 154.67 26.325 154.88 26.395 ;
    RECT 154.67 26.685 154.88 26.755 ;
    RECT 150.89 25.965 151.1 26.035 ;
    RECT 150.89 26.325 151.1 26.395 ;
    RECT 150.89 26.685 151.1 26.755 ;
    RECT 151.35 25.965 151.56 26.035 ;
    RECT 151.35 26.325 151.56 26.395 ;
    RECT 151.35 26.685 151.56 26.755 ;
    RECT 147.57 25.965 147.78 26.035 ;
    RECT 147.57 26.325 147.78 26.395 ;
    RECT 147.57 26.685 147.78 26.755 ;
    RECT 148.03 25.965 148.24 26.035 ;
    RECT 148.03 26.325 148.24 26.395 ;
    RECT 148.03 26.685 148.24 26.755 ;
    RECT 144.25 25.965 144.46 26.035 ;
    RECT 144.25 26.325 144.46 26.395 ;
    RECT 144.25 26.685 144.46 26.755 ;
    RECT 144.71 25.965 144.92 26.035 ;
    RECT 144.71 26.325 144.92 26.395 ;
    RECT 144.71 26.685 144.92 26.755 ;
    RECT 140.93 25.965 141.14 26.035 ;
    RECT 140.93 26.325 141.14 26.395 ;
    RECT 140.93 26.685 141.14 26.755 ;
    RECT 141.39 25.965 141.6 26.035 ;
    RECT 141.39 26.325 141.6 26.395 ;
    RECT 141.39 26.685 141.6 26.755 ;
    RECT 137.61 25.965 137.82 26.035 ;
    RECT 137.61 26.325 137.82 26.395 ;
    RECT 137.61 26.685 137.82 26.755 ;
    RECT 138.07 25.965 138.28 26.035 ;
    RECT 138.07 26.325 138.28 26.395 ;
    RECT 138.07 26.685 138.28 26.755 ;
    RECT 134.29 25.965 134.5 26.035 ;
    RECT 134.29 26.325 134.5 26.395 ;
    RECT 134.29 26.685 134.5 26.755 ;
    RECT 134.75 25.965 134.96 26.035 ;
    RECT 134.75 26.325 134.96 26.395 ;
    RECT 134.75 26.685 134.96 26.755 ;
    RECT 64.57 25.965 64.78 26.035 ;
    RECT 64.57 26.325 64.78 26.395 ;
    RECT 64.57 26.685 64.78 26.755 ;
    RECT 65.03 25.965 65.24 26.035 ;
    RECT 65.03 26.325 65.24 26.395 ;
    RECT 65.03 26.685 65.24 26.755 ;
    RECT 61.25 25.245 61.46 25.315 ;
    RECT 61.25 25.605 61.46 25.675 ;
    RECT 61.25 25.965 61.46 26.035 ;
    RECT 61.71 25.245 61.92 25.315 ;
    RECT 61.71 25.605 61.92 25.675 ;
    RECT 61.71 25.965 61.92 26.035 ;
    RECT 57.93 25.245 58.14 25.315 ;
    RECT 57.93 25.605 58.14 25.675 ;
    RECT 57.93 25.965 58.14 26.035 ;
    RECT 58.39 25.245 58.6 25.315 ;
    RECT 58.39 25.605 58.6 25.675 ;
    RECT 58.39 25.965 58.6 26.035 ;
    RECT 54.61 25.245 54.82 25.315 ;
    RECT 54.61 25.605 54.82 25.675 ;
    RECT 54.61 25.965 54.82 26.035 ;
    RECT 55.07 25.245 55.28 25.315 ;
    RECT 55.07 25.605 55.28 25.675 ;
    RECT 55.07 25.965 55.28 26.035 ;
    RECT 51.29 25.245 51.5 25.315 ;
    RECT 51.29 25.605 51.5 25.675 ;
    RECT 51.29 25.965 51.5 26.035 ;
    RECT 51.75 25.245 51.96 25.315 ;
    RECT 51.75 25.605 51.96 25.675 ;
    RECT 51.75 25.965 51.96 26.035 ;
    RECT 47.97 25.245 48.18 25.315 ;
    RECT 47.97 25.605 48.18 25.675 ;
    RECT 47.97 25.965 48.18 26.035 ;
    RECT 48.43 25.245 48.64 25.315 ;
    RECT 48.43 25.605 48.64 25.675 ;
    RECT 48.43 25.965 48.64 26.035 ;
    RECT 44.65 25.245 44.86 25.315 ;
    RECT 44.65 25.605 44.86 25.675 ;
    RECT 44.65 25.965 44.86 26.035 ;
    RECT 45.11 25.245 45.32 25.315 ;
    RECT 45.11 25.605 45.32 25.675 ;
    RECT 45.11 25.965 45.32 26.035 ;
    RECT 41.33 25.245 41.54 25.315 ;
    RECT 41.33 25.605 41.54 25.675 ;
    RECT 41.33 25.965 41.54 26.035 ;
    RECT 41.79 25.245 42.0 25.315 ;
    RECT 41.79 25.605 42.0 25.675 ;
    RECT 41.79 25.965 42.0 26.035 ;
    RECT 38.01 25.245 38.22 25.315 ;
    RECT 38.01 25.605 38.22 25.675 ;
    RECT 38.01 25.965 38.22 26.035 ;
    RECT 38.47 25.245 38.68 25.315 ;
    RECT 38.47 25.605 38.68 25.675 ;
    RECT 38.47 25.965 38.68 26.035 ;
    RECT 34.69 25.245 34.9 25.315 ;
    RECT 34.69 25.605 34.9 25.675 ;
    RECT 34.69 25.965 34.9 26.035 ;
    RECT 35.15 25.245 35.36 25.315 ;
    RECT 35.15 25.605 35.36 25.675 ;
    RECT 35.15 25.965 35.36 26.035 ;
    RECT 173.945 25.605 174.015 25.675 ;
    RECT 130.97 25.245 131.18 25.315 ;
    RECT 130.97 25.605 131.18 25.675 ;
    RECT 130.97 25.965 131.18 26.035 ;
    RECT 131.43 25.245 131.64 25.315 ;
    RECT 131.43 25.605 131.64 25.675 ;
    RECT 131.43 25.965 131.64 26.035 ;
    RECT 127.65 25.245 127.86 25.315 ;
    RECT 127.65 25.605 127.86 25.675 ;
    RECT 127.65 25.965 127.86 26.035 ;
    RECT 128.11 25.245 128.32 25.315 ;
    RECT 128.11 25.605 128.32 25.675 ;
    RECT 128.11 25.965 128.32 26.035 ;
    RECT 124.33 25.245 124.54 25.315 ;
    RECT 124.33 25.605 124.54 25.675 ;
    RECT 124.33 25.965 124.54 26.035 ;
    RECT 124.79 25.245 125.0 25.315 ;
    RECT 124.79 25.605 125.0 25.675 ;
    RECT 124.79 25.965 125.0 26.035 ;
    RECT 121.01 25.245 121.22 25.315 ;
    RECT 121.01 25.605 121.22 25.675 ;
    RECT 121.01 25.965 121.22 26.035 ;
    RECT 121.47 25.245 121.68 25.315 ;
    RECT 121.47 25.605 121.68 25.675 ;
    RECT 121.47 25.965 121.68 26.035 ;
    RECT 117.69 25.245 117.9 25.315 ;
    RECT 117.69 25.605 117.9 25.675 ;
    RECT 117.69 25.965 117.9 26.035 ;
    RECT 118.15 25.245 118.36 25.315 ;
    RECT 118.15 25.605 118.36 25.675 ;
    RECT 118.15 25.965 118.36 26.035 ;
    RECT 114.37 25.245 114.58 25.315 ;
    RECT 114.37 25.605 114.58 25.675 ;
    RECT 114.37 25.965 114.58 26.035 ;
    RECT 114.83 25.245 115.04 25.315 ;
    RECT 114.83 25.605 115.04 25.675 ;
    RECT 114.83 25.965 115.04 26.035 ;
    RECT 111.05 25.245 111.26 25.315 ;
    RECT 111.05 25.605 111.26 25.675 ;
    RECT 111.05 25.965 111.26 26.035 ;
    RECT 111.51 25.245 111.72 25.315 ;
    RECT 111.51 25.605 111.72 25.675 ;
    RECT 111.51 25.965 111.72 26.035 ;
    RECT 107.73 25.245 107.94 25.315 ;
    RECT 107.73 25.605 107.94 25.675 ;
    RECT 107.73 25.965 107.94 26.035 ;
    RECT 108.19 25.245 108.4 25.315 ;
    RECT 108.19 25.605 108.4 25.675 ;
    RECT 108.19 25.965 108.4 26.035 ;
    RECT 104.41 25.245 104.62 25.315 ;
    RECT 104.41 25.605 104.62 25.675 ;
    RECT 104.41 25.965 104.62 26.035 ;
    RECT 104.87 25.245 105.08 25.315 ;
    RECT 104.87 25.605 105.08 25.675 ;
    RECT 104.87 25.965 105.08 26.035 ;
    RECT 101.09 25.245 101.3 25.315 ;
    RECT 101.09 25.605 101.3 25.675 ;
    RECT 101.09 25.965 101.3 26.035 ;
    RECT 101.55 25.245 101.76 25.315 ;
    RECT 101.55 25.605 101.76 25.675 ;
    RECT 101.55 25.965 101.76 26.035 ;
    RECT 0.4 25.605 0.47 25.675 ;
    RECT 170.81 25.245 171.02 25.315 ;
    RECT 170.81 25.605 171.02 25.675 ;
    RECT 170.81 25.965 171.02 26.035 ;
    RECT 171.27 25.245 171.48 25.315 ;
    RECT 171.27 25.605 171.48 25.675 ;
    RECT 171.27 25.965 171.48 26.035 ;
    RECT 167.49 25.245 167.7 25.315 ;
    RECT 167.49 25.605 167.7 25.675 ;
    RECT 167.49 25.965 167.7 26.035 ;
    RECT 167.95 25.245 168.16 25.315 ;
    RECT 167.95 25.605 168.16 25.675 ;
    RECT 167.95 25.965 168.16 26.035 ;
    RECT 97.77 25.245 97.98 25.315 ;
    RECT 97.77 25.605 97.98 25.675 ;
    RECT 97.77 25.965 97.98 26.035 ;
    RECT 98.23 25.245 98.44 25.315 ;
    RECT 98.23 25.605 98.44 25.675 ;
    RECT 98.23 25.965 98.44 26.035 ;
    RECT 94.45 25.245 94.66 25.315 ;
    RECT 94.45 25.605 94.66 25.675 ;
    RECT 94.45 25.965 94.66 26.035 ;
    RECT 94.91 25.245 95.12 25.315 ;
    RECT 94.91 25.605 95.12 25.675 ;
    RECT 94.91 25.965 95.12 26.035 ;
    RECT 91.13 25.245 91.34 25.315 ;
    RECT 91.13 25.605 91.34 25.675 ;
    RECT 91.13 25.965 91.34 26.035 ;
    RECT 91.59 25.245 91.8 25.315 ;
    RECT 91.59 25.605 91.8 25.675 ;
    RECT 91.59 25.965 91.8 26.035 ;
    RECT 87.81 25.245 88.02 25.315 ;
    RECT 87.81 25.605 88.02 25.675 ;
    RECT 87.81 25.965 88.02 26.035 ;
    RECT 88.27 25.245 88.48 25.315 ;
    RECT 88.27 25.605 88.48 25.675 ;
    RECT 88.27 25.965 88.48 26.035 ;
    RECT 84.49 25.245 84.7 25.315 ;
    RECT 84.49 25.605 84.7 25.675 ;
    RECT 84.49 25.965 84.7 26.035 ;
    RECT 84.95 25.245 85.16 25.315 ;
    RECT 84.95 25.605 85.16 25.675 ;
    RECT 84.95 25.965 85.16 26.035 ;
    RECT 81.17 25.245 81.38 25.315 ;
    RECT 81.17 25.605 81.38 25.675 ;
    RECT 81.17 25.965 81.38 26.035 ;
    RECT 81.63 25.245 81.84 25.315 ;
    RECT 81.63 25.605 81.84 25.675 ;
    RECT 81.63 25.965 81.84 26.035 ;
    RECT 77.85 25.245 78.06 25.315 ;
    RECT 77.85 25.605 78.06 25.675 ;
    RECT 77.85 25.965 78.06 26.035 ;
    RECT 78.31 25.245 78.52 25.315 ;
    RECT 78.31 25.605 78.52 25.675 ;
    RECT 78.31 25.965 78.52 26.035 ;
    RECT 74.53 25.245 74.74 25.315 ;
    RECT 74.53 25.605 74.74 25.675 ;
    RECT 74.53 25.965 74.74 26.035 ;
    RECT 74.99 25.245 75.2 25.315 ;
    RECT 74.99 25.605 75.2 25.675 ;
    RECT 74.99 25.965 75.2 26.035 ;
    RECT 71.21 25.245 71.42 25.315 ;
    RECT 71.21 25.605 71.42 25.675 ;
    RECT 71.21 25.965 71.42 26.035 ;
    RECT 71.67 25.245 71.88 25.315 ;
    RECT 71.67 25.605 71.88 25.675 ;
    RECT 71.67 25.965 71.88 26.035 ;
    RECT 31.37 25.245 31.58 25.315 ;
    RECT 31.37 25.605 31.58 25.675 ;
    RECT 31.37 25.965 31.58 26.035 ;
    RECT 31.83 25.245 32.04 25.315 ;
    RECT 31.83 25.605 32.04 25.675 ;
    RECT 31.83 25.965 32.04 26.035 ;
    RECT 67.89 25.245 68.1 25.315 ;
    RECT 67.89 25.605 68.1 25.675 ;
    RECT 67.89 25.965 68.1 26.035 ;
    RECT 68.35 25.245 68.56 25.315 ;
    RECT 68.35 25.605 68.56 25.675 ;
    RECT 68.35 25.965 68.56 26.035 ;
    RECT 28.05 25.245 28.26 25.315 ;
    RECT 28.05 25.605 28.26 25.675 ;
    RECT 28.05 25.965 28.26 26.035 ;
    RECT 28.51 25.245 28.72 25.315 ;
    RECT 28.51 25.605 28.72 25.675 ;
    RECT 28.51 25.965 28.72 26.035 ;
    RECT 24.73 25.245 24.94 25.315 ;
    RECT 24.73 25.605 24.94 25.675 ;
    RECT 24.73 25.965 24.94 26.035 ;
    RECT 25.19 25.245 25.4 25.315 ;
    RECT 25.19 25.605 25.4 25.675 ;
    RECT 25.19 25.965 25.4 26.035 ;
    RECT 21.41 25.245 21.62 25.315 ;
    RECT 21.41 25.605 21.62 25.675 ;
    RECT 21.41 25.965 21.62 26.035 ;
    RECT 21.87 25.245 22.08 25.315 ;
    RECT 21.87 25.605 22.08 25.675 ;
    RECT 21.87 25.965 22.08 26.035 ;
    RECT 18.09 25.245 18.3 25.315 ;
    RECT 18.09 25.605 18.3 25.675 ;
    RECT 18.09 25.965 18.3 26.035 ;
    RECT 18.55 25.245 18.76 25.315 ;
    RECT 18.55 25.605 18.76 25.675 ;
    RECT 18.55 25.965 18.76 26.035 ;
    RECT 14.77 25.245 14.98 25.315 ;
    RECT 14.77 25.605 14.98 25.675 ;
    RECT 14.77 25.965 14.98 26.035 ;
    RECT 15.23 25.245 15.44 25.315 ;
    RECT 15.23 25.605 15.44 25.675 ;
    RECT 15.23 25.965 15.44 26.035 ;
    RECT 11.45 25.245 11.66 25.315 ;
    RECT 11.45 25.605 11.66 25.675 ;
    RECT 11.45 25.965 11.66 26.035 ;
    RECT 11.91 25.245 12.12 25.315 ;
    RECT 11.91 25.605 12.12 25.675 ;
    RECT 11.91 25.965 12.12 26.035 ;
    RECT 8.13 25.245 8.34 25.315 ;
    RECT 8.13 25.605 8.34 25.675 ;
    RECT 8.13 25.965 8.34 26.035 ;
    RECT 8.59 25.245 8.8 25.315 ;
    RECT 8.59 25.605 8.8 25.675 ;
    RECT 8.59 25.965 8.8 26.035 ;
    RECT 4.81 25.245 5.02 25.315 ;
    RECT 4.81 25.605 5.02 25.675 ;
    RECT 4.81 25.965 5.02 26.035 ;
    RECT 5.27 25.245 5.48 25.315 ;
    RECT 5.27 25.605 5.48 25.675 ;
    RECT 5.27 25.965 5.48 26.035 ;
    RECT 164.17 25.245 164.38 25.315 ;
    RECT 164.17 25.605 164.38 25.675 ;
    RECT 164.17 25.965 164.38 26.035 ;
    RECT 164.63 25.245 164.84 25.315 ;
    RECT 164.63 25.605 164.84 25.675 ;
    RECT 164.63 25.965 164.84 26.035 ;
    RECT 1.49 25.245 1.7 25.315 ;
    RECT 1.49 25.605 1.7 25.675 ;
    RECT 1.49 25.965 1.7 26.035 ;
    RECT 1.95 25.245 2.16 25.315 ;
    RECT 1.95 25.605 2.16 25.675 ;
    RECT 1.95 25.965 2.16 26.035 ;
    RECT 160.85 25.245 161.06 25.315 ;
    RECT 160.85 25.605 161.06 25.675 ;
    RECT 160.85 25.965 161.06 26.035 ;
    RECT 161.31 25.245 161.52 25.315 ;
    RECT 161.31 25.605 161.52 25.675 ;
    RECT 161.31 25.965 161.52 26.035 ;
    RECT 157.53 25.245 157.74 25.315 ;
    RECT 157.53 25.605 157.74 25.675 ;
    RECT 157.53 25.965 157.74 26.035 ;
    RECT 157.99 25.245 158.2 25.315 ;
    RECT 157.99 25.605 158.2 25.675 ;
    RECT 157.99 25.965 158.2 26.035 ;
    RECT 154.21 25.245 154.42 25.315 ;
    RECT 154.21 25.605 154.42 25.675 ;
    RECT 154.21 25.965 154.42 26.035 ;
    RECT 154.67 25.245 154.88 25.315 ;
    RECT 154.67 25.605 154.88 25.675 ;
    RECT 154.67 25.965 154.88 26.035 ;
    RECT 150.89 25.245 151.1 25.315 ;
    RECT 150.89 25.605 151.1 25.675 ;
    RECT 150.89 25.965 151.1 26.035 ;
    RECT 151.35 25.245 151.56 25.315 ;
    RECT 151.35 25.605 151.56 25.675 ;
    RECT 151.35 25.965 151.56 26.035 ;
    RECT 147.57 25.245 147.78 25.315 ;
    RECT 147.57 25.605 147.78 25.675 ;
    RECT 147.57 25.965 147.78 26.035 ;
    RECT 148.03 25.245 148.24 25.315 ;
    RECT 148.03 25.605 148.24 25.675 ;
    RECT 148.03 25.965 148.24 26.035 ;
    RECT 144.25 25.245 144.46 25.315 ;
    RECT 144.25 25.605 144.46 25.675 ;
    RECT 144.25 25.965 144.46 26.035 ;
    RECT 144.71 25.245 144.92 25.315 ;
    RECT 144.71 25.605 144.92 25.675 ;
    RECT 144.71 25.965 144.92 26.035 ;
    RECT 140.93 25.245 141.14 25.315 ;
    RECT 140.93 25.605 141.14 25.675 ;
    RECT 140.93 25.965 141.14 26.035 ;
    RECT 141.39 25.245 141.6 25.315 ;
    RECT 141.39 25.605 141.6 25.675 ;
    RECT 141.39 25.965 141.6 26.035 ;
    RECT 137.61 25.245 137.82 25.315 ;
    RECT 137.61 25.605 137.82 25.675 ;
    RECT 137.61 25.965 137.82 26.035 ;
    RECT 138.07 25.245 138.28 25.315 ;
    RECT 138.07 25.605 138.28 25.675 ;
    RECT 138.07 25.965 138.28 26.035 ;
    RECT 134.29 25.245 134.5 25.315 ;
    RECT 134.29 25.605 134.5 25.675 ;
    RECT 134.29 25.965 134.5 26.035 ;
    RECT 134.75 25.245 134.96 25.315 ;
    RECT 134.75 25.605 134.96 25.675 ;
    RECT 134.75 25.965 134.96 26.035 ;
    RECT 64.57 25.245 64.78 25.315 ;
    RECT 64.57 25.605 64.78 25.675 ;
    RECT 64.57 25.965 64.78 26.035 ;
    RECT 65.03 25.245 65.24 25.315 ;
    RECT 65.03 25.605 65.24 25.675 ;
    RECT 65.03 25.965 65.24 26.035 ;
    RECT 61.25 24.525 61.46 24.595 ;
    RECT 61.25 24.885 61.46 24.955 ;
    RECT 61.25 25.245 61.46 25.315 ;
    RECT 61.71 24.525 61.92 24.595 ;
    RECT 61.71 24.885 61.92 24.955 ;
    RECT 61.71 25.245 61.92 25.315 ;
    RECT 57.93 24.525 58.14 24.595 ;
    RECT 57.93 24.885 58.14 24.955 ;
    RECT 57.93 25.245 58.14 25.315 ;
    RECT 58.39 24.525 58.6 24.595 ;
    RECT 58.39 24.885 58.6 24.955 ;
    RECT 58.39 25.245 58.6 25.315 ;
    RECT 54.61 24.525 54.82 24.595 ;
    RECT 54.61 24.885 54.82 24.955 ;
    RECT 54.61 25.245 54.82 25.315 ;
    RECT 55.07 24.525 55.28 24.595 ;
    RECT 55.07 24.885 55.28 24.955 ;
    RECT 55.07 25.245 55.28 25.315 ;
    RECT 51.29 24.525 51.5 24.595 ;
    RECT 51.29 24.885 51.5 24.955 ;
    RECT 51.29 25.245 51.5 25.315 ;
    RECT 51.75 24.525 51.96 24.595 ;
    RECT 51.75 24.885 51.96 24.955 ;
    RECT 51.75 25.245 51.96 25.315 ;
    RECT 47.97 24.525 48.18 24.595 ;
    RECT 47.97 24.885 48.18 24.955 ;
    RECT 47.97 25.245 48.18 25.315 ;
    RECT 48.43 24.525 48.64 24.595 ;
    RECT 48.43 24.885 48.64 24.955 ;
    RECT 48.43 25.245 48.64 25.315 ;
    RECT 44.65 24.525 44.86 24.595 ;
    RECT 44.65 24.885 44.86 24.955 ;
    RECT 44.65 25.245 44.86 25.315 ;
    RECT 45.11 24.525 45.32 24.595 ;
    RECT 45.11 24.885 45.32 24.955 ;
    RECT 45.11 25.245 45.32 25.315 ;
    RECT 41.33 24.525 41.54 24.595 ;
    RECT 41.33 24.885 41.54 24.955 ;
    RECT 41.33 25.245 41.54 25.315 ;
    RECT 41.79 24.525 42.0 24.595 ;
    RECT 41.79 24.885 42.0 24.955 ;
    RECT 41.79 25.245 42.0 25.315 ;
    RECT 38.01 24.525 38.22 24.595 ;
    RECT 38.01 24.885 38.22 24.955 ;
    RECT 38.01 25.245 38.22 25.315 ;
    RECT 38.47 24.525 38.68 24.595 ;
    RECT 38.47 24.885 38.68 24.955 ;
    RECT 38.47 25.245 38.68 25.315 ;
    RECT 34.69 24.525 34.9 24.595 ;
    RECT 34.69 24.885 34.9 24.955 ;
    RECT 34.69 25.245 34.9 25.315 ;
    RECT 35.15 24.525 35.36 24.595 ;
    RECT 35.15 24.885 35.36 24.955 ;
    RECT 35.15 25.245 35.36 25.315 ;
    RECT 173.945 24.885 174.015 24.955 ;
    RECT 130.97 24.525 131.18 24.595 ;
    RECT 130.97 24.885 131.18 24.955 ;
    RECT 130.97 25.245 131.18 25.315 ;
    RECT 131.43 24.525 131.64 24.595 ;
    RECT 131.43 24.885 131.64 24.955 ;
    RECT 131.43 25.245 131.64 25.315 ;
    RECT 127.65 24.525 127.86 24.595 ;
    RECT 127.65 24.885 127.86 24.955 ;
    RECT 127.65 25.245 127.86 25.315 ;
    RECT 128.11 24.525 128.32 24.595 ;
    RECT 128.11 24.885 128.32 24.955 ;
    RECT 128.11 25.245 128.32 25.315 ;
    RECT 124.33 24.525 124.54 24.595 ;
    RECT 124.33 24.885 124.54 24.955 ;
    RECT 124.33 25.245 124.54 25.315 ;
    RECT 124.79 24.525 125.0 24.595 ;
    RECT 124.79 24.885 125.0 24.955 ;
    RECT 124.79 25.245 125.0 25.315 ;
    RECT 121.01 24.525 121.22 24.595 ;
    RECT 121.01 24.885 121.22 24.955 ;
    RECT 121.01 25.245 121.22 25.315 ;
    RECT 121.47 24.525 121.68 24.595 ;
    RECT 121.47 24.885 121.68 24.955 ;
    RECT 121.47 25.245 121.68 25.315 ;
    RECT 117.69 24.525 117.9 24.595 ;
    RECT 117.69 24.885 117.9 24.955 ;
    RECT 117.69 25.245 117.9 25.315 ;
    RECT 118.15 24.525 118.36 24.595 ;
    RECT 118.15 24.885 118.36 24.955 ;
    RECT 118.15 25.245 118.36 25.315 ;
    RECT 114.37 24.525 114.58 24.595 ;
    RECT 114.37 24.885 114.58 24.955 ;
    RECT 114.37 25.245 114.58 25.315 ;
    RECT 114.83 24.525 115.04 24.595 ;
    RECT 114.83 24.885 115.04 24.955 ;
    RECT 114.83 25.245 115.04 25.315 ;
    RECT 111.05 24.525 111.26 24.595 ;
    RECT 111.05 24.885 111.26 24.955 ;
    RECT 111.05 25.245 111.26 25.315 ;
    RECT 111.51 24.525 111.72 24.595 ;
    RECT 111.51 24.885 111.72 24.955 ;
    RECT 111.51 25.245 111.72 25.315 ;
    RECT 107.73 24.525 107.94 24.595 ;
    RECT 107.73 24.885 107.94 24.955 ;
    RECT 107.73 25.245 107.94 25.315 ;
    RECT 108.19 24.525 108.4 24.595 ;
    RECT 108.19 24.885 108.4 24.955 ;
    RECT 108.19 25.245 108.4 25.315 ;
    RECT 104.41 24.525 104.62 24.595 ;
    RECT 104.41 24.885 104.62 24.955 ;
    RECT 104.41 25.245 104.62 25.315 ;
    RECT 104.87 24.525 105.08 24.595 ;
    RECT 104.87 24.885 105.08 24.955 ;
    RECT 104.87 25.245 105.08 25.315 ;
    RECT 101.09 24.525 101.3 24.595 ;
    RECT 101.09 24.885 101.3 24.955 ;
    RECT 101.09 25.245 101.3 25.315 ;
    RECT 101.55 24.525 101.76 24.595 ;
    RECT 101.55 24.885 101.76 24.955 ;
    RECT 101.55 25.245 101.76 25.315 ;
    RECT 0.4 24.885 0.47 24.955 ;
    RECT 170.81 24.525 171.02 24.595 ;
    RECT 170.81 24.885 171.02 24.955 ;
    RECT 170.81 25.245 171.02 25.315 ;
    RECT 171.27 24.525 171.48 24.595 ;
    RECT 171.27 24.885 171.48 24.955 ;
    RECT 171.27 25.245 171.48 25.315 ;
    RECT 167.49 24.525 167.7 24.595 ;
    RECT 167.49 24.885 167.7 24.955 ;
    RECT 167.49 25.245 167.7 25.315 ;
    RECT 167.95 24.525 168.16 24.595 ;
    RECT 167.95 24.885 168.16 24.955 ;
    RECT 167.95 25.245 168.16 25.315 ;
    RECT 97.77 24.525 97.98 24.595 ;
    RECT 97.77 24.885 97.98 24.955 ;
    RECT 97.77 25.245 97.98 25.315 ;
    RECT 98.23 24.525 98.44 24.595 ;
    RECT 98.23 24.885 98.44 24.955 ;
    RECT 98.23 25.245 98.44 25.315 ;
    RECT 94.45 24.525 94.66 24.595 ;
    RECT 94.45 24.885 94.66 24.955 ;
    RECT 94.45 25.245 94.66 25.315 ;
    RECT 94.91 24.525 95.12 24.595 ;
    RECT 94.91 24.885 95.12 24.955 ;
    RECT 94.91 25.245 95.12 25.315 ;
    RECT 91.13 24.525 91.34 24.595 ;
    RECT 91.13 24.885 91.34 24.955 ;
    RECT 91.13 25.245 91.34 25.315 ;
    RECT 91.59 24.525 91.8 24.595 ;
    RECT 91.59 24.885 91.8 24.955 ;
    RECT 91.59 25.245 91.8 25.315 ;
    RECT 87.81 24.525 88.02 24.595 ;
    RECT 87.81 24.885 88.02 24.955 ;
    RECT 87.81 25.245 88.02 25.315 ;
    RECT 88.27 24.525 88.48 24.595 ;
    RECT 88.27 24.885 88.48 24.955 ;
    RECT 88.27 25.245 88.48 25.315 ;
    RECT 84.49 24.525 84.7 24.595 ;
    RECT 84.49 24.885 84.7 24.955 ;
    RECT 84.49 25.245 84.7 25.315 ;
    RECT 84.95 24.525 85.16 24.595 ;
    RECT 84.95 24.885 85.16 24.955 ;
    RECT 84.95 25.245 85.16 25.315 ;
    RECT 81.17 24.525 81.38 24.595 ;
    RECT 81.17 24.885 81.38 24.955 ;
    RECT 81.17 25.245 81.38 25.315 ;
    RECT 81.63 24.525 81.84 24.595 ;
    RECT 81.63 24.885 81.84 24.955 ;
    RECT 81.63 25.245 81.84 25.315 ;
    RECT 77.85 24.525 78.06 24.595 ;
    RECT 77.85 24.885 78.06 24.955 ;
    RECT 77.85 25.245 78.06 25.315 ;
    RECT 78.31 24.525 78.52 24.595 ;
    RECT 78.31 24.885 78.52 24.955 ;
    RECT 78.31 25.245 78.52 25.315 ;
    RECT 74.53 24.525 74.74 24.595 ;
    RECT 74.53 24.885 74.74 24.955 ;
    RECT 74.53 25.245 74.74 25.315 ;
    RECT 74.99 24.525 75.2 24.595 ;
    RECT 74.99 24.885 75.2 24.955 ;
    RECT 74.99 25.245 75.2 25.315 ;
    RECT 71.21 24.525 71.42 24.595 ;
    RECT 71.21 24.885 71.42 24.955 ;
    RECT 71.21 25.245 71.42 25.315 ;
    RECT 71.67 24.525 71.88 24.595 ;
    RECT 71.67 24.885 71.88 24.955 ;
    RECT 71.67 25.245 71.88 25.315 ;
    RECT 31.37 24.525 31.58 24.595 ;
    RECT 31.37 24.885 31.58 24.955 ;
    RECT 31.37 25.245 31.58 25.315 ;
    RECT 31.83 24.525 32.04 24.595 ;
    RECT 31.83 24.885 32.04 24.955 ;
    RECT 31.83 25.245 32.04 25.315 ;
    RECT 67.89 24.525 68.1 24.595 ;
    RECT 67.89 24.885 68.1 24.955 ;
    RECT 67.89 25.245 68.1 25.315 ;
    RECT 68.35 24.525 68.56 24.595 ;
    RECT 68.35 24.885 68.56 24.955 ;
    RECT 68.35 25.245 68.56 25.315 ;
    RECT 28.05 24.525 28.26 24.595 ;
    RECT 28.05 24.885 28.26 24.955 ;
    RECT 28.05 25.245 28.26 25.315 ;
    RECT 28.51 24.525 28.72 24.595 ;
    RECT 28.51 24.885 28.72 24.955 ;
    RECT 28.51 25.245 28.72 25.315 ;
    RECT 24.73 24.525 24.94 24.595 ;
    RECT 24.73 24.885 24.94 24.955 ;
    RECT 24.73 25.245 24.94 25.315 ;
    RECT 25.19 24.525 25.4 24.595 ;
    RECT 25.19 24.885 25.4 24.955 ;
    RECT 25.19 25.245 25.4 25.315 ;
    RECT 21.41 24.525 21.62 24.595 ;
    RECT 21.41 24.885 21.62 24.955 ;
    RECT 21.41 25.245 21.62 25.315 ;
    RECT 21.87 24.525 22.08 24.595 ;
    RECT 21.87 24.885 22.08 24.955 ;
    RECT 21.87 25.245 22.08 25.315 ;
    RECT 18.09 24.525 18.3 24.595 ;
    RECT 18.09 24.885 18.3 24.955 ;
    RECT 18.09 25.245 18.3 25.315 ;
    RECT 18.55 24.525 18.76 24.595 ;
    RECT 18.55 24.885 18.76 24.955 ;
    RECT 18.55 25.245 18.76 25.315 ;
    RECT 14.77 24.525 14.98 24.595 ;
    RECT 14.77 24.885 14.98 24.955 ;
    RECT 14.77 25.245 14.98 25.315 ;
    RECT 15.23 24.525 15.44 24.595 ;
    RECT 15.23 24.885 15.44 24.955 ;
    RECT 15.23 25.245 15.44 25.315 ;
    RECT 11.45 24.525 11.66 24.595 ;
    RECT 11.45 24.885 11.66 24.955 ;
    RECT 11.45 25.245 11.66 25.315 ;
    RECT 11.91 24.525 12.12 24.595 ;
    RECT 11.91 24.885 12.12 24.955 ;
    RECT 11.91 25.245 12.12 25.315 ;
    RECT 8.13 24.525 8.34 24.595 ;
    RECT 8.13 24.885 8.34 24.955 ;
    RECT 8.13 25.245 8.34 25.315 ;
    RECT 8.59 24.525 8.8 24.595 ;
    RECT 8.59 24.885 8.8 24.955 ;
    RECT 8.59 25.245 8.8 25.315 ;
    RECT 4.81 24.525 5.02 24.595 ;
    RECT 4.81 24.885 5.02 24.955 ;
    RECT 4.81 25.245 5.02 25.315 ;
    RECT 5.27 24.525 5.48 24.595 ;
    RECT 5.27 24.885 5.48 24.955 ;
    RECT 5.27 25.245 5.48 25.315 ;
    RECT 164.17 24.525 164.38 24.595 ;
    RECT 164.17 24.885 164.38 24.955 ;
    RECT 164.17 25.245 164.38 25.315 ;
    RECT 164.63 24.525 164.84 24.595 ;
    RECT 164.63 24.885 164.84 24.955 ;
    RECT 164.63 25.245 164.84 25.315 ;
    RECT 1.49 24.525 1.7 24.595 ;
    RECT 1.49 24.885 1.7 24.955 ;
    RECT 1.49 25.245 1.7 25.315 ;
    RECT 1.95 24.525 2.16 24.595 ;
    RECT 1.95 24.885 2.16 24.955 ;
    RECT 1.95 25.245 2.16 25.315 ;
    RECT 160.85 24.525 161.06 24.595 ;
    RECT 160.85 24.885 161.06 24.955 ;
    RECT 160.85 25.245 161.06 25.315 ;
    RECT 161.31 24.525 161.52 24.595 ;
    RECT 161.31 24.885 161.52 24.955 ;
    RECT 161.31 25.245 161.52 25.315 ;
    RECT 157.53 24.525 157.74 24.595 ;
    RECT 157.53 24.885 157.74 24.955 ;
    RECT 157.53 25.245 157.74 25.315 ;
    RECT 157.99 24.525 158.2 24.595 ;
    RECT 157.99 24.885 158.2 24.955 ;
    RECT 157.99 25.245 158.2 25.315 ;
    RECT 154.21 24.525 154.42 24.595 ;
    RECT 154.21 24.885 154.42 24.955 ;
    RECT 154.21 25.245 154.42 25.315 ;
    RECT 154.67 24.525 154.88 24.595 ;
    RECT 154.67 24.885 154.88 24.955 ;
    RECT 154.67 25.245 154.88 25.315 ;
    RECT 150.89 24.525 151.1 24.595 ;
    RECT 150.89 24.885 151.1 24.955 ;
    RECT 150.89 25.245 151.1 25.315 ;
    RECT 151.35 24.525 151.56 24.595 ;
    RECT 151.35 24.885 151.56 24.955 ;
    RECT 151.35 25.245 151.56 25.315 ;
    RECT 147.57 24.525 147.78 24.595 ;
    RECT 147.57 24.885 147.78 24.955 ;
    RECT 147.57 25.245 147.78 25.315 ;
    RECT 148.03 24.525 148.24 24.595 ;
    RECT 148.03 24.885 148.24 24.955 ;
    RECT 148.03 25.245 148.24 25.315 ;
    RECT 144.25 24.525 144.46 24.595 ;
    RECT 144.25 24.885 144.46 24.955 ;
    RECT 144.25 25.245 144.46 25.315 ;
    RECT 144.71 24.525 144.92 24.595 ;
    RECT 144.71 24.885 144.92 24.955 ;
    RECT 144.71 25.245 144.92 25.315 ;
    RECT 140.93 24.525 141.14 24.595 ;
    RECT 140.93 24.885 141.14 24.955 ;
    RECT 140.93 25.245 141.14 25.315 ;
    RECT 141.39 24.525 141.6 24.595 ;
    RECT 141.39 24.885 141.6 24.955 ;
    RECT 141.39 25.245 141.6 25.315 ;
    RECT 137.61 24.525 137.82 24.595 ;
    RECT 137.61 24.885 137.82 24.955 ;
    RECT 137.61 25.245 137.82 25.315 ;
    RECT 138.07 24.525 138.28 24.595 ;
    RECT 138.07 24.885 138.28 24.955 ;
    RECT 138.07 25.245 138.28 25.315 ;
    RECT 134.29 24.525 134.5 24.595 ;
    RECT 134.29 24.885 134.5 24.955 ;
    RECT 134.29 25.245 134.5 25.315 ;
    RECT 134.75 24.525 134.96 24.595 ;
    RECT 134.75 24.885 134.96 24.955 ;
    RECT 134.75 25.245 134.96 25.315 ;
    RECT 64.57 24.525 64.78 24.595 ;
    RECT 64.57 24.885 64.78 24.955 ;
    RECT 64.57 25.245 64.78 25.315 ;
    RECT 65.03 24.525 65.24 24.595 ;
    RECT 65.03 24.885 65.24 24.955 ;
    RECT 65.03 25.245 65.24 25.315 ;
    RECT 61.25 23.805 61.46 23.875 ;
    RECT 61.25 24.165 61.46 24.235 ;
    RECT 61.25 24.525 61.46 24.595 ;
    RECT 61.71 23.805 61.92 23.875 ;
    RECT 61.71 24.165 61.92 24.235 ;
    RECT 61.71 24.525 61.92 24.595 ;
    RECT 57.93 23.805 58.14 23.875 ;
    RECT 57.93 24.165 58.14 24.235 ;
    RECT 57.93 24.525 58.14 24.595 ;
    RECT 58.39 23.805 58.6 23.875 ;
    RECT 58.39 24.165 58.6 24.235 ;
    RECT 58.39 24.525 58.6 24.595 ;
    RECT 54.61 23.805 54.82 23.875 ;
    RECT 54.61 24.165 54.82 24.235 ;
    RECT 54.61 24.525 54.82 24.595 ;
    RECT 55.07 23.805 55.28 23.875 ;
    RECT 55.07 24.165 55.28 24.235 ;
    RECT 55.07 24.525 55.28 24.595 ;
    RECT 51.29 23.805 51.5 23.875 ;
    RECT 51.29 24.165 51.5 24.235 ;
    RECT 51.29 24.525 51.5 24.595 ;
    RECT 51.75 23.805 51.96 23.875 ;
    RECT 51.75 24.165 51.96 24.235 ;
    RECT 51.75 24.525 51.96 24.595 ;
    RECT 47.97 23.805 48.18 23.875 ;
    RECT 47.97 24.165 48.18 24.235 ;
    RECT 47.97 24.525 48.18 24.595 ;
    RECT 48.43 23.805 48.64 23.875 ;
    RECT 48.43 24.165 48.64 24.235 ;
    RECT 48.43 24.525 48.64 24.595 ;
    RECT 44.65 23.805 44.86 23.875 ;
    RECT 44.65 24.165 44.86 24.235 ;
    RECT 44.65 24.525 44.86 24.595 ;
    RECT 45.11 23.805 45.32 23.875 ;
    RECT 45.11 24.165 45.32 24.235 ;
    RECT 45.11 24.525 45.32 24.595 ;
    RECT 41.33 23.805 41.54 23.875 ;
    RECT 41.33 24.165 41.54 24.235 ;
    RECT 41.33 24.525 41.54 24.595 ;
    RECT 41.79 23.805 42.0 23.875 ;
    RECT 41.79 24.165 42.0 24.235 ;
    RECT 41.79 24.525 42.0 24.595 ;
    RECT 38.01 23.805 38.22 23.875 ;
    RECT 38.01 24.165 38.22 24.235 ;
    RECT 38.01 24.525 38.22 24.595 ;
    RECT 38.47 23.805 38.68 23.875 ;
    RECT 38.47 24.165 38.68 24.235 ;
    RECT 38.47 24.525 38.68 24.595 ;
    RECT 34.69 23.805 34.9 23.875 ;
    RECT 34.69 24.165 34.9 24.235 ;
    RECT 34.69 24.525 34.9 24.595 ;
    RECT 35.15 23.805 35.36 23.875 ;
    RECT 35.15 24.165 35.36 24.235 ;
    RECT 35.15 24.525 35.36 24.595 ;
    RECT 173.945 24.165 174.015 24.235 ;
    RECT 130.97 23.805 131.18 23.875 ;
    RECT 130.97 24.165 131.18 24.235 ;
    RECT 130.97 24.525 131.18 24.595 ;
    RECT 131.43 23.805 131.64 23.875 ;
    RECT 131.43 24.165 131.64 24.235 ;
    RECT 131.43 24.525 131.64 24.595 ;
    RECT 127.65 23.805 127.86 23.875 ;
    RECT 127.65 24.165 127.86 24.235 ;
    RECT 127.65 24.525 127.86 24.595 ;
    RECT 128.11 23.805 128.32 23.875 ;
    RECT 128.11 24.165 128.32 24.235 ;
    RECT 128.11 24.525 128.32 24.595 ;
    RECT 124.33 23.805 124.54 23.875 ;
    RECT 124.33 24.165 124.54 24.235 ;
    RECT 124.33 24.525 124.54 24.595 ;
    RECT 124.79 23.805 125.0 23.875 ;
    RECT 124.79 24.165 125.0 24.235 ;
    RECT 124.79 24.525 125.0 24.595 ;
    RECT 121.01 23.805 121.22 23.875 ;
    RECT 121.01 24.165 121.22 24.235 ;
    RECT 121.01 24.525 121.22 24.595 ;
    RECT 121.47 23.805 121.68 23.875 ;
    RECT 121.47 24.165 121.68 24.235 ;
    RECT 121.47 24.525 121.68 24.595 ;
    RECT 117.69 23.805 117.9 23.875 ;
    RECT 117.69 24.165 117.9 24.235 ;
    RECT 117.69 24.525 117.9 24.595 ;
    RECT 118.15 23.805 118.36 23.875 ;
    RECT 118.15 24.165 118.36 24.235 ;
    RECT 118.15 24.525 118.36 24.595 ;
    RECT 114.37 23.805 114.58 23.875 ;
    RECT 114.37 24.165 114.58 24.235 ;
    RECT 114.37 24.525 114.58 24.595 ;
    RECT 114.83 23.805 115.04 23.875 ;
    RECT 114.83 24.165 115.04 24.235 ;
    RECT 114.83 24.525 115.04 24.595 ;
    RECT 111.05 23.805 111.26 23.875 ;
    RECT 111.05 24.165 111.26 24.235 ;
    RECT 111.05 24.525 111.26 24.595 ;
    RECT 111.51 23.805 111.72 23.875 ;
    RECT 111.51 24.165 111.72 24.235 ;
    RECT 111.51 24.525 111.72 24.595 ;
    RECT 107.73 23.805 107.94 23.875 ;
    RECT 107.73 24.165 107.94 24.235 ;
    RECT 107.73 24.525 107.94 24.595 ;
    RECT 108.19 23.805 108.4 23.875 ;
    RECT 108.19 24.165 108.4 24.235 ;
    RECT 108.19 24.525 108.4 24.595 ;
    RECT 104.41 23.805 104.62 23.875 ;
    RECT 104.41 24.165 104.62 24.235 ;
    RECT 104.41 24.525 104.62 24.595 ;
    RECT 104.87 23.805 105.08 23.875 ;
    RECT 104.87 24.165 105.08 24.235 ;
    RECT 104.87 24.525 105.08 24.595 ;
    RECT 101.09 23.805 101.3 23.875 ;
    RECT 101.09 24.165 101.3 24.235 ;
    RECT 101.09 24.525 101.3 24.595 ;
    RECT 101.55 23.805 101.76 23.875 ;
    RECT 101.55 24.165 101.76 24.235 ;
    RECT 101.55 24.525 101.76 24.595 ;
    RECT 0.4 24.165 0.47 24.235 ;
    RECT 170.81 23.805 171.02 23.875 ;
    RECT 170.81 24.165 171.02 24.235 ;
    RECT 170.81 24.525 171.02 24.595 ;
    RECT 171.27 23.805 171.48 23.875 ;
    RECT 171.27 24.165 171.48 24.235 ;
    RECT 171.27 24.525 171.48 24.595 ;
    RECT 167.49 23.805 167.7 23.875 ;
    RECT 167.49 24.165 167.7 24.235 ;
    RECT 167.49 24.525 167.7 24.595 ;
    RECT 167.95 23.805 168.16 23.875 ;
    RECT 167.95 24.165 168.16 24.235 ;
    RECT 167.95 24.525 168.16 24.595 ;
    RECT 97.77 23.805 97.98 23.875 ;
    RECT 97.77 24.165 97.98 24.235 ;
    RECT 97.77 24.525 97.98 24.595 ;
    RECT 98.23 23.805 98.44 23.875 ;
    RECT 98.23 24.165 98.44 24.235 ;
    RECT 98.23 24.525 98.44 24.595 ;
    RECT 94.45 23.805 94.66 23.875 ;
    RECT 94.45 24.165 94.66 24.235 ;
    RECT 94.45 24.525 94.66 24.595 ;
    RECT 94.91 23.805 95.12 23.875 ;
    RECT 94.91 24.165 95.12 24.235 ;
    RECT 94.91 24.525 95.12 24.595 ;
    RECT 91.13 23.805 91.34 23.875 ;
    RECT 91.13 24.165 91.34 24.235 ;
    RECT 91.13 24.525 91.34 24.595 ;
    RECT 91.59 23.805 91.8 23.875 ;
    RECT 91.59 24.165 91.8 24.235 ;
    RECT 91.59 24.525 91.8 24.595 ;
    RECT 87.81 23.805 88.02 23.875 ;
    RECT 87.81 24.165 88.02 24.235 ;
    RECT 87.81 24.525 88.02 24.595 ;
    RECT 88.27 23.805 88.48 23.875 ;
    RECT 88.27 24.165 88.48 24.235 ;
    RECT 88.27 24.525 88.48 24.595 ;
    RECT 84.49 23.805 84.7 23.875 ;
    RECT 84.49 24.165 84.7 24.235 ;
    RECT 84.49 24.525 84.7 24.595 ;
    RECT 84.95 23.805 85.16 23.875 ;
    RECT 84.95 24.165 85.16 24.235 ;
    RECT 84.95 24.525 85.16 24.595 ;
    RECT 81.17 23.805 81.38 23.875 ;
    RECT 81.17 24.165 81.38 24.235 ;
    RECT 81.17 24.525 81.38 24.595 ;
    RECT 81.63 23.805 81.84 23.875 ;
    RECT 81.63 24.165 81.84 24.235 ;
    RECT 81.63 24.525 81.84 24.595 ;
    RECT 77.85 23.805 78.06 23.875 ;
    RECT 77.85 24.165 78.06 24.235 ;
    RECT 77.85 24.525 78.06 24.595 ;
    RECT 78.31 23.805 78.52 23.875 ;
    RECT 78.31 24.165 78.52 24.235 ;
    RECT 78.31 24.525 78.52 24.595 ;
    RECT 74.53 23.805 74.74 23.875 ;
    RECT 74.53 24.165 74.74 24.235 ;
    RECT 74.53 24.525 74.74 24.595 ;
    RECT 74.99 23.805 75.2 23.875 ;
    RECT 74.99 24.165 75.2 24.235 ;
    RECT 74.99 24.525 75.2 24.595 ;
    RECT 71.21 23.805 71.42 23.875 ;
    RECT 71.21 24.165 71.42 24.235 ;
    RECT 71.21 24.525 71.42 24.595 ;
    RECT 71.67 23.805 71.88 23.875 ;
    RECT 71.67 24.165 71.88 24.235 ;
    RECT 71.67 24.525 71.88 24.595 ;
    RECT 31.37 23.805 31.58 23.875 ;
    RECT 31.37 24.165 31.58 24.235 ;
    RECT 31.37 24.525 31.58 24.595 ;
    RECT 31.83 23.805 32.04 23.875 ;
    RECT 31.83 24.165 32.04 24.235 ;
    RECT 31.83 24.525 32.04 24.595 ;
    RECT 67.89 23.805 68.1 23.875 ;
    RECT 67.89 24.165 68.1 24.235 ;
    RECT 67.89 24.525 68.1 24.595 ;
    RECT 68.35 23.805 68.56 23.875 ;
    RECT 68.35 24.165 68.56 24.235 ;
    RECT 68.35 24.525 68.56 24.595 ;
    RECT 28.05 23.805 28.26 23.875 ;
    RECT 28.05 24.165 28.26 24.235 ;
    RECT 28.05 24.525 28.26 24.595 ;
    RECT 28.51 23.805 28.72 23.875 ;
    RECT 28.51 24.165 28.72 24.235 ;
    RECT 28.51 24.525 28.72 24.595 ;
    RECT 24.73 23.805 24.94 23.875 ;
    RECT 24.73 24.165 24.94 24.235 ;
    RECT 24.73 24.525 24.94 24.595 ;
    RECT 25.19 23.805 25.4 23.875 ;
    RECT 25.19 24.165 25.4 24.235 ;
    RECT 25.19 24.525 25.4 24.595 ;
    RECT 21.41 23.805 21.62 23.875 ;
    RECT 21.41 24.165 21.62 24.235 ;
    RECT 21.41 24.525 21.62 24.595 ;
    RECT 21.87 23.805 22.08 23.875 ;
    RECT 21.87 24.165 22.08 24.235 ;
    RECT 21.87 24.525 22.08 24.595 ;
    RECT 18.09 23.805 18.3 23.875 ;
    RECT 18.09 24.165 18.3 24.235 ;
    RECT 18.09 24.525 18.3 24.595 ;
    RECT 18.55 23.805 18.76 23.875 ;
    RECT 18.55 24.165 18.76 24.235 ;
    RECT 18.55 24.525 18.76 24.595 ;
    RECT 14.77 23.805 14.98 23.875 ;
    RECT 14.77 24.165 14.98 24.235 ;
    RECT 14.77 24.525 14.98 24.595 ;
    RECT 15.23 23.805 15.44 23.875 ;
    RECT 15.23 24.165 15.44 24.235 ;
    RECT 15.23 24.525 15.44 24.595 ;
    RECT 11.45 23.805 11.66 23.875 ;
    RECT 11.45 24.165 11.66 24.235 ;
    RECT 11.45 24.525 11.66 24.595 ;
    RECT 11.91 23.805 12.12 23.875 ;
    RECT 11.91 24.165 12.12 24.235 ;
    RECT 11.91 24.525 12.12 24.595 ;
    RECT 8.13 23.805 8.34 23.875 ;
    RECT 8.13 24.165 8.34 24.235 ;
    RECT 8.13 24.525 8.34 24.595 ;
    RECT 8.59 23.805 8.8 23.875 ;
    RECT 8.59 24.165 8.8 24.235 ;
    RECT 8.59 24.525 8.8 24.595 ;
    RECT 4.81 23.805 5.02 23.875 ;
    RECT 4.81 24.165 5.02 24.235 ;
    RECT 4.81 24.525 5.02 24.595 ;
    RECT 5.27 23.805 5.48 23.875 ;
    RECT 5.27 24.165 5.48 24.235 ;
    RECT 5.27 24.525 5.48 24.595 ;
    RECT 164.17 23.805 164.38 23.875 ;
    RECT 164.17 24.165 164.38 24.235 ;
    RECT 164.17 24.525 164.38 24.595 ;
    RECT 164.63 23.805 164.84 23.875 ;
    RECT 164.63 24.165 164.84 24.235 ;
    RECT 164.63 24.525 164.84 24.595 ;
    RECT 1.49 23.805 1.7 23.875 ;
    RECT 1.49 24.165 1.7 24.235 ;
    RECT 1.49 24.525 1.7 24.595 ;
    RECT 1.95 23.805 2.16 23.875 ;
    RECT 1.95 24.165 2.16 24.235 ;
    RECT 1.95 24.525 2.16 24.595 ;
    RECT 160.85 23.805 161.06 23.875 ;
    RECT 160.85 24.165 161.06 24.235 ;
    RECT 160.85 24.525 161.06 24.595 ;
    RECT 161.31 23.805 161.52 23.875 ;
    RECT 161.31 24.165 161.52 24.235 ;
    RECT 161.31 24.525 161.52 24.595 ;
    RECT 157.53 23.805 157.74 23.875 ;
    RECT 157.53 24.165 157.74 24.235 ;
    RECT 157.53 24.525 157.74 24.595 ;
    RECT 157.99 23.805 158.2 23.875 ;
    RECT 157.99 24.165 158.2 24.235 ;
    RECT 157.99 24.525 158.2 24.595 ;
    RECT 154.21 23.805 154.42 23.875 ;
    RECT 154.21 24.165 154.42 24.235 ;
    RECT 154.21 24.525 154.42 24.595 ;
    RECT 154.67 23.805 154.88 23.875 ;
    RECT 154.67 24.165 154.88 24.235 ;
    RECT 154.67 24.525 154.88 24.595 ;
    RECT 150.89 23.805 151.1 23.875 ;
    RECT 150.89 24.165 151.1 24.235 ;
    RECT 150.89 24.525 151.1 24.595 ;
    RECT 151.35 23.805 151.56 23.875 ;
    RECT 151.35 24.165 151.56 24.235 ;
    RECT 151.35 24.525 151.56 24.595 ;
    RECT 147.57 23.805 147.78 23.875 ;
    RECT 147.57 24.165 147.78 24.235 ;
    RECT 147.57 24.525 147.78 24.595 ;
    RECT 148.03 23.805 148.24 23.875 ;
    RECT 148.03 24.165 148.24 24.235 ;
    RECT 148.03 24.525 148.24 24.595 ;
    RECT 144.25 23.805 144.46 23.875 ;
    RECT 144.25 24.165 144.46 24.235 ;
    RECT 144.25 24.525 144.46 24.595 ;
    RECT 144.71 23.805 144.92 23.875 ;
    RECT 144.71 24.165 144.92 24.235 ;
    RECT 144.71 24.525 144.92 24.595 ;
    RECT 140.93 23.805 141.14 23.875 ;
    RECT 140.93 24.165 141.14 24.235 ;
    RECT 140.93 24.525 141.14 24.595 ;
    RECT 141.39 23.805 141.6 23.875 ;
    RECT 141.39 24.165 141.6 24.235 ;
    RECT 141.39 24.525 141.6 24.595 ;
    RECT 137.61 23.805 137.82 23.875 ;
    RECT 137.61 24.165 137.82 24.235 ;
    RECT 137.61 24.525 137.82 24.595 ;
    RECT 138.07 23.805 138.28 23.875 ;
    RECT 138.07 24.165 138.28 24.235 ;
    RECT 138.07 24.525 138.28 24.595 ;
    RECT 134.29 23.805 134.5 23.875 ;
    RECT 134.29 24.165 134.5 24.235 ;
    RECT 134.29 24.525 134.5 24.595 ;
    RECT 134.75 23.805 134.96 23.875 ;
    RECT 134.75 24.165 134.96 24.235 ;
    RECT 134.75 24.525 134.96 24.595 ;
    RECT 64.57 23.805 64.78 23.875 ;
    RECT 64.57 24.165 64.78 24.235 ;
    RECT 64.57 24.525 64.78 24.595 ;
    RECT 65.03 23.805 65.24 23.875 ;
    RECT 65.03 24.165 65.24 24.235 ;
    RECT 65.03 24.525 65.24 24.595 ;
    RECT 61.25 23.085 61.46 23.155 ;
    RECT 61.25 23.445 61.46 23.515 ;
    RECT 61.25 23.805 61.46 23.875 ;
    RECT 61.71 23.085 61.92 23.155 ;
    RECT 61.71 23.445 61.92 23.515 ;
    RECT 61.71 23.805 61.92 23.875 ;
    RECT 57.93 23.085 58.14 23.155 ;
    RECT 57.93 23.445 58.14 23.515 ;
    RECT 57.93 23.805 58.14 23.875 ;
    RECT 58.39 23.085 58.6 23.155 ;
    RECT 58.39 23.445 58.6 23.515 ;
    RECT 58.39 23.805 58.6 23.875 ;
    RECT 54.61 23.085 54.82 23.155 ;
    RECT 54.61 23.445 54.82 23.515 ;
    RECT 54.61 23.805 54.82 23.875 ;
    RECT 55.07 23.085 55.28 23.155 ;
    RECT 55.07 23.445 55.28 23.515 ;
    RECT 55.07 23.805 55.28 23.875 ;
    RECT 51.29 23.085 51.5 23.155 ;
    RECT 51.29 23.445 51.5 23.515 ;
    RECT 51.29 23.805 51.5 23.875 ;
    RECT 51.75 23.085 51.96 23.155 ;
    RECT 51.75 23.445 51.96 23.515 ;
    RECT 51.75 23.805 51.96 23.875 ;
    RECT 47.97 23.085 48.18 23.155 ;
    RECT 47.97 23.445 48.18 23.515 ;
    RECT 47.97 23.805 48.18 23.875 ;
    RECT 48.43 23.085 48.64 23.155 ;
    RECT 48.43 23.445 48.64 23.515 ;
    RECT 48.43 23.805 48.64 23.875 ;
    RECT 44.65 23.085 44.86 23.155 ;
    RECT 44.65 23.445 44.86 23.515 ;
    RECT 44.65 23.805 44.86 23.875 ;
    RECT 45.11 23.085 45.32 23.155 ;
    RECT 45.11 23.445 45.32 23.515 ;
    RECT 45.11 23.805 45.32 23.875 ;
    RECT 41.33 23.085 41.54 23.155 ;
    RECT 41.33 23.445 41.54 23.515 ;
    RECT 41.33 23.805 41.54 23.875 ;
    RECT 41.79 23.085 42.0 23.155 ;
    RECT 41.79 23.445 42.0 23.515 ;
    RECT 41.79 23.805 42.0 23.875 ;
    RECT 38.01 23.085 38.22 23.155 ;
    RECT 38.01 23.445 38.22 23.515 ;
    RECT 38.01 23.805 38.22 23.875 ;
    RECT 38.47 23.085 38.68 23.155 ;
    RECT 38.47 23.445 38.68 23.515 ;
    RECT 38.47 23.805 38.68 23.875 ;
    RECT 34.69 23.085 34.9 23.155 ;
    RECT 34.69 23.445 34.9 23.515 ;
    RECT 34.69 23.805 34.9 23.875 ;
    RECT 35.15 23.085 35.36 23.155 ;
    RECT 35.15 23.445 35.36 23.515 ;
    RECT 35.15 23.805 35.36 23.875 ;
    RECT 173.945 23.445 174.015 23.515 ;
    RECT 130.97 23.085 131.18 23.155 ;
    RECT 130.97 23.445 131.18 23.515 ;
    RECT 130.97 23.805 131.18 23.875 ;
    RECT 131.43 23.085 131.64 23.155 ;
    RECT 131.43 23.445 131.64 23.515 ;
    RECT 131.43 23.805 131.64 23.875 ;
    RECT 127.65 23.085 127.86 23.155 ;
    RECT 127.65 23.445 127.86 23.515 ;
    RECT 127.65 23.805 127.86 23.875 ;
    RECT 128.11 23.085 128.32 23.155 ;
    RECT 128.11 23.445 128.32 23.515 ;
    RECT 128.11 23.805 128.32 23.875 ;
    RECT 124.33 23.085 124.54 23.155 ;
    RECT 124.33 23.445 124.54 23.515 ;
    RECT 124.33 23.805 124.54 23.875 ;
    RECT 124.79 23.085 125.0 23.155 ;
    RECT 124.79 23.445 125.0 23.515 ;
    RECT 124.79 23.805 125.0 23.875 ;
    RECT 121.01 23.085 121.22 23.155 ;
    RECT 121.01 23.445 121.22 23.515 ;
    RECT 121.01 23.805 121.22 23.875 ;
    RECT 121.47 23.085 121.68 23.155 ;
    RECT 121.47 23.445 121.68 23.515 ;
    RECT 121.47 23.805 121.68 23.875 ;
    RECT 117.69 23.085 117.9 23.155 ;
    RECT 117.69 23.445 117.9 23.515 ;
    RECT 117.69 23.805 117.9 23.875 ;
    RECT 118.15 23.085 118.36 23.155 ;
    RECT 118.15 23.445 118.36 23.515 ;
    RECT 118.15 23.805 118.36 23.875 ;
    RECT 114.37 23.085 114.58 23.155 ;
    RECT 114.37 23.445 114.58 23.515 ;
    RECT 114.37 23.805 114.58 23.875 ;
    RECT 114.83 23.085 115.04 23.155 ;
    RECT 114.83 23.445 115.04 23.515 ;
    RECT 114.83 23.805 115.04 23.875 ;
    RECT 111.05 23.085 111.26 23.155 ;
    RECT 111.05 23.445 111.26 23.515 ;
    RECT 111.05 23.805 111.26 23.875 ;
    RECT 111.51 23.085 111.72 23.155 ;
    RECT 111.51 23.445 111.72 23.515 ;
    RECT 111.51 23.805 111.72 23.875 ;
    RECT 107.73 23.085 107.94 23.155 ;
    RECT 107.73 23.445 107.94 23.515 ;
    RECT 107.73 23.805 107.94 23.875 ;
    RECT 108.19 23.085 108.4 23.155 ;
    RECT 108.19 23.445 108.4 23.515 ;
    RECT 108.19 23.805 108.4 23.875 ;
    RECT 104.41 23.085 104.62 23.155 ;
    RECT 104.41 23.445 104.62 23.515 ;
    RECT 104.41 23.805 104.62 23.875 ;
    RECT 104.87 23.085 105.08 23.155 ;
    RECT 104.87 23.445 105.08 23.515 ;
    RECT 104.87 23.805 105.08 23.875 ;
    RECT 101.09 23.085 101.3 23.155 ;
    RECT 101.09 23.445 101.3 23.515 ;
    RECT 101.09 23.805 101.3 23.875 ;
    RECT 101.55 23.085 101.76 23.155 ;
    RECT 101.55 23.445 101.76 23.515 ;
    RECT 101.55 23.805 101.76 23.875 ;
    RECT 0.4 23.445 0.47 23.515 ;
    RECT 170.81 23.085 171.02 23.155 ;
    RECT 170.81 23.445 171.02 23.515 ;
    RECT 170.81 23.805 171.02 23.875 ;
    RECT 171.27 23.085 171.48 23.155 ;
    RECT 171.27 23.445 171.48 23.515 ;
    RECT 171.27 23.805 171.48 23.875 ;
    RECT 167.49 23.085 167.7 23.155 ;
    RECT 167.49 23.445 167.7 23.515 ;
    RECT 167.49 23.805 167.7 23.875 ;
    RECT 167.95 23.085 168.16 23.155 ;
    RECT 167.95 23.445 168.16 23.515 ;
    RECT 167.95 23.805 168.16 23.875 ;
    RECT 97.77 23.085 97.98 23.155 ;
    RECT 97.77 23.445 97.98 23.515 ;
    RECT 97.77 23.805 97.98 23.875 ;
    RECT 98.23 23.085 98.44 23.155 ;
    RECT 98.23 23.445 98.44 23.515 ;
    RECT 98.23 23.805 98.44 23.875 ;
    RECT 94.45 23.085 94.66 23.155 ;
    RECT 94.45 23.445 94.66 23.515 ;
    RECT 94.45 23.805 94.66 23.875 ;
    RECT 94.91 23.085 95.12 23.155 ;
    RECT 94.91 23.445 95.12 23.515 ;
    RECT 94.91 23.805 95.12 23.875 ;
    RECT 91.13 23.085 91.34 23.155 ;
    RECT 91.13 23.445 91.34 23.515 ;
    RECT 91.13 23.805 91.34 23.875 ;
    RECT 91.59 23.085 91.8 23.155 ;
    RECT 91.59 23.445 91.8 23.515 ;
    RECT 91.59 23.805 91.8 23.875 ;
    RECT 87.81 23.085 88.02 23.155 ;
    RECT 87.81 23.445 88.02 23.515 ;
    RECT 87.81 23.805 88.02 23.875 ;
    RECT 88.27 23.085 88.48 23.155 ;
    RECT 88.27 23.445 88.48 23.515 ;
    RECT 88.27 23.805 88.48 23.875 ;
    RECT 84.49 23.085 84.7 23.155 ;
    RECT 84.49 23.445 84.7 23.515 ;
    RECT 84.49 23.805 84.7 23.875 ;
    RECT 84.95 23.085 85.16 23.155 ;
    RECT 84.95 23.445 85.16 23.515 ;
    RECT 84.95 23.805 85.16 23.875 ;
    RECT 81.17 23.085 81.38 23.155 ;
    RECT 81.17 23.445 81.38 23.515 ;
    RECT 81.17 23.805 81.38 23.875 ;
    RECT 81.63 23.085 81.84 23.155 ;
    RECT 81.63 23.445 81.84 23.515 ;
    RECT 81.63 23.805 81.84 23.875 ;
    RECT 77.85 23.085 78.06 23.155 ;
    RECT 77.85 23.445 78.06 23.515 ;
    RECT 77.85 23.805 78.06 23.875 ;
    RECT 78.31 23.085 78.52 23.155 ;
    RECT 78.31 23.445 78.52 23.515 ;
    RECT 78.31 23.805 78.52 23.875 ;
    RECT 74.53 23.085 74.74 23.155 ;
    RECT 74.53 23.445 74.74 23.515 ;
    RECT 74.53 23.805 74.74 23.875 ;
    RECT 74.99 23.085 75.2 23.155 ;
    RECT 74.99 23.445 75.2 23.515 ;
    RECT 74.99 23.805 75.2 23.875 ;
    RECT 71.21 23.085 71.42 23.155 ;
    RECT 71.21 23.445 71.42 23.515 ;
    RECT 71.21 23.805 71.42 23.875 ;
    RECT 71.67 23.085 71.88 23.155 ;
    RECT 71.67 23.445 71.88 23.515 ;
    RECT 71.67 23.805 71.88 23.875 ;
    RECT 31.37 23.085 31.58 23.155 ;
    RECT 31.37 23.445 31.58 23.515 ;
    RECT 31.37 23.805 31.58 23.875 ;
    RECT 31.83 23.085 32.04 23.155 ;
    RECT 31.83 23.445 32.04 23.515 ;
    RECT 31.83 23.805 32.04 23.875 ;
    RECT 67.89 23.085 68.1 23.155 ;
    RECT 67.89 23.445 68.1 23.515 ;
    RECT 67.89 23.805 68.1 23.875 ;
    RECT 68.35 23.085 68.56 23.155 ;
    RECT 68.35 23.445 68.56 23.515 ;
    RECT 68.35 23.805 68.56 23.875 ;
    RECT 28.05 23.085 28.26 23.155 ;
    RECT 28.05 23.445 28.26 23.515 ;
    RECT 28.05 23.805 28.26 23.875 ;
    RECT 28.51 23.085 28.72 23.155 ;
    RECT 28.51 23.445 28.72 23.515 ;
    RECT 28.51 23.805 28.72 23.875 ;
    RECT 24.73 23.085 24.94 23.155 ;
    RECT 24.73 23.445 24.94 23.515 ;
    RECT 24.73 23.805 24.94 23.875 ;
    RECT 25.19 23.085 25.4 23.155 ;
    RECT 25.19 23.445 25.4 23.515 ;
    RECT 25.19 23.805 25.4 23.875 ;
    RECT 21.41 23.085 21.62 23.155 ;
    RECT 21.41 23.445 21.62 23.515 ;
    RECT 21.41 23.805 21.62 23.875 ;
    RECT 21.87 23.085 22.08 23.155 ;
    RECT 21.87 23.445 22.08 23.515 ;
    RECT 21.87 23.805 22.08 23.875 ;
    RECT 18.09 23.085 18.3 23.155 ;
    RECT 18.09 23.445 18.3 23.515 ;
    RECT 18.09 23.805 18.3 23.875 ;
    RECT 18.55 23.085 18.76 23.155 ;
    RECT 18.55 23.445 18.76 23.515 ;
    RECT 18.55 23.805 18.76 23.875 ;
    RECT 14.77 23.085 14.98 23.155 ;
    RECT 14.77 23.445 14.98 23.515 ;
    RECT 14.77 23.805 14.98 23.875 ;
    RECT 15.23 23.085 15.44 23.155 ;
    RECT 15.23 23.445 15.44 23.515 ;
    RECT 15.23 23.805 15.44 23.875 ;
    RECT 11.45 23.085 11.66 23.155 ;
    RECT 11.45 23.445 11.66 23.515 ;
    RECT 11.45 23.805 11.66 23.875 ;
    RECT 11.91 23.085 12.12 23.155 ;
    RECT 11.91 23.445 12.12 23.515 ;
    RECT 11.91 23.805 12.12 23.875 ;
    RECT 8.13 23.085 8.34 23.155 ;
    RECT 8.13 23.445 8.34 23.515 ;
    RECT 8.13 23.805 8.34 23.875 ;
    RECT 8.59 23.085 8.8 23.155 ;
    RECT 8.59 23.445 8.8 23.515 ;
    RECT 8.59 23.805 8.8 23.875 ;
    RECT 4.81 23.085 5.02 23.155 ;
    RECT 4.81 23.445 5.02 23.515 ;
    RECT 4.81 23.805 5.02 23.875 ;
    RECT 5.27 23.085 5.48 23.155 ;
    RECT 5.27 23.445 5.48 23.515 ;
    RECT 5.27 23.805 5.48 23.875 ;
    RECT 164.17 23.085 164.38 23.155 ;
    RECT 164.17 23.445 164.38 23.515 ;
    RECT 164.17 23.805 164.38 23.875 ;
    RECT 164.63 23.085 164.84 23.155 ;
    RECT 164.63 23.445 164.84 23.515 ;
    RECT 164.63 23.805 164.84 23.875 ;
    RECT 1.49 23.085 1.7 23.155 ;
    RECT 1.49 23.445 1.7 23.515 ;
    RECT 1.49 23.805 1.7 23.875 ;
    RECT 1.95 23.085 2.16 23.155 ;
    RECT 1.95 23.445 2.16 23.515 ;
    RECT 1.95 23.805 2.16 23.875 ;
    RECT 160.85 23.085 161.06 23.155 ;
    RECT 160.85 23.445 161.06 23.515 ;
    RECT 160.85 23.805 161.06 23.875 ;
    RECT 161.31 23.085 161.52 23.155 ;
    RECT 161.31 23.445 161.52 23.515 ;
    RECT 161.31 23.805 161.52 23.875 ;
    RECT 157.53 23.085 157.74 23.155 ;
    RECT 157.53 23.445 157.74 23.515 ;
    RECT 157.53 23.805 157.74 23.875 ;
    RECT 157.99 23.085 158.2 23.155 ;
    RECT 157.99 23.445 158.2 23.515 ;
    RECT 157.99 23.805 158.2 23.875 ;
    RECT 154.21 23.085 154.42 23.155 ;
    RECT 154.21 23.445 154.42 23.515 ;
    RECT 154.21 23.805 154.42 23.875 ;
    RECT 154.67 23.085 154.88 23.155 ;
    RECT 154.67 23.445 154.88 23.515 ;
    RECT 154.67 23.805 154.88 23.875 ;
    RECT 150.89 23.085 151.1 23.155 ;
    RECT 150.89 23.445 151.1 23.515 ;
    RECT 150.89 23.805 151.1 23.875 ;
    RECT 151.35 23.085 151.56 23.155 ;
    RECT 151.35 23.445 151.56 23.515 ;
    RECT 151.35 23.805 151.56 23.875 ;
    RECT 147.57 23.085 147.78 23.155 ;
    RECT 147.57 23.445 147.78 23.515 ;
    RECT 147.57 23.805 147.78 23.875 ;
    RECT 148.03 23.085 148.24 23.155 ;
    RECT 148.03 23.445 148.24 23.515 ;
    RECT 148.03 23.805 148.24 23.875 ;
    RECT 144.25 23.085 144.46 23.155 ;
    RECT 144.25 23.445 144.46 23.515 ;
    RECT 144.25 23.805 144.46 23.875 ;
    RECT 144.71 23.085 144.92 23.155 ;
    RECT 144.71 23.445 144.92 23.515 ;
    RECT 144.71 23.805 144.92 23.875 ;
    RECT 140.93 23.085 141.14 23.155 ;
    RECT 140.93 23.445 141.14 23.515 ;
    RECT 140.93 23.805 141.14 23.875 ;
    RECT 141.39 23.085 141.6 23.155 ;
    RECT 141.39 23.445 141.6 23.515 ;
    RECT 141.39 23.805 141.6 23.875 ;
    RECT 137.61 23.085 137.82 23.155 ;
    RECT 137.61 23.445 137.82 23.515 ;
    RECT 137.61 23.805 137.82 23.875 ;
    RECT 138.07 23.085 138.28 23.155 ;
    RECT 138.07 23.445 138.28 23.515 ;
    RECT 138.07 23.805 138.28 23.875 ;
    RECT 134.29 23.085 134.5 23.155 ;
    RECT 134.29 23.445 134.5 23.515 ;
    RECT 134.29 23.805 134.5 23.875 ;
    RECT 134.75 23.085 134.96 23.155 ;
    RECT 134.75 23.445 134.96 23.515 ;
    RECT 134.75 23.805 134.96 23.875 ;
    RECT 64.57 23.085 64.78 23.155 ;
    RECT 64.57 23.445 64.78 23.515 ;
    RECT 64.57 23.805 64.78 23.875 ;
    RECT 65.03 23.085 65.24 23.155 ;
    RECT 65.03 23.445 65.24 23.515 ;
    RECT 65.03 23.805 65.24 23.875 ;
    RECT 61.25 22.365 61.46 22.435 ;
    RECT 61.25 22.725 61.46 22.795 ;
    RECT 61.25 23.085 61.46 23.155 ;
    RECT 61.71 22.365 61.92 22.435 ;
    RECT 61.71 22.725 61.92 22.795 ;
    RECT 61.71 23.085 61.92 23.155 ;
    RECT 57.93 22.365 58.14 22.435 ;
    RECT 57.93 22.725 58.14 22.795 ;
    RECT 57.93 23.085 58.14 23.155 ;
    RECT 58.39 22.365 58.6 22.435 ;
    RECT 58.39 22.725 58.6 22.795 ;
    RECT 58.39 23.085 58.6 23.155 ;
    RECT 54.61 22.365 54.82 22.435 ;
    RECT 54.61 22.725 54.82 22.795 ;
    RECT 54.61 23.085 54.82 23.155 ;
    RECT 55.07 22.365 55.28 22.435 ;
    RECT 55.07 22.725 55.28 22.795 ;
    RECT 55.07 23.085 55.28 23.155 ;
    RECT 51.29 22.365 51.5 22.435 ;
    RECT 51.29 22.725 51.5 22.795 ;
    RECT 51.29 23.085 51.5 23.155 ;
    RECT 51.75 22.365 51.96 22.435 ;
    RECT 51.75 22.725 51.96 22.795 ;
    RECT 51.75 23.085 51.96 23.155 ;
    RECT 47.97 22.365 48.18 22.435 ;
    RECT 47.97 22.725 48.18 22.795 ;
    RECT 47.97 23.085 48.18 23.155 ;
    RECT 48.43 22.365 48.64 22.435 ;
    RECT 48.43 22.725 48.64 22.795 ;
    RECT 48.43 23.085 48.64 23.155 ;
    RECT 44.65 22.365 44.86 22.435 ;
    RECT 44.65 22.725 44.86 22.795 ;
    RECT 44.65 23.085 44.86 23.155 ;
    RECT 45.11 22.365 45.32 22.435 ;
    RECT 45.11 22.725 45.32 22.795 ;
    RECT 45.11 23.085 45.32 23.155 ;
    RECT 41.33 22.365 41.54 22.435 ;
    RECT 41.33 22.725 41.54 22.795 ;
    RECT 41.33 23.085 41.54 23.155 ;
    RECT 41.79 22.365 42.0 22.435 ;
    RECT 41.79 22.725 42.0 22.795 ;
    RECT 41.79 23.085 42.0 23.155 ;
    RECT 38.01 22.365 38.22 22.435 ;
    RECT 38.01 22.725 38.22 22.795 ;
    RECT 38.01 23.085 38.22 23.155 ;
    RECT 38.47 22.365 38.68 22.435 ;
    RECT 38.47 22.725 38.68 22.795 ;
    RECT 38.47 23.085 38.68 23.155 ;
    RECT 34.69 22.365 34.9 22.435 ;
    RECT 34.69 22.725 34.9 22.795 ;
    RECT 34.69 23.085 34.9 23.155 ;
    RECT 35.15 22.365 35.36 22.435 ;
    RECT 35.15 22.725 35.36 22.795 ;
    RECT 35.15 23.085 35.36 23.155 ;
    RECT 173.945 22.725 174.015 22.795 ;
    RECT 130.97 22.365 131.18 22.435 ;
    RECT 130.97 22.725 131.18 22.795 ;
    RECT 130.97 23.085 131.18 23.155 ;
    RECT 131.43 22.365 131.64 22.435 ;
    RECT 131.43 22.725 131.64 22.795 ;
    RECT 131.43 23.085 131.64 23.155 ;
    RECT 127.65 22.365 127.86 22.435 ;
    RECT 127.65 22.725 127.86 22.795 ;
    RECT 127.65 23.085 127.86 23.155 ;
    RECT 128.11 22.365 128.32 22.435 ;
    RECT 128.11 22.725 128.32 22.795 ;
    RECT 128.11 23.085 128.32 23.155 ;
    RECT 124.33 22.365 124.54 22.435 ;
    RECT 124.33 22.725 124.54 22.795 ;
    RECT 124.33 23.085 124.54 23.155 ;
    RECT 124.79 22.365 125.0 22.435 ;
    RECT 124.79 22.725 125.0 22.795 ;
    RECT 124.79 23.085 125.0 23.155 ;
    RECT 121.01 22.365 121.22 22.435 ;
    RECT 121.01 22.725 121.22 22.795 ;
    RECT 121.01 23.085 121.22 23.155 ;
    RECT 121.47 22.365 121.68 22.435 ;
    RECT 121.47 22.725 121.68 22.795 ;
    RECT 121.47 23.085 121.68 23.155 ;
    RECT 117.69 22.365 117.9 22.435 ;
    RECT 117.69 22.725 117.9 22.795 ;
    RECT 117.69 23.085 117.9 23.155 ;
    RECT 118.15 22.365 118.36 22.435 ;
    RECT 118.15 22.725 118.36 22.795 ;
    RECT 118.15 23.085 118.36 23.155 ;
    RECT 114.37 22.365 114.58 22.435 ;
    RECT 114.37 22.725 114.58 22.795 ;
    RECT 114.37 23.085 114.58 23.155 ;
    RECT 114.83 22.365 115.04 22.435 ;
    RECT 114.83 22.725 115.04 22.795 ;
    RECT 114.83 23.085 115.04 23.155 ;
    RECT 111.05 22.365 111.26 22.435 ;
    RECT 111.05 22.725 111.26 22.795 ;
    RECT 111.05 23.085 111.26 23.155 ;
    RECT 111.51 22.365 111.72 22.435 ;
    RECT 111.51 22.725 111.72 22.795 ;
    RECT 111.51 23.085 111.72 23.155 ;
    RECT 107.73 22.365 107.94 22.435 ;
    RECT 107.73 22.725 107.94 22.795 ;
    RECT 107.73 23.085 107.94 23.155 ;
    RECT 108.19 22.365 108.4 22.435 ;
    RECT 108.19 22.725 108.4 22.795 ;
    RECT 108.19 23.085 108.4 23.155 ;
    RECT 104.41 22.365 104.62 22.435 ;
    RECT 104.41 22.725 104.62 22.795 ;
    RECT 104.41 23.085 104.62 23.155 ;
    RECT 104.87 22.365 105.08 22.435 ;
    RECT 104.87 22.725 105.08 22.795 ;
    RECT 104.87 23.085 105.08 23.155 ;
    RECT 101.09 22.365 101.3 22.435 ;
    RECT 101.09 22.725 101.3 22.795 ;
    RECT 101.09 23.085 101.3 23.155 ;
    RECT 101.55 22.365 101.76 22.435 ;
    RECT 101.55 22.725 101.76 22.795 ;
    RECT 101.55 23.085 101.76 23.155 ;
    RECT 0.4 22.725 0.47 22.795 ;
    RECT 170.81 22.365 171.02 22.435 ;
    RECT 170.81 22.725 171.02 22.795 ;
    RECT 170.81 23.085 171.02 23.155 ;
    RECT 171.27 22.365 171.48 22.435 ;
    RECT 171.27 22.725 171.48 22.795 ;
    RECT 171.27 23.085 171.48 23.155 ;
    RECT 167.49 22.365 167.7 22.435 ;
    RECT 167.49 22.725 167.7 22.795 ;
    RECT 167.49 23.085 167.7 23.155 ;
    RECT 167.95 22.365 168.16 22.435 ;
    RECT 167.95 22.725 168.16 22.795 ;
    RECT 167.95 23.085 168.16 23.155 ;
    RECT 97.77 22.365 97.98 22.435 ;
    RECT 97.77 22.725 97.98 22.795 ;
    RECT 97.77 23.085 97.98 23.155 ;
    RECT 98.23 22.365 98.44 22.435 ;
    RECT 98.23 22.725 98.44 22.795 ;
    RECT 98.23 23.085 98.44 23.155 ;
    RECT 94.45 22.365 94.66 22.435 ;
    RECT 94.45 22.725 94.66 22.795 ;
    RECT 94.45 23.085 94.66 23.155 ;
    RECT 94.91 22.365 95.12 22.435 ;
    RECT 94.91 22.725 95.12 22.795 ;
    RECT 94.91 23.085 95.12 23.155 ;
    RECT 91.13 22.365 91.34 22.435 ;
    RECT 91.13 22.725 91.34 22.795 ;
    RECT 91.13 23.085 91.34 23.155 ;
    RECT 91.59 22.365 91.8 22.435 ;
    RECT 91.59 22.725 91.8 22.795 ;
    RECT 91.59 23.085 91.8 23.155 ;
    RECT 87.81 22.365 88.02 22.435 ;
    RECT 87.81 22.725 88.02 22.795 ;
    RECT 87.81 23.085 88.02 23.155 ;
    RECT 88.27 22.365 88.48 22.435 ;
    RECT 88.27 22.725 88.48 22.795 ;
    RECT 88.27 23.085 88.48 23.155 ;
    RECT 84.49 22.365 84.7 22.435 ;
    RECT 84.49 22.725 84.7 22.795 ;
    RECT 84.49 23.085 84.7 23.155 ;
    RECT 84.95 22.365 85.16 22.435 ;
    RECT 84.95 22.725 85.16 22.795 ;
    RECT 84.95 23.085 85.16 23.155 ;
    RECT 81.17 22.365 81.38 22.435 ;
    RECT 81.17 22.725 81.38 22.795 ;
    RECT 81.17 23.085 81.38 23.155 ;
    RECT 81.63 22.365 81.84 22.435 ;
    RECT 81.63 22.725 81.84 22.795 ;
    RECT 81.63 23.085 81.84 23.155 ;
    RECT 77.85 22.365 78.06 22.435 ;
    RECT 77.85 22.725 78.06 22.795 ;
    RECT 77.85 23.085 78.06 23.155 ;
    RECT 78.31 22.365 78.52 22.435 ;
    RECT 78.31 22.725 78.52 22.795 ;
    RECT 78.31 23.085 78.52 23.155 ;
    RECT 74.53 22.365 74.74 22.435 ;
    RECT 74.53 22.725 74.74 22.795 ;
    RECT 74.53 23.085 74.74 23.155 ;
    RECT 74.99 22.365 75.2 22.435 ;
    RECT 74.99 22.725 75.2 22.795 ;
    RECT 74.99 23.085 75.2 23.155 ;
    RECT 71.21 22.365 71.42 22.435 ;
    RECT 71.21 22.725 71.42 22.795 ;
    RECT 71.21 23.085 71.42 23.155 ;
    RECT 71.67 22.365 71.88 22.435 ;
    RECT 71.67 22.725 71.88 22.795 ;
    RECT 71.67 23.085 71.88 23.155 ;
    RECT 31.37 22.365 31.58 22.435 ;
    RECT 31.37 22.725 31.58 22.795 ;
    RECT 31.37 23.085 31.58 23.155 ;
    RECT 31.83 22.365 32.04 22.435 ;
    RECT 31.83 22.725 32.04 22.795 ;
    RECT 31.83 23.085 32.04 23.155 ;
    RECT 67.89 22.365 68.1 22.435 ;
    RECT 67.89 22.725 68.1 22.795 ;
    RECT 67.89 23.085 68.1 23.155 ;
    RECT 68.35 22.365 68.56 22.435 ;
    RECT 68.35 22.725 68.56 22.795 ;
    RECT 68.35 23.085 68.56 23.155 ;
    RECT 28.05 22.365 28.26 22.435 ;
    RECT 28.05 22.725 28.26 22.795 ;
    RECT 28.05 23.085 28.26 23.155 ;
    RECT 28.51 22.365 28.72 22.435 ;
    RECT 28.51 22.725 28.72 22.795 ;
    RECT 28.51 23.085 28.72 23.155 ;
    RECT 24.73 22.365 24.94 22.435 ;
    RECT 24.73 22.725 24.94 22.795 ;
    RECT 24.73 23.085 24.94 23.155 ;
    RECT 25.19 22.365 25.4 22.435 ;
    RECT 25.19 22.725 25.4 22.795 ;
    RECT 25.19 23.085 25.4 23.155 ;
    RECT 21.41 22.365 21.62 22.435 ;
    RECT 21.41 22.725 21.62 22.795 ;
    RECT 21.41 23.085 21.62 23.155 ;
    RECT 21.87 22.365 22.08 22.435 ;
    RECT 21.87 22.725 22.08 22.795 ;
    RECT 21.87 23.085 22.08 23.155 ;
    RECT 18.09 22.365 18.3 22.435 ;
    RECT 18.09 22.725 18.3 22.795 ;
    RECT 18.09 23.085 18.3 23.155 ;
    RECT 18.55 22.365 18.76 22.435 ;
    RECT 18.55 22.725 18.76 22.795 ;
    RECT 18.55 23.085 18.76 23.155 ;
    RECT 14.77 22.365 14.98 22.435 ;
    RECT 14.77 22.725 14.98 22.795 ;
    RECT 14.77 23.085 14.98 23.155 ;
    RECT 15.23 22.365 15.44 22.435 ;
    RECT 15.23 22.725 15.44 22.795 ;
    RECT 15.23 23.085 15.44 23.155 ;
    RECT 11.45 22.365 11.66 22.435 ;
    RECT 11.45 22.725 11.66 22.795 ;
    RECT 11.45 23.085 11.66 23.155 ;
    RECT 11.91 22.365 12.12 22.435 ;
    RECT 11.91 22.725 12.12 22.795 ;
    RECT 11.91 23.085 12.12 23.155 ;
    RECT 8.13 22.365 8.34 22.435 ;
    RECT 8.13 22.725 8.34 22.795 ;
    RECT 8.13 23.085 8.34 23.155 ;
    RECT 8.59 22.365 8.8 22.435 ;
    RECT 8.59 22.725 8.8 22.795 ;
    RECT 8.59 23.085 8.8 23.155 ;
    RECT 4.81 22.365 5.02 22.435 ;
    RECT 4.81 22.725 5.02 22.795 ;
    RECT 4.81 23.085 5.02 23.155 ;
    RECT 5.27 22.365 5.48 22.435 ;
    RECT 5.27 22.725 5.48 22.795 ;
    RECT 5.27 23.085 5.48 23.155 ;
    RECT 164.17 22.365 164.38 22.435 ;
    RECT 164.17 22.725 164.38 22.795 ;
    RECT 164.17 23.085 164.38 23.155 ;
    RECT 164.63 22.365 164.84 22.435 ;
    RECT 164.63 22.725 164.84 22.795 ;
    RECT 164.63 23.085 164.84 23.155 ;
    RECT 1.49 22.365 1.7 22.435 ;
    RECT 1.49 22.725 1.7 22.795 ;
    RECT 1.49 23.085 1.7 23.155 ;
    RECT 1.95 22.365 2.16 22.435 ;
    RECT 1.95 22.725 2.16 22.795 ;
    RECT 1.95 23.085 2.16 23.155 ;
    RECT 160.85 22.365 161.06 22.435 ;
    RECT 160.85 22.725 161.06 22.795 ;
    RECT 160.85 23.085 161.06 23.155 ;
    RECT 161.31 22.365 161.52 22.435 ;
    RECT 161.31 22.725 161.52 22.795 ;
    RECT 161.31 23.085 161.52 23.155 ;
    RECT 157.53 22.365 157.74 22.435 ;
    RECT 157.53 22.725 157.74 22.795 ;
    RECT 157.53 23.085 157.74 23.155 ;
    RECT 157.99 22.365 158.2 22.435 ;
    RECT 157.99 22.725 158.2 22.795 ;
    RECT 157.99 23.085 158.2 23.155 ;
    RECT 154.21 22.365 154.42 22.435 ;
    RECT 154.21 22.725 154.42 22.795 ;
    RECT 154.21 23.085 154.42 23.155 ;
    RECT 154.67 22.365 154.88 22.435 ;
    RECT 154.67 22.725 154.88 22.795 ;
    RECT 154.67 23.085 154.88 23.155 ;
    RECT 150.89 22.365 151.1 22.435 ;
    RECT 150.89 22.725 151.1 22.795 ;
    RECT 150.89 23.085 151.1 23.155 ;
    RECT 151.35 22.365 151.56 22.435 ;
    RECT 151.35 22.725 151.56 22.795 ;
    RECT 151.35 23.085 151.56 23.155 ;
    RECT 147.57 22.365 147.78 22.435 ;
    RECT 147.57 22.725 147.78 22.795 ;
    RECT 147.57 23.085 147.78 23.155 ;
    RECT 148.03 22.365 148.24 22.435 ;
    RECT 148.03 22.725 148.24 22.795 ;
    RECT 148.03 23.085 148.24 23.155 ;
    RECT 144.25 22.365 144.46 22.435 ;
    RECT 144.25 22.725 144.46 22.795 ;
    RECT 144.25 23.085 144.46 23.155 ;
    RECT 144.71 22.365 144.92 22.435 ;
    RECT 144.71 22.725 144.92 22.795 ;
    RECT 144.71 23.085 144.92 23.155 ;
    RECT 140.93 22.365 141.14 22.435 ;
    RECT 140.93 22.725 141.14 22.795 ;
    RECT 140.93 23.085 141.14 23.155 ;
    RECT 141.39 22.365 141.6 22.435 ;
    RECT 141.39 22.725 141.6 22.795 ;
    RECT 141.39 23.085 141.6 23.155 ;
    RECT 137.61 22.365 137.82 22.435 ;
    RECT 137.61 22.725 137.82 22.795 ;
    RECT 137.61 23.085 137.82 23.155 ;
    RECT 138.07 22.365 138.28 22.435 ;
    RECT 138.07 22.725 138.28 22.795 ;
    RECT 138.07 23.085 138.28 23.155 ;
    RECT 134.29 22.365 134.5 22.435 ;
    RECT 134.29 22.725 134.5 22.795 ;
    RECT 134.29 23.085 134.5 23.155 ;
    RECT 134.75 22.365 134.96 22.435 ;
    RECT 134.75 22.725 134.96 22.795 ;
    RECT 134.75 23.085 134.96 23.155 ;
    RECT 64.57 22.365 64.78 22.435 ;
    RECT 64.57 22.725 64.78 22.795 ;
    RECT 64.57 23.085 64.78 23.155 ;
    RECT 65.03 22.365 65.24 22.435 ;
    RECT 65.03 22.725 65.24 22.795 ;
    RECT 65.03 23.085 65.24 23.155 ;
    RECT 61.25 35.325 61.46 35.395 ;
    RECT 61.25 35.685 61.46 35.755 ;
    RECT 61.25 36.045 61.46 36.115 ;
    RECT 61.71 35.325 61.92 35.395 ;
    RECT 61.71 35.685 61.92 35.755 ;
    RECT 61.71 36.045 61.92 36.115 ;
    RECT 57.93 35.325 58.14 35.395 ;
    RECT 57.93 35.685 58.14 35.755 ;
    RECT 57.93 36.045 58.14 36.115 ;
    RECT 58.39 35.325 58.6 35.395 ;
    RECT 58.39 35.685 58.6 35.755 ;
    RECT 58.39 36.045 58.6 36.115 ;
    RECT 54.61 35.325 54.82 35.395 ;
    RECT 54.61 35.685 54.82 35.755 ;
    RECT 54.61 36.045 54.82 36.115 ;
    RECT 55.07 35.325 55.28 35.395 ;
    RECT 55.07 35.685 55.28 35.755 ;
    RECT 55.07 36.045 55.28 36.115 ;
    RECT 51.29 35.325 51.5 35.395 ;
    RECT 51.29 35.685 51.5 35.755 ;
    RECT 51.29 36.045 51.5 36.115 ;
    RECT 51.75 35.325 51.96 35.395 ;
    RECT 51.75 35.685 51.96 35.755 ;
    RECT 51.75 36.045 51.96 36.115 ;
    RECT 47.97 35.325 48.18 35.395 ;
    RECT 47.97 35.685 48.18 35.755 ;
    RECT 47.97 36.045 48.18 36.115 ;
    RECT 48.43 35.325 48.64 35.395 ;
    RECT 48.43 35.685 48.64 35.755 ;
    RECT 48.43 36.045 48.64 36.115 ;
    RECT 44.65 35.325 44.86 35.395 ;
    RECT 44.65 35.685 44.86 35.755 ;
    RECT 44.65 36.045 44.86 36.115 ;
    RECT 45.11 35.325 45.32 35.395 ;
    RECT 45.11 35.685 45.32 35.755 ;
    RECT 45.11 36.045 45.32 36.115 ;
    RECT 41.33 35.325 41.54 35.395 ;
    RECT 41.33 35.685 41.54 35.755 ;
    RECT 41.33 36.045 41.54 36.115 ;
    RECT 41.79 35.325 42.0 35.395 ;
    RECT 41.79 35.685 42.0 35.755 ;
    RECT 41.79 36.045 42.0 36.115 ;
    RECT 38.01 35.325 38.22 35.395 ;
    RECT 38.01 35.685 38.22 35.755 ;
    RECT 38.01 36.045 38.22 36.115 ;
    RECT 38.47 35.325 38.68 35.395 ;
    RECT 38.47 35.685 38.68 35.755 ;
    RECT 38.47 36.045 38.68 36.115 ;
    RECT 34.69 35.325 34.9 35.395 ;
    RECT 34.69 35.685 34.9 35.755 ;
    RECT 34.69 36.045 34.9 36.115 ;
    RECT 35.15 35.325 35.36 35.395 ;
    RECT 35.15 35.685 35.36 35.755 ;
    RECT 35.15 36.045 35.36 36.115 ;
    RECT 130.97 35.325 131.18 35.395 ;
    RECT 130.97 35.685 131.18 35.755 ;
    RECT 130.97 36.045 131.18 36.115 ;
    RECT 131.43 35.325 131.64 35.395 ;
    RECT 131.43 35.685 131.64 35.755 ;
    RECT 131.43 36.045 131.64 36.115 ;
    RECT 127.65 35.325 127.86 35.395 ;
    RECT 127.65 35.685 127.86 35.755 ;
    RECT 127.65 36.045 127.86 36.115 ;
    RECT 128.11 35.325 128.32 35.395 ;
    RECT 128.11 35.685 128.32 35.755 ;
    RECT 128.11 36.045 128.32 36.115 ;
    RECT 124.33 35.325 124.54 35.395 ;
    RECT 124.33 35.685 124.54 35.755 ;
    RECT 124.33 36.045 124.54 36.115 ;
    RECT 124.79 35.325 125.0 35.395 ;
    RECT 124.79 35.685 125.0 35.755 ;
    RECT 124.79 36.045 125.0 36.115 ;
    RECT 121.01 35.325 121.22 35.395 ;
    RECT 121.01 35.685 121.22 35.755 ;
    RECT 121.01 36.045 121.22 36.115 ;
    RECT 121.47 35.325 121.68 35.395 ;
    RECT 121.47 35.685 121.68 35.755 ;
    RECT 121.47 36.045 121.68 36.115 ;
    RECT 117.69 35.325 117.9 35.395 ;
    RECT 117.69 35.685 117.9 35.755 ;
    RECT 117.69 36.045 117.9 36.115 ;
    RECT 118.15 35.325 118.36 35.395 ;
    RECT 118.15 35.685 118.36 35.755 ;
    RECT 118.15 36.045 118.36 36.115 ;
    RECT 114.37 35.325 114.58 35.395 ;
    RECT 114.37 35.685 114.58 35.755 ;
    RECT 114.37 36.045 114.58 36.115 ;
    RECT 114.83 35.325 115.04 35.395 ;
    RECT 114.83 35.685 115.04 35.755 ;
    RECT 114.83 36.045 115.04 36.115 ;
    RECT 111.05 35.325 111.26 35.395 ;
    RECT 111.05 35.685 111.26 35.755 ;
    RECT 111.05 36.045 111.26 36.115 ;
    RECT 111.51 35.325 111.72 35.395 ;
    RECT 111.51 35.685 111.72 35.755 ;
    RECT 111.51 36.045 111.72 36.115 ;
    RECT 107.73 35.325 107.94 35.395 ;
    RECT 107.73 35.685 107.94 35.755 ;
    RECT 107.73 36.045 107.94 36.115 ;
    RECT 108.19 35.325 108.4 35.395 ;
    RECT 108.19 35.685 108.4 35.755 ;
    RECT 108.19 36.045 108.4 36.115 ;
    RECT 104.41 35.325 104.62 35.395 ;
    RECT 104.41 35.685 104.62 35.755 ;
    RECT 104.41 36.045 104.62 36.115 ;
    RECT 104.87 35.325 105.08 35.395 ;
    RECT 104.87 35.685 105.08 35.755 ;
    RECT 104.87 36.045 105.08 36.115 ;
    RECT 101.09 35.325 101.3 35.395 ;
    RECT 101.09 35.685 101.3 35.755 ;
    RECT 101.09 36.045 101.3 36.115 ;
    RECT 101.55 35.325 101.76 35.395 ;
    RECT 101.55 35.685 101.76 35.755 ;
    RECT 101.55 36.045 101.76 36.115 ;
    RECT 0.4 35.685 0.47 35.755 ;
    RECT 170.81 35.325 171.02 35.395 ;
    RECT 170.81 35.685 171.02 35.755 ;
    RECT 170.81 36.045 171.02 36.115 ;
    RECT 171.27 35.325 171.48 35.395 ;
    RECT 171.27 35.685 171.48 35.755 ;
    RECT 171.27 36.045 171.48 36.115 ;
    RECT 167.49 35.325 167.7 35.395 ;
    RECT 167.49 35.685 167.7 35.755 ;
    RECT 167.49 36.045 167.7 36.115 ;
    RECT 167.95 35.325 168.16 35.395 ;
    RECT 167.95 35.685 168.16 35.755 ;
    RECT 167.95 36.045 168.16 36.115 ;
    RECT 97.77 35.325 97.98 35.395 ;
    RECT 97.77 35.685 97.98 35.755 ;
    RECT 97.77 36.045 97.98 36.115 ;
    RECT 98.23 35.325 98.44 35.395 ;
    RECT 98.23 35.685 98.44 35.755 ;
    RECT 98.23 36.045 98.44 36.115 ;
    RECT 94.45 35.325 94.66 35.395 ;
    RECT 94.45 35.685 94.66 35.755 ;
    RECT 94.45 36.045 94.66 36.115 ;
    RECT 94.91 35.325 95.12 35.395 ;
    RECT 94.91 35.685 95.12 35.755 ;
    RECT 94.91 36.045 95.12 36.115 ;
    RECT 91.13 35.325 91.34 35.395 ;
    RECT 91.13 35.685 91.34 35.755 ;
    RECT 91.13 36.045 91.34 36.115 ;
    RECT 91.59 35.325 91.8 35.395 ;
    RECT 91.59 35.685 91.8 35.755 ;
    RECT 91.59 36.045 91.8 36.115 ;
    RECT 87.81 35.325 88.02 35.395 ;
    RECT 87.81 35.685 88.02 35.755 ;
    RECT 87.81 36.045 88.02 36.115 ;
    RECT 88.27 35.325 88.48 35.395 ;
    RECT 88.27 35.685 88.48 35.755 ;
    RECT 88.27 36.045 88.48 36.115 ;
    RECT 84.49 35.325 84.7 35.395 ;
    RECT 84.49 35.685 84.7 35.755 ;
    RECT 84.49 36.045 84.7 36.115 ;
    RECT 84.95 35.325 85.16 35.395 ;
    RECT 84.95 35.685 85.16 35.755 ;
    RECT 84.95 36.045 85.16 36.115 ;
    RECT 81.17 35.325 81.38 35.395 ;
    RECT 81.17 35.685 81.38 35.755 ;
    RECT 81.17 36.045 81.38 36.115 ;
    RECT 81.63 35.325 81.84 35.395 ;
    RECT 81.63 35.685 81.84 35.755 ;
    RECT 81.63 36.045 81.84 36.115 ;
    RECT 77.85 35.325 78.06 35.395 ;
    RECT 77.85 35.685 78.06 35.755 ;
    RECT 77.85 36.045 78.06 36.115 ;
    RECT 78.31 35.325 78.52 35.395 ;
    RECT 78.31 35.685 78.52 35.755 ;
    RECT 78.31 36.045 78.52 36.115 ;
    RECT 74.53 35.325 74.74 35.395 ;
    RECT 74.53 35.685 74.74 35.755 ;
    RECT 74.53 36.045 74.74 36.115 ;
    RECT 74.99 35.325 75.2 35.395 ;
    RECT 74.99 35.685 75.2 35.755 ;
    RECT 74.99 36.045 75.2 36.115 ;
    RECT 71.21 35.325 71.42 35.395 ;
    RECT 71.21 35.685 71.42 35.755 ;
    RECT 71.21 36.045 71.42 36.115 ;
    RECT 71.67 35.325 71.88 35.395 ;
    RECT 71.67 35.685 71.88 35.755 ;
    RECT 71.67 36.045 71.88 36.115 ;
    RECT 31.37 35.325 31.58 35.395 ;
    RECT 31.37 35.685 31.58 35.755 ;
    RECT 31.37 36.045 31.58 36.115 ;
    RECT 31.83 35.325 32.04 35.395 ;
    RECT 31.83 35.685 32.04 35.755 ;
    RECT 31.83 36.045 32.04 36.115 ;
    RECT 67.89 35.325 68.1 35.395 ;
    RECT 67.89 35.685 68.1 35.755 ;
    RECT 67.89 36.045 68.1 36.115 ;
    RECT 68.35 35.325 68.56 35.395 ;
    RECT 68.35 35.685 68.56 35.755 ;
    RECT 68.35 36.045 68.56 36.115 ;
    RECT 28.05 35.325 28.26 35.395 ;
    RECT 28.05 35.685 28.26 35.755 ;
    RECT 28.05 36.045 28.26 36.115 ;
    RECT 28.51 35.325 28.72 35.395 ;
    RECT 28.51 35.685 28.72 35.755 ;
    RECT 28.51 36.045 28.72 36.115 ;
    RECT 24.73 35.325 24.94 35.395 ;
    RECT 24.73 35.685 24.94 35.755 ;
    RECT 24.73 36.045 24.94 36.115 ;
    RECT 25.19 35.325 25.4 35.395 ;
    RECT 25.19 35.685 25.4 35.755 ;
    RECT 25.19 36.045 25.4 36.115 ;
    RECT 21.41 35.325 21.62 35.395 ;
    RECT 21.41 35.685 21.62 35.755 ;
    RECT 21.41 36.045 21.62 36.115 ;
    RECT 21.87 35.325 22.08 35.395 ;
    RECT 21.87 35.685 22.08 35.755 ;
    RECT 21.87 36.045 22.08 36.115 ;
    RECT 18.09 35.325 18.3 35.395 ;
    RECT 18.09 35.685 18.3 35.755 ;
    RECT 18.09 36.045 18.3 36.115 ;
    RECT 18.55 35.325 18.76 35.395 ;
    RECT 18.55 35.685 18.76 35.755 ;
    RECT 18.55 36.045 18.76 36.115 ;
    RECT 14.77 35.325 14.98 35.395 ;
    RECT 14.77 35.685 14.98 35.755 ;
    RECT 14.77 36.045 14.98 36.115 ;
    RECT 15.23 35.325 15.44 35.395 ;
    RECT 15.23 35.685 15.44 35.755 ;
    RECT 15.23 36.045 15.44 36.115 ;
    RECT 11.45 35.325 11.66 35.395 ;
    RECT 11.45 35.685 11.66 35.755 ;
    RECT 11.45 36.045 11.66 36.115 ;
    RECT 11.91 35.325 12.12 35.395 ;
    RECT 11.91 35.685 12.12 35.755 ;
    RECT 11.91 36.045 12.12 36.115 ;
    RECT 173.945 35.685 174.015 35.755 ;
    RECT 8.13 35.325 8.34 35.395 ;
    RECT 8.13 35.685 8.34 35.755 ;
    RECT 8.13 36.045 8.34 36.115 ;
    RECT 8.59 35.325 8.8 35.395 ;
    RECT 8.59 35.685 8.8 35.755 ;
    RECT 8.59 36.045 8.8 36.115 ;
    RECT 4.81 35.325 5.02 35.395 ;
    RECT 4.81 35.685 5.02 35.755 ;
    RECT 4.81 36.045 5.02 36.115 ;
    RECT 5.27 35.325 5.48 35.395 ;
    RECT 5.27 35.685 5.48 35.755 ;
    RECT 5.27 36.045 5.48 36.115 ;
    RECT 164.17 35.325 164.38 35.395 ;
    RECT 164.17 35.685 164.38 35.755 ;
    RECT 164.17 36.045 164.38 36.115 ;
    RECT 164.63 35.325 164.84 35.395 ;
    RECT 164.63 35.685 164.84 35.755 ;
    RECT 164.63 36.045 164.84 36.115 ;
    RECT 1.49 35.325 1.7 35.395 ;
    RECT 1.49 35.685 1.7 35.755 ;
    RECT 1.49 36.045 1.7 36.115 ;
    RECT 1.95 35.325 2.16 35.395 ;
    RECT 1.95 35.685 2.16 35.755 ;
    RECT 1.95 36.045 2.16 36.115 ;
    RECT 160.85 35.325 161.06 35.395 ;
    RECT 160.85 35.685 161.06 35.755 ;
    RECT 160.85 36.045 161.06 36.115 ;
    RECT 161.31 35.325 161.52 35.395 ;
    RECT 161.31 35.685 161.52 35.755 ;
    RECT 161.31 36.045 161.52 36.115 ;
    RECT 157.53 35.325 157.74 35.395 ;
    RECT 157.53 35.685 157.74 35.755 ;
    RECT 157.53 36.045 157.74 36.115 ;
    RECT 157.99 35.325 158.2 35.395 ;
    RECT 157.99 35.685 158.2 35.755 ;
    RECT 157.99 36.045 158.2 36.115 ;
    RECT 154.21 35.325 154.42 35.395 ;
    RECT 154.21 35.685 154.42 35.755 ;
    RECT 154.21 36.045 154.42 36.115 ;
    RECT 154.67 35.325 154.88 35.395 ;
    RECT 154.67 35.685 154.88 35.755 ;
    RECT 154.67 36.045 154.88 36.115 ;
    RECT 150.89 35.325 151.1 35.395 ;
    RECT 150.89 35.685 151.1 35.755 ;
    RECT 150.89 36.045 151.1 36.115 ;
    RECT 151.35 35.325 151.56 35.395 ;
    RECT 151.35 35.685 151.56 35.755 ;
    RECT 151.35 36.045 151.56 36.115 ;
    RECT 147.57 35.325 147.78 35.395 ;
    RECT 147.57 35.685 147.78 35.755 ;
    RECT 147.57 36.045 147.78 36.115 ;
    RECT 148.03 35.325 148.24 35.395 ;
    RECT 148.03 35.685 148.24 35.755 ;
    RECT 148.03 36.045 148.24 36.115 ;
    RECT 144.25 35.325 144.46 35.395 ;
    RECT 144.25 35.685 144.46 35.755 ;
    RECT 144.25 36.045 144.46 36.115 ;
    RECT 144.71 35.325 144.92 35.395 ;
    RECT 144.71 35.685 144.92 35.755 ;
    RECT 144.71 36.045 144.92 36.115 ;
    RECT 140.93 35.325 141.14 35.395 ;
    RECT 140.93 35.685 141.14 35.755 ;
    RECT 140.93 36.045 141.14 36.115 ;
    RECT 141.39 35.325 141.6 35.395 ;
    RECT 141.39 35.685 141.6 35.755 ;
    RECT 141.39 36.045 141.6 36.115 ;
    RECT 137.61 35.325 137.82 35.395 ;
    RECT 137.61 35.685 137.82 35.755 ;
    RECT 137.61 36.045 137.82 36.115 ;
    RECT 138.07 35.325 138.28 35.395 ;
    RECT 138.07 35.685 138.28 35.755 ;
    RECT 138.07 36.045 138.28 36.115 ;
    RECT 134.29 35.325 134.5 35.395 ;
    RECT 134.29 35.685 134.5 35.755 ;
    RECT 134.29 36.045 134.5 36.115 ;
    RECT 134.75 35.325 134.96 35.395 ;
    RECT 134.75 35.685 134.96 35.755 ;
    RECT 134.75 36.045 134.96 36.115 ;
    RECT 64.57 35.325 64.78 35.395 ;
    RECT 64.57 35.685 64.78 35.755 ;
    RECT 64.57 36.045 64.78 36.115 ;
    RECT 65.03 35.325 65.24 35.395 ;
    RECT 65.03 35.685 65.24 35.755 ;
    RECT 65.03 36.045 65.24 36.115 ;
    RECT 61.25 21.645 61.46 21.715 ;
    RECT 61.25 22.005 61.46 22.075 ;
    RECT 61.25 22.365 61.46 22.435 ;
    RECT 61.71 21.645 61.92 21.715 ;
    RECT 61.71 22.005 61.92 22.075 ;
    RECT 61.71 22.365 61.92 22.435 ;
    RECT 57.93 21.645 58.14 21.715 ;
    RECT 57.93 22.005 58.14 22.075 ;
    RECT 57.93 22.365 58.14 22.435 ;
    RECT 58.39 21.645 58.6 21.715 ;
    RECT 58.39 22.005 58.6 22.075 ;
    RECT 58.39 22.365 58.6 22.435 ;
    RECT 54.61 21.645 54.82 21.715 ;
    RECT 54.61 22.005 54.82 22.075 ;
    RECT 54.61 22.365 54.82 22.435 ;
    RECT 55.07 21.645 55.28 21.715 ;
    RECT 55.07 22.005 55.28 22.075 ;
    RECT 55.07 22.365 55.28 22.435 ;
    RECT 51.29 21.645 51.5 21.715 ;
    RECT 51.29 22.005 51.5 22.075 ;
    RECT 51.29 22.365 51.5 22.435 ;
    RECT 51.75 21.645 51.96 21.715 ;
    RECT 51.75 22.005 51.96 22.075 ;
    RECT 51.75 22.365 51.96 22.435 ;
    RECT 47.97 21.645 48.18 21.715 ;
    RECT 47.97 22.005 48.18 22.075 ;
    RECT 47.97 22.365 48.18 22.435 ;
    RECT 48.43 21.645 48.64 21.715 ;
    RECT 48.43 22.005 48.64 22.075 ;
    RECT 48.43 22.365 48.64 22.435 ;
    RECT 44.65 21.645 44.86 21.715 ;
    RECT 44.65 22.005 44.86 22.075 ;
    RECT 44.65 22.365 44.86 22.435 ;
    RECT 45.11 21.645 45.32 21.715 ;
    RECT 45.11 22.005 45.32 22.075 ;
    RECT 45.11 22.365 45.32 22.435 ;
    RECT 41.33 21.645 41.54 21.715 ;
    RECT 41.33 22.005 41.54 22.075 ;
    RECT 41.33 22.365 41.54 22.435 ;
    RECT 41.79 21.645 42.0 21.715 ;
    RECT 41.79 22.005 42.0 22.075 ;
    RECT 41.79 22.365 42.0 22.435 ;
    RECT 38.01 21.645 38.22 21.715 ;
    RECT 38.01 22.005 38.22 22.075 ;
    RECT 38.01 22.365 38.22 22.435 ;
    RECT 38.47 21.645 38.68 21.715 ;
    RECT 38.47 22.005 38.68 22.075 ;
    RECT 38.47 22.365 38.68 22.435 ;
    RECT 34.69 21.645 34.9 21.715 ;
    RECT 34.69 22.005 34.9 22.075 ;
    RECT 34.69 22.365 34.9 22.435 ;
    RECT 35.15 21.645 35.36 21.715 ;
    RECT 35.15 22.005 35.36 22.075 ;
    RECT 35.15 22.365 35.36 22.435 ;
    RECT 173.945 22.005 174.015 22.075 ;
    RECT 130.97 21.645 131.18 21.715 ;
    RECT 130.97 22.005 131.18 22.075 ;
    RECT 130.97 22.365 131.18 22.435 ;
    RECT 131.43 21.645 131.64 21.715 ;
    RECT 131.43 22.005 131.64 22.075 ;
    RECT 131.43 22.365 131.64 22.435 ;
    RECT 127.65 21.645 127.86 21.715 ;
    RECT 127.65 22.005 127.86 22.075 ;
    RECT 127.65 22.365 127.86 22.435 ;
    RECT 128.11 21.645 128.32 21.715 ;
    RECT 128.11 22.005 128.32 22.075 ;
    RECT 128.11 22.365 128.32 22.435 ;
    RECT 124.33 21.645 124.54 21.715 ;
    RECT 124.33 22.005 124.54 22.075 ;
    RECT 124.33 22.365 124.54 22.435 ;
    RECT 124.79 21.645 125.0 21.715 ;
    RECT 124.79 22.005 125.0 22.075 ;
    RECT 124.79 22.365 125.0 22.435 ;
    RECT 121.01 21.645 121.22 21.715 ;
    RECT 121.01 22.005 121.22 22.075 ;
    RECT 121.01 22.365 121.22 22.435 ;
    RECT 121.47 21.645 121.68 21.715 ;
    RECT 121.47 22.005 121.68 22.075 ;
    RECT 121.47 22.365 121.68 22.435 ;
    RECT 117.69 21.645 117.9 21.715 ;
    RECT 117.69 22.005 117.9 22.075 ;
    RECT 117.69 22.365 117.9 22.435 ;
    RECT 118.15 21.645 118.36 21.715 ;
    RECT 118.15 22.005 118.36 22.075 ;
    RECT 118.15 22.365 118.36 22.435 ;
    RECT 114.37 21.645 114.58 21.715 ;
    RECT 114.37 22.005 114.58 22.075 ;
    RECT 114.37 22.365 114.58 22.435 ;
    RECT 114.83 21.645 115.04 21.715 ;
    RECT 114.83 22.005 115.04 22.075 ;
    RECT 114.83 22.365 115.04 22.435 ;
    RECT 111.05 21.645 111.26 21.715 ;
    RECT 111.05 22.005 111.26 22.075 ;
    RECT 111.05 22.365 111.26 22.435 ;
    RECT 111.51 21.645 111.72 21.715 ;
    RECT 111.51 22.005 111.72 22.075 ;
    RECT 111.51 22.365 111.72 22.435 ;
    RECT 107.73 21.645 107.94 21.715 ;
    RECT 107.73 22.005 107.94 22.075 ;
    RECT 107.73 22.365 107.94 22.435 ;
    RECT 108.19 21.645 108.4 21.715 ;
    RECT 108.19 22.005 108.4 22.075 ;
    RECT 108.19 22.365 108.4 22.435 ;
    RECT 104.41 21.645 104.62 21.715 ;
    RECT 104.41 22.005 104.62 22.075 ;
    RECT 104.41 22.365 104.62 22.435 ;
    RECT 104.87 21.645 105.08 21.715 ;
    RECT 104.87 22.005 105.08 22.075 ;
    RECT 104.87 22.365 105.08 22.435 ;
    RECT 101.09 21.645 101.3 21.715 ;
    RECT 101.09 22.005 101.3 22.075 ;
    RECT 101.09 22.365 101.3 22.435 ;
    RECT 101.55 21.645 101.76 21.715 ;
    RECT 101.55 22.005 101.76 22.075 ;
    RECT 101.55 22.365 101.76 22.435 ;
    RECT 0.4 22.005 0.47 22.075 ;
    RECT 170.81 21.645 171.02 21.715 ;
    RECT 170.81 22.005 171.02 22.075 ;
    RECT 170.81 22.365 171.02 22.435 ;
    RECT 171.27 21.645 171.48 21.715 ;
    RECT 171.27 22.005 171.48 22.075 ;
    RECT 171.27 22.365 171.48 22.435 ;
    RECT 167.49 21.645 167.7 21.715 ;
    RECT 167.49 22.005 167.7 22.075 ;
    RECT 167.49 22.365 167.7 22.435 ;
    RECT 167.95 21.645 168.16 21.715 ;
    RECT 167.95 22.005 168.16 22.075 ;
    RECT 167.95 22.365 168.16 22.435 ;
    RECT 97.77 21.645 97.98 21.715 ;
    RECT 97.77 22.005 97.98 22.075 ;
    RECT 97.77 22.365 97.98 22.435 ;
    RECT 98.23 21.645 98.44 21.715 ;
    RECT 98.23 22.005 98.44 22.075 ;
    RECT 98.23 22.365 98.44 22.435 ;
    RECT 94.45 21.645 94.66 21.715 ;
    RECT 94.45 22.005 94.66 22.075 ;
    RECT 94.45 22.365 94.66 22.435 ;
    RECT 94.91 21.645 95.12 21.715 ;
    RECT 94.91 22.005 95.12 22.075 ;
    RECT 94.91 22.365 95.12 22.435 ;
    RECT 91.13 21.645 91.34 21.715 ;
    RECT 91.13 22.005 91.34 22.075 ;
    RECT 91.13 22.365 91.34 22.435 ;
    RECT 91.59 21.645 91.8 21.715 ;
    RECT 91.59 22.005 91.8 22.075 ;
    RECT 91.59 22.365 91.8 22.435 ;
    RECT 87.81 21.645 88.02 21.715 ;
    RECT 87.81 22.005 88.02 22.075 ;
    RECT 87.81 22.365 88.02 22.435 ;
    RECT 88.27 21.645 88.48 21.715 ;
    RECT 88.27 22.005 88.48 22.075 ;
    RECT 88.27 22.365 88.48 22.435 ;
    RECT 84.49 21.645 84.7 21.715 ;
    RECT 84.49 22.005 84.7 22.075 ;
    RECT 84.49 22.365 84.7 22.435 ;
    RECT 84.95 21.645 85.16 21.715 ;
    RECT 84.95 22.005 85.16 22.075 ;
    RECT 84.95 22.365 85.16 22.435 ;
    RECT 81.17 21.645 81.38 21.715 ;
    RECT 81.17 22.005 81.38 22.075 ;
    RECT 81.17 22.365 81.38 22.435 ;
    RECT 81.63 21.645 81.84 21.715 ;
    RECT 81.63 22.005 81.84 22.075 ;
    RECT 81.63 22.365 81.84 22.435 ;
    RECT 77.85 21.645 78.06 21.715 ;
    RECT 77.85 22.005 78.06 22.075 ;
    RECT 77.85 22.365 78.06 22.435 ;
    RECT 78.31 21.645 78.52 21.715 ;
    RECT 78.31 22.005 78.52 22.075 ;
    RECT 78.31 22.365 78.52 22.435 ;
    RECT 74.53 21.645 74.74 21.715 ;
    RECT 74.53 22.005 74.74 22.075 ;
    RECT 74.53 22.365 74.74 22.435 ;
    RECT 74.99 21.645 75.2 21.715 ;
    RECT 74.99 22.005 75.2 22.075 ;
    RECT 74.99 22.365 75.2 22.435 ;
    RECT 71.21 21.645 71.42 21.715 ;
    RECT 71.21 22.005 71.42 22.075 ;
    RECT 71.21 22.365 71.42 22.435 ;
    RECT 71.67 21.645 71.88 21.715 ;
    RECT 71.67 22.005 71.88 22.075 ;
    RECT 71.67 22.365 71.88 22.435 ;
    RECT 31.37 21.645 31.58 21.715 ;
    RECT 31.37 22.005 31.58 22.075 ;
    RECT 31.37 22.365 31.58 22.435 ;
    RECT 31.83 21.645 32.04 21.715 ;
    RECT 31.83 22.005 32.04 22.075 ;
    RECT 31.83 22.365 32.04 22.435 ;
    RECT 67.89 21.645 68.1 21.715 ;
    RECT 67.89 22.005 68.1 22.075 ;
    RECT 67.89 22.365 68.1 22.435 ;
    RECT 68.35 21.645 68.56 21.715 ;
    RECT 68.35 22.005 68.56 22.075 ;
    RECT 68.35 22.365 68.56 22.435 ;
    RECT 28.05 21.645 28.26 21.715 ;
    RECT 28.05 22.005 28.26 22.075 ;
    RECT 28.05 22.365 28.26 22.435 ;
    RECT 28.51 21.645 28.72 21.715 ;
    RECT 28.51 22.005 28.72 22.075 ;
    RECT 28.51 22.365 28.72 22.435 ;
    RECT 24.73 21.645 24.94 21.715 ;
    RECT 24.73 22.005 24.94 22.075 ;
    RECT 24.73 22.365 24.94 22.435 ;
    RECT 25.19 21.645 25.4 21.715 ;
    RECT 25.19 22.005 25.4 22.075 ;
    RECT 25.19 22.365 25.4 22.435 ;
    RECT 21.41 21.645 21.62 21.715 ;
    RECT 21.41 22.005 21.62 22.075 ;
    RECT 21.41 22.365 21.62 22.435 ;
    RECT 21.87 21.645 22.08 21.715 ;
    RECT 21.87 22.005 22.08 22.075 ;
    RECT 21.87 22.365 22.08 22.435 ;
    RECT 18.09 21.645 18.3 21.715 ;
    RECT 18.09 22.005 18.3 22.075 ;
    RECT 18.09 22.365 18.3 22.435 ;
    RECT 18.55 21.645 18.76 21.715 ;
    RECT 18.55 22.005 18.76 22.075 ;
    RECT 18.55 22.365 18.76 22.435 ;
    RECT 14.77 21.645 14.98 21.715 ;
    RECT 14.77 22.005 14.98 22.075 ;
    RECT 14.77 22.365 14.98 22.435 ;
    RECT 15.23 21.645 15.44 21.715 ;
    RECT 15.23 22.005 15.44 22.075 ;
    RECT 15.23 22.365 15.44 22.435 ;
    RECT 11.45 21.645 11.66 21.715 ;
    RECT 11.45 22.005 11.66 22.075 ;
    RECT 11.45 22.365 11.66 22.435 ;
    RECT 11.91 21.645 12.12 21.715 ;
    RECT 11.91 22.005 12.12 22.075 ;
    RECT 11.91 22.365 12.12 22.435 ;
    RECT 8.13 21.645 8.34 21.715 ;
    RECT 8.13 22.005 8.34 22.075 ;
    RECT 8.13 22.365 8.34 22.435 ;
    RECT 8.59 21.645 8.8 21.715 ;
    RECT 8.59 22.005 8.8 22.075 ;
    RECT 8.59 22.365 8.8 22.435 ;
    RECT 4.81 21.645 5.02 21.715 ;
    RECT 4.81 22.005 5.02 22.075 ;
    RECT 4.81 22.365 5.02 22.435 ;
    RECT 5.27 21.645 5.48 21.715 ;
    RECT 5.27 22.005 5.48 22.075 ;
    RECT 5.27 22.365 5.48 22.435 ;
    RECT 164.17 21.645 164.38 21.715 ;
    RECT 164.17 22.005 164.38 22.075 ;
    RECT 164.17 22.365 164.38 22.435 ;
    RECT 164.63 21.645 164.84 21.715 ;
    RECT 164.63 22.005 164.84 22.075 ;
    RECT 164.63 22.365 164.84 22.435 ;
    RECT 1.49 21.645 1.7 21.715 ;
    RECT 1.49 22.005 1.7 22.075 ;
    RECT 1.49 22.365 1.7 22.435 ;
    RECT 1.95 21.645 2.16 21.715 ;
    RECT 1.95 22.005 2.16 22.075 ;
    RECT 1.95 22.365 2.16 22.435 ;
    RECT 160.85 21.645 161.06 21.715 ;
    RECT 160.85 22.005 161.06 22.075 ;
    RECT 160.85 22.365 161.06 22.435 ;
    RECT 161.31 21.645 161.52 21.715 ;
    RECT 161.31 22.005 161.52 22.075 ;
    RECT 161.31 22.365 161.52 22.435 ;
    RECT 157.53 21.645 157.74 21.715 ;
    RECT 157.53 22.005 157.74 22.075 ;
    RECT 157.53 22.365 157.74 22.435 ;
    RECT 157.99 21.645 158.2 21.715 ;
    RECT 157.99 22.005 158.2 22.075 ;
    RECT 157.99 22.365 158.2 22.435 ;
    RECT 154.21 21.645 154.42 21.715 ;
    RECT 154.21 22.005 154.42 22.075 ;
    RECT 154.21 22.365 154.42 22.435 ;
    RECT 154.67 21.645 154.88 21.715 ;
    RECT 154.67 22.005 154.88 22.075 ;
    RECT 154.67 22.365 154.88 22.435 ;
    RECT 150.89 21.645 151.1 21.715 ;
    RECT 150.89 22.005 151.1 22.075 ;
    RECT 150.89 22.365 151.1 22.435 ;
    RECT 151.35 21.645 151.56 21.715 ;
    RECT 151.35 22.005 151.56 22.075 ;
    RECT 151.35 22.365 151.56 22.435 ;
    RECT 147.57 21.645 147.78 21.715 ;
    RECT 147.57 22.005 147.78 22.075 ;
    RECT 147.57 22.365 147.78 22.435 ;
    RECT 148.03 21.645 148.24 21.715 ;
    RECT 148.03 22.005 148.24 22.075 ;
    RECT 148.03 22.365 148.24 22.435 ;
    RECT 144.25 21.645 144.46 21.715 ;
    RECT 144.25 22.005 144.46 22.075 ;
    RECT 144.25 22.365 144.46 22.435 ;
    RECT 144.71 21.645 144.92 21.715 ;
    RECT 144.71 22.005 144.92 22.075 ;
    RECT 144.71 22.365 144.92 22.435 ;
    RECT 140.93 21.645 141.14 21.715 ;
    RECT 140.93 22.005 141.14 22.075 ;
    RECT 140.93 22.365 141.14 22.435 ;
    RECT 141.39 21.645 141.6 21.715 ;
    RECT 141.39 22.005 141.6 22.075 ;
    RECT 141.39 22.365 141.6 22.435 ;
    RECT 137.61 21.645 137.82 21.715 ;
    RECT 137.61 22.005 137.82 22.075 ;
    RECT 137.61 22.365 137.82 22.435 ;
    RECT 138.07 21.645 138.28 21.715 ;
    RECT 138.07 22.005 138.28 22.075 ;
    RECT 138.07 22.365 138.28 22.435 ;
    RECT 134.29 21.645 134.5 21.715 ;
    RECT 134.29 22.005 134.5 22.075 ;
    RECT 134.29 22.365 134.5 22.435 ;
    RECT 134.75 21.645 134.96 21.715 ;
    RECT 134.75 22.005 134.96 22.075 ;
    RECT 134.75 22.365 134.96 22.435 ;
    RECT 64.57 21.645 64.78 21.715 ;
    RECT 64.57 22.005 64.78 22.075 ;
    RECT 64.57 22.365 64.78 22.435 ;
    RECT 65.03 21.645 65.24 21.715 ;
    RECT 65.03 22.005 65.24 22.075 ;
    RECT 65.03 22.365 65.24 22.435 ;
    RECT 61.25 20.925 61.46 20.995 ;
    RECT 61.25 21.285 61.46 21.355 ;
    RECT 61.25 21.645 61.46 21.715 ;
    RECT 61.71 20.925 61.92 20.995 ;
    RECT 61.71 21.285 61.92 21.355 ;
    RECT 61.71 21.645 61.92 21.715 ;
    RECT 57.93 20.925 58.14 20.995 ;
    RECT 57.93 21.285 58.14 21.355 ;
    RECT 57.93 21.645 58.14 21.715 ;
    RECT 58.39 20.925 58.6 20.995 ;
    RECT 58.39 21.285 58.6 21.355 ;
    RECT 58.39 21.645 58.6 21.715 ;
    RECT 54.61 20.925 54.82 20.995 ;
    RECT 54.61 21.285 54.82 21.355 ;
    RECT 54.61 21.645 54.82 21.715 ;
    RECT 55.07 20.925 55.28 20.995 ;
    RECT 55.07 21.285 55.28 21.355 ;
    RECT 55.07 21.645 55.28 21.715 ;
    RECT 51.29 20.925 51.5 20.995 ;
    RECT 51.29 21.285 51.5 21.355 ;
    RECT 51.29 21.645 51.5 21.715 ;
    RECT 51.75 20.925 51.96 20.995 ;
    RECT 51.75 21.285 51.96 21.355 ;
    RECT 51.75 21.645 51.96 21.715 ;
    RECT 47.97 20.925 48.18 20.995 ;
    RECT 47.97 21.285 48.18 21.355 ;
    RECT 47.97 21.645 48.18 21.715 ;
    RECT 48.43 20.925 48.64 20.995 ;
    RECT 48.43 21.285 48.64 21.355 ;
    RECT 48.43 21.645 48.64 21.715 ;
    RECT 44.65 20.925 44.86 20.995 ;
    RECT 44.65 21.285 44.86 21.355 ;
    RECT 44.65 21.645 44.86 21.715 ;
    RECT 45.11 20.925 45.32 20.995 ;
    RECT 45.11 21.285 45.32 21.355 ;
    RECT 45.11 21.645 45.32 21.715 ;
    RECT 41.33 20.925 41.54 20.995 ;
    RECT 41.33 21.285 41.54 21.355 ;
    RECT 41.33 21.645 41.54 21.715 ;
    RECT 41.79 20.925 42.0 20.995 ;
    RECT 41.79 21.285 42.0 21.355 ;
    RECT 41.79 21.645 42.0 21.715 ;
    RECT 38.01 20.925 38.22 20.995 ;
    RECT 38.01 21.285 38.22 21.355 ;
    RECT 38.01 21.645 38.22 21.715 ;
    RECT 38.47 20.925 38.68 20.995 ;
    RECT 38.47 21.285 38.68 21.355 ;
    RECT 38.47 21.645 38.68 21.715 ;
    RECT 34.69 20.925 34.9 20.995 ;
    RECT 34.69 21.285 34.9 21.355 ;
    RECT 34.69 21.645 34.9 21.715 ;
    RECT 35.15 20.925 35.36 20.995 ;
    RECT 35.15 21.285 35.36 21.355 ;
    RECT 35.15 21.645 35.36 21.715 ;
    RECT 173.945 21.285 174.015 21.355 ;
    RECT 130.97 20.925 131.18 20.995 ;
    RECT 130.97 21.285 131.18 21.355 ;
    RECT 130.97 21.645 131.18 21.715 ;
    RECT 131.43 20.925 131.64 20.995 ;
    RECT 131.43 21.285 131.64 21.355 ;
    RECT 131.43 21.645 131.64 21.715 ;
    RECT 127.65 20.925 127.86 20.995 ;
    RECT 127.65 21.285 127.86 21.355 ;
    RECT 127.65 21.645 127.86 21.715 ;
    RECT 128.11 20.925 128.32 20.995 ;
    RECT 128.11 21.285 128.32 21.355 ;
    RECT 128.11 21.645 128.32 21.715 ;
    RECT 124.33 20.925 124.54 20.995 ;
    RECT 124.33 21.285 124.54 21.355 ;
    RECT 124.33 21.645 124.54 21.715 ;
    RECT 124.79 20.925 125.0 20.995 ;
    RECT 124.79 21.285 125.0 21.355 ;
    RECT 124.79 21.645 125.0 21.715 ;
    RECT 121.01 20.925 121.22 20.995 ;
    RECT 121.01 21.285 121.22 21.355 ;
    RECT 121.01 21.645 121.22 21.715 ;
    RECT 121.47 20.925 121.68 20.995 ;
    RECT 121.47 21.285 121.68 21.355 ;
    RECT 121.47 21.645 121.68 21.715 ;
    RECT 117.69 20.925 117.9 20.995 ;
    RECT 117.69 21.285 117.9 21.355 ;
    RECT 117.69 21.645 117.9 21.715 ;
    RECT 118.15 20.925 118.36 20.995 ;
    RECT 118.15 21.285 118.36 21.355 ;
    RECT 118.15 21.645 118.36 21.715 ;
    RECT 114.37 20.925 114.58 20.995 ;
    RECT 114.37 21.285 114.58 21.355 ;
    RECT 114.37 21.645 114.58 21.715 ;
    RECT 114.83 20.925 115.04 20.995 ;
    RECT 114.83 21.285 115.04 21.355 ;
    RECT 114.83 21.645 115.04 21.715 ;
    RECT 111.05 20.925 111.26 20.995 ;
    RECT 111.05 21.285 111.26 21.355 ;
    RECT 111.05 21.645 111.26 21.715 ;
    RECT 111.51 20.925 111.72 20.995 ;
    RECT 111.51 21.285 111.72 21.355 ;
    RECT 111.51 21.645 111.72 21.715 ;
    RECT 107.73 20.925 107.94 20.995 ;
    RECT 107.73 21.285 107.94 21.355 ;
    RECT 107.73 21.645 107.94 21.715 ;
    RECT 108.19 20.925 108.4 20.995 ;
    RECT 108.19 21.285 108.4 21.355 ;
    RECT 108.19 21.645 108.4 21.715 ;
    RECT 104.41 20.925 104.62 20.995 ;
    RECT 104.41 21.285 104.62 21.355 ;
    RECT 104.41 21.645 104.62 21.715 ;
    RECT 104.87 20.925 105.08 20.995 ;
    RECT 104.87 21.285 105.08 21.355 ;
    RECT 104.87 21.645 105.08 21.715 ;
    RECT 101.09 20.925 101.3 20.995 ;
    RECT 101.09 21.285 101.3 21.355 ;
    RECT 101.09 21.645 101.3 21.715 ;
    RECT 101.55 20.925 101.76 20.995 ;
    RECT 101.55 21.285 101.76 21.355 ;
    RECT 101.55 21.645 101.76 21.715 ;
    RECT 0.4 21.285 0.47 21.355 ;
    RECT 170.81 20.925 171.02 20.995 ;
    RECT 170.81 21.285 171.02 21.355 ;
    RECT 170.81 21.645 171.02 21.715 ;
    RECT 171.27 20.925 171.48 20.995 ;
    RECT 171.27 21.285 171.48 21.355 ;
    RECT 171.27 21.645 171.48 21.715 ;
    RECT 167.49 20.925 167.7 20.995 ;
    RECT 167.49 21.285 167.7 21.355 ;
    RECT 167.49 21.645 167.7 21.715 ;
    RECT 167.95 20.925 168.16 20.995 ;
    RECT 167.95 21.285 168.16 21.355 ;
    RECT 167.95 21.645 168.16 21.715 ;
    RECT 97.77 20.925 97.98 20.995 ;
    RECT 97.77 21.285 97.98 21.355 ;
    RECT 97.77 21.645 97.98 21.715 ;
    RECT 98.23 20.925 98.44 20.995 ;
    RECT 98.23 21.285 98.44 21.355 ;
    RECT 98.23 21.645 98.44 21.715 ;
    RECT 94.45 20.925 94.66 20.995 ;
    RECT 94.45 21.285 94.66 21.355 ;
    RECT 94.45 21.645 94.66 21.715 ;
    RECT 94.91 20.925 95.12 20.995 ;
    RECT 94.91 21.285 95.12 21.355 ;
    RECT 94.91 21.645 95.12 21.715 ;
    RECT 91.13 20.925 91.34 20.995 ;
    RECT 91.13 21.285 91.34 21.355 ;
    RECT 91.13 21.645 91.34 21.715 ;
    RECT 91.59 20.925 91.8 20.995 ;
    RECT 91.59 21.285 91.8 21.355 ;
    RECT 91.59 21.645 91.8 21.715 ;
    RECT 87.81 20.925 88.02 20.995 ;
    RECT 87.81 21.285 88.02 21.355 ;
    RECT 87.81 21.645 88.02 21.715 ;
    RECT 88.27 20.925 88.48 20.995 ;
    RECT 88.27 21.285 88.48 21.355 ;
    RECT 88.27 21.645 88.48 21.715 ;
    RECT 84.49 20.925 84.7 20.995 ;
    RECT 84.49 21.285 84.7 21.355 ;
    RECT 84.49 21.645 84.7 21.715 ;
    RECT 84.95 20.925 85.16 20.995 ;
    RECT 84.95 21.285 85.16 21.355 ;
    RECT 84.95 21.645 85.16 21.715 ;
    RECT 81.17 20.925 81.38 20.995 ;
    RECT 81.17 21.285 81.38 21.355 ;
    RECT 81.17 21.645 81.38 21.715 ;
    RECT 81.63 20.925 81.84 20.995 ;
    RECT 81.63 21.285 81.84 21.355 ;
    RECT 81.63 21.645 81.84 21.715 ;
    RECT 77.85 20.925 78.06 20.995 ;
    RECT 77.85 21.285 78.06 21.355 ;
    RECT 77.85 21.645 78.06 21.715 ;
    RECT 78.31 20.925 78.52 20.995 ;
    RECT 78.31 21.285 78.52 21.355 ;
    RECT 78.31 21.645 78.52 21.715 ;
    RECT 74.53 20.925 74.74 20.995 ;
    RECT 74.53 21.285 74.74 21.355 ;
    RECT 74.53 21.645 74.74 21.715 ;
    RECT 74.99 20.925 75.2 20.995 ;
    RECT 74.99 21.285 75.2 21.355 ;
    RECT 74.99 21.645 75.2 21.715 ;
    RECT 71.21 20.925 71.42 20.995 ;
    RECT 71.21 21.285 71.42 21.355 ;
    RECT 71.21 21.645 71.42 21.715 ;
    RECT 71.67 20.925 71.88 20.995 ;
    RECT 71.67 21.285 71.88 21.355 ;
    RECT 71.67 21.645 71.88 21.715 ;
    RECT 31.37 20.925 31.58 20.995 ;
    RECT 31.37 21.285 31.58 21.355 ;
    RECT 31.37 21.645 31.58 21.715 ;
    RECT 31.83 20.925 32.04 20.995 ;
    RECT 31.83 21.285 32.04 21.355 ;
    RECT 31.83 21.645 32.04 21.715 ;
    RECT 67.89 20.925 68.1 20.995 ;
    RECT 67.89 21.285 68.1 21.355 ;
    RECT 67.89 21.645 68.1 21.715 ;
    RECT 68.35 20.925 68.56 20.995 ;
    RECT 68.35 21.285 68.56 21.355 ;
    RECT 68.35 21.645 68.56 21.715 ;
    RECT 28.05 20.925 28.26 20.995 ;
    RECT 28.05 21.285 28.26 21.355 ;
    RECT 28.05 21.645 28.26 21.715 ;
    RECT 28.51 20.925 28.72 20.995 ;
    RECT 28.51 21.285 28.72 21.355 ;
    RECT 28.51 21.645 28.72 21.715 ;
    RECT 24.73 20.925 24.94 20.995 ;
    RECT 24.73 21.285 24.94 21.355 ;
    RECT 24.73 21.645 24.94 21.715 ;
    RECT 25.19 20.925 25.4 20.995 ;
    RECT 25.19 21.285 25.4 21.355 ;
    RECT 25.19 21.645 25.4 21.715 ;
    RECT 21.41 20.925 21.62 20.995 ;
    RECT 21.41 21.285 21.62 21.355 ;
    RECT 21.41 21.645 21.62 21.715 ;
    RECT 21.87 20.925 22.08 20.995 ;
    RECT 21.87 21.285 22.08 21.355 ;
    RECT 21.87 21.645 22.08 21.715 ;
    RECT 18.09 20.925 18.3 20.995 ;
    RECT 18.09 21.285 18.3 21.355 ;
    RECT 18.09 21.645 18.3 21.715 ;
    RECT 18.55 20.925 18.76 20.995 ;
    RECT 18.55 21.285 18.76 21.355 ;
    RECT 18.55 21.645 18.76 21.715 ;
    RECT 14.77 20.925 14.98 20.995 ;
    RECT 14.77 21.285 14.98 21.355 ;
    RECT 14.77 21.645 14.98 21.715 ;
    RECT 15.23 20.925 15.44 20.995 ;
    RECT 15.23 21.285 15.44 21.355 ;
    RECT 15.23 21.645 15.44 21.715 ;
    RECT 11.45 20.925 11.66 20.995 ;
    RECT 11.45 21.285 11.66 21.355 ;
    RECT 11.45 21.645 11.66 21.715 ;
    RECT 11.91 20.925 12.12 20.995 ;
    RECT 11.91 21.285 12.12 21.355 ;
    RECT 11.91 21.645 12.12 21.715 ;
    RECT 8.13 20.925 8.34 20.995 ;
    RECT 8.13 21.285 8.34 21.355 ;
    RECT 8.13 21.645 8.34 21.715 ;
    RECT 8.59 20.925 8.8 20.995 ;
    RECT 8.59 21.285 8.8 21.355 ;
    RECT 8.59 21.645 8.8 21.715 ;
    RECT 4.81 20.925 5.02 20.995 ;
    RECT 4.81 21.285 5.02 21.355 ;
    RECT 4.81 21.645 5.02 21.715 ;
    RECT 5.27 20.925 5.48 20.995 ;
    RECT 5.27 21.285 5.48 21.355 ;
    RECT 5.27 21.645 5.48 21.715 ;
    RECT 164.17 20.925 164.38 20.995 ;
    RECT 164.17 21.285 164.38 21.355 ;
    RECT 164.17 21.645 164.38 21.715 ;
    RECT 164.63 20.925 164.84 20.995 ;
    RECT 164.63 21.285 164.84 21.355 ;
    RECT 164.63 21.645 164.84 21.715 ;
    RECT 1.49 20.925 1.7 20.995 ;
    RECT 1.49 21.285 1.7 21.355 ;
    RECT 1.49 21.645 1.7 21.715 ;
    RECT 1.95 20.925 2.16 20.995 ;
    RECT 1.95 21.285 2.16 21.355 ;
    RECT 1.95 21.645 2.16 21.715 ;
    RECT 160.85 20.925 161.06 20.995 ;
    RECT 160.85 21.285 161.06 21.355 ;
    RECT 160.85 21.645 161.06 21.715 ;
    RECT 161.31 20.925 161.52 20.995 ;
    RECT 161.31 21.285 161.52 21.355 ;
    RECT 161.31 21.645 161.52 21.715 ;
    RECT 157.53 20.925 157.74 20.995 ;
    RECT 157.53 21.285 157.74 21.355 ;
    RECT 157.53 21.645 157.74 21.715 ;
    RECT 157.99 20.925 158.2 20.995 ;
    RECT 157.99 21.285 158.2 21.355 ;
    RECT 157.99 21.645 158.2 21.715 ;
    RECT 154.21 20.925 154.42 20.995 ;
    RECT 154.21 21.285 154.42 21.355 ;
    RECT 154.21 21.645 154.42 21.715 ;
    RECT 154.67 20.925 154.88 20.995 ;
    RECT 154.67 21.285 154.88 21.355 ;
    RECT 154.67 21.645 154.88 21.715 ;
    RECT 150.89 20.925 151.1 20.995 ;
    RECT 150.89 21.285 151.1 21.355 ;
    RECT 150.89 21.645 151.1 21.715 ;
    RECT 151.35 20.925 151.56 20.995 ;
    RECT 151.35 21.285 151.56 21.355 ;
    RECT 151.35 21.645 151.56 21.715 ;
    RECT 147.57 20.925 147.78 20.995 ;
    RECT 147.57 21.285 147.78 21.355 ;
    RECT 147.57 21.645 147.78 21.715 ;
    RECT 148.03 20.925 148.24 20.995 ;
    RECT 148.03 21.285 148.24 21.355 ;
    RECT 148.03 21.645 148.24 21.715 ;
    RECT 144.25 20.925 144.46 20.995 ;
    RECT 144.25 21.285 144.46 21.355 ;
    RECT 144.25 21.645 144.46 21.715 ;
    RECT 144.71 20.925 144.92 20.995 ;
    RECT 144.71 21.285 144.92 21.355 ;
    RECT 144.71 21.645 144.92 21.715 ;
    RECT 140.93 20.925 141.14 20.995 ;
    RECT 140.93 21.285 141.14 21.355 ;
    RECT 140.93 21.645 141.14 21.715 ;
    RECT 141.39 20.925 141.6 20.995 ;
    RECT 141.39 21.285 141.6 21.355 ;
    RECT 141.39 21.645 141.6 21.715 ;
    RECT 137.61 20.925 137.82 20.995 ;
    RECT 137.61 21.285 137.82 21.355 ;
    RECT 137.61 21.645 137.82 21.715 ;
    RECT 138.07 20.925 138.28 20.995 ;
    RECT 138.07 21.285 138.28 21.355 ;
    RECT 138.07 21.645 138.28 21.715 ;
    RECT 134.29 20.925 134.5 20.995 ;
    RECT 134.29 21.285 134.5 21.355 ;
    RECT 134.29 21.645 134.5 21.715 ;
    RECT 134.75 20.925 134.96 20.995 ;
    RECT 134.75 21.285 134.96 21.355 ;
    RECT 134.75 21.645 134.96 21.715 ;
    RECT 64.57 20.925 64.78 20.995 ;
    RECT 64.57 21.285 64.78 21.355 ;
    RECT 64.57 21.645 64.78 21.715 ;
    RECT 65.03 20.925 65.24 20.995 ;
    RECT 65.03 21.285 65.24 21.355 ;
    RECT 65.03 21.645 65.24 21.715 ;
    RECT 61.25 20.205 61.46 20.275 ;
    RECT 61.25 20.565 61.46 20.635 ;
    RECT 61.25 20.925 61.46 20.995 ;
    RECT 61.71 20.205 61.92 20.275 ;
    RECT 61.71 20.565 61.92 20.635 ;
    RECT 61.71 20.925 61.92 20.995 ;
    RECT 57.93 20.205 58.14 20.275 ;
    RECT 57.93 20.565 58.14 20.635 ;
    RECT 57.93 20.925 58.14 20.995 ;
    RECT 58.39 20.205 58.6 20.275 ;
    RECT 58.39 20.565 58.6 20.635 ;
    RECT 58.39 20.925 58.6 20.995 ;
    RECT 54.61 20.205 54.82 20.275 ;
    RECT 54.61 20.565 54.82 20.635 ;
    RECT 54.61 20.925 54.82 20.995 ;
    RECT 55.07 20.205 55.28 20.275 ;
    RECT 55.07 20.565 55.28 20.635 ;
    RECT 55.07 20.925 55.28 20.995 ;
    RECT 51.29 20.205 51.5 20.275 ;
    RECT 51.29 20.565 51.5 20.635 ;
    RECT 51.29 20.925 51.5 20.995 ;
    RECT 51.75 20.205 51.96 20.275 ;
    RECT 51.75 20.565 51.96 20.635 ;
    RECT 51.75 20.925 51.96 20.995 ;
    RECT 47.97 20.205 48.18 20.275 ;
    RECT 47.97 20.565 48.18 20.635 ;
    RECT 47.97 20.925 48.18 20.995 ;
    RECT 48.43 20.205 48.64 20.275 ;
    RECT 48.43 20.565 48.64 20.635 ;
    RECT 48.43 20.925 48.64 20.995 ;
    RECT 44.65 20.205 44.86 20.275 ;
    RECT 44.65 20.565 44.86 20.635 ;
    RECT 44.65 20.925 44.86 20.995 ;
    RECT 45.11 20.205 45.32 20.275 ;
    RECT 45.11 20.565 45.32 20.635 ;
    RECT 45.11 20.925 45.32 20.995 ;
    RECT 41.33 20.205 41.54 20.275 ;
    RECT 41.33 20.565 41.54 20.635 ;
    RECT 41.33 20.925 41.54 20.995 ;
    RECT 41.79 20.205 42.0 20.275 ;
    RECT 41.79 20.565 42.0 20.635 ;
    RECT 41.79 20.925 42.0 20.995 ;
    RECT 38.01 20.205 38.22 20.275 ;
    RECT 38.01 20.565 38.22 20.635 ;
    RECT 38.01 20.925 38.22 20.995 ;
    RECT 38.47 20.205 38.68 20.275 ;
    RECT 38.47 20.565 38.68 20.635 ;
    RECT 38.47 20.925 38.68 20.995 ;
    RECT 34.69 20.205 34.9 20.275 ;
    RECT 34.69 20.565 34.9 20.635 ;
    RECT 34.69 20.925 34.9 20.995 ;
    RECT 35.15 20.205 35.36 20.275 ;
    RECT 35.15 20.565 35.36 20.635 ;
    RECT 35.15 20.925 35.36 20.995 ;
    RECT 173.945 20.565 174.015 20.635 ;
    RECT 130.97 20.205 131.18 20.275 ;
    RECT 130.97 20.565 131.18 20.635 ;
    RECT 130.97 20.925 131.18 20.995 ;
    RECT 131.43 20.205 131.64 20.275 ;
    RECT 131.43 20.565 131.64 20.635 ;
    RECT 131.43 20.925 131.64 20.995 ;
    RECT 127.65 20.205 127.86 20.275 ;
    RECT 127.65 20.565 127.86 20.635 ;
    RECT 127.65 20.925 127.86 20.995 ;
    RECT 128.11 20.205 128.32 20.275 ;
    RECT 128.11 20.565 128.32 20.635 ;
    RECT 128.11 20.925 128.32 20.995 ;
    RECT 124.33 20.205 124.54 20.275 ;
    RECT 124.33 20.565 124.54 20.635 ;
    RECT 124.33 20.925 124.54 20.995 ;
    RECT 124.79 20.205 125.0 20.275 ;
    RECT 124.79 20.565 125.0 20.635 ;
    RECT 124.79 20.925 125.0 20.995 ;
    RECT 121.01 20.205 121.22 20.275 ;
    RECT 121.01 20.565 121.22 20.635 ;
    RECT 121.01 20.925 121.22 20.995 ;
    RECT 121.47 20.205 121.68 20.275 ;
    RECT 121.47 20.565 121.68 20.635 ;
    RECT 121.47 20.925 121.68 20.995 ;
    RECT 117.69 20.205 117.9 20.275 ;
    RECT 117.69 20.565 117.9 20.635 ;
    RECT 117.69 20.925 117.9 20.995 ;
    RECT 118.15 20.205 118.36 20.275 ;
    RECT 118.15 20.565 118.36 20.635 ;
    RECT 118.15 20.925 118.36 20.995 ;
    RECT 114.37 20.205 114.58 20.275 ;
    RECT 114.37 20.565 114.58 20.635 ;
    RECT 114.37 20.925 114.58 20.995 ;
    RECT 114.83 20.205 115.04 20.275 ;
    RECT 114.83 20.565 115.04 20.635 ;
    RECT 114.83 20.925 115.04 20.995 ;
    RECT 111.05 20.205 111.26 20.275 ;
    RECT 111.05 20.565 111.26 20.635 ;
    RECT 111.05 20.925 111.26 20.995 ;
    RECT 111.51 20.205 111.72 20.275 ;
    RECT 111.51 20.565 111.72 20.635 ;
    RECT 111.51 20.925 111.72 20.995 ;
    RECT 107.73 20.205 107.94 20.275 ;
    RECT 107.73 20.565 107.94 20.635 ;
    RECT 107.73 20.925 107.94 20.995 ;
    RECT 108.19 20.205 108.4 20.275 ;
    RECT 108.19 20.565 108.4 20.635 ;
    RECT 108.19 20.925 108.4 20.995 ;
    RECT 104.41 20.205 104.62 20.275 ;
    RECT 104.41 20.565 104.62 20.635 ;
    RECT 104.41 20.925 104.62 20.995 ;
    RECT 104.87 20.205 105.08 20.275 ;
    RECT 104.87 20.565 105.08 20.635 ;
    RECT 104.87 20.925 105.08 20.995 ;
    RECT 101.09 20.205 101.3 20.275 ;
    RECT 101.09 20.565 101.3 20.635 ;
    RECT 101.09 20.925 101.3 20.995 ;
    RECT 101.55 20.205 101.76 20.275 ;
    RECT 101.55 20.565 101.76 20.635 ;
    RECT 101.55 20.925 101.76 20.995 ;
    RECT 0.4 20.565 0.47 20.635 ;
    RECT 170.81 20.205 171.02 20.275 ;
    RECT 170.81 20.565 171.02 20.635 ;
    RECT 170.81 20.925 171.02 20.995 ;
    RECT 171.27 20.205 171.48 20.275 ;
    RECT 171.27 20.565 171.48 20.635 ;
    RECT 171.27 20.925 171.48 20.995 ;
    RECT 167.49 20.205 167.7 20.275 ;
    RECT 167.49 20.565 167.7 20.635 ;
    RECT 167.49 20.925 167.7 20.995 ;
    RECT 167.95 20.205 168.16 20.275 ;
    RECT 167.95 20.565 168.16 20.635 ;
    RECT 167.95 20.925 168.16 20.995 ;
    RECT 97.77 20.205 97.98 20.275 ;
    RECT 97.77 20.565 97.98 20.635 ;
    RECT 97.77 20.925 97.98 20.995 ;
    RECT 98.23 20.205 98.44 20.275 ;
    RECT 98.23 20.565 98.44 20.635 ;
    RECT 98.23 20.925 98.44 20.995 ;
    RECT 94.45 20.205 94.66 20.275 ;
    RECT 94.45 20.565 94.66 20.635 ;
    RECT 94.45 20.925 94.66 20.995 ;
    RECT 94.91 20.205 95.12 20.275 ;
    RECT 94.91 20.565 95.12 20.635 ;
    RECT 94.91 20.925 95.12 20.995 ;
    RECT 91.13 20.205 91.34 20.275 ;
    RECT 91.13 20.565 91.34 20.635 ;
    RECT 91.13 20.925 91.34 20.995 ;
    RECT 91.59 20.205 91.8 20.275 ;
    RECT 91.59 20.565 91.8 20.635 ;
    RECT 91.59 20.925 91.8 20.995 ;
    RECT 87.81 20.205 88.02 20.275 ;
    RECT 87.81 20.565 88.02 20.635 ;
    RECT 87.81 20.925 88.02 20.995 ;
    RECT 88.27 20.205 88.48 20.275 ;
    RECT 88.27 20.565 88.48 20.635 ;
    RECT 88.27 20.925 88.48 20.995 ;
    RECT 84.49 20.205 84.7 20.275 ;
    RECT 84.49 20.565 84.7 20.635 ;
    RECT 84.49 20.925 84.7 20.995 ;
    RECT 84.95 20.205 85.16 20.275 ;
    RECT 84.95 20.565 85.16 20.635 ;
    RECT 84.95 20.925 85.16 20.995 ;
    RECT 81.17 20.205 81.38 20.275 ;
    RECT 81.17 20.565 81.38 20.635 ;
    RECT 81.17 20.925 81.38 20.995 ;
    RECT 81.63 20.205 81.84 20.275 ;
    RECT 81.63 20.565 81.84 20.635 ;
    RECT 81.63 20.925 81.84 20.995 ;
    RECT 77.85 20.205 78.06 20.275 ;
    RECT 77.85 20.565 78.06 20.635 ;
    RECT 77.85 20.925 78.06 20.995 ;
    RECT 78.31 20.205 78.52 20.275 ;
    RECT 78.31 20.565 78.52 20.635 ;
    RECT 78.31 20.925 78.52 20.995 ;
    RECT 74.53 20.205 74.74 20.275 ;
    RECT 74.53 20.565 74.74 20.635 ;
    RECT 74.53 20.925 74.74 20.995 ;
    RECT 74.99 20.205 75.2 20.275 ;
    RECT 74.99 20.565 75.2 20.635 ;
    RECT 74.99 20.925 75.2 20.995 ;
    RECT 71.21 20.205 71.42 20.275 ;
    RECT 71.21 20.565 71.42 20.635 ;
    RECT 71.21 20.925 71.42 20.995 ;
    RECT 71.67 20.205 71.88 20.275 ;
    RECT 71.67 20.565 71.88 20.635 ;
    RECT 71.67 20.925 71.88 20.995 ;
    RECT 31.37 20.205 31.58 20.275 ;
    RECT 31.37 20.565 31.58 20.635 ;
    RECT 31.37 20.925 31.58 20.995 ;
    RECT 31.83 20.205 32.04 20.275 ;
    RECT 31.83 20.565 32.04 20.635 ;
    RECT 31.83 20.925 32.04 20.995 ;
    RECT 67.89 20.205 68.1 20.275 ;
    RECT 67.89 20.565 68.1 20.635 ;
    RECT 67.89 20.925 68.1 20.995 ;
    RECT 68.35 20.205 68.56 20.275 ;
    RECT 68.35 20.565 68.56 20.635 ;
    RECT 68.35 20.925 68.56 20.995 ;
    RECT 28.05 20.205 28.26 20.275 ;
    RECT 28.05 20.565 28.26 20.635 ;
    RECT 28.05 20.925 28.26 20.995 ;
    RECT 28.51 20.205 28.72 20.275 ;
    RECT 28.51 20.565 28.72 20.635 ;
    RECT 28.51 20.925 28.72 20.995 ;
    RECT 24.73 20.205 24.94 20.275 ;
    RECT 24.73 20.565 24.94 20.635 ;
    RECT 24.73 20.925 24.94 20.995 ;
    RECT 25.19 20.205 25.4 20.275 ;
    RECT 25.19 20.565 25.4 20.635 ;
    RECT 25.19 20.925 25.4 20.995 ;
    RECT 21.41 20.205 21.62 20.275 ;
    RECT 21.41 20.565 21.62 20.635 ;
    RECT 21.41 20.925 21.62 20.995 ;
    RECT 21.87 20.205 22.08 20.275 ;
    RECT 21.87 20.565 22.08 20.635 ;
    RECT 21.87 20.925 22.08 20.995 ;
    RECT 18.09 20.205 18.3 20.275 ;
    RECT 18.09 20.565 18.3 20.635 ;
    RECT 18.09 20.925 18.3 20.995 ;
    RECT 18.55 20.205 18.76 20.275 ;
    RECT 18.55 20.565 18.76 20.635 ;
    RECT 18.55 20.925 18.76 20.995 ;
    RECT 14.77 20.205 14.98 20.275 ;
    RECT 14.77 20.565 14.98 20.635 ;
    RECT 14.77 20.925 14.98 20.995 ;
    RECT 15.23 20.205 15.44 20.275 ;
    RECT 15.23 20.565 15.44 20.635 ;
    RECT 15.23 20.925 15.44 20.995 ;
    RECT 11.45 20.205 11.66 20.275 ;
    RECT 11.45 20.565 11.66 20.635 ;
    RECT 11.45 20.925 11.66 20.995 ;
    RECT 11.91 20.205 12.12 20.275 ;
    RECT 11.91 20.565 12.12 20.635 ;
    RECT 11.91 20.925 12.12 20.995 ;
    RECT 8.13 20.205 8.34 20.275 ;
    RECT 8.13 20.565 8.34 20.635 ;
    RECT 8.13 20.925 8.34 20.995 ;
    RECT 8.59 20.205 8.8 20.275 ;
    RECT 8.59 20.565 8.8 20.635 ;
    RECT 8.59 20.925 8.8 20.995 ;
    RECT 4.81 20.205 5.02 20.275 ;
    RECT 4.81 20.565 5.02 20.635 ;
    RECT 4.81 20.925 5.02 20.995 ;
    RECT 5.27 20.205 5.48 20.275 ;
    RECT 5.27 20.565 5.48 20.635 ;
    RECT 5.27 20.925 5.48 20.995 ;
    RECT 164.17 20.205 164.38 20.275 ;
    RECT 164.17 20.565 164.38 20.635 ;
    RECT 164.17 20.925 164.38 20.995 ;
    RECT 164.63 20.205 164.84 20.275 ;
    RECT 164.63 20.565 164.84 20.635 ;
    RECT 164.63 20.925 164.84 20.995 ;
    RECT 1.49 20.205 1.7 20.275 ;
    RECT 1.49 20.565 1.7 20.635 ;
    RECT 1.49 20.925 1.7 20.995 ;
    RECT 1.95 20.205 2.16 20.275 ;
    RECT 1.95 20.565 2.16 20.635 ;
    RECT 1.95 20.925 2.16 20.995 ;
    RECT 160.85 20.205 161.06 20.275 ;
    RECT 160.85 20.565 161.06 20.635 ;
    RECT 160.85 20.925 161.06 20.995 ;
    RECT 161.31 20.205 161.52 20.275 ;
    RECT 161.31 20.565 161.52 20.635 ;
    RECT 161.31 20.925 161.52 20.995 ;
    RECT 157.53 20.205 157.74 20.275 ;
    RECT 157.53 20.565 157.74 20.635 ;
    RECT 157.53 20.925 157.74 20.995 ;
    RECT 157.99 20.205 158.2 20.275 ;
    RECT 157.99 20.565 158.2 20.635 ;
    RECT 157.99 20.925 158.2 20.995 ;
    RECT 154.21 20.205 154.42 20.275 ;
    RECT 154.21 20.565 154.42 20.635 ;
    RECT 154.21 20.925 154.42 20.995 ;
    RECT 154.67 20.205 154.88 20.275 ;
    RECT 154.67 20.565 154.88 20.635 ;
    RECT 154.67 20.925 154.88 20.995 ;
    RECT 150.89 20.205 151.1 20.275 ;
    RECT 150.89 20.565 151.1 20.635 ;
    RECT 150.89 20.925 151.1 20.995 ;
    RECT 151.35 20.205 151.56 20.275 ;
    RECT 151.35 20.565 151.56 20.635 ;
    RECT 151.35 20.925 151.56 20.995 ;
    RECT 147.57 20.205 147.78 20.275 ;
    RECT 147.57 20.565 147.78 20.635 ;
    RECT 147.57 20.925 147.78 20.995 ;
    RECT 148.03 20.205 148.24 20.275 ;
    RECT 148.03 20.565 148.24 20.635 ;
    RECT 148.03 20.925 148.24 20.995 ;
    RECT 144.25 20.205 144.46 20.275 ;
    RECT 144.25 20.565 144.46 20.635 ;
    RECT 144.25 20.925 144.46 20.995 ;
    RECT 144.71 20.205 144.92 20.275 ;
    RECT 144.71 20.565 144.92 20.635 ;
    RECT 144.71 20.925 144.92 20.995 ;
    RECT 140.93 20.205 141.14 20.275 ;
    RECT 140.93 20.565 141.14 20.635 ;
    RECT 140.93 20.925 141.14 20.995 ;
    RECT 141.39 20.205 141.6 20.275 ;
    RECT 141.39 20.565 141.6 20.635 ;
    RECT 141.39 20.925 141.6 20.995 ;
    RECT 137.61 20.205 137.82 20.275 ;
    RECT 137.61 20.565 137.82 20.635 ;
    RECT 137.61 20.925 137.82 20.995 ;
    RECT 138.07 20.205 138.28 20.275 ;
    RECT 138.07 20.565 138.28 20.635 ;
    RECT 138.07 20.925 138.28 20.995 ;
    RECT 134.29 20.205 134.5 20.275 ;
    RECT 134.29 20.565 134.5 20.635 ;
    RECT 134.29 20.925 134.5 20.995 ;
    RECT 134.75 20.205 134.96 20.275 ;
    RECT 134.75 20.565 134.96 20.635 ;
    RECT 134.75 20.925 134.96 20.995 ;
    RECT 64.57 20.205 64.78 20.275 ;
    RECT 64.57 20.565 64.78 20.635 ;
    RECT 64.57 20.925 64.78 20.995 ;
    RECT 65.03 20.205 65.24 20.275 ;
    RECT 65.03 20.565 65.24 20.635 ;
    RECT 65.03 20.925 65.24 20.995 ;
    RECT 61.25 19.485 61.46 19.555 ;
    RECT 61.25 19.845 61.46 19.915 ;
    RECT 61.25 20.205 61.46 20.275 ;
    RECT 61.71 19.485 61.92 19.555 ;
    RECT 61.71 19.845 61.92 19.915 ;
    RECT 61.71 20.205 61.92 20.275 ;
    RECT 57.93 19.485 58.14 19.555 ;
    RECT 57.93 19.845 58.14 19.915 ;
    RECT 57.93 20.205 58.14 20.275 ;
    RECT 58.39 19.485 58.6 19.555 ;
    RECT 58.39 19.845 58.6 19.915 ;
    RECT 58.39 20.205 58.6 20.275 ;
    RECT 54.61 19.485 54.82 19.555 ;
    RECT 54.61 19.845 54.82 19.915 ;
    RECT 54.61 20.205 54.82 20.275 ;
    RECT 55.07 19.485 55.28 19.555 ;
    RECT 55.07 19.845 55.28 19.915 ;
    RECT 55.07 20.205 55.28 20.275 ;
    RECT 51.29 19.485 51.5 19.555 ;
    RECT 51.29 19.845 51.5 19.915 ;
    RECT 51.29 20.205 51.5 20.275 ;
    RECT 51.75 19.485 51.96 19.555 ;
    RECT 51.75 19.845 51.96 19.915 ;
    RECT 51.75 20.205 51.96 20.275 ;
    RECT 47.97 19.485 48.18 19.555 ;
    RECT 47.97 19.845 48.18 19.915 ;
    RECT 47.97 20.205 48.18 20.275 ;
    RECT 48.43 19.485 48.64 19.555 ;
    RECT 48.43 19.845 48.64 19.915 ;
    RECT 48.43 20.205 48.64 20.275 ;
    RECT 44.65 19.485 44.86 19.555 ;
    RECT 44.65 19.845 44.86 19.915 ;
    RECT 44.65 20.205 44.86 20.275 ;
    RECT 45.11 19.485 45.32 19.555 ;
    RECT 45.11 19.845 45.32 19.915 ;
    RECT 45.11 20.205 45.32 20.275 ;
    RECT 41.33 19.485 41.54 19.555 ;
    RECT 41.33 19.845 41.54 19.915 ;
    RECT 41.33 20.205 41.54 20.275 ;
    RECT 41.79 19.485 42.0 19.555 ;
    RECT 41.79 19.845 42.0 19.915 ;
    RECT 41.79 20.205 42.0 20.275 ;
    RECT 38.01 19.485 38.22 19.555 ;
    RECT 38.01 19.845 38.22 19.915 ;
    RECT 38.01 20.205 38.22 20.275 ;
    RECT 38.47 19.485 38.68 19.555 ;
    RECT 38.47 19.845 38.68 19.915 ;
    RECT 38.47 20.205 38.68 20.275 ;
    RECT 34.69 19.485 34.9 19.555 ;
    RECT 34.69 19.845 34.9 19.915 ;
    RECT 34.69 20.205 34.9 20.275 ;
    RECT 35.15 19.485 35.36 19.555 ;
    RECT 35.15 19.845 35.36 19.915 ;
    RECT 35.15 20.205 35.36 20.275 ;
    RECT 173.945 19.845 174.015 19.915 ;
    RECT 130.97 19.485 131.18 19.555 ;
    RECT 130.97 19.845 131.18 19.915 ;
    RECT 130.97 20.205 131.18 20.275 ;
    RECT 131.43 19.485 131.64 19.555 ;
    RECT 131.43 19.845 131.64 19.915 ;
    RECT 131.43 20.205 131.64 20.275 ;
    RECT 127.65 19.485 127.86 19.555 ;
    RECT 127.65 19.845 127.86 19.915 ;
    RECT 127.65 20.205 127.86 20.275 ;
    RECT 128.11 19.485 128.32 19.555 ;
    RECT 128.11 19.845 128.32 19.915 ;
    RECT 128.11 20.205 128.32 20.275 ;
    RECT 124.33 19.485 124.54 19.555 ;
    RECT 124.33 19.845 124.54 19.915 ;
    RECT 124.33 20.205 124.54 20.275 ;
    RECT 124.79 19.485 125.0 19.555 ;
    RECT 124.79 19.845 125.0 19.915 ;
    RECT 124.79 20.205 125.0 20.275 ;
    RECT 121.01 19.485 121.22 19.555 ;
    RECT 121.01 19.845 121.22 19.915 ;
    RECT 121.01 20.205 121.22 20.275 ;
    RECT 121.47 19.485 121.68 19.555 ;
    RECT 121.47 19.845 121.68 19.915 ;
    RECT 121.47 20.205 121.68 20.275 ;
    RECT 117.69 19.485 117.9 19.555 ;
    RECT 117.69 19.845 117.9 19.915 ;
    RECT 117.69 20.205 117.9 20.275 ;
    RECT 118.15 19.485 118.36 19.555 ;
    RECT 118.15 19.845 118.36 19.915 ;
    RECT 118.15 20.205 118.36 20.275 ;
    RECT 114.37 19.485 114.58 19.555 ;
    RECT 114.37 19.845 114.58 19.915 ;
    RECT 114.37 20.205 114.58 20.275 ;
    RECT 114.83 19.485 115.04 19.555 ;
    RECT 114.83 19.845 115.04 19.915 ;
    RECT 114.83 20.205 115.04 20.275 ;
    RECT 111.05 19.485 111.26 19.555 ;
    RECT 111.05 19.845 111.26 19.915 ;
    RECT 111.05 20.205 111.26 20.275 ;
    RECT 111.51 19.485 111.72 19.555 ;
    RECT 111.51 19.845 111.72 19.915 ;
    RECT 111.51 20.205 111.72 20.275 ;
    RECT 107.73 19.485 107.94 19.555 ;
    RECT 107.73 19.845 107.94 19.915 ;
    RECT 107.73 20.205 107.94 20.275 ;
    RECT 108.19 19.485 108.4 19.555 ;
    RECT 108.19 19.845 108.4 19.915 ;
    RECT 108.19 20.205 108.4 20.275 ;
    RECT 104.41 19.485 104.62 19.555 ;
    RECT 104.41 19.845 104.62 19.915 ;
    RECT 104.41 20.205 104.62 20.275 ;
    RECT 104.87 19.485 105.08 19.555 ;
    RECT 104.87 19.845 105.08 19.915 ;
    RECT 104.87 20.205 105.08 20.275 ;
    RECT 101.09 19.485 101.3 19.555 ;
    RECT 101.09 19.845 101.3 19.915 ;
    RECT 101.09 20.205 101.3 20.275 ;
    RECT 101.55 19.485 101.76 19.555 ;
    RECT 101.55 19.845 101.76 19.915 ;
    RECT 101.55 20.205 101.76 20.275 ;
    RECT 0.4 19.845 0.47 19.915 ;
    RECT 170.81 19.485 171.02 19.555 ;
    RECT 170.81 19.845 171.02 19.915 ;
    RECT 170.81 20.205 171.02 20.275 ;
    RECT 171.27 19.485 171.48 19.555 ;
    RECT 171.27 19.845 171.48 19.915 ;
    RECT 171.27 20.205 171.48 20.275 ;
    RECT 167.49 19.485 167.7 19.555 ;
    RECT 167.49 19.845 167.7 19.915 ;
    RECT 167.49 20.205 167.7 20.275 ;
    RECT 167.95 19.485 168.16 19.555 ;
    RECT 167.95 19.845 168.16 19.915 ;
    RECT 167.95 20.205 168.16 20.275 ;
    RECT 97.77 19.485 97.98 19.555 ;
    RECT 97.77 19.845 97.98 19.915 ;
    RECT 97.77 20.205 97.98 20.275 ;
    RECT 98.23 19.485 98.44 19.555 ;
    RECT 98.23 19.845 98.44 19.915 ;
    RECT 98.23 20.205 98.44 20.275 ;
    RECT 94.45 19.485 94.66 19.555 ;
    RECT 94.45 19.845 94.66 19.915 ;
    RECT 94.45 20.205 94.66 20.275 ;
    RECT 94.91 19.485 95.12 19.555 ;
    RECT 94.91 19.845 95.12 19.915 ;
    RECT 94.91 20.205 95.12 20.275 ;
    RECT 91.13 19.485 91.34 19.555 ;
    RECT 91.13 19.845 91.34 19.915 ;
    RECT 91.13 20.205 91.34 20.275 ;
    RECT 91.59 19.485 91.8 19.555 ;
    RECT 91.59 19.845 91.8 19.915 ;
    RECT 91.59 20.205 91.8 20.275 ;
    RECT 87.81 19.485 88.02 19.555 ;
    RECT 87.81 19.845 88.02 19.915 ;
    RECT 87.81 20.205 88.02 20.275 ;
    RECT 88.27 19.485 88.48 19.555 ;
    RECT 88.27 19.845 88.48 19.915 ;
    RECT 88.27 20.205 88.48 20.275 ;
    RECT 84.49 19.485 84.7 19.555 ;
    RECT 84.49 19.845 84.7 19.915 ;
    RECT 84.49 20.205 84.7 20.275 ;
    RECT 84.95 19.485 85.16 19.555 ;
    RECT 84.95 19.845 85.16 19.915 ;
    RECT 84.95 20.205 85.16 20.275 ;
    RECT 81.17 19.485 81.38 19.555 ;
    RECT 81.17 19.845 81.38 19.915 ;
    RECT 81.17 20.205 81.38 20.275 ;
    RECT 81.63 19.485 81.84 19.555 ;
    RECT 81.63 19.845 81.84 19.915 ;
    RECT 81.63 20.205 81.84 20.275 ;
    RECT 77.85 19.485 78.06 19.555 ;
    RECT 77.85 19.845 78.06 19.915 ;
    RECT 77.85 20.205 78.06 20.275 ;
    RECT 78.31 19.485 78.52 19.555 ;
    RECT 78.31 19.845 78.52 19.915 ;
    RECT 78.31 20.205 78.52 20.275 ;
    RECT 74.53 19.485 74.74 19.555 ;
    RECT 74.53 19.845 74.74 19.915 ;
    RECT 74.53 20.205 74.74 20.275 ;
    RECT 74.99 19.485 75.2 19.555 ;
    RECT 74.99 19.845 75.2 19.915 ;
    RECT 74.99 20.205 75.2 20.275 ;
    RECT 71.21 19.485 71.42 19.555 ;
    RECT 71.21 19.845 71.42 19.915 ;
    RECT 71.21 20.205 71.42 20.275 ;
    RECT 71.67 19.485 71.88 19.555 ;
    RECT 71.67 19.845 71.88 19.915 ;
    RECT 71.67 20.205 71.88 20.275 ;
    RECT 31.37 19.485 31.58 19.555 ;
    RECT 31.37 19.845 31.58 19.915 ;
    RECT 31.37 20.205 31.58 20.275 ;
    RECT 31.83 19.485 32.04 19.555 ;
    RECT 31.83 19.845 32.04 19.915 ;
    RECT 31.83 20.205 32.04 20.275 ;
    RECT 67.89 19.485 68.1 19.555 ;
    RECT 67.89 19.845 68.1 19.915 ;
    RECT 67.89 20.205 68.1 20.275 ;
    RECT 68.35 19.485 68.56 19.555 ;
    RECT 68.35 19.845 68.56 19.915 ;
    RECT 68.35 20.205 68.56 20.275 ;
    RECT 28.05 19.485 28.26 19.555 ;
    RECT 28.05 19.845 28.26 19.915 ;
    RECT 28.05 20.205 28.26 20.275 ;
    RECT 28.51 19.485 28.72 19.555 ;
    RECT 28.51 19.845 28.72 19.915 ;
    RECT 28.51 20.205 28.72 20.275 ;
    RECT 24.73 19.485 24.94 19.555 ;
    RECT 24.73 19.845 24.94 19.915 ;
    RECT 24.73 20.205 24.94 20.275 ;
    RECT 25.19 19.485 25.4 19.555 ;
    RECT 25.19 19.845 25.4 19.915 ;
    RECT 25.19 20.205 25.4 20.275 ;
    RECT 21.41 19.485 21.62 19.555 ;
    RECT 21.41 19.845 21.62 19.915 ;
    RECT 21.41 20.205 21.62 20.275 ;
    RECT 21.87 19.485 22.08 19.555 ;
    RECT 21.87 19.845 22.08 19.915 ;
    RECT 21.87 20.205 22.08 20.275 ;
    RECT 18.09 19.485 18.3 19.555 ;
    RECT 18.09 19.845 18.3 19.915 ;
    RECT 18.09 20.205 18.3 20.275 ;
    RECT 18.55 19.485 18.76 19.555 ;
    RECT 18.55 19.845 18.76 19.915 ;
    RECT 18.55 20.205 18.76 20.275 ;
    RECT 14.77 19.485 14.98 19.555 ;
    RECT 14.77 19.845 14.98 19.915 ;
    RECT 14.77 20.205 14.98 20.275 ;
    RECT 15.23 19.485 15.44 19.555 ;
    RECT 15.23 19.845 15.44 19.915 ;
    RECT 15.23 20.205 15.44 20.275 ;
    RECT 11.45 19.485 11.66 19.555 ;
    RECT 11.45 19.845 11.66 19.915 ;
    RECT 11.45 20.205 11.66 20.275 ;
    RECT 11.91 19.485 12.12 19.555 ;
    RECT 11.91 19.845 12.12 19.915 ;
    RECT 11.91 20.205 12.12 20.275 ;
    RECT 8.13 19.485 8.34 19.555 ;
    RECT 8.13 19.845 8.34 19.915 ;
    RECT 8.13 20.205 8.34 20.275 ;
    RECT 8.59 19.485 8.8 19.555 ;
    RECT 8.59 19.845 8.8 19.915 ;
    RECT 8.59 20.205 8.8 20.275 ;
    RECT 4.81 19.485 5.02 19.555 ;
    RECT 4.81 19.845 5.02 19.915 ;
    RECT 4.81 20.205 5.02 20.275 ;
    RECT 5.27 19.485 5.48 19.555 ;
    RECT 5.27 19.845 5.48 19.915 ;
    RECT 5.27 20.205 5.48 20.275 ;
    RECT 164.17 19.485 164.38 19.555 ;
    RECT 164.17 19.845 164.38 19.915 ;
    RECT 164.17 20.205 164.38 20.275 ;
    RECT 164.63 19.485 164.84 19.555 ;
    RECT 164.63 19.845 164.84 19.915 ;
    RECT 164.63 20.205 164.84 20.275 ;
    RECT 1.49 19.485 1.7 19.555 ;
    RECT 1.49 19.845 1.7 19.915 ;
    RECT 1.49 20.205 1.7 20.275 ;
    RECT 1.95 19.485 2.16 19.555 ;
    RECT 1.95 19.845 2.16 19.915 ;
    RECT 1.95 20.205 2.16 20.275 ;
    RECT 160.85 19.485 161.06 19.555 ;
    RECT 160.85 19.845 161.06 19.915 ;
    RECT 160.85 20.205 161.06 20.275 ;
    RECT 161.31 19.485 161.52 19.555 ;
    RECT 161.31 19.845 161.52 19.915 ;
    RECT 161.31 20.205 161.52 20.275 ;
    RECT 157.53 19.485 157.74 19.555 ;
    RECT 157.53 19.845 157.74 19.915 ;
    RECT 157.53 20.205 157.74 20.275 ;
    RECT 157.99 19.485 158.2 19.555 ;
    RECT 157.99 19.845 158.2 19.915 ;
    RECT 157.99 20.205 158.2 20.275 ;
    RECT 154.21 19.485 154.42 19.555 ;
    RECT 154.21 19.845 154.42 19.915 ;
    RECT 154.21 20.205 154.42 20.275 ;
    RECT 154.67 19.485 154.88 19.555 ;
    RECT 154.67 19.845 154.88 19.915 ;
    RECT 154.67 20.205 154.88 20.275 ;
    RECT 150.89 19.485 151.1 19.555 ;
    RECT 150.89 19.845 151.1 19.915 ;
    RECT 150.89 20.205 151.1 20.275 ;
    RECT 151.35 19.485 151.56 19.555 ;
    RECT 151.35 19.845 151.56 19.915 ;
    RECT 151.35 20.205 151.56 20.275 ;
    RECT 147.57 19.485 147.78 19.555 ;
    RECT 147.57 19.845 147.78 19.915 ;
    RECT 147.57 20.205 147.78 20.275 ;
    RECT 148.03 19.485 148.24 19.555 ;
    RECT 148.03 19.845 148.24 19.915 ;
    RECT 148.03 20.205 148.24 20.275 ;
    RECT 144.25 19.485 144.46 19.555 ;
    RECT 144.25 19.845 144.46 19.915 ;
    RECT 144.25 20.205 144.46 20.275 ;
    RECT 144.71 19.485 144.92 19.555 ;
    RECT 144.71 19.845 144.92 19.915 ;
    RECT 144.71 20.205 144.92 20.275 ;
    RECT 140.93 19.485 141.14 19.555 ;
    RECT 140.93 19.845 141.14 19.915 ;
    RECT 140.93 20.205 141.14 20.275 ;
    RECT 141.39 19.485 141.6 19.555 ;
    RECT 141.39 19.845 141.6 19.915 ;
    RECT 141.39 20.205 141.6 20.275 ;
    RECT 137.61 19.485 137.82 19.555 ;
    RECT 137.61 19.845 137.82 19.915 ;
    RECT 137.61 20.205 137.82 20.275 ;
    RECT 138.07 19.485 138.28 19.555 ;
    RECT 138.07 19.845 138.28 19.915 ;
    RECT 138.07 20.205 138.28 20.275 ;
    RECT 134.29 19.485 134.5 19.555 ;
    RECT 134.29 19.845 134.5 19.915 ;
    RECT 134.29 20.205 134.5 20.275 ;
    RECT 134.75 19.485 134.96 19.555 ;
    RECT 134.75 19.845 134.96 19.915 ;
    RECT 134.75 20.205 134.96 20.275 ;
    RECT 64.57 19.485 64.78 19.555 ;
    RECT 64.57 19.845 64.78 19.915 ;
    RECT 64.57 20.205 64.78 20.275 ;
    RECT 65.03 19.485 65.24 19.555 ;
    RECT 65.03 19.845 65.24 19.915 ;
    RECT 65.03 20.205 65.24 20.275 ;
    RECT 61.25 18.765 61.46 18.835 ;
    RECT 61.25 19.125 61.46 19.195 ;
    RECT 61.25 19.485 61.46 19.555 ;
    RECT 61.71 18.765 61.92 18.835 ;
    RECT 61.71 19.125 61.92 19.195 ;
    RECT 61.71 19.485 61.92 19.555 ;
    RECT 57.93 18.765 58.14 18.835 ;
    RECT 57.93 19.125 58.14 19.195 ;
    RECT 57.93 19.485 58.14 19.555 ;
    RECT 58.39 18.765 58.6 18.835 ;
    RECT 58.39 19.125 58.6 19.195 ;
    RECT 58.39 19.485 58.6 19.555 ;
    RECT 54.61 18.765 54.82 18.835 ;
    RECT 54.61 19.125 54.82 19.195 ;
    RECT 54.61 19.485 54.82 19.555 ;
    RECT 55.07 18.765 55.28 18.835 ;
    RECT 55.07 19.125 55.28 19.195 ;
    RECT 55.07 19.485 55.28 19.555 ;
    RECT 51.29 18.765 51.5 18.835 ;
    RECT 51.29 19.125 51.5 19.195 ;
    RECT 51.29 19.485 51.5 19.555 ;
    RECT 51.75 18.765 51.96 18.835 ;
    RECT 51.75 19.125 51.96 19.195 ;
    RECT 51.75 19.485 51.96 19.555 ;
    RECT 47.97 18.765 48.18 18.835 ;
    RECT 47.97 19.125 48.18 19.195 ;
    RECT 47.97 19.485 48.18 19.555 ;
    RECT 48.43 18.765 48.64 18.835 ;
    RECT 48.43 19.125 48.64 19.195 ;
    RECT 48.43 19.485 48.64 19.555 ;
    RECT 44.65 18.765 44.86 18.835 ;
    RECT 44.65 19.125 44.86 19.195 ;
    RECT 44.65 19.485 44.86 19.555 ;
    RECT 45.11 18.765 45.32 18.835 ;
    RECT 45.11 19.125 45.32 19.195 ;
    RECT 45.11 19.485 45.32 19.555 ;
    RECT 41.33 18.765 41.54 18.835 ;
    RECT 41.33 19.125 41.54 19.195 ;
    RECT 41.33 19.485 41.54 19.555 ;
    RECT 41.79 18.765 42.0 18.835 ;
    RECT 41.79 19.125 42.0 19.195 ;
    RECT 41.79 19.485 42.0 19.555 ;
    RECT 38.01 18.765 38.22 18.835 ;
    RECT 38.01 19.125 38.22 19.195 ;
    RECT 38.01 19.485 38.22 19.555 ;
    RECT 38.47 18.765 38.68 18.835 ;
    RECT 38.47 19.125 38.68 19.195 ;
    RECT 38.47 19.485 38.68 19.555 ;
    RECT 34.69 18.765 34.9 18.835 ;
    RECT 34.69 19.125 34.9 19.195 ;
    RECT 34.69 19.485 34.9 19.555 ;
    RECT 35.15 18.765 35.36 18.835 ;
    RECT 35.15 19.125 35.36 19.195 ;
    RECT 35.15 19.485 35.36 19.555 ;
    RECT 173.945 19.125 174.015 19.195 ;
    RECT 130.97 18.765 131.18 18.835 ;
    RECT 130.97 19.125 131.18 19.195 ;
    RECT 130.97 19.485 131.18 19.555 ;
    RECT 131.43 18.765 131.64 18.835 ;
    RECT 131.43 19.125 131.64 19.195 ;
    RECT 131.43 19.485 131.64 19.555 ;
    RECT 127.65 18.765 127.86 18.835 ;
    RECT 127.65 19.125 127.86 19.195 ;
    RECT 127.65 19.485 127.86 19.555 ;
    RECT 128.11 18.765 128.32 18.835 ;
    RECT 128.11 19.125 128.32 19.195 ;
    RECT 128.11 19.485 128.32 19.555 ;
    RECT 124.33 18.765 124.54 18.835 ;
    RECT 124.33 19.125 124.54 19.195 ;
    RECT 124.33 19.485 124.54 19.555 ;
    RECT 124.79 18.765 125.0 18.835 ;
    RECT 124.79 19.125 125.0 19.195 ;
    RECT 124.79 19.485 125.0 19.555 ;
    RECT 121.01 18.765 121.22 18.835 ;
    RECT 121.01 19.125 121.22 19.195 ;
    RECT 121.01 19.485 121.22 19.555 ;
    RECT 121.47 18.765 121.68 18.835 ;
    RECT 121.47 19.125 121.68 19.195 ;
    RECT 121.47 19.485 121.68 19.555 ;
    RECT 117.69 18.765 117.9 18.835 ;
    RECT 117.69 19.125 117.9 19.195 ;
    RECT 117.69 19.485 117.9 19.555 ;
    RECT 118.15 18.765 118.36 18.835 ;
    RECT 118.15 19.125 118.36 19.195 ;
    RECT 118.15 19.485 118.36 19.555 ;
    RECT 114.37 18.765 114.58 18.835 ;
    RECT 114.37 19.125 114.58 19.195 ;
    RECT 114.37 19.485 114.58 19.555 ;
    RECT 114.83 18.765 115.04 18.835 ;
    RECT 114.83 19.125 115.04 19.195 ;
    RECT 114.83 19.485 115.04 19.555 ;
    RECT 111.05 18.765 111.26 18.835 ;
    RECT 111.05 19.125 111.26 19.195 ;
    RECT 111.05 19.485 111.26 19.555 ;
    RECT 111.51 18.765 111.72 18.835 ;
    RECT 111.51 19.125 111.72 19.195 ;
    RECT 111.51 19.485 111.72 19.555 ;
    RECT 107.73 18.765 107.94 18.835 ;
    RECT 107.73 19.125 107.94 19.195 ;
    RECT 107.73 19.485 107.94 19.555 ;
    RECT 108.19 18.765 108.4 18.835 ;
    RECT 108.19 19.125 108.4 19.195 ;
    RECT 108.19 19.485 108.4 19.555 ;
    RECT 104.41 18.765 104.62 18.835 ;
    RECT 104.41 19.125 104.62 19.195 ;
    RECT 104.41 19.485 104.62 19.555 ;
    RECT 104.87 18.765 105.08 18.835 ;
    RECT 104.87 19.125 105.08 19.195 ;
    RECT 104.87 19.485 105.08 19.555 ;
    RECT 101.09 18.765 101.3 18.835 ;
    RECT 101.09 19.125 101.3 19.195 ;
    RECT 101.09 19.485 101.3 19.555 ;
    RECT 101.55 18.765 101.76 18.835 ;
    RECT 101.55 19.125 101.76 19.195 ;
    RECT 101.55 19.485 101.76 19.555 ;
    RECT 0.4 19.125 0.47 19.195 ;
    RECT 170.81 18.765 171.02 18.835 ;
    RECT 170.81 19.125 171.02 19.195 ;
    RECT 170.81 19.485 171.02 19.555 ;
    RECT 171.27 18.765 171.48 18.835 ;
    RECT 171.27 19.125 171.48 19.195 ;
    RECT 171.27 19.485 171.48 19.555 ;
    RECT 167.49 18.765 167.7 18.835 ;
    RECT 167.49 19.125 167.7 19.195 ;
    RECT 167.49 19.485 167.7 19.555 ;
    RECT 167.95 18.765 168.16 18.835 ;
    RECT 167.95 19.125 168.16 19.195 ;
    RECT 167.95 19.485 168.16 19.555 ;
    RECT 97.77 18.765 97.98 18.835 ;
    RECT 97.77 19.125 97.98 19.195 ;
    RECT 97.77 19.485 97.98 19.555 ;
    RECT 98.23 18.765 98.44 18.835 ;
    RECT 98.23 19.125 98.44 19.195 ;
    RECT 98.23 19.485 98.44 19.555 ;
    RECT 94.45 18.765 94.66 18.835 ;
    RECT 94.45 19.125 94.66 19.195 ;
    RECT 94.45 19.485 94.66 19.555 ;
    RECT 94.91 18.765 95.12 18.835 ;
    RECT 94.91 19.125 95.12 19.195 ;
    RECT 94.91 19.485 95.12 19.555 ;
    RECT 91.13 18.765 91.34 18.835 ;
    RECT 91.13 19.125 91.34 19.195 ;
    RECT 91.13 19.485 91.34 19.555 ;
    RECT 91.59 18.765 91.8 18.835 ;
    RECT 91.59 19.125 91.8 19.195 ;
    RECT 91.59 19.485 91.8 19.555 ;
    RECT 87.81 18.765 88.02 18.835 ;
    RECT 87.81 19.125 88.02 19.195 ;
    RECT 87.81 19.485 88.02 19.555 ;
    RECT 88.27 18.765 88.48 18.835 ;
    RECT 88.27 19.125 88.48 19.195 ;
    RECT 88.27 19.485 88.48 19.555 ;
    RECT 84.49 18.765 84.7 18.835 ;
    RECT 84.49 19.125 84.7 19.195 ;
    RECT 84.49 19.485 84.7 19.555 ;
    RECT 84.95 18.765 85.16 18.835 ;
    RECT 84.95 19.125 85.16 19.195 ;
    RECT 84.95 19.485 85.16 19.555 ;
    RECT 81.17 18.765 81.38 18.835 ;
    RECT 81.17 19.125 81.38 19.195 ;
    RECT 81.17 19.485 81.38 19.555 ;
    RECT 81.63 18.765 81.84 18.835 ;
    RECT 81.63 19.125 81.84 19.195 ;
    RECT 81.63 19.485 81.84 19.555 ;
    RECT 77.85 18.765 78.06 18.835 ;
    RECT 77.85 19.125 78.06 19.195 ;
    RECT 77.85 19.485 78.06 19.555 ;
    RECT 78.31 18.765 78.52 18.835 ;
    RECT 78.31 19.125 78.52 19.195 ;
    RECT 78.31 19.485 78.52 19.555 ;
    RECT 74.53 18.765 74.74 18.835 ;
    RECT 74.53 19.125 74.74 19.195 ;
    RECT 74.53 19.485 74.74 19.555 ;
    RECT 74.99 18.765 75.2 18.835 ;
    RECT 74.99 19.125 75.2 19.195 ;
    RECT 74.99 19.485 75.2 19.555 ;
    RECT 71.21 18.765 71.42 18.835 ;
    RECT 71.21 19.125 71.42 19.195 ;
    RECT 71.21 19.485 71.42 19.555 ;
    RECT 71.67 18.765 71.88 18.835 ;
    RECT 71.67 19.125 71.88 19.195 ;
    RECT 71.67 19.485 71.88 19.555 ;
    RECT 31.37 18.765 31.58 18.835 ;
    RECT 31.37 19.125 31.58 19.195 ;
    RECT 31.37 19.485 31.58 19.555 ;
    RECT 31.83 18.765 32.04 18.835 ;
    RECT 31.83 19.125 32.04 19.195 ;
    RECT 31.83 19.485 32.04 19.555 ;
    RECT 67.89 18.765 68.1 18.835 ;
    RECT 67.89 19.125 68.1 19.195 ;
    RECT 67.89 19.485 68.1 19.555 ;
    RECT 68.35 18.765 68.56 18.835 ;
    RECT 68.35 19.125 68.56 19.195 ;
    RECT 68.35 19.485 68.56 19.555 ;
    RECT 28.05 18.765 28.26 18.835 ;
    RECT 28.05 19.125 28.26 19.195 ;
    RECT 28.05 19.485 28.26 19.555 ;
    RECT 28.51 18.765 28.72 18.835 ;
    RECT 28.51 19.125 28.72 19.195 ;
    RECT 28.51 19.485 28.72 19.555 ;
    RECT 24.73 18.765 24.94 18.835 ;
    RECT 24.73 19.125 24.94 19.195 ;
    RECT 24.73 19.485 24.94 19.555 ;
    RECT 25.19 18.765 25.4 18.835 ;
    RECT 25.19 19.125 25.4 19.195 ;
    RECT 25.19 19.485 25.4 19.555 ;
    RECT 21.41 18.765 21.62 18.835 ;
    RECT 21.41 19.125 21.62 19.195 ;
    RECT 21.41 19.485 21.62 19.555 ;
    RECT 21.87 18.765 22.08 18.835 ;
    RECT 21.87 19.125 22.08 19.195 ;
    RECT 21.87 19.485 22.08 19.555 ;
    RECT 18.09 18.765 18.3 18.835 ;
    RECT 18.09 19.125 18.3 19.195 ;
    RECT 18.09 19.485 18.3 19.555 ;
    RECT 18.55 18.765 18.76 18.835 ;
    RECT 18.55 19.125 18.76 19.195 ;
    RECT 18.55 19.485 18.76 19.555 ;
    RECT 14.77 18.765 14.98 18.835 ;
    RECT 14.77 19.125 14.98 19.195 ;
    RECT 14.77 19.485 14.98 19.555 ;
    RECT 15.23 18.765 15.44 18.835 ;
    RECT 15.23 19.125 15.44 19.195 ;
    RECT 15.23 19.485 15.44 19.555 ;
    RECT 11.45 18.765 11.66 18.835 ;
    RECT 11.45 19.125 11.66 19.195 ;
    RECT 11.45 19.485 11.66 19.555 ;
    RECT 11.91 18.765 12.12 18.835 ;
    RECT 11.91 19.125 12.12 19.195 ;
    RECT 11.91 19.485 12.12 19.555 ;
    RECT 8.13 18.765 8.34 18.835 ;
    RECT 8.13 19.125 8.34 19.195 ;
    RECT 8.13 19.485 8.34 19.555 ;
    RECT 8.59 18.765 8.8 18.835 ;
    RECT 8.59 19.125 8.8 19.195 ;
    RECT 8.59 19.485 8.8 19.555 ;
    RECT 4.81 18.765 5.02 18.835 ;
    RECT 4.81 19.125 5.02 19.195 ;
    RECT 4.81 19.485 5.02 19.555 ;
    RECT 5.27 18.765 5.48 18.835 ;
    RECT 5.27 19.125 5.48 19.195 ;
    RECT 5.27 19.485 5.48 19.555 ;
    RECT 164.17 18.765 164.38 18.835 ;
    RECT 164.17 19.125 164.38 19.195 ;
    RECT 164.17 19.485 164.38 19.555 ;
    RECT 164.63 18.765 164.84 18.835 ;
    RECT 164.63 19.125 164.84 19.195 ;
    RECT 164.63 19.485 164.84 19.555 ;
    RECT 1.49 18.765 1.7 18.835 ;
    RECT 1.49 19.125 1.7 19.195 ;
    RECT 1.49 19.485 1.7 19.555 ;
    RECT 1.95 18.765 2.16 18.835 ;
    RECT 1.95 19.125 2.16 19.195 ;
    RECT 1.95 19.485 2.16 19.555 ;
    RECT 160.85 18.765 161.06 18.835 ;
    RECT 160.85 19.125 161.06 19.195 ;
    RECT 160.85 19.485 161.06 19.555 ;
    RECT 161.31 18.765 161.52 18.835 ;
    RECT 161.31 19.125 161.52 19.195 ;
    RECT 161.31 19.485 161.52 19.555 ;
    RECT 157.53 18.765 157.74 18.835 ;
    RECT 157.53 19.125 157.74 19.195 ;
    RECT 157.53 19.485 157.74 19.555 ;
    RECT 157.99 18.765 158.2 18.835 ;
    RECT 157.99 19.125 158.2 19.195 ;
    RECT 157.99 19.485 158.2 19.555 ;
    RECT 154.21 18.765 154.42 18.835 ;
    RECT 154.21 19.125 154.42 19.195 ;
    RECT 154.21 19.485 154.42 19.555 ;
    RECT 154.67 18.765 154.88 18.835 ;
    RECT 154.67 19.125 154.88 19.195 ;
    RECT 154.67 19.485 154.88 19.555 ;
    RECT 150.89 18.765 151.1 18.835 ;
    RECT 150.89 19.125 151.1 19.195 ;
    RECT 150.89 19.485 151.1 19.555 ;
    RECT 151.35 18.765 151.56 18.835 ;
    RECT 151.35 19.125 151.56 19.195 ;
    RECT 151.35 19.485 151.56 19.555 ;
    RECT 147.57 18.765 147.78 18.835 ;
    RECT 147.57 19.125 147.78 19.195 ;
    RECT 147.57 19.485 147.78 19.555 ;
    RECT 148.03 18.765 148.24 18.835 ;
    RECT 148.03 19.125 148.24 19.195 ;
    RECT 148.03 19.485 148.24 19.555 ;
    RECT 144.25 18.765 144.46 18.835 ;
    RECT 144.25 19.125 144.46 19.195 ;
    RECT 144.25 19.485 144.46 19.555 ;
    RECT 144.71 18.765 144.92 18.835 ;
    RECT 144.71 19.125 144.92 19.195 ;
    RECT 144.71 19.485 144.92 19.555 ;
    RECT 140.93 18.765 141.14 18.835 ;
    RECT 140.93 19.125 141.14 19.195 ;
    RECT 140.93 19.485 141.14 19.555 ;
    RECT 141.39 18.765 141.6 18.835 ;
    RECT 141.39 19.125 141.6 19.195 ;
    RECT 141.39 19.485 141.6 19.555 ;
    RECT 137.61 18.765 137.82 18.835 ;
    RECT 137.61 19.125 137.82 19.195 ;
    RECT 137.61 19.485 137.82 19.555 ;
    RECT 138.07 18.765 138.28 18.835 ;
    RECT 138.07 19.125 138.28 19.195 ;
    RECT 138.07 19.485 138.28 19.555 ;
    RECT 134.29 18.765 134.5 18.835 ;
    RECT 134.29 19.125 134.5 19.195 ;
    RECT 134.29 19.485 134.5 19.555 ;
    RECT 134.75 18.765 134.96 18.835 ;
    RECT 134.75 19.125 134.96 19.195 ;
    RECT 134.75 19.485 134.96 19.555 ;
    RECT 64.57 18.765 64.78 18.835 ;
    RECT 64.57 19.125 64.78 19.195 ;
    RECT 64.57 19.485 64.78 19.555 ;
    RECT 65.03 18.765 65.24 18.835 ;
    RECT 65.03 19.125 65.24 19.195 ;
    RECT 65.03 19.485 65.24 19.555 ;
    RECT 61.71 58.145 61.92 58.215 ;
    RECT 65.52 57.885 65.73 57.955 ;
    RECT 61.25 58.145 61.46 58.215 ;
    RECT 131.43 58.145 131.64 58.215 ;
    RECT 130.97 58.145 131.18 58.215 ;
    RECT 84.95 58.145 85.16 58.215 ;
    RECT 84.49 58.145 84.7 58.215 ;
    RECT 154.67 58.145 154.88 58.215 ;
    RECT 154.21 58.145 154.42 58.215 ;
    RECT 131.92 57.885 132.13 57.955 ;
    RECT 151.84 57.885 152.05 57.955 ;
    RECT 1.95 58.145 2.16 58.215 ;
    RECT 1.49 58.145 1.7 58.215 ;
    RECT 24.73 58.145 24.94 58.215 ;
    RECT 38.47 58.145 38.68 58.215 ;
    RECT 121.47 58.145 121.68 58.215 ;
    RECT 167.95 58.145 168.16 58.215 ;
    RECT 38.01 58.145 38.22 58.215 ;
    RECT 121.01 58.145 121.22 58.215 ;
    RECT 167.49 58.145 167.7 58.215 ;
    RECT 35.64 57.885 35.85 57.955 ;
    RECT 5.76 57.885 5.97 57.955 ;
    RECT 88.76 57.885 88.97 57.955 ;
    RECT 102.04 57.885 102.25 57.955 ;
    RECT 58.88 57.885 59.09 57.955 ;
    RECT 29.0 57.885 29.21 57.955 ;
    RECT 124.79 58.145 125.0 58.215 ;
    RECT 78.31 58.145 78.52 58.215 ;
    RECT 125.28 57.885 125.49 57.955 ;
    RECT 145.2 57.885 145.41 57.955 ;
    RECT 77.85 58.145 78.06 58.215 ;
    RECT 148.03 58.145 148.24 58.215 ;
    RECT 147.57 58.145 147.78 58.215 ;
    RECT 18.55 58.145 18.76 58.215 ;
    RECT 18.09 58.145 18.3 58.215 ;
    RECT 168.44 57.885 168.65 57.955 ;
    RECT 114.83 58.145 115.04 58.215 ;
    RECT 114.37 58.145 114.58 58.215 ;
    RECT 55.07 58.145 55.28 58.215 ;
    RECT 54.61 58.145 54.82 58.215 ;
    RECT 82.12 57.885 82.33 57.955 ;
    RECT 72.16 57.885 72.37 57.955 ;
    RECT 138.56 57.885 138.77 57.955 ;
    RECT 94.91 58.145 95.12 58.215 ;
    RECT 141.39 58.145 141.6 58.215 ;
    RECT 94.45 58.145 94.66 58.215 ;
    RECT 164.63 58.145 164.84 58.215 ;
    RECT 164.17 58.145 164.38 58.215 ;
    RECT 11.91 58.145 12.12 58.215 ;
    RECT 11.45 58.145 11.66 58.215 ;
    RECT 161.8 57.885 162.01 57.955 ;
    RECT 174.155 57.885 174.225 57.955 ;
    RECT 173.945 58.145 174.015 58.215 ;
    RECT 52.24 57.885 52.45 57.955 ;
    RECT 22.36 57.885 22.57 57.955 ;
    RECT 108.19 58.145 108.4 58.215 ;
    RECT 0.19 57.885 0.26 57.955 ;
    RECT 0.4 58.145 0.47 58.215 ;
    RECT 48.43 58.145 48.64 58.215 ;
    RECT 47.97 58.145 48.18 58.215 ;
    RECT 98.72 57.885 98.93 57.955 ;
    RECT 118.64 57.885 118.85 57.955 ;
    RECT 71.67 58.145 71.88 58.215 ;
    RECT 71.21 58.145 71.42 58.215 ;
    RECT 140.93 58.145 141.14 58.215 ;
    RECT 107.73 58.145 107.94 58.215 ;
    RECT 157.99 58.145 158.2 58.215 ;
    RECT 28.51 58.145 28.72 58.215 ;
    RECT 28.05 58.145 28.26 58.215 ;
    RECT 45.6 57.885 45.81 57.955 ;
    RECT 15.72 57.885 15.93 57.955 ;
    RECT 41.79 58.145 42.0 58.215 ;
    RECT 112.0 57.885 112.21 57.955 ;
    RECT 65.03 58.145 65.24 58.215 ;
    RECT 92.08 57.885 92.29 57.955 ;
    RECT 64.57 58.145 64.78 58.215 ;
    RECT 88.27 58.145 88.48 58.215 ;
    RECT 134.75 58.145 134.96 58.215 ;
    RECT 87.81 58.145 88.02 58.215 ;
    RECT 134.29 58.145 134.5 58.215 ;
    RECT 157.53 58.145 157.74 58.215 ;
    RECT 155.16 57.885 155.37 57.955 ;
    RECT 5.27 58.145 5.48 58.215 ;
    RECT 4.81 58.145 5.02 58.215 ;
    RECT 101.55 58.145 101.76 58.215 ;
    RECT 101.09 58.145 101.3 58.215 ;
    RECT 171.27 58.145 171.48 58.215 ;
    RECT 41.33 58.145 41.54 58.215 ;
    RECT 124.33 58.145 124.54 58.215 ;
    RECT 170.81 58.145 171.02 58.215 ;
    RECT 38.96 57.885 39.17 57.955 ;
    RECT 9.08 57.885 9.29 57.955 ;
    RECT 105.36 57.885 105.57 57.955 ;
    RECT 62.2 57.885 62.41 57.955 ;
    RECT 32.32 57.885 32.53 57.955 ;
    RECT 58.39 58.145 58.6 58.215 ;
    RECT 128.11 58.145 128.32 58.215 ;
    RECT 127.65 58.145 127.86 58.215 ;
    RECT 81.63 58.145 81.84 58.215 ;
    RECT 81.17 58.145 81.38 58.215 ;
    RECT 128.6 57.885 128.81 57.955 ;
    RECT 148.52 57.885 148.73 57.955 ;
    RECT 151.35 58.145 151.56 58.215 ;
    RECT 150.89 58.145 151.1 58.215 ;
    RECT 21.87 58.145 22.08 58.215 ;
    RECT 21.41 58.145 21.62 58.215 ;
    RECT 35.15 58.145 35.36 58.215 ;
    RECT 118.15 58.145 118.36 58.215 ;
    RECT 171.76 57.885 171.97 57.955 ;
    RECT 34.69 58.145 34.9 58.215 ;
    RECT 117.69 58.145 117.9 58.215 ;
    RECT 57.93 58.145 58.14 58.215 ;
    RECT 2.44 57.885 2.65 57.955 ;
    RECT 85.44 57.885 85.65 57.955 ;
    RECT 75.48 57.885 75.69 57.955 ;
    RECT 25.68 57.885 25.89 57.955 ;
    RECT 141.88 57.885 142.09 57.955 ;
    RECT 74.99 58.145 75.2 58.215 ;
    RECT 98.23 58.145 98.44 58.215 ;
    RECT 144.71 58.145 144.92 58.215 ;
    RECT 97.77 58.145 97.98 58.215 ;
    RECT 144.25 58.145 144.46 58.215 ;
    RECT 15.23 58.145 15.44 58.215 ;
    RECT 14.77 58.145 14.98 58.215 ;
    RECT 165.12 57.885 165.33 57.955 ;
    RECT 55.56 57.885 55.77 57.955 ;
    RECT 111.51 58.145 111.72 58.215 ;
    RECT 111.05 58.145 111.26 58.215 ;
    RECT 51.75 58.145 51.96 58.215 ;
    RECT 51.29 58.145 51.5 58.215 ;
    RECT 121.96 57.885 122.17 57.955 ;
    RECT 74.53 58.145 74.74 58.215 ;
    RECT 78.8 57.885 79.01 57.955 ;
    RECT 68.84 57.885 69.05 57.955 ;
    RECT 135.24 57.885 135.45 57.955 ;
    RECT 91.59 58.145 91.8 58.215 ;
    RECT 161.31 58.145 161.52 58.215 ;
    RECT 160.85 58.145 161.06 58.215 ;
    RECT 8.59 58.145 8.8 58.215 ;
    RECT 158.48 57.885 158.69 57.955 ;
    RECT 31.83 58.145 32.04 58.215 ;
    RECT 31.37 58.145 31.58 58.215 ;
    RECT 48.92 57.885 49.13 57.955 ;
    RECT 19.04 57.885 19.25 57.955 ;
    RECT 45.11 58.145 45.32 58.215 ;
    RECT 44.65 58.145 44.86 58.215 ;
    RECT 95.4 57.885 95.61 57.955 ;
    RECT 115.32 57.885 115.53 57.955 ;
    RECT 68.35 58.145 68.56 58.215 ;
    RECT 67.89 58.145 68.1 58.215 ;
    RECT 138.07 58.145 138.28 58.215 ;
    RECT 91.13 58.145 91.34 58.215 ;
    RECT 137.61 58.145 137.82 58.215 ;
    RECT 8.13 58.145 8.34 58.215 ;
    RECT 104.87 58.145 105.08 58.215 ;
    RECT 104.41 58.145 104.62 58.215 ;
    RECT 25.19 58.145 25.4 58.215 ;
    RECT 42.28 57.885 42.49 57.955 ;
    RECT 12.4 57.885 12.61 57.955 ;
    RECT 108.68 57.885 108.89 57.955 ;
    RECT 61.25 56.925 61.46 56.995 ;
    RECT 61.25 57.285 61.46 57.355 ;
    RECT 61.25 57.645 61.46 57.715 ;
    RECT 61.71 56.925 61.92 56.995 ;
    RECT 61.71 57.285 61.92 57.355 ;
    RECT 61.71 57.645 61.92 57.715 ;
    RECT 57.93 56.925 58.14 56.995 ;
    RECT 57.93 57.285 58.14 57.355 ;
    RECT 57.93 57.645 58.14 57.715 ;
    RECT 58.39 56.925 58.6 56.995 ;
    RECT 58.39 57.285 58.6 57.355 ;
    RECT 58.39 57.645 58.6 57.715 ;
    RECT 54.61 56.925 54.82 56.995 ;
    RECT 54.61 57.285 54.82 57.355 ;
    RECT 54.61 57.645 54.82 57.715 ;
    RECT 55.07 56.925 55.28 56.995 ;
    RECT 55.07 57.285 55.28 57.355 ;
    RECT 55.07 57.645 55.28 57.715 ;
    RECT 51.29 56.925 51.5 56.995 ;
    RECT 51.29 57.285 51.5 57.355 ;
    RECT 51.29 57.645 51.5 57.715 ;
    RECT 51.75 56.925 51.96 56.995 ;
    RECT 51.75 57.285 51.96 57.355 ;
    RECT 51.75 57.645 51.96 57.715 ;
    RECT 47.97 56.925 48.18 56.995 ;
    RECT 47.97 57.285 48.18 57.355 ;
    RECT 47.97 57.645 48.18 57.715 ;
    RECT 48.43 56.925 48.64 56.995 ;
    RECT 48.43 57.285 48.64 57.355 ;
    RECT 48.43 57.645 48.64 57.715 ;
    RECT 44.65 56.925 44.86 56.995 ;
    RECT 44.65 57.285 44.86 57.355 ;
    RECT 44.65 57.645 44.86 57.715 ;
    RECT 45.11 56.925 45.32 56.995 ;
    RECT 45.11 57.285 45.32 57.355 ;
    RECT 45.11 57.645 45.32 57.715 ;
    RECT 41.33 56.925 41.54 56.995 ;
    RECT 41.33 57.285 41.54 57.355 ;
    RECT 41.33 57.645 41.54 57.715 ;
    RECT 41.79 56.925 42.0 56.995 ;
    RECT 41.79 57.285 42.0 57.355 ;
    RECT 41.79 57.645 42.0 57.715 ;
    RECT 38.01 56.925 38.22 56.995 ;
    RECT 38.01 57.285 38.22 57.355 ;
    RECT 38.01 57.645 38.22 57.715 ;
    RECT 38.47 56.925 38.68 56.995 ;
    RECT 38.47 57.285 38.68 57.355 ;
    RECT 38.47 57.645 38.68 57.715 ;
    RECT 34.69 56.925 34.9 56.995 ;
    RECT 34.69 57.285 34.9 57.355 ;
    RECT 34.69 57.645 34.9 57.715 ;
    RECT 35.15 56.925 35.36 56.995 ;
    RECT 35.15 57.285 35.36 57.355 ;
    RECT 35.15 57.645 35.36 57.715 ;
    RECT 173.945 57.285 174.015 57.355 ;
    RECT 130.97 56.925 131.18 56.995 ;
    RECT 130.97 57.285 131.18 57.355 ;
    RECT 130.97 57.645 131.18 57.715 ;
    RECT 131.43 56.925 131.64 56.995 ;
    RECT 131.43 57.285 131.64 57.355 ;
    RECT 131.43 57.645 131.64 57.715 ;
    RECT 127.65 56.925 127.86 56.995 ;
    RECT 127.65 57.285 127.86 57.355 ;
    RECT 127.65 57.645 127.86 57.715 ;
    RECT 128.11 56.925 128.32 56.995 ;
    RECT 128.11 57.285 128.32 57.355 ;
    RECT 128.11 57.645 128.32 57.715 ;
    RECT 124.33 56.925 124.54 56.995 ;
    RECT 124.33 57.285 124.54 57.355 ;
    RECT 124.33 57.645 124.54 57.715 ;
    RECT 124.79 56.925 125.0 56.995 ;
    RECT 124.79 57.285 125.0 57.355 ;
    RECT 124.79 57.645 125.0 57.715 ;
    RECT 121.01 56.925 121.22 56.995 ;
    RECT 121.01 57.285 121.22 57.355 ;
    RECT 121.01 57.645 121.22 57.715 ;
    RECT 121.47 56.925 121.68 56.995 ;
    RECT 121.47 57.285 121.68 57.355 ;
    RECT 121.47 57.645 121.68 57.715 ;
    RECT 117.69 56.925 117.9 56.995 ;
    RECT 117.69 57.285 117.9 57.355 ;
    RECT 117.69 57.645 117.9 57.715 ;
    RECT 118.15 56.925 118.36 56.995 ;
    RECT 118.15 57.285 118.36 57.355 ;
    RECT 118.15 57.645 118.36 57.715 ;
    RECT 114.37 56.925 114.58 56.995 ;
    RECT 114.37 57.285 114.58 57.355 ;
    RECT 114.37 57.645 114.58 57.715 ;
    RECT 114.83 56.925 115.04 56.995 ;
    RECT 114.83 57.285 115.04 57.355 ;
    RECT 114.83 57.645 115.04 57.715 ;
    RECT 111.05 56.925 111.26 56.995 ;
    RECT 111.05 57.285 111.26 57.355 ;
    RECT 111.05 57.645 111.26 57.715 ;
    RECT 111.51 56.925 111.72 56.995 ;
    RECT 111.51 57.285 111.72 57.355 ;
    RECT 111.51 57.645 111.72 57.715 ;
    RECT 107.73 56.925 107.94 56.995 ;
    RECT 107.73 57.285 107.94 57.355 ;
    RECT 107.73 57.645 107.94 57.715 ;
    RECT 108.19 56.925 108.4 56.995 ;
    RECT 108.19 57.285 108.4 57.355 ;
    RECT 108.19 57.645 108.4 57.715 ;
    RECT 104.41 56.925 104.62 56.995 ;
    RECT 104.41 57.285 104.62 57.355 ;
    RECT 104.41 57.645 104.62 57.715 ;
    RECT 104.87 56.925 105.08 56.995 ;
    RECT 104.87 57.285 105.08 57.355 ;
    RECT 104.87 57.645 105.08 57.715 ;
    RECT 101.09 56.925 101.3 56.995 ;
    RECT 101.09 57.285 101.3 57.355 ;
    RECT 101.09 57.645 101.3 57.715 ;
    RECT 101.55 56.925 101.76 56.995 ;
    RECT 101.55 57.285 101.76 57.355 ;
    RECT 101.55 57.645 101.76 57.715 ;
    RECT 0.4 57.285 0.47 57.355 ;
    RECT 170.81 56.925 171.02 56.995 ;
    RECT 170.81 57.285 171.02 57.355 ;
    RECT 170.81 57.645 171.02 57.715 ;
    RECT 171.27 56.925 171.48 56.995 ;
    RECT 171.27 57.285 171.48 57.355 ;
    RECT 171.27 57.645 171.48 57.715 ;
    RECT 167.49 56.925 167.7 56.995 ;
    RECT 167.49 57.285 167.7 57.355 ;
    RECT 167.49 57.645 167.7 57.715 ;
    RECT 167.95 56.925 168.16 56.995 ;
    RECT 167.95 57.285 168.16 57.355 ;
    RECT 167.95 57.645 168.16 57.715 ;
    RECT 97.77 56.925 97.98 56.995 ;
    RECT 97.77 57.285 97.98 57.355 ;
    RECT 97.77 57.645 97.98 57.715 ;
    RECT 98.23 56.925 98.44 56.995 ;
    RECT 98.23 57.285 98.44 57.355 ;
    RECT 98.23 57.645 98.44 57.715 ;
    RECT 94.45 56.925 94.66 56.995 ;
    RECT 94.45 57.285 94.66 57.355 ;
    RECT 94.45 57.645 94.66 57.715 ;
    RECT 94.91 56.925 95.12 56.995 ;
    RECT 94.91 57.285 95.12 57.355 ;
    RECT 94.91 57.645 95.12 57.715 ;
    RECT 91.13 56.925 91.34 56.995 ;
    RECT 91.13 57.285 91.34 57.355 ;
    RECT 91.13 57.645 91.34 57.715 ;
    RECT 91.59 56.925 91.8 56.995 ;
    RECT 91.59 57.285 91.8 57.355 ;
    RECT 91.59 57.645 91.8 57.715 ;
    RECT 87.81 56.925 88.02 56.995 ;
    RECT 87.81 57.285 88.02 57.355 ;
    RECT 87.81 57.645 88.02 57.715 ;
    RECT 88.27 56.925 88.48 56.995 ;
    RECT 88.27 57.285 88.48 57.355 ;
    RECT 88.27 57.645 88.48 57.715 ;
    RECT 84.49 56.925 84.7 56.995 ;
    RECT 84.49 57.285 84.7 57.355 ;
    RECT 84.49 57.645 84.7 57.715 ;
    RECT 84.95 56.925 85.16 56.995 ;
    RECT 84.95 57.285 85.16 57.355 ;
    RECT 84.95 57.645 85.16 57.715 ;
    RECT 81.17 56.925 81.38 56.995 ;
    RECT 81.17 57.285 81.38 57.355 ;
    RECT 81.17 57.645 81.38 57.715 ;
    RECT 81.63 56.925 81.84 56.995 ;
    RECT 81.63 57.285 81.84 57.355 ;
    RECT 81.63 57.645 81.84 57.715 ;
    RECT 77.85 56.925 78.06 56.995 ;
    RECT 77.85 57.285 78.06 57.355 ;
    RECT 77.85 57.645 78.06 57.715 ;
    RECT 78.31 56.925 78.52 56.995 ;
    RECT 78.31 57.285 78.52 57.355 ;
    RECT 78.31 57.645 78.52 57.715 ;
    RECT 74.53 56.925 74.74 56.995 ;
    RECT 74.53 57.285 74.74 57.355 ;
    RECT 74.53 57.645 74.74 57.715 ;
    RECT 74.99 56.925 75.2 56.995 ;
    RECT 74.99 57.285 75.2 57.355 ;
    RECT 74.99 57.645 75.2 57.715 ;
    RECT 71.21 56.925 71.42 56.995 ;
    RECT 71.21 57.285 71.42 57.355 ;
    RECT 71.21 57.645 71.42 57.715 ;
    RECT 71.67 56.925 71.88 56.995 ;
    RECT 71.67 57.285 71.88 57.355 ;
    RECT 71.67 57.645 71.88 57.715 ;
    RECT 31.37 56.925 31.58 56.995 ;
    RECT 31.37 57.285 31.58 57.355 ;
    RECT 31.37 57.645 31.58 57.715 ;
    RECT 31.83 56.925 32.04 56.995 ;
    RECT 31.83 57.285 32.04 57.355 ;
    RECT 31.83 57.645 32.04 57.715 ;
    RECT 67.89 56.925 68.1 56.995 ;
    RECT 67.89 57.285 68.1 57.355 ;
    RECT 67.89 57.645 68.1 57.715 ;
    RECT 68.35 56.925 68.56 56.995 ;
    RECT 68.35 57.285 68.56 57.355 ;
    RECT 68.35 57.645 68.56 57.715 ;
    RECT 28.05 56.925 28.26 56.995 ;
    RECT 28.05 57.285 28.26 57.355 ;
    RECT 28.05 57.645 28.26 57.715 ;
    RECT 28.51 56.925 28.72 56.995 ;
    RECT 28.51 57.285 28.72 57.355 ;
    RECT 28.51 57.645 28.72 57.715 ;
    RECT 24.73 56.925 24.94 56.995 ;
    RECT 24.73 57.285 24.94 57.355 ;
    RECT 24.73 57.645 24.94 57.715 ;
    RECT 25.19 56.925 25.4 56.995 ;
    RECT 25.19 57.285 25.4 57.355 ;
    RECT 25.19 57.645 25.4 57.715 ;
    RECT 21.41 56.925 21.62 56.995 ;
    RECT 21.41 57.285 21.62 57.355 ;
    RECT 21.41 57.645 21.62 57.715 ;
    RECT 21.87 56.925 22.08 56.995 ;
    RECT 21.87 57.285 22.08 57.355 ;
    RECT 21.87 57.645 22.08 57.715 ;
    RECT 18.09 56.925 18.3 56.995 ;
    RECT 18.09 57.285 18.3 57.355 ;
    RECT 18.09 57.645 18.3 57.715 ;
    RECT 18.55 56.925 18.76 56.995 ;
    RECT 18.55 57.285 18.76 57.355 ;
    RECT 18.55 57.645 18.76 57.715 ;
    RECT 14.77 56.925 14.98 56.995 ;
    RECT 14.77 57.285 14.98 57.355 ;
    RECT 14.77 57.645 14.98 57.715 ;
    RECT 15.23 56.925 15.44 56.995 ;
    RECT 15.23 57.285 15.44 57.355 ;
    RECT 15.23 57.645 15.44 57.715 ;
    RECT 11.45 56.925 11.66 56.995 ;
    RECT 11.45 57.285 11.66 57.355 ;
    RECT 11.45 57.645 11.66 57.715 ;
    RECT 11.91 56.925 12.12 56.995 ;
    RECT 11.91 57.285 12.12 57.355 ;
    RECT 11.91 57.645 12.12 57.715 ;
    RECT 8.13 56.925 8.34 56.995 ;
    RECT 8.13 57.285 8.34 57.355 ;
    RECT 8.13 57.645 8.34 57.715 ;
    RECT 8.59 56.925 8.8 56.995 ;
    RECT 8.59 57.285 8.8 57.355 ;
    RECT 8.59 57.645 8.8 57.715 ;
    RECT 4.81 56.925 5.02 56.995 ;
    RECT 4.81 57.285 5.02 57.355 ;
    RECT 4.81 57.645 5.02 57.715 ;
    RECT 5.27 56.925 5.48 56.995 ;
    RECT 5.27 57.285 5.48 57.355 ;
    RECT 5.27 57.645 5.48 57.715 ;
    RECT 164.17 56.925 164.38 56.995 ;
    RECT 164.17 57.285 164.38 57.355 ;
    RECT 164.17 57.645 164.38 57.715 ;
    RECT 164.63 56.925 164.84 56.995 ;
    RECT 164.63 57.285 164.84 57.355 ;
    RECT 164.63 57.645 164.84 57.715 ;
    RECT 1.49 56.925 1.7 56.995 ;
    RECT 1.49 57.285 1.7 57.355 ;
    RECT 1.49 57.645 1.7 57.715 ;
    RECT 1.95 56.925 2.16 56.995 ;
    RECT 1.95 57.285 2.16 57.355 ;
    RECT 1.95 57.645 2.16 57.715 ;
    RECT 160.85 56.925 161.06 56.995 ;
    RECT 160.85 57.285 161.06 57.355 ;
    RECT 160.85 57.645 161.06 57.715 ;
    RECT 161.31 56.925 161.52 56.995 ;
    RECT 161.31 57.285 161.52 57.355 ;
    RECT 161.31 57.645 161.52 57.715 ;
    RECT 157.53 56.925 157.74 56.995 ;
    RECT 157.53 57.285 157.74 57.355 ;
    RECT 157.53 57.645 157.74 57.715 ;
    RECT 157.99 56.925 158.2 56.995 ;
    RECT 157.99 57.285 158.2 57.355 ;
    RECT 157.99 57.645 158.2 57.715 ;
    RECT 154.21 56.925 154.42 56.995 ;
    RECT 154.21 57.285 154.42 57.355 ;
    RECT 154.21 57.645 154.42 57.715 ;
    RECT 154.67 56.925 154.88 56.995 ;
    RECT 154.67 57.285 154.88 57.355 ;
    RECT 154.67 57.645 154.88 57.715 ;
    RECT 150.89 56.925 151.1 56.995 ;
    RECT 150.89 57.285 151.1 57.355 ;
    RECT 150.89 57.645 151.1 57.715 ;
    RECT 151.35 56.925 151.56 56.995 ;
    RECT 151.35 57.285 151.56 57.355 ;
    RECT 151.35 57.645 151.56 57.715 ;
    RECT 147.57 56.925 147.78 56.995 ;
    RECT 147.57 57.285 147.78 57.355 ;
    RECT 147.57 57.645 147.78 57.715 ;
    RECT 148.03 56.925 148.24 56.995 ;
    RECT 148.03 57.285 148.24 57.355 ;
    RECT 148.03 57.645 148.24 57.715 ;
    RECT 144.25 56.925 144.46 56.995 ;
    RECT 144.25 57.285 144.46 57.355 ;
    RECT 144.25 57.645 144.46 57.715 ;
    RECT 144.71 56.925 144.92 56.995 ;
    RECT 144.71 57.285 144.92 57.355 ;
    RECT 144.71 57.645 144.92 57.715 ;
    RECT 140.93 56.925 141.14 56.995 ;
    RECT 140.93 57.285 141.14 57.355 ;
    RECT 140.93 57.645 141.14 57.715 ;
    RECT 141.39 56.925 141.6 56.995 ;
    RECT 141.39 57.285 141.6 57.355 ;
    RECT 141.39 57.645 141.6 57.715 ;
    RECT 137.61 56.925 137.82 56.995 ;
    RECT 137.61 57.285 137.82 57.355 ;
    RECT 137.61 57.645 137.82 57.715 ;
    RECT 138.07 56.925 138.28 56.995 ;
    RECT 138.07 57.285 138.28 57.355 ;
    RECT 138.07 57.645 138.28 57.715 ;
    RECT 134.29 56.925 134.5 56.995 ;
    RECT 134.29 57.285 134.5 57.355 ;
    RECT 134.29 57.645 134.5 57.715 ;
    RECT 134.75 56.925 134.96 56.995 ;
    RECT 134.75 57.285 134.96 57.355 ;
    RECT 134.75 57.645 134.96 57.715 ;
    RECT 64.57 56.925 64.78 56.995 ;
    RECT 64.57 57.285 64.78 57.355 ;
    RECT 64.57 57.645 64.78 57.715 ;
    RECT 65.03 56.925 65.24 56.995 ;
    RECT 65.03 57.285 65.24 57.355 ;
    RECT 65.03 57.645 65.24 57.715 ;
    RECT 61.25 56.205 61.46 56.275 ;
    RECT 61.25 56.565 61.46 56.635 ;
    RECT 61.25 56.925 61.46 56.995 ;
    RECT 61.71 56.205 61.92 56.275 ;
    RECT 61.71 56.565 61.92 56.635 ;
    RECT 61.71 56.925 61.92 56.995 ;
    RECT 57.93 56.205 58.14 56.275 ;
    RECT 57.93 56.565 58.14 56.635 ;
    RECT 57.93 56.925 58.14 56.995 ;
    RECT 58.39 56.205 58.6 56.275 ;
    RECT 58.39 56.565 58.6 56.635 ;
    RECT 58.39 56.925 58.6 56.995 ;
    RECT 54.61 56.205 54.82 56.275 ;
    RECT 54.61 56.565 54.82 56.635 ;
    RECT 54.61 56.925 54.82 56.995 ;
    RECT 55.07 56.205 55.28 56.275 ;
    RECT 55.07 56.565 55.28 56.635 ;
    RECT 55.07 56.925 55.28 56.995 ;
    RECT 51.29 56.205 51.5 56.275 ;
    RECT 51.29 56.565 51.5 56.635 ;
    RECT 51.29 56.925 51.5 56.995 ;
    RECT 51.75 56.205 51.96 56.275 ;
    RECT 51.75 56.565 51.96 56.635 ;
    RECT 51.75 56.925 51.96 56.995 ;
    RECT 47.97 56.205 48.18 56.275 ;
    RECT 47.97 56.565 48.18 56.635 ;
    RECT 47.97 56.925 48.18 56.995 ;
    RECT 48.43 56.205 48.64 56.275 ;
    RECT 48.43 56.565 48.64 56.635 ;
    RECT 48.43 56.925 48.64 56.995 ;
    RECT 44.65 56.205 44.86 56.275 ;
    RECT 44.65 56.565 44.86 56.635 ;
    RECT 44.65 56.925 44.86 56.995 ;
    RECT 45.11 56.205 45.32 56.275 ;
    RECT 45.11 56.565 45.32 56.635 ;
    RECT 45.11 56.925 45.32 56.995 ;
    RECT 41.33 56.205 41.54 56.275 ;
    RECT 41.33 56.565 41.54 56.635 ;
    RECT 41.33 56.925 41.54 56.995 ;
    RECT 41.79 56.205 42.0 56.275 ;
    RECT 41.79 56.565 42.0 56.635 ;
    RECT 41.79 56.925 42.0 56.995 ;
    RECT 38.01 56.205 38.22 56.275 ;
    RECT 38.01 56.565 38.22 56.635 ;
    RECT 38.01 56.925 38.22 56.995 ;
    RECT 38.47 56.205 38.68 56.275 ;
    RECT 38.47 56.565 38.68 56.635 ;
    RECT 38.47 56.925 38.68 56.995 ;
    RECT 34.69 56.205 34.9 56.275 ;
    RECT 34.69 56.565 34.9 56.635 ;
    RECT 34.69 56.925 34.9 56.995 ;
    RECT 35.15 56.205 35.36 56.275 ;
    RECT 35.15 56.565 35.36 56.635 ;
    RECT 35.15 56.925 35.36 56.995 ;
    RECT 173.945 56.565 174.015 56.635 ;
    RECT 130.97 56.205 131.18 56.275 ;
    RECT 130.97 56.565 131.18 56.635 ;
    RECT 130.97 56.925 131.18 56.995 ;
    RECT 131.43 56.205 131.64 56.275 ;
    RECT 131.43 56.565 131.64 56.635 ;
    RECT 131.43 56.925 131.64 56.995 ;
    RECT 127.65 56.205 127.86 56.275 ;
    RECT 127.65 56.565 127.86 56.635 ;
    RECT 127.65 56.925 127.86 56.995 ;
    RECT 128.11 56.205 128.32 56.275 ;
    RECT 128.11 56.565 128.32 56.635 ;
    RECT 128.11 56.925 128.32 56.995 ;
    RECT 124.33 56.205 124.54 56.275 ;
    RECT 124.33 56.565 124.54 56.635 ;
    RECT 124.33 56.925 124.54 56.995 ;
    RECT 124.79 56.205 125.0 56.275 ;
    RECT 124.79 56.565 125.0 56.635 ;
    RECT 124.79 56.925 125.0 56.995 ;
    RECT 121.01 56.205 121.22 56.275 ;
    RECT 121.01 56.565 121.22 56.635 ;
    RECT 121.01 56.925 121.22 56.995 ;
    RECT 121.47 56.205 121.68 56.275 ;
    RECT 121.47 56.565 121.68 56.635 ;
    RECT 121.47 56.925 121.68 56.995 ;
    RECT 117.69 56.205 117.9 56.275 ;
    RECT 117.69 56.565 117.9 56.635 ;
    RECT 117.69 56.925 117.9 56.995 ;
    RECT 118.15 56.205 118.36 56.275 ;
    RECT 118.15 56.565 118.36 56.635 ;
    RECT 118.15 56.925 118.36 56.995 ;
    RECT 114.37 56.205 114.58 56.275 ;
    RECT 114.37 56.565 114.58 56.635 ;
    RECT 114.37 56.925 114.58 56.995 ;
    RECT 114.83 56.205 115.04 56.275 ;
    RECT 114.83 56.565 115.04 56.635 ;
    RECT 114.83 56.925 115.04 56.995 ;
    RECT 111.05 56.205 111.26 56.275 ;
    RECT 111.05 56.565 111.26 56.635 ;
    RECT 111.05 56.925 111.26 56.995 ;
    RECT 111.51 56.205 111.72 56.275 ;
    RECT 111.51 56.565 111.72 56.635 ;
    RECT 111.51 56.925 111.72 56.995 ;
    RECT 107.73 56.205 107.94 56.275 ;
    RECT 107.73 56.565 107.94 56.635 ;
    RECT 107.73 56.925 107.94 56.995 ;
    RECT 108.19 56.205 108.4 56.275 ;
    RECT 108.19 56.565 108.4 56.635 ;
    RECT 108.19 56.925 108.4 56.995 ;
    RECT 104.41 56.205 104.62 56.275 ;
    RECT 104.41 56.565 104.62 56.635 ;
    RECT 104.41 56.925 104.62 56.995 ;
    RECT 104.87 56.205 105.08 56.275 ;
    RECT 104.87 56.565 105.08 56.635 ;
    RECT 104.87 56.925 105.08 56.995 ;
    RECT 101.09 56.205 101.3 56.275 ;
    RECT 101.09 56.565 101.3 56.635 ;
    RECT 101.09 56.925 101.3 56.995 ;
    RECT 101.55 56.205 101.76 56.275 ;
    RECT 101.55 56.565 101.76 56.635 ;
    RECT 101.55 56.925 101.76 56.995 ;
    RECT 0.4 56.565 0.47 56.635 ;
    RECT 170.81 56.205 171.02 56.275 ;
    RECT 170.81 56.565 171.02 56.635 ;
    RECT 170.81 56.925 171.02 56.995 ;
    RECT 171.27 56.205 171.48 56.275 ;
    RECT 171.27 56.565 171.48 56.635 ;
    RECT 171.27 56.925 171.48 56.995 ;
    RECT 167.49 56.205 167.7 56.275 ;
    RECT 167.49 56.565 167.7 56.635 ;
    RECT 167.49 56.925 167.7 56.995 ;
    RECT 167.95 56.205 168.16 56.275 ;
    RECT 167.95 56.565 168.16 56.635 ;
    RECT 167.95 56.925 168.16 56.995 ;
    RECT 97.77 56.205 97.98 56.275 ;
    RECT 97.77 56.565 97.98 56.635 ;
    RECT 97.77 56.925 97.98 56.995 ;
    RECT 98.23 56.205 98.44 56.275 ;
    RECT 98.23 56.565 98.44 56.635 ;
    RECT 98.23 56.925 98.44 56.995 ;
    RECT 94.45 56.205 94.66 56.275 ;
    RECT 94.45 56.565 94.66 56.635 ;
    RECT 94.45 56.925 94.66 56.995 ;
    RECT 94.91 56.205 95.12 56.275 ;
    RECT 94.91 56.565 95.12 56.635 ;
    RECT 94.91 56.925 95.12 56.995 ;
    RECT 91.13 56.205 91.34 56.275 ;
    RECT 91.13 56.565 91.34 56.635 ;
    RECT 91.13 56.925 91.34 56.995 ;
    RECT 91.59 56.205 91.8 56.275 ;
    RECT 91.59 56.565 91.8 56.635 ;
    RECT 91.59 56.925 91.8 56.995 ;
    RECT 87.81 56.205 88.02 56.275 ;
    RECT 87.81 56.565 88.02 56.635 ;
    RECT 87.81 56.925 88.02 56.995 ;
    RECT 88.27 56.205 88.48 56.275 ;
    RECT 88.27 56.565 88.48 56.635 ;
    RECT 88.27 56.925 88.48 56.995 ;
    RECT 84.49 56.205 84.7 56.275 ;
    RECT 84.49 56.565 84.7 56.635 ;
    RECT 84.49 56.925 84.7 56.995 ;
    RECT 84.95 56.205 85.16 56.275 ;
    RECT 84.95 56.565 85.16 56.635 ;
    RECT 84.95 56.925 85.16 56.995 ;
    RECT 81.17 56.205 81.38 56.275 ;
    RECT 81.17 56.565 81.38 56.635 ;
    RECT 81.17 56.925 81.38 56.995 ;
    RECT 81.63 56.205 81.84 56.275 ;
    RECT 81.63 56.565 81.84 56.635 ;
    RECT 81.63 56.925 81.84 56.995 ;
    RECT 77.85 56.205 78.06 56.275 ;
    RECT 77.85 56.565 78.06 56.635 ;
    RECT 77.85 56.925 78.06 56.995 ;
    RECT 78.31 56.205 78.52 56.275 ;
    RECT 78.31 56.565 78.52 56.635 ;
    RECT 78.31 56.925 78.52 56.995 ;
    RECT 74.53 56.205 74.74 56.275 ;
    RECT 74.53 56.565 74.74 56.635 ;
    RECT 74.53 56.925 74.74 56.995 ;
    RECT 74.99 56.205 75.2 56.275 ;
    RECT 74.99 56.565 75.2 56.635 ;
    RECT 74.99 56.925 75.2 56.995 ;
    RECT 71.21 56.205 71.42 56.275 ;
    RECT 71.21 56.565 71.42 56.635 ;
    RECT 71.21 56.925 71.42 56.995 ;
    RECT 71.67 56.205 71.88 56.275 ;
    RECT 71.67 56.565 71.88 56.635 ;
    RECT 71.67 56.925 71.88 56.995 ;
    RECT 31.37 56.205 31.58 56.275 ;
    RECT 31.37 56.565 31.58 56.635 ;
    RECT 31.37 56.925 31.58 56.995 ;
    RECT 31.83 56.205 32.04 56.275 ;
    RECT 31.83 56.565 32.04 56.635 ;
    RECT 31.83 56.925 32.04 56.995 ;
    RECT 67.89 56.205 68.1 56.275 ;
    RECT 67.89 56.565 68.1 56.635 ;
    RECT 67.89 56.925 68.1 56.995 ;
    RECT 68.35 56.205 68.56 56.275 ;
    RECT 68.35 56.565 68.56 56.635 ;
    RECT 68.35 56.925 68.56 56.995 ;
    RECT 28.05 56.205 28.26 56.275 ;
    RECT 28.05 56.565 28.26 56.635 ;
    RECT 28.05 56.925 28.26 56.995 ;
    RECT 28.51 56.205 28.72 56.275 ;
    RECT 28.51 56.565 28.72 56.635 ;
    RECT 28.51 56.925 28.72 56.995 ;
    RECT 24.73 56.205 24.94 56.275 ;
    RECT 24.73 56.565 24.94 56.635 ;
    RECT 24.73 56.925 24.94 56.995 ;
    RECT 25.19 56.205 25.4 56.275 ;
    RECT 25.19 56.565 25.4 56.635 ;
    RECT 25.19 56.925 25.4 56.995 ;
    RECT 21.41 56.205 21.62 56.275 ;
    RECT 21.41 56.565 21.62 56.635 ;
    RECT 21.41 56.925 21.62 56.995 ;
    RECT 21.87 56.205 22.08 56.275 ;
    RECT 21.87 56.565 22.08 56.635 ;
    RECT 21.87 56.925 22.08 56.995 ;
    RECT 18.09 56.205 18.3 56.275 ;
    RECT 18.09 56.565 18.3 56.635 ;
    RECT 18.09 56.925 18.3 56.995 ;
    RECT 18.55 56.205 18.76 56.275 ;
    RECT 18.55 56.565 18.76 56.635 ;
    RECT 18.55 56.925 18.76 56.995 ;
    RECT 14.77 56.205 14.98 56.275 ;
    RECT 14.77 56.565 14.98 56.635 ;
    RECT 14.77 56.925 14.98 56.995 ;
    RECT 15.23 56.205 15.44 56.275 ;
    RECT 15.23 56.565 15.44 56.635 ;
    RECT 15.23 56.925 15.44 56.995 ;
    RECT 11.45 56.205 11.66 56.275 ;
    RECT 11.45 56.565 11.66 56.635 ;
    RECT 11.45 56.925 11.66 56.995 ;
    RECT 11.91 56.205 12.12 56.275 ;
    RECT 11.91 56.565 12.12 56.635 ;
    RECT 11.91 56.925 12.12 56.995 ;
    RECT 8.13 56.205 8.34 56.275 ;
    RECT 8.13 56.565 8.34 56.635 ;
    RECT 8.13 56.925 8.34 56.995 ;
    RECT 8.59 56.205 8.8 56.275 ;
    RECT 8.59 56.565 8.8 56.635 ;
    RECT 8.59 56.925 8.8 56.995 ;
    RECT 4.81 56.205 5.02 56.275 ;
    RECT 4.81 56.565 5.02 56.635 ;
    RECT 4.81 56.925 5.02 56.995 ;
    RECT 5.27 56.205 5.48 56.275 ;
    RECT 5.27 56.565 5.48 56.635 ;
    RECT 5.27 56.925 5.48 56.995 ;
    RECT 164.17 56.205 164.38 56.275 ;
    RECT 164.17 56.565 164.38 56.635 ;
    RECT 164.17 56.925 164.38 56.995 ;
    RECT 164.63 56.205 164.84 56.275 ;
    RECT 164.63 56.565 164.84 56.635 ;
    RECT 164.63 56.925 164.84 56.995 ;
    RECT 1.49 56.205 1.7 56.275 ;
    RECT 1.49 56.565 1.7 56.635 ;
    RECT 1.49 56.925 1.7 56.995 ;
    RECT 1.95 56.205 2.16 56.275 ;
    RECT 1.95 56.565 2.16 56.635 ;
    RECT 1.95 56.925 2.16 56.995 ;
    RECT 160.85 56.205 161.06 56.275 ;
    RECT 160.85 56.565 161.06 56.635 ;
    RECT 160.85 56.925 161.06 56.995 ;
    RECT 161.31 56.205 161.52 56.275 ;
    RECT 161.31 56.565 161.52 56.635 ;
    RECT 161.31 56.925 161.52 56.995 ;
    RECT 157.53 56.205 157.74 56.275 ;
    RECT 157.53 56.565 157.74 56.635 ;
    RECT 157.53 56.925 157.74 56.995 ;
    RECT 157.99 56.205 158.2 56.275 ;
    RECT 157.99 56.565 158.2 56.635 ;
    RECT 157.99 56.925 158.2 56.995 ;
    RECT 154.21 56.205 154.42 56.275 ;
    RECT 154.21 56.565 154.42 56.635 ;
    RECT 154.21 56.925 154.42 56.995 ;
    RECT 154.67 56.205 154.88 56.275 ;
    RECT 154.67 56.565 154.88 56.635 ;
    RECT 154.67 56.925 154.88 56.995 ;
    RECT 150.89 56.205 151.1 56.275 ;
    RECT 150.89 56.565 151.1 56.635 ;
    RECT 150.89 56.925 151.1 56.995 ;
    RECT 151.35 56.205 151.56 56.275 ;
    RECT 151.35 56.565 151.56 56.635 ;
    RECT 151.35 56.925 151.56 56.995 ;
    RECT 147.57 56.205 147.78 56.275 ;
    RECT 147.57 56.565 147.78 56.635 ;
    RECT 147.57 56.925 147.78 56.995 ;
    RECT 148.03 56.205 148.24 56.275 ;
    RECT 148.03 56.565 148.24 56.635 ;
    RECT 148.03 56.925 148.24 56.995 ;
    RECT 144.25 56.205 144.46 56.275 ;
    RECT 144.25 56.565 144.46 56.635 ;
    RECT 144.25 56.925 144.46 56.995 ;
    RECT 144.71 56.205 144.92 56.275 ;
    RECT 144.71 56.565 144.92 56.635 ;
    RECT 144.71 56.925 144.92 56.995 ;
    RECT 140.93 56.205 141.14 56.275 ;
    RECT 140.93 56.565 141.14 56.635 ;
    RECT 140.93 56.925 141.14 56.995 ;
    RECT 141.39 56.205 141.6 56.275 ;
    RECT 141.39 56.565 141.6 56.635 ;
    RECT 141.39 56.925 141.6 56.995 ;
    RECT 137.61 56.205 137.82 56.275 ;
    RECT 137.61 56.565 137.82 56.635 ;
    RECT 137.61 56.925 137.82 56.995 ;
    RECT 138.07 56.205 138.28 56.275 ;
    RECT 138.07 56.565 138.28 56.635 ;
    RECT 138.07 56.925 138.28 56.995 ;
    RECT 134.29 56.205 134.5 56.275 ;
    RECT 134.29 56.565 134.5 56.635 ;
    RECT 134.29 56.925 134.5 56.995 ;
    RECT 134.75 56.205 134.96 56.275 ;
    RECT 134.75 56.565 134.96 56.635 ;
    RECT 134.75 56.925 134.96 56.995 ;
    RECT 64.57 56.205 64.78 56.275 ;
    RECT 64.57 56.565 64.78 56.635 ;
    RECT 64.57 56.925 64.78 56.995 ;
    RECT 65.03 56.205 65.24 56.275 ;
    RECT 65.03 56.565 65.24 56.635 ;
    RECT 65.03 56.925 65.24 56.995 ;
    RECT 61.25 55.485 61.46 55.555 ;
    RECT 61.25 55.845 61.46 55.915 ;
    RECT 61.25 56.205 61.46 56.275 ;
    RECT 61.71 55.485 61.92 55.555 ;
    RECT 61.71 55.845 61.92 55.915 ;
    RECT 61.71 56.205 61.92 56.275 ;
    RECT 57.93 55.485 58.14 55.555 ;
    RECT 57.93 55.845 58.14 55.915 ;
    RECT 57.93 56.205 58.14 56.275 ;
    RECT 58.39 55.485 58.6 55.555 ;
    RECT 58.39 55.845 58.6 55.915 ;
    RECT 58.39 56.205 58.6 56.275 ;
    RECT 54.61 55.485 54.82 55.555 ;
    RECT 54.61 55.845 54.82 55.915 ;
    RECT 54.61 56.205 54.82 56.275 ;
    RECT 55.07 55.485 55.28 55.555 ;
    RECT 55.07 55.845 55.28 55.915 ;
    RECT 55.07 56.205 55.28 56.275 ;
    RECT 51.29 55.485 51.5 55.555 ;
    RECT 51.29 55.845 51.5 55.915 ;
    RECT 51.29 56.205 51.5 56.275 ;
    RECT 51.75 55.485 51.96 55.555 ;
    RECT 51.75 55.845 51.96 55.915 ;
    RECT 51.75 56.205 51.96 56.275 ;
    RECT 47.97 55.485 48.18 55.555 ;
    RECT 47.97 55.845 48.18 55.915 ;
    RECT 47.97 56.205 48.18 56.275 ;
    RECT 48.43 55.485 48.64 55.555 ;
    RECT 48.43 55.845 48.64 55.915 ;
    RECT 48.43 56.205 48.64 56.275 ;
    RECT 44.65 55.485 44.86 55.555 ;
    RECT 44.65 55.845 44.86 55.915 ;
    RECT 44.65 56.205 44.86 56.275 ;
    RECT 45.11 55.485 45.32 55.555 ;
    RECT 45.11 55.845 45.32 55.915 ;
    RECT 45.11 56.205 45.32 56.275 ;
    RECT 41.33 55.485 41.54 55.555 ;
    RECT 41.33 55.845 41.54 55.915 ;
    RECT 41.33 56.205 41.54 56.275 ;
    RECT 41.79 55.485 42.0 55.555 ;
    RECT 41.79 55.845 42.0 55.915 ;
    RECT 41.79 56.205 42.0 56.275 ;
    RECT 38.01 55.485 38.22 55.555 ;
    RECT 38.01 55.845 38.22 55.915 ;
    RECT 38.01 56.205 38.22 56.275 ;
    RECT 38.47 55.485 38.68 55.555 ;
    RECT 38.47 55.845 38.68 55.915 ;
    RECT 38.47 56.205 38.68 56.275 ;
    RECT 34.69 55.485 34.9 55.555 ;
    RECT 34.69 55.845 34.9 55.915 ;
    RECT 34.69 56.205 34.9 56.275 ;
    RECT 35.15 55.485 35.36 55.555 ;
    RECT 35.15 55.845 35.36 55.915 ;
    RECT 35.15 56.205 35.36 56.275 ;
    RECT 173.945 55.845 174.015 55.915 ;
    RECT 130.97 55.485 131.18 55.555 ;
    RECT 130.97 55.845 131.18 55.915 ;
    RECT 130.97 56.205 131.18 56.275 ;
    RECT 131.43 55.485 131.64 55.555 ;
    RECT 131.43 55.845 131.64 55.915 ;
    RECT 131.43 56.205 131.64 56.275 ;
    RECT 127.65 55.485 127.86 55.555 ;
    RECT 127.65 55.845 127.86 55.915 ;
    RECT 127.65 56.205 127.86 56.275 ;
    RECT 128.11 55.485 128.32 55.555 ;
    RECT 128.11 55.845 128.32 55.915 ;
    RECT 128.11 56.205 128.32 56.275 ;
    RECT 124.33 55.485 124.54 55.555 ;
    RECT 124.33 55.845 124.54 55.915 ;
    RECT 124.33 56.205 124.54 56.275 ;
    RECT 124.79 55.485 125.0 55.555 ;
    RECT 124.79 55.845 125.0 55.915 ;
    RECT 124.79 56.205 125.0 56.275 ;
    RECT 121.01 55.485 121.22 55.555 ;
    RECT 121.01 55.845 121.22 55.915 ;
    RECT 121.01 56.205 121.22 56.275 ;
    RECT 121.47 55.485 121.68 55.555 ;
    RECT 121.47 55.845 121.68 55.915 ;
    RECT 121.47 56.205 121.68 56.275 ;
    RECT 117.69 55.485 117.9 55.555 ;
    RECT 117.69 55.845 117.9 55.915 ;
    RECT 117.69 56.205 117.9 56.275 ;
    RECT 118.15 55.485 118.36 55.555 ;
    RECT 118.15 55.845 118.36 55.915 ;
    RECT 118.15 56.205 118.36 56.275 ;
    RECT 114.37 55.485 114.58 55.555 ;
    RECT 114.37 55.845 114.58 55.915 ;
    RECT 114.37 56.205 114.58 56.275 ;
    RECT 114.83 55.485 115.04 55.555 ;
    RECT 114.83 55.845 115.04 55.915 ;
    RECT 114.83 56.205 115.04 56.275 ;
    RECT 111.05 55.485 111.26 55.555 ;
    RECT 111.05 55.845 111.26 55.915 ;
    RECT 111.05 56.205 111.26 56.275 ;
    RECT 111.51 55.485 111.72 55.555 ;
    RECT 111.51 55.845 111.72 55.915 ;
    RECT 111.51 56.205 111.72 56.275 ;
    RECT 107.73 55.485 107.94 55.555 ;
    RECT 107.73 55.845 107.94 55.915 ;
    RECT 107.73 56.205 107.94 56.275 ;
    RECT 108.19 55.485 108.4 55.555 ;
    RECT 108.19 55.845 108.4 55.915 ;
    RECT 108.19 56.205 108.4 56.275 ;
    RECT 104.41 55.485 104.62 55.555 ;
    RECT 104.41 55.845 104.62 55.915 ;
    RECT 104.41 56.205 104.62 56.275 ;
    RECT 104.87 55.485 105.08 55.555 ;
    RECT 104.87 55.845 105.08 55.915 ;
    RECT 104.87 56.205 105.08 56.275 ;
    RECT 101.09 55.485 101.3 55.555 ;
    RECT 101.09 55.845 101.3 55.915 ;
    RECT 101.09 56.205 101.3 56.275 ;
    RECT 101.55 55.485 101.76 55.555 ;
    RECT 101.55 55.845 101.76 55.915 ;
    RECT 101.55 56.205 101.76 56.275 ;
    RECT 0.4 55.845 0.47 55.915 ;
    RECT 170.81 55.485 171.02 55.555 ;
    RECT 170.81 55.845 171.02 55.915 ;
    RECT 170.81 56.205 171.02 56.275 ;
    RECT 171.27 55.485 171.48 55.555 ;
    RECT 171.27 55.845 171.48 55.915 ;
    RECT 171.27 56.205 171.48 56.275 ;
    RECT 167.49 55.485 167.7 55.555 ;
    RECT 167.49 55.845 167.7 55.915 ;
    RECT 167.49 56.205 167.7 56.275 ;
    RECT 167.95 55.485 168.16 55.555 ;
    RECT 167.95 55.845 168.16 55.915 ;
    RECT 167.95 56.205 168.16 56.275 ;
    RECT 97.77 55.485 97.98 55.555 ;
    RECT 97.77 55.845 97.98 55.915 ;
    RECT 97.77 56.205 97.98 56.275 ;
    RECT 98.23 55.485 98.44 55.555 ;
    RECT 98.23 55.845 98.44 55.915 ;
    RECT 98.23 56.205 98.44 56.275 ;
    RECT 94.45 55.485 94.66 55.555 ;
    RECT 94.45 55.845 94.66 55.915 ;
    RECT 94.45 56.205 94.66 56.275 ;
    RECT 94.91 55.485 95.12 55.555 ;
    RECT 94.91 55.845 95.12 55.915 ;
    RECT 94.91 56.205 95.12 56.275 ;
    RECT 91.13 55.485 91.34 55.555 ;
    RECT 91.13 55.845 91.34 55.915 ;
    RECT 91.13 56.205 91.34 56.275 ;
    RECT 91.59 55.485 91.8 55.555 ;
    RECT 91.59 55.845 91.8 55.915 ;
    RECT 91.59 56.205 91.8 56.275 ;
    RECT 87.81 55.485 88.02 55.555 ;
    RECT 87.81 55.845 88.02 55.915 ;
    RECT 87.81 56.205 88.02 56.275 ;
    RECT 88.27 55.485 88.48 55.555 ;
    RECT 88.27 55.845 88.48 55.915 ;
    RECT 88.27 56.205 88.48 56.275 ;
    RECT 84.49 55.485 84.7 55.555 ;
    RECT 84.49 55.845 84.7 55.915 ;
    RECT 84.49 56.205 84.7 56.275 ;
    RECT 84.95 55.485 85.16 55.555 ;
    RECT 84.95 55.845 85.16 55.915 ;
    RECT 84.95 56.205 85.16 56.275 ;
    RECT 81.17 55.485 81.38 55.555 ;
    RECT 81.17 55.845 81.38 55.915 ;
    RECT 81.17 56.205 81.38 56.275 ;
    RECT 81.63 55.485 81.84 55.555 ;
    RECT 81.63 55.845 81.84 55.915 ;
    RECT 81.63 56.205 81.84 56.275 ;
    RECT 77.85 55.485 78.06 55.555 ;
    RECT 77.85 55.845 78.06 55.915 ;
    RECT 77.85 56.205 78.06 56.275 ;
    RECT 78.31 55.485 78.52 55.555 ;
    RECT 78.31 55.845 78.52 55.915 ;
    RECT 78.31 56.205 78.52 56.275 ;
    RECT 74.53 55.485 74.74 55.555 ;
    RECT 74.53 55.845 74.74 55.915 ;
    RECT 74.53 56.205 74.74 56.275 ;
    RECT 74.99 55.485 75.2 55.555 ;
    RECT 74.99 55.845 75.2 55.915 ;
    RECT 74.99 56.205 75.2 56.275 ;
    RECT 71.21 55.485 71.42 55.555 ;
    RECT 71.21 55.845 71.42 55.915 ;
    RECT 71.21 56.205 71.42 56.275 ;
    RECT 71.67 55.485 71.88 55.555 ;
    RECT 71.67 55.845 71.88 55.915 ;
    RECT 71.67 56.205 71.88 56.275 ;
    RECT 31.37 55.485 31.58 55.555 ;
    RECT 31.37 55.845 31.58 55.915 ;
    RECT 31.37 56.205 31.58 56.275 ;
    RECT 31.83 55.485 32.04 55.555 ;
    RECT 31.83 55.845 32.04 55.915 ;
    RECT 31.83 56.205 32.04 56.275 ;
    RECT 67.89 55.485 68.1 55.555 ;
    RECT 67.89 55.845 68.1 55.915 ;
    RECT 67.89 56.205 68.1 56.275 ;
    RECT 68.35 55.485 68.56 55.555 ;
    RECT 68.35 55.845 68.56 55.915 ;
    RECT 68.35 56.205 68.56 56.275 ;
    RECT 28.05 55.485 28.26 55.555 ;
    RECT 28.05 55.845 28.26 55.915 ;
    RECT 28.05 56.205 28.26 56.275 ;
    RECT 28.51 55.485 28.72 55.555 ;
    RECT 28.51 55.845 28.72 55.915 ;
    RECT 28.51 56.205 28.72 56.275 ;
    RECT 24.73 55.485 24.94 55.555 ;
    RECT 24.73 55.845 24.94 55.915 ;
    RECT 24.73 56.205 24.94 56.275 ;
    RECT 25.19 55.485 25.4 55.555 ;
    RECT 25.19 55.845 25.4 55.915 ;
    RECT 25.19 56.205 25.4 56.275 ;
    RECT 21.41 55.485 21.62 55.555 ;
    RECT 21.41 55.845 21.62 55.915 ;
    RECT 21.41 56.205 21.62 56.275 ;
    RECT 21.87 55.485 22.08 55.555 ;
    RECT 21.87 55.845 22.08 55.915 ;
    RECT 21.87 56.205 22.08 56.275 ;
    RECT 18.09 55.485 18.3 55.555 ;
    RECT 18.09 55.845 18.3 55.915 ;
    RECT 18.09 56.205 18.3 56.275 ;
    RECT 18.55 55.485 18.76 55.555 ;
    RECT 18.55 55.845 18.76 55.915 ;
    RECT 18.55 56.205 18.76 56.275 ;
    RECT 14.77 55.485 14.98 55.555 ;
    RECT 14.77 55.845 14.98 55.915 ;
    RECT 14.77 56.205 14.98 56.275 ;
    RECT 15.23 55.485 15.44 55.555 ;
    RECT 15.23 55.845 15.44 55.915 ;
    RECT 15.23 56.205 15.44 56.275 ;
    RECT 11.45 55.485 11.66 55.555 ;
    RECT 11.45 55.845 11.66 55.915 ;
    RECT 11.45 56.205 11.66 56.275 ;
    RECT 11.91 55.485 12.12 55.555 ;
    RECT 11.91 55.845 12.12 55.915 ;
    RECT 11.91 56.205 12.12 56.275 ;
    RECT 8.13 55.485 8.34 55.555 ;
    RECT 8.13 55.845 8.34 55.915 ;
    RECT 8.13 56.205 8.34 56.275 ;
    RECT 8.59 55.485 8.8 55.555 ;
    RECT 8.59 55.845 8.8 55.915 ;
    RECT 8.59 56.205 8.8 56.275 ;
    RECT 4.81 55.485 5.02 55.555 ;
    RECT 4.81 55.845 5.02 55.915 ;
    RECT 4.81 56.205 5.02 56.275 ;
    RECT 5.27 55.485 5.48 55.555 ;
    RECT 5.27 55.845 5.48 55.915 ;
    RECT 5.27 56.205 5.48 56.275 ;
    RECT 164.17 55.485 164.38 55.555 ;
    RECT 164.17 55.845 164.38 55.915 ;
    RECT 164.17 56.205 164.38 56.275 ;
    RECT 164.63 55.485 164.84 55.555 ;
    RECT 164.63 55.845 164.84 55.915 ;
    RECT 164.63 56.205 164.84 56.275 ;
    RECT 1.49 55.485 1.7 55.555 ;
    RECT 1.49 55.845 1.7 55.915 ;
    RECT 1.49 56.205 1.7 56.275 ;
    RECT 1.95 55.485 2.16 55.555 ;
    RECT 1.95 55.845 2.16 55.915 ;
    RECT 1.95 56.205 2.16 56.275 ;
    RECT 160.85 55.485 161.06 55.555 ;
    RECT 160.85 55.845 161.06 55.915 ;
    RECT 160.85 56.205 161.06 56.275 ;
    RECT 161.31 55.485 161.52 55.555 ;
    RECT 161.31 55.845 161.52 55.915 ;
    RECT 161.31 56.205 161.52 56.275 ;
    RECT 157.53 55.485 157.74 55.555 ;
    RECT 157.53 55.845 157.74 55.915 ;
    RECT 157.53 56.205 157.74 56.275 ;
    RECT 157.99 55.485 158.2 55.555 ;
    RECT 157.99 55.845 158.2 55.915 ;
    RECT 157.99 56.205 158.2 56.275 ;
    RECT 154.21 55.485 154.42 55.555 ;
    RECT 154.21 55.845 154.42 55.915 ;
    RECT 154.21 56.205 154.42 56.275 ;
    RECT 154.67 55.485 154.88 55.555 ;
    RECT 154.67 55.845 154.88 55.915 ;
    RECT 154.67 56.205 154.88 56.275 ;
    RECT 150.89 55.485 151.1 55.555 ;
    RECT 150.89 55.845 151.1 55.915 ;
    RECT 150.89 56.205 151.1 56.275 ;
    RECT 151.35 55.485 151.56 55.555 ;
    RECT 151.35 55.845 151.56 55.915 ;
    RECT 151.35 56.205 151.56 56.275 ;
    RECT 147.57 55.485 147.78 55.555 ;
    RECT 147.57 55.845 147.78 55.915 ;
    RECT 147.57 56.205 147.78 56.275 ;
    RECT 148.03 55.485 148.24 55.555 ;
    RECT 148.03 55.845 148.24 55.915 ;
    RECT 148.03 56.205 148.24 56.275 ;
    RECT 144.25 55.485 144.46 55.555 ;
    RECT 144.25 55.845 144.46 55.915 ;
    RECT 144.25 56.205 144.46 56.275 ;
    RECT 144.71 55.485 144.92 55.555 ;
    RECT 144.71 55.845 144.92 55.915 ;
    RECT 144.71 56.205 144.92 56.275 ;
    RECT 140.93 55.485 141.14 55.555 ;
    RECT 140.93 55.845 141.14 55.915 ;
    RECT 140.93 56.205 141.14 56.275 ;
    RECT 141.39 55.485 141.6 55.555 ;
    RECT 141.39 55.845 141.6 55.915 ;
    RECT 141.39 56.205 141.6 56.275 ;
    RECT 137.61 55.485 137.82 55.555 ;
    RECT 137.61 55.845 137.82 55.915 ;
    RECT 137.61 56.205 137.82 56.275 ;
    RECT 138.07 55.485 138.28 55.555 ;
    RECT 138.07 55.845 138.28 55.915 ;
    RECT 138.07 56.205 138.28 56.275 ;
    RECT 134.29 55.485 134.5 55.555 ;
    RECT 134.29 55.845 134.5 55.915 ;
    RECT 134.29 56.205 134.5 56.275 ;
    RECT 134.75 55.485 134.96 55.555 ;
    RECT 134.75 55.845 134.96 55.915 ;
    RECT 134.75 56.205 134.96 56.275 ;
    RECT 64.57 55.485 64.78 55.555 ;
    RECT 64.57 55.845 64.78 55.915 ;
    RECT 64.57 56.205 64.78 56.275 ;
    RECT 65.03 55.485 65.24 55.555 ;
    RECT 65.03 55.845 65.24 55.915 ;
    RECT 65.03 56.205 65.24 56.275 ;
    RECT 61.25 54.765 61.46 54.835 ;
    RECT 61.25 55.125 61.46 55.195 ;
    RECT 61.25 55.485 61.46 55.555 ;
    RECT 61.71 54.765 61.92 54.835 ;
    RECT 61.71 55.125 61.92 55.195 ;
    RECT 61.71 55.485 61.92 55.555 ;
    RECT 57.93 54.765 58.14 54.835 ;
    RECT 57.93 55.125 58.14 55.195 ;
    RECT 57.93 55.485 58.14 55.555 ;
    RECT 58.39 54.765 58.6 54.835 ;
    RECT 58.39 55.125 58.6 55.195 ;
    RECT 58.39 55.485 58.6 55.555 ;
    RECT 54.61 54.765 54.82 54.835 ;
    RECT 54.61 55.125 54.82 55.195 ;
    RECT 54.61 55.485 54.82 55.555 ;
    RECT 55.07 54.765 55.28 54.835 ;
    RECT 55.07 55.125 55.28 55.195 ;
    RECT 55.07 55.485 55.28 55.555 ;
    RECT 51.29 54.765 51.5 54.835 ;
    RECT 51.29 55.125 51.5 55.195 ;
    RECT 51.29 55.485 51.5 55.555 ;
    RECT 51.75 54.765 51.96 54.835 ;
    RECT 51.75 55.125 51.96 55.195 ;
    RECT 51.75 55.485 51.96 55.555 ;
    RECT 47.97 54.765 48.18 54.835 ;
    RECT 47.97 55.125 48.18 55.195 ;
    RECT 47.97 55.485 48.18 55.555 ;
    RECT 48.43 54.765 48.64 54.835 ;
    RECT 48.43 55.125 48.64 55.195 ;
    RECT 48.43 55.485 48.64 55.555 ;
    RECT 44.65 54.765 44.86 54.835 ;
    RECT 44.65 55.125 44.86 55.195 ;
    RECT 44.65 55.485 44.86 55.555 ;
    RECT 45.11 54.765 45.32 54.835 ;
    RECT 45.11 55.125 45.32 55.195 ;
    RECT 45.11 55.485 45.32 55.555 ;
    RECT 41.33 54.765 41.54 54.835 ;
    RECT 41.33 55.125 41.54 55.195 ;
    RECT 41.33 55.485 41.54 55.555 ;
    RECT 41.79 54.765 42.0 54.835 ;
    RECT 41.79 55.125 42.0 55.195 ;
    RECT 41.79 55.485 42.0 55.555 ;
    RECT 38.01 54.765 38.22 54.835 ;
    RECT 38.01 55.125 38.22 55.195 ;
    RECT 38.01 55.485 38.22 55.555 ;
    RECT 38.47 54.765 38.68 54.835 ;
    RECT 38.47 55.125 38.68 55.195 ;
    RECT 38.47 55.485 38.68 55.555 ;
    RECT 34.69 54.765 34.9 54.835 ;
    RECT 34.69 55.125 34.9 55.195 ;
    RECT 34.69 55.485 34.9 55.555 ;
    RECT 35.15 54.765 35.36 54.835 ;
    RECT 35.15 55.125 35.36 55.195 ;
    RECT 35.15 55.485 35.36 55.555 ;
    RECT 173.945 55.125 174.015 55.195 ;
    RECT 130.97 54.765 131.18 54.835 ;
    RECT 130.97 55.125 131.18 55.195 ;
    RECT 130.97 55.485 131.18 55.555 ;
    RECT 131.43 54.765 131.64 54.835 ;
    RECT 131.43 55.125 131.64 55.195 ;
    RECT 131.43 55.485 131.64 55.555 ;
    RECT 127.65 54.765 127.86 54.835 ;
    RECT 127.65 55.125 127.86 55.195 ;
    RECT 127.65 55.485 127.86 55.555 ;
    RECT 128.11 54.765 128.32 54.835 ;
    RECT 128.11 55.125 128.32 55.195 ;
    RECT 128.11 55.485 128.32 55.555 ;
    RECT 124.33 54.765 124.54 54.835 ;
    RECT 124.33 55.125 124.54 55.195 ;
    RECT 124.33 55.485 124.54 55.555 ;
    RECT 124.79 54.765 125.0 54.835 ;
    RECT 124.79 55.125 125.0 55.195 ;
    RECT 124.79 55.485 125.0 55.555 ;
    RECT 121.01 54.765 121.22 54.835 ;
    RECT 121.01 55.125 121.22 55.195 ;
    RECT 121.01 55.485 121.22 55.555 ;
    RECT 121.47 54.765 121.68 54.835 ;
    RECT 121.47 55.125 121.68 55.195 ;
    RECT 121.47 55.485 121.68 55.555 ;
    RECT 117.69 54.765 117.9 54.835 ;
    RECT 117.69 55.125 117.9 55.195 ;
    RECT 117.69 55.485 117.9 55.555 ;
    RECT 118.15 54.765 118.36 54.835 ;
    RECT 118.15 55.125 118.36 55.195 ;
    RECT 118.15 55.485 118.36 55.555 ;
    RECT 114.37 54.765 114.58 54.835 ;
    RECT 114.37 55.125 114.58 55.195 ;
    RECT 114.37 55.485 114.58 55.555 ;
    RECT 114.83 54.765 115.04 54.835 ;
    RECT 114.83 55.125 115.04 55.195 ;
    RECT 114.83 55.485 115.04 55.555 ;
    RECT 111.05 54.765 111.26 54.835 ;
    RECT 111.05 55.125 111.26 55.195 ;
    RECT 111.05 55.485 111.26 55.555 ;
    RECT 111.51 54.765 111.72 54.835 ;
    RECT 111.51 55.125 111.72 55.195 ;
    RECT 111.51 55.485 111.72 55.555 ;
    RECT 107.73 54.765 107.94 54.835 ;
    RECT 107.73 55.125 107.94 55.195 ;
    RECT 107.73 55.485 107.94 55.555 ;
    RECT 108.19 54.765 108.4 54.835 ;
    RECT 108.19 55.125 108.4 55.195 ;
    RECT 108.19 55.485 108.4 55.555 ;
    RECT 104.41 54.765 104.62 54.835 ;
    RECT 104.41 55.125 104.62 55.195 ;
    RECT 104.41 55.485 104.62 55.555 ;
    RECT 104.87 54.765 105.08 54.835 ;
    RECT 104.87 55.125 105.08 55.195 ;
    RECT 104.87 55.485 105.08 55.555 ;
    RECT 101.09 54.765 101.3 54.835 ;
    RECT 101.09 55.125 101.3 55.195 ;
    RECT 101.09 55.485 101.3 55.555 ;
    RECT 101.55 54.765 101.76 54.835 ;
    RECT 101.55 55.125 101.76 55.195 ;
    RECT 101.55 55.485 101.76 55.555 ;
    RECT 0.4 55.125 0.47 55.195 ;
    RECT 170.81 54.765 171.02 54.835 ;
    RECT 170.81 55.125 171.02 55.195 ;
    RECT 170.81 55.485 171.02 55.555 ;
    RECT 171.27 54.765 171.48 54.835 ;
    RECT 171.27 55.125 171.48 55.195 ;
    RECT 171.27 55.485 171.48 55.555 ;
    RECT 167.49 54.765 167.7 54.835 ;
    RECT 167.49 55.125 167.7 55.195 ;
    RECT 167.49 55.485 167.7 55.555 ;
    RECT 167.95 54.765 168.16 54.835 ;
    RECT 167.95 55.125 168.16 55.195 ;
    RECT 167.95 55.485 168.16 55.555 ;
    RECT 97.77 54.765 97.98 54.835 ;
    RECT 97.77 55.125 97.98 55.195 ;
    RECT 97.77 55.485 97.98 55.555 ;
    RECT 98.23 54.765 98.44 54.835 ;
    RECT 98.23 55.125 98.44 55.195 ;
    RECT 98.23 55.485 98.44 55.555 ;
    RECT 94.45 54.765 94.66 54.835 ;
    RECT 94.45 55.125 94.66 55.195 ;
    RECT 94.45 55.485 94.66 55.555 ;
    RECT 94.91 54.765 95.12 54.835 ;
    RECT 94.91 55.125 95.12 55.195 ;
    RECT 94.91 55.485 95.12 55.555 ;
    RECT 91.13 54.765 91.34 54.835 ;
    RECT 91.13 55.125 91.34 55.195 ;
    RECT 91.13 55.485 91.34 55.555 ;
    RECT 91.59 54.765 91.8 54.835 ;
    RECT 91.59 55.125 91.8 55.195 ;
    RECT 91.59 55.485 91.8 55.555 ;
    RECT 87.81 54.765 88.02 54.835 ;
    RECT 87.81 55.125 88.02 55.195 ;
    RECT 87.81 55.485 88.02 55.555 ;
    RECT 88.27 54.765 88.48 54.835 ;
    RECT 88.27 55.125 88.48 55.195 ;
    RECT 88.27 55.485 88.48 55.555 ;
    RECT 84.49 54.765 84.7 54.835 ;
    RECT 84.49 55.125 84.7 55.195 ;
    RECT 84.49 55.485 84.7 55.555 ;
    RECT 84.95 54.765 85.16 54.835 ;
    RECT 84.95 55.125 85.16 55.195 ;
    RECT 84.95 55.485 85.16 55.555 ;
    RECT 81.17 54.765 81.38 54.835 ;
    RECT 81.17 55.125 81.38 55.195 ;
    RECT 81.17 55.485 81.38 55.555 ;
    RECT 81.63 54.765 81.84 54.835 ;
    RECT 81.63 55.125 81.84 55.195 ;
    RECT 81.63 55.485 81.84 55.555 ;
    RECT 77.85 54.765 78.06 54.835 ;
    RECT 77.85 55.125 78.06 55.195 ;
    RECT 77.85 55.485 78.06 55.555 ;
    RECT 78.31 54.765 78.52 54.835 ;
    RECT 78.31 55.125 78.52 55.195 ;
    RECT 78.31 55.485 78.52 55.555 ;
    RECT 74.53 54.765 74.74 54.835 ;
    RECT 74.53 55.125 74.74 55.195 ;
    RECT 74.53 55.485 74.74 55.555 ;
    RECT 74.99 54.765 75.2 54.835 ;
    RECT 74.99 55.125 75.2 55.195 ;
    RECT 74.99 55.485 75.2 55.555 ;
    RECT 71.21 54.765 71.42 54.835 ;
    RECT 71.21 55.125 71.42 55.195 ;
    RECT 71.21 55.485 71.42 55.555 ;
    RECT 71.67 54.765 71.88 54.835 ;
    RECT 71.67 55.125 71.88 55.195 ;
    RECT 71.67 55.485 71.88 55.555 ;
    RECT 31.37 54.765 31.58 54.835 ;
    RECT 31.37 55.125 31.58 55.195 ;
    RECT 31.37 55.485 31.58 55.555 ;
    RECT 31.83 54.765 32.04 54.835 ;
    RECT 31.83 55.125 32.04 55.195 ;
    RECT 31.83 55.485 32.04 55.555 ;
    RECT 67.89 54.765 68.1 54.835 ;
    RECT 67.89 55.125 68.1 55.195 ;
    RECT 67.89 55.485 68.1 55.555 ;
    RECT 68.35 54.765 68.56 54.835 ;
    RECT 68.35 55.125 68.56 55.195 ;
    RECT 68.35 55.485 68.56 55.555 ;
    RECT 28.05 54.765 28.26 54.835 ;
    RECT 28.05 55.125 28.26 55.195 ;
    RECT 28.05 55.485 28.26 55.555 ;
    RECT 28.51 54.765 28.72 54.835 ;
    RECT 28.51 55.125 28.72 55.195 ;
    RECT 28.51 55.485 28.72 55.555 ;
    RECT 24.73 54.765 24.94 54.835 ;
    RECT 24.73 55.125 24.94 55.195 ;
    RECT 24.73 55.485 24.94 55.555 ;
    RECT 25.19 54.765 25.4 54.835 ;
    RECT 25.19 55.125 25.4 55.195 ;
    RECT 25.19 55.485 25.4 55.555 ;
    RECT 21.41 54.765 21.62 54.835 ;
    RECT 21.41 55.125 21.62 55.195 ;
    RECT 21.41 55.485 21.62 55.555 ;
    RECT 21.87 54.765 22.08 54.835 ;
    RECT 21.87 55.125 22.08 55.195 ;
    RECT 21.87 55.485 22.08 55.555 ;
    RECT 18.09 54.765 18.3 54.835 ;
    RECT 18.09 55.125 18.3 55.195 ;
    RECT 18.09 55.485 18.3 55.555 ;
    RECT 18.55 54.765 18.76 54.835 ;
    RECT 18.55 55.125 18.76 55.195 ;
    RECT 18.55 55.485 18.76 55.555 ;
    RECT 14.77 54.765 14.98 54.835 ;
    RECT 14.77 55.125 14.98 55.195 ;
    RECT 14.77 55.485 14.98 55.555 ;
    RECT 15.23 54.765 15.44 54.835 ;
    RECT 15.23 55.125 15.44 55.195 ;
    RECT 15.23 55.485 15.44 55.555 ;
    RECT 11.45 54.765 11.66 54.835 ;
    RECT 11.45 55.125 11.66 55.195 ;
    RECT 11.45 55.485 11.66 55.555 ;
    RECT 11.91 54.765 12.12 54.835 ;
    RECT 11.91 55.125 12.12 55.195 ;
    RECT 11.91 55.485 12.12 55.555 ;
    RECT 8.13 54.765 8.34 54.835 ;
    RECT 8.13 55.125 8.34 55.195 ;
    RECT 8.13 55.485 8.34 55.555 ;
    RECT 8.59 54.765 8.8 54.835 ;
    RECT 8.59 55.125 8.8 55.195 ;
    RECT 8.59 55.485 8.8 55.555 ;
    RECT 4.81 54.765 5.02 54.835 ;
    RECT 4.81 55.125 5.02 55.195 ;
    RECT 4.81 55.485 5.02 55.555 ;
    RECT 5.27 54.765 5.48 54.835 ;
    RECT 5.27 55.125 5.48 55.195 ;
    RECT 5.27 55.485 5.48 55.555 ;
    RECT 164.17 54.765 164.38 54.835 ;
    RECT 164.17 55.125 164.38 55.195 ;
    RECT 164.17 55.485 164.38 55.555 ;
    RECT 164.63 54.765 164.84 54.835 ;
    RECT 164.63 55.125 164.84 55.195 ;
    RECT 164.63 55.485 164.84 55.555 ;
    RECT 1.49 54.765 1.7 54.835 ;
    RECT 1.49 55.125 1.7 55.195 ;
    RECT 1.49 55.485 1.7 55.555 ;
    RECT 1.95 54.765 2.16 54.835 ;
    RECT 1.95 55.125 2.16 55.195 ;
    RECT 1.95 55.485 2.16 55.555 ;
    RECT 160.85 54.765 161.06 54.835 ;
    RECT 160.85 55.125 161.06 55.195 ;
    RECT 160.85 55.485 161.06 55.555 ;
    RECT 161.31 54.765 161.52 54.835 ;
    RECT 161.31 55.125 161.52 55.195 ;
    RECT 161.31 55.485 161.52 55.555 ;
    RECT 157.53 54.765 157.74 54.835 ;
    RECT 157.53 55.125 157.74 55.195 ;
    RECT 157.53 55.485 157.74 55.555 ;
    RECT 157.99 54.765 158.2 54.835 ;
    RECT 157.99 55.125 158.2 55.195 ;
    RECT 157.99 55.485 158.2 55.555 ;
    RECT 154.21 54.765 154.42 54.835 ;
    RECT 154.21 55.125 154.42 55.195 ;
    RECT 154.21 55.485 154.42 55.555 ;
    RECT 154.67 54.765 154.88 54.835 ;
    RECT 154.67 55.125 154.88 55.195 ;
    RECT 154.67 55.485 154.88 55.555 ;
    RECT 150.89 54.765 151.1 54.835 ;
    RECT 150.89 55.125 151.1 55.195 ;
    RECT 150.89 55.485 151.1 55.555 ;
    RECT 151.35 54.765 151.56 54.835 ;
    RECT 151.35 55.125 151.56 55.195 ;
    RECT 151.35 55.485 151.56 55.555 ;
    RECT 147.57 54.765 147.78 54.835 ;
    RECT 147.57 55.125 147.78 55.195 ;
    RECT 147.57 55.485 147.78 55.555 ;
    RECT 148.03 54.765 148.24 54.835 ;
    RECT 148.03 55.125 148.24 55.195 ;
    RECT 148.03 55.485 148.24 55.555 ;
    RECT 144.25 54.765 144.46 54.835 ;
    RECT 144.25 55.125 144.46 55.195 ;
    RECT 144.25 55.485 144.46 55.555 ;
    RECT 144.71 54.765 144.92 54.835 ;
    RECT 144.71 55.125 144.92 55.195 ;
    RECT 144.71 55.485 144.92 55.555 ;
    RECT 140.93 54.765 141.14 54.835 ;
    RECT 140.93 55.125 141.14 55.195 ;
    RECT 140.93 55.485 141.14 55.555 ;
    RECT 141.39 54.765 141.6 54.835 ;
    RECT 141.39 55.125 141.6 55.195 ;
    RECT 141.39 55.485 141.6 55.555 ;
    RECT 137.61 54.765 137.82 54.835 ;
    RECT 137.61 55.125 137.82 55.195 ;
    RECT 137.61 55.485 137.82 55.555 ;
    RECT 138.07 54.765 138.28 54.835 ;
    RECT 138.07 55.125 138.28 55.195 ;
    RECT 138.07 55.485 138.28 55.555 ;
    RECT 134.29 54.765 134.5 54.835 ;
    RECT 134.29 55.125 134.5 55.195 ;
    RECT 134.29 55.485 134.5 55.555 ;
    RECT 134.75 54.765 134.96 54.835 ;
    RECT 134.75 55.125 134.96 55.195 ;
    RECT 134.75 55.485 134.96 55.555 ;
    RECT 64.57 54.765 64.78 54.835 ;
    RECT 64.57 55.125 64.78 55.195 ;
    RECT 64.57 55.485 64.78 55.555 ;
    RECT 65.03 54.765 65.24 54.835 ;
    RECT 65.03 55.125 65.24 55.195 ;
    RECT 65.03 55.485 65.24 55.555 ;
    RECT 19.04 59.865 19.25 59.935 ;
    RECT 131.92 59.865 132.13 59.935 ;
    RECT 104.87 59.345 105.08 59.415 ;
    RECT 104.41 59.345 104.62 59.415 ;
    RECT 141.88 59.605 142.09 59.675 ;
    RECT 48.43 59.345 48.64 59.415 ;
    RECT 47.97 59.345 48.18 59.415 ;
    RECT 98.72 59.605 98.93 59.675 ;
    RECT 164.63 59.345 164.84 59.415 ;
    RECT 164.17 59.345 164.38 59.415 ;
    RECT 15.72 59.865 15.93 59.935 ;
    RECT 128.6 59.865 128.81 59.935 ;
    RECT 101.55 59.345 101.76 59.415 ;
    RECT 101.09 59.345 101.3 59.415 ;
    RECT 138.56 59.605 138.77 59.675 ;
    RECT 45.11 59.345 45.32 59.415 ;
    RECT 44.65 59.345 44.86 59.415 ;
    RECT 95.4 59.605 95.61 59.675 ;
    RECT 161.31 59.345 161.52 59.415 ;
    RECT 160.85 59.345 161.06 59.415 ;
    RECT 12.4 59.865 12.61 59.935 ;
    RECT 65.52 59.865 65.73 59.935 ;
    RECT 135.24 59.605 135.45 59.675 ;
    RECT 75.48 59.605 75.69 59.675 ;
    RECT 41.79 59.345 42.0 59.415 ;
    RECT 41.33 59.345 41.54 59.415 ;
    RECT 92.08 59.605 92.29 59.675 ;
    RECT 125.28 59.865 125.49 59.935 ;
    RECT 157.99 59.345 158.2 59.415 ;
    RECT 157.53 59.345 157.74 59.415 ;
    RECT 9.08 59.865 9.29 59.935 ;
    RECT 62.2 59.865 62.41 59.935 ;
    RECT 31.83 59.345 32.04 59.415 ;
    RECT 31.37 59.345 31.58 59.415 ;
    RECT 72.16 59.605 72.37 59.675 ;
    RECT 88.76 59.605 88.97 59.675 ;
    RECT 121.96 59.865 122.17 59.935 ;
    RECT 5.76 59.865 5.97 59.935 ;
    RECT 38.47 59.345 38.68 59.415 ;
    RECT 38.01 59.345 38.22 59.415 ;
    RECT 28.51 59.345 28.72 59.415 ;
    RECT 28.05 59.345 28.26 59.415 ;
    RECT 154.67 59.345 154.88 59.415 ;
    RECT 68.84 59.605 69.05 59.675 ;
    RECT 154.21 59.345 154.42 59.415 ;
    RECT 98.23 59.345 98.44 59.415 ;
    RECT 97.77 59.345 97.98 59.415 ;
    RECT 85.44 59.605 85.65 59.675 ;
    RECT 118.64 59.865 118.85 59.935 ;
    RECT 58.88 59.865 59.09 59.935 ;
    RECT 2.44 59.865 2.65 59.935 ;
    RECT 35.15 59.345 35.36 59.415 ;
    RECT 34.69 59.345 34.9 59.415 ;
    RECT 25.19 59.345 25.4 59.415 ;
    RECT 30.905 60.125 31.125 60.195 ;
    RECT 24.73 59.345 24.94 59.415 ;
    RECT 27.585 60.125 27.805 60.195 ;
    RECT 24.265 60.125 24.485 60.195 ;
    RECT 151.35 59.345 151.56 59.415 ;
    RECT 20.945 60.125 21.165 60.195 ;
    RECT 150.89 59.345 151.1 59.415 ;
    RECT 17.625 60.125 17.845 60.195 ;
    RECT 14.305 60.125 14.525 60.195 ;
    RECT 10.985 60.125 11.205 60.195 ;
    RECT 94.91 59.345 95.12 59.415 ;
    RECT 7.665 60.125 7.885 60.195 ;
    RECT 94.45 59.345 94.66 59.415 ;
    RECT 165.12 59.865 165.33 59.935 ;
    RECT 4.345 60.125 4.565 60.195 ;
    RECT 82.12 59.605 82.33 59.675 ;
    RECT 1.025 60.125 1.245 60.195 ;
    RECT 115.32 59.865 115.53 59.935 ;
    RECT 55.56 59.865 55.77 59.935 ;
    RECT 131.92 59.605 132.13 59.675 ;
    RECT 32.32 59.605 32.53 59.675 ;
    RECT 148.03 59.345 148.24 59.415 ;
    RECT 147.57 59.345 147.78 59.415 ;
    RECT 91.59 59.345 91.8 59.415 ;
    RECT 161.8 59.865 162.01 59.935 ;
    RECT 91.13 59.345 91.34 59.415 ;
    RECT 78.8 59.605 79.01 59.675 ;
    RECT 171.76 59.865 171.97 59.935 ;
    RECT 112.0 59.865 112.21 59.935 ;
    RECT 52.24 59.865 52.45 59.935 ;
    RECT 170.345 60.125 170.565 60.195 ;
    RECT 167.025 60.125 167.245 60.195 ;
    RECT 128.6 59.605 128.81 59.675 ;
    RECT 29.0 59.605 29.21 59.675 ;
    RECT 21.87 59.345 22.08 59.415 ;
    RECT 21.41 59.345 21.62 59.415 ;
    RECT 163.705 60.125 163.925 60.195 ;
    RECT 160.385 60.125 160.605 60.195 ;
    RECT 157.065 60.125 157.285 60.195 ;
    RECT 153.745 60.125 153.965 60.195 ;
    RECT 150.425 60.125 150.645 60.195 ;
    RECT 144.71 59.345 144.92 59.415 ;
    RECT 147.105 60.125 147.325 60.195 ;
    RECT 144.25 59.345 144.46 59.415 ;
    RECT 143.785 60.125 144.005 60.195 ;
    RECT 140.465 60.125 140.685 60.195 ;
    RECT 137.145 60.125 137.365 60.195 ;
    RECT 98.72 59.865 98.93 59.935 ;
    RECT 168.44 59.865 168.65 59.935 ;
    RECT 133.825 60.125 134.045 60.195 ;
    RECT 108.68 59.865 108.89 59.935 ;
    RECT 48.92 59.865 49.13 59.935 ;
    RECT 125.28 59.605 125.49 59.675 ;
    RECT 65.52 59.605 65.73 59.675 ;
    RECT 158.48 59.865 158.69 59.935 ;
    RECT 88.27 59.345 88.48 59.415 ;
    RECT 87.81 59.345 88.02 59.415 ;
    RECT 130.505 60.125 130.725 60.195 ;
    RECT 25.68 59.605 25.89 59.675 ;
    RECT 127.185 60.125 127.405 60.195 ;
    RECT 123.865 60.125 124.085 60.195 ;
    RECT 120.545 60.125 120.765 60.195 ;
    RECT 18.55 59.345 18.76 59.415 ;
    RECT 117.225 60.125 117.445 60.195 ;
    RECT 18.09 59.345 18.3 59.415 ;
    RECT 113.905 60.125 114.125 60.195 ;
    RECT 110.585 60.125 110.805 60.195 ;
    RECT 107.265 60.125 107.485 60.195 ;
    RECT 103.945 60.125 104.165 60.195 ;
    RECT 100.625 60.125 100.845 60.195 ;
    RECT 141.39 59.345 141.6 59.415 ;
    RECT 140.93 59.345 141.14 59.415 ;
    RECT 95.4 59.865 95.61 59.935 ;
    RECT 105.36 59.865 105.57 59.935 ;
    RECT 45.6 59.865 45.81 59.935 ;
    RECT 121.96 59.605 122.17 59.675 ;
    RECT 97.305 60.125 97.525 60.195 ;
    RECT 131.43 59.345 131.64 59.415 ;
    RECT 62.2 59.605 62.41 59.675 ;
    RECT 93.985 60.125 94.205 60.195 ;
    RECT 130.97 59.345 131.18 59.415 ;
    RECT 155.16 59.865 155.37 59.935 ;
    RECT 90.665 60.125 90.885 60.195 ;
    RECT 87.345 60.125 87.565 60.195 ;
    RECT 84.95 59.345 85.16 59.415 ;
    RECT 84.025 60.125 84.245 60.195 ;
    RECT 84.49 59.345 84.7 59.415 ;
    RECT 22.36 59.605 22.57 59.675 ;
    RECT 80.705 60.125 80.925 60.195 ;
    RECT 77.385 60.125 77.605 60.195 ;
    RECT 74.065 60.125 74.285 60.195 ;
    RECT 70.745 60.125 70.965 60.195 ;
    RECT 15.23 59.345 15.44 59.415 ;
    RECT 67.425 60.125 67.645 60.195 ;
    RECT 14.77 59.345 14.98 59.415 ;
    RECT 102.04 59.865 102.25 59.935 ;
    RECT 42.28 59.865 42.49 59.935 ;
    RECT 64.105 60.125 64.325 60.195 ;
    RECT 60.785 60.125 61.005 60.195 ;
    RECT 57.465 60.125 57.685 60.195 ;
    RECT 54.145 60.125 54.365 60.195 ;
    RECT 118.64 59.605 118.85 59.675 ;
    RECT 50.825 60.125 51.045 60.195 ;
    RECT 138.07 59.345 138.28 59.415 ;
    RECT 58.88 59.605 59.09 59.675 ;
    RECT 47.505 60.125 47.725 60.195 ;
    RECT 137.61 59.345 137.82 59.415 ;
    RECT 128.11 59.345 128.32 59.415 ;
    RECT 151.84 59.865 152.05 59.935 ;
    RECT 44.185 60.125 44.405 60.195 ;
    RECT 127.65 59.345 127.86 59.415 ;
    RECT 92.08 59.865 92.29 59.935 ;
    RECT 40.865 60.125 41.085 60.195 ;
    RECT 37.545 60.125 37.765 60.195 ;
    RECT 81.63 59.345 81.84 59.415 ;
    RECT 19.04 59.605 19.25 59.675 ;
    RECT 34.225 60.125 34.445 60.195 ;
    RECT 81.17 59.345 81.38 59.415 ;
    RECT 11.91 59.345 12.12 59.415 ;
    RECT 11.45 59.345 11.66 59.415 ;
    RECT 38.96 59.865 39.17 59.935 ;
    RECT 115.32 59.605 115.53 59.675 ;
    RECT 55.56 59.605 55.77 59.675 ;
    RECT 134.75 59.345 134.96 59.415 ;
    RECT 148.52 59.865 148.73 59.935 ;
    RECT 124.79 59.345 125.0 59.415 ;
    RECT 134.29 59.345 134.5 59.415 ;
    RECT 88.76 59.865 88.97 59.935 ;
    RECT 124.33 59.345 124.54 59.415 ;
    RECT 15.72 59.605 15.93 59.675 ;
    RECT 78.31 59.345 78.52 59.415 ;
    RECT 77.85 59.345 78.06 59.415 ;
    RECT 8.59 59.345 8.8 59.415 ;
    RECT 8.13 59.345 8.34 59.415 ;
    RECT 165.12 59.605 165.33 59.675 ;
    RECT 35.64 59.865 35.85 59.935 ;
    RECT 171.76 59.605 171.97 59.675 ;
    RECT 112.0 59.605 112.21 59.675 ;
    RECT 52.24 59.605 52.45 59.675 ;
    RECT 145.2 59.865 145.41 59.935 ;
    RECT 85.44 59.865 85.65 59.935 ;
    RECT 12.4 59.605 12.61 59.675 ;
    RECT 74.99 59.345 75.2 59.415 ;
    RECT 74.53 59.345 74.74 59.415 ;
    RECT 161.8 59.605 162.01 59.675 ;
    RECT 121.47 59.345 121.68 59.415 ;
    RECT 121.01 59.345 121.22 59.415 ;
    RECT 65.03 59.345 65.24 59.415 ;
    RECT 64.57 59.345 64.78 59.415 ;
    RECT 168.44 59.605 168.65 59.675 ;
    RECT 5.27 59.345 5.48 59.415 ;
    RECT 108.68 59.605 108.89 59.675 ;
    RECT 4.81 59.345 5.02 59.415 ;
    RECT 48.92 59.605 49.13 59.675 ;
    RECT 141.88 59.865 142.09 59.935 ;
    RECT 82.12 59.865 82.33 59.935 ;
    RECT 9.08 59.605 9.29 59.675 ;
    RECT 32.32 59.865 32.53 59.935 ;
    RECT 158.48 59.605 158.69 59.675 ;
    RECT 118.15 59.345 118.36 59.415 ;
    RECT 117.69 59.345 117.9 59.415 ;
    RECT 71.67 59.345 71.88 59.415 ;
    RECT 61.71 59.345 61.92 59.415 ;
    RECT 71.21 59.345 71.42 59.415 ;
    RECT 61.25 59.345 61.46 59.415 ;
    RECT 105.36 59.605 105.57 59.675 ;
    RECT 1.95 59.345 2.16 59.415 ;
    RECT 45.6 59.605 45.81 59.675 ;
    RECT 1.49 59.345 1.7 59.415 ;
    RECT 138.56 59.865 138.77 59.935 ;
    RECT 78.8 59.865 79.01 59.935 ;
    RECT 5.76 59.605 5.97 59.675 ;
    RECT 29.0 59.865 29.21 59.935 ;
    RECT 155.16 59.605 155.37 59.675 ;
    RECT 171.27 59.345 171.48 59.415 ;
    RECT 170.81 59.345 171.02 59.415 ;
    RECT 114.83 59.345 115.04 59.415 ;
    RECT 114.37 59.345 114.58 59.415 ;
    RECT 68.35 59.345 68.56 59.415 ;
    RECT 58.39 59.345 58.6 59.415 ;
    RECT 67.89 59.345 68.1 59.415 ;
    RECT 57.93 59.345 58.14 59.415 ;
    RECT 102.04 59.605 102.25 59.675 ;
    RECT 42.28 59.605 42.49 59.675 ;
    RECT 135.24 59.865 135.45 59.935 ;
    RECT 75.48 59.865 75.69 59.935 ;
    RECT 2.44 59.605 2.65 59.675 ;
    RECT 151.84 59.605 152.05 59.675 ;
    RECT 167.95 59.345 168.16 59.415 ;
    RECT 167.49 59.345 167.7 59.415 ;
    RECT 111.51 59.345 111.72 59.415 ;
    RECT 111.05 59.345 111.26 59.415 ;
    RECT 38.96 59.605 39.17 59.675 ;
    RECT 25.68 59.865 25.89 59.935 ;
    RECT 72.16 59.865 72.37 59.935 ;
    RECT 174.155 59.605 174.225 59.675 ;
    RECT 173.945 59.345 174.015 59.415 ;
    RECT 55.07 59.345 55.28 59.415 ;
    RECT 148.52 59.605 148.73 59.675 ;
    RECT 54.61 59.345 54.82 59.415 ;
    RECT 0.19 59.605 0.26 59.675 ;
    RECT 0.4 59.345 0.47 59.415 ;
    RECT 108.19 59.345 108.4 59.415 ;
    RECT 107.73 59.345 107.94 59.415 ;
    RECT 35.64 59.605 35.85 59.675 ;
    RECT 22.36 59.865 22.57 59.935 ;
    RECT 68.84 59.865 69.05 59.935 ;
    RECT 145.2 59.605 145.41 59.675 ;
    RECT 51.75 59.345 51.96 59.415 ;
    RECT 51.29 59.345 51.5 59.415 ;
    RECT 61.25 33.885 61.46 33.955 ;
    RECT 61.25 34.245 61.46 34.315 ;
    RECT 61.25 34.605 61.46 34.675 ;
    RECT 61.71 33.885 61.92 33.955 ;
    RECT 61.71 34.245 61.92 34.315 ;
    RECT 61.71 34.605 61.92 34.675 ;
    RECT 57.93 33.885 58.14 33.955 ;
    RECT 57.93 34.245 58.14 34.315 ;
    RECT 57.93 34.605 58.14 34.675 ;
    RECT 58.39 33.885 58.6 33.955 ;
    RECT 58.39 34.245 58.6 34.315 ;
    RECT 58.39 34.605 58.6 34.675 ;
    RECT 54.61 33.885 54.82 33.955 ;
    RECT 54.61 34.245 54.82 34.315 ;
    RECT 54.61 34.605 54.82 34.675 ;
    RECT 55.07 33.885 55.28 33.955 ;
    RECT 55.07 34.245 55.28 34.315 ;
    RECT 55.07 34.605 55.28 34.675 ;
    RECT 51.29 33.885 51.5 33.955 ;
    RECT 51.29 34.245 51.5 34.315 ;
    RECT 51.29 34.605 51.5 34.675 ;
    RECT 51.75 33.885 51.96 33.955 ;
    RECT 51.75 34.245 51.96 34.315 ;
    RECT 51.75 34.605 51.96 34.675 ;
    RECT 47.97 33.885 48.18 33.955 ;
    RECT 47.97 34.245 48.18 34.315 ;
    RECT 47.97 34.605 48.18 34.675 ;
    RECT 48.43 33.885 48.64 33.955 ;
    RECT 48.43 34.245 48.64 34.315 ;
    RECT 48.43 34.605 48.64 34.675 ;
    RECT 44.65 33.885 44.86 33.955 ;
    RECT 44.65 34.245 44.86 34.315 ;
    RECT 44.65 34.605 44.86 34.675 ;
    RECT 45.11 33.885 45.32 33.955 ;
    RECT 45.11 34.245 45.32 34.315 ;
    RECT 45.11 34.605 45.32 34.675 ;
    RECT 41.33 33.885 41.54 33.955 ;
    RECT 41.33 34.245 41.54 34.315 ;
    RECT 41.33 34.605 41.54 34.675 ;
    RECT 41.79 33.885 42.0 33.955 ;
    RECT 41.79 34.245 42.0 34.315 ;
    RECT 41.79 34.605 42.0 34.675 ;
    RECT 38.01 33.885 38.22 33.955 ;
    RECT 38.01 34.245 38.22 34.315 ;
    RECT 38.01 34.605 38.22 34.675 ;
    RECT 38.47 33.885 38.68 33.955 ;
    RECT 38.47 34.245 38.68 34.315 ;
    RECT 38.47 34.605 38.68 34.675 ;
    RECT 34.69 33.885 34.9 33.955 ;
    RECT 34.69 34.245 34.9 34.315 ;
    RECT 34.69 34.605 34.9 34.675 ;
    RECT 35.15 33.885 35.36 33.955 ;
    RECT 35.15 34.245 35.36 34.315 ;
    RECT 35.15 34.605 35.36 34.675 ;
    RECT 173.945 34.245 174.015 34.315 ;
    RECT 130.97 33.885 131.18 33.955 ;
    RECT 130.97 34.245 131.18 34.315 ;
    RECT 130.97 34.605 131.18 34.675 ;
    RECT 131.43 33.885 131.64 33.955 ;
    RECT 131.43 34.245 131.64 34.315 ;
    RECT 131.43 34.605 131.64 34.675 ;
    RECT 127.65 33.885 127.86 33.955 ;
    RECT 127.65 34.245 127.86 34.315 ;
    RECT 127.65 34.605 127.86 34.675 ;
    RECT 128.11 33.885 128.32 33.955 ;
    RECT 128.11 34.245 128.32 34.315 ;
    RECT 128.11 34.605 128.32 34.675 ;
    RECT 124.33 33.885 124.54 33.955 ;
    RECT 124.33 34.245 124.54 34.315 ;
    RECT 124.33 34.605 124.54 34.675 ;
    RECT 124.79 33.885 125.0 33.955 ;
    RECT 124.79 34.245 125.0 34.315 ;
    RECT 124.79 34.605 125.0 34.675 ;
    RECT 121.01 33.885 121.22 33.955 ;
    RECT 121.01 34.245 121.22 34.315 ;
    RECT 121.01 34.605 121.22 34.675 ;
    RECT 121.47 33.885 121.68 33.955 ;
    RECT 121.47 34.245 121.68 34.315 ;
    RECT 121.47 34.605 121.68 34.675 ;
    RECT 117.69 33.885 117.9 33.955 ;
    RECT 117.69 34.245 117.9 34.315 ;
    RECT 117.69 34.605 117.9 34.675 ;
    RECT 118.15 33.885 118.36 33.955 ;
    RECT 118.15 34.245 118.36 34.315 ;
    RECT 118.15 34.605 118.36 34.675 ;
    RECT 114.37 33.885 114.58 33.955 ;
    RECT 114.37 34.245 114.58 34.315 ;
    RECT 114.37 34.605 114.58 34.675 ;
    RECT 114.83 33.885 115.04 33.955 ;
    RECT 114.83 34.245 115.04 34.315 ;
    RECT 114.83 34.605 115.04 34.675 ;
    RECT 111.05 33.885 111.26 33.955 ;
    RECT 111.05 34.245 111.26 34.315 ;
    RECT 111.05 34.605 111.26 34.675 ;
    RECT 111.51 33.885 111.72 33.955 ;
    RECT 111.51 34.245 111.72 34.315 ;
    RECT 111.51 34.605 111.72 34.675 ;
    RECT 107.73 33.885 107.94 33.955 ;
    RECT 107.73 34.245 107.94 34.315 ;
    RECT 107.73 34.605 107.94 34.675 ;
    RECT 108.19 33.885 108.4 33.955 ;
    RECT 108.19 34.245 108.4 34.315 ;
    RECT 108.19 34.605 108.4 34.675 ;
    RECT 104.41 33.885 104.62 33.955 ;
    RECT 104.41 34.245 104.62 34.315 ;
    RECT 104.41 34.605 104.62 34.675 ;
    RECT 104.87 33.885 105.08 33.955 ;
    RECT 104.87 34.245 105.08 34.315 ;
    RECT 104.87 34.605 105.08 34.675 ;
    RECT 101.09 33.885 101.3 33.955 ;
    RECT 101.09 34.245 101.3 34.315 ;
    RECT 101.09 34.605 101.3 34.675 ;
    RECT 101.55 33.885 101.76 33.955 ;
    RECT 101.55 34.245 101.76 34.315 ;
    RECT 101.55 34.605 101.76 34.675 ;
    RECT 0.4 34.245 0.47 34.315 ;
    RECT 170.81 33.885 171.02 33.955 ;
    RECT 170.81 34.245 171.02 34.315 ;
    RECT 170.81 34.605 171.02 34.675 ;
    RECT 171.27 33.885 171.48 33.955 ;
    RECT 171.27 34.245 171.48 34.315 ;
    RECT 171.27 34.605 171.48 34.675 ;
    RECT 167.49 33.885 167.7 33.955 ;
    RECT 167.49 34.245 167.7 34.315 ;
    RECT 167.49 34.605 167.7 34.675 ;
    RECT 167.95 33.885 168.16 33.955 ;
    RECT 167.95 34.245 168.16 34.315 ;
    RECT 167.95 34.605 168.16 34.675 ;
    RECT 97.77 33.885 97.98 33.955 ;
    RECT 97.77 34.245 97.98 34.315 ;
    RECT 97.77 34.605 97.98 34.675 ;
    RECT 98.23 33.885 98.44 33.955 ;
    RECT 98.23 34.245 98.44 34.315 ;
    RECT 98.23 34.605 98.44 34.675 ;
    RECT 94.45 33.885 94.66 33.955 ;
    RECT 94.45 34.245 94.66 34.315 ;
    RECT 94.45 34.605 94.66 34.675 ;
    RECT 94.91 33.885 95.12 33.955 ;
    RECT 94.91 34.245 95.12 34.315 ;
    RECT 94.91 34.605 95.12 34.675 ;
    RECT 91.13 33.885 91.34 33.955 ;
    RECT 91.13 34.245 91.34 34.315 ;
    RECT 91.13 34.605 91.34 34.675 ;
    RECT 91.59 33.885 91.8 33.955 ;
    RECT 91.59 34.245 91.8 34.315 ;
    RECT 91.59 34.605 91.8 34.675 ;
    RECT 87.81 33.885 88.02 33.955 ;
    RECT 87.81 34.245 88.02 34.315 ;
    RECT 87.81 34.605 88.02 34.675 ;
    RECT 88.27 33.885 88.48 33.955 ;
    RECT 88.27 34.245 88.48 34.315 ;
    RECT 88.27 34.605 88.48 34.675 ;
    RECT 84.49 33.885 84.7 33.955 ;
    RECT 84.49 34.245 84.7 34.315 ;
    RECT 84.49 34.605 84.7 34.675 ;
    RECT 84.95 33.885 85.16 33.955 ;
    RECT 84.95 34.245 85.16 34.315 ;
    RECT 84.95 34.605 85.16 34.675 ;
    RECT 81.17 33.885 81.38 33.955 ;
    RECT 81.17 34.245 81.38 34.315 ;
    RECT 81.17 34.605 81.38 34.675 ;
    RECT 81.63 33.885 81.84 33.955 ;
    RECT 81.63 34.245 81.84 34.315 ;
    RECT 81.63 34.605 81.84 34.675 ;
    RECT 77.85 33.885 78.06 33.955 ;
    RECT 77.85 34.245 78.06 34.315 ;
    RECT 77.85 34.605 78.06 34.675 ;
    RECT 78.31 33.885 78.52 33.955 ;
    RECT 78.31 34.245 78.52 34.315 ;
    RECT 78.31 34.605 78.52 34.675 ;
    RECT 74.53 33.885 74.74 33.955 ;
    RECT 74.53 34.245 74.74 34.315 ;
    RECT 74.53 34.605 74.74 34.675 ;
    RECT 74.99 33.885 75.2 33.955 ;
    RECT 74.99 34.245 75.2 34.315 ;
    RECT 74.99 34.605 75.2 34.675 ;
    RECT 71.21 33.885 71.42 33.955 ;
    RECT 71.21 34.245 71.42 34.315 ;
    RECT 71.21 34.605 71.42 34.675 ;
    RECT 71.67 33.885 71.88 33.955 ;
    RECT 71.67 34.245 71.88 34.315 ;
    RECT 71.67 34.605 71.88 34.675 ;
    RECT 31.37 33.885 31.58 33.955 ;
    RECT 31.37 34.245 31.58 34.315 ;
    RECT 31.37 34.605 31.58 34.675 ;
    RECT 31.83 33.885 32.04 33.955 ;
    RECT 31.83 34.245 32.04 34.315 ;
    RECT 31.83 34.605 32.04 34.675 ;
    RECT 67.89 33.885 68.1 33.955 ;
    RECT 67.89 34.245 68.1 34.315 ;
    RECT 67.89 34.605 68.1 34.675 ;
    RECT 68.35 33.885 68.56 33.955 ;
    RECT 68.35 34.245 68.56 34.315 ;
    RECT 68.35 34.605 68.56 34.675 ;
    RECT 28.05 33.885 28.26 33.955 ;
    RECT 28.05 34.245 28.26 34.315 ;
    RECT 28.05 34.605 28.26 34.675 ;
    RECT 28.51 33.885 28.72 33.955 ;
    RECT 28.51 34.245 28.72 34.315 ;
    RECT 28.51 34.605 28.72 34.675 ;
    RECT 24.73 33.885 24.94 33.955 ;
    RECT 24.73 34.245 24.94 34.315 ;
    RECT 24.73 34.605 24.94 34.675 ;
    RECT 25.19 33.885 25.4 33.955 ;
    RECT 25.19 34.245 25.4 34.315 ;
    RECT 25.19 34.605 25.4 34.675 ;
    RECT 21.41 33.885 21.62 33.955 ;
    RECT 21.41 34.245 21.62 34.315 ;
    RECT 21.41 34.605 21.62 34.675 ;
    RECT 21.87 33.885 22.08 33.955 ;
    RECT 21.87 34.245 22.08 34.315 ;
    RECT 21.87 34.605 22.08 34.675 ;
    RECT 18.09 33.885 18.3 33.955 ;
    RECT 18.09 34.245 18.3 34.315 ;
    RECT 18.09 34.605 18.3 34.675 ;
    RECT 18.55 33.885 18.76 33.955 ;
    RECT 18.55 34.245 18.76 34.315 ;
    RECT 18.55 34.605 18.76 34.675 ;
    RECT 14.77 33.885 14.98 33.955 ;
    RECT 14.77 34.245 14.98 34.315 ;
    RECT 14.77 34.605 14.98 34.675 ;
    RECT 15.23 33.885 15.44 33.955 ;
    RECT 15.23 34.245 15.44 34.315 ;
    RECT 15.23 34.605 15.44 34.675 ;
    RECT 11.45 33.885 11.66 33.955 ;
    RECT 11.45 34.245 11.66 34.315 ;
    RECT 11.45 34.605 11.66 34.675 ;
    RECT 11.91 33.885 12.12 33.955 ;
    RECT 11.91 34.245 12.12 34.315 ;
    RECT 11.91 34.605 12.12 34.675 ;
    RECT 8.13 33.885 8.34 33.955 ;
    RECT 8.13 34.245 8.34 34.315 ;
    RECT 8.13 34.605 8.34 34.675 ;
    RECT 8.59 33.885 8.8 33.955 ;
    RECT 8.59 34.245 8.8 34.315 ;
    RECT 8.59 34.605 8.8 34.675 ;
    RECT 4.81 33.885 5.02 33.955 ;
    RECT 4.81 34.245 5.02 34.315 ;
    RECT 4.81 34.605 5.02 34.675 ;
    RECT 5.27 33.885 5.48 33.955 ;
    RECT 5.27 34.245 5.48 34.315 ;
    RECT 5.27 34.605 5.48 34.675 ;
    RECT 164.17 33.885 164.38 33.955 ;
    RECT 164.17 34.245 164.38 34.315 ;
    RECT 164.17 34.605 164.38 34.675 ;
    RECT 164.63 33.885 164.84 33.955 ;
    RECT 164.63 34.245 164.84 34.315 ;
    RECT 164.63 34.605 164.84 34.675 ;
    RECT 1.49 33.885 1.7 33.955 ;
    RECT 1.49 34.245 1.7 34.315 ;
    RECT 1.49 34.605 1.7 34.675 ;
    RECT 1.95 33.885 2.16 33.955 ;
    RECT 1.95 34.245 2.16 34.315 ;
    RECT 1.95 34.605 2.16 34.675 ;
    RECT 160.85 33.885 161.06 33.955 ;
    RECT 160.85 34.245 161.06 34.315 ;
    RECT 160.85 34.605 161.06 34.675 ;
    RECT 161.31 33.885 161.52 33.955 ;
    RECT 161.31 34.245 161.52 34.315 ;
    RECT 161.31 34.605 161.52 34.675 ;
    RECT 157.53 33.885 157.74 33.955 ;
    RECT 157.53 34.245 157.74 34.315 ;
    RECT 157.53 34.605 157.74 34.675 ;
    RECT 157.99 33.885 158.2 33.955 ;
    RECT 157.99 34.245 158.2 34.315 ;
    RECT 157.99 34.605 158.2 34.675 ;
    RECT 154.21 33.885 154.42 33.955 ;
    RECT 154.21 34.245 154.42 34.315 ;
    RECT 154.21 34.605 154.42 34.675 ;
    RECT 154.67 33.885 154.88 33.955 ;
    RECT 154.67 34.245 154.88 34.315 ;
    RECT 154.67 34.605 154.88 34.675 ;
    RECT 150.89 33.885 151.1 33.955 ;
    RECT 150.89 34.245 151.1 34.315 ;
    RECT 150.89 34.605 151.1 34.675 ;
    RECT 151.35 33.885 151.56 33.955 ;
    RECT 151.35 34.245 151.56 34.315 ;
    RECT 151.35 34.605 151.56 34.675 ;
    RECT 147.57 33.885 147.78 33.955 ;
    RECT 147.57 34.245 147.78 34.315 ;
    RECT 147.57 34.605 147.78 34.675 ;
    RECT 148.03 33.885 148.24 33.955 ;
    RECT 148.03 34.245 148.24 34.315 ;
    RECT 148.03 34.605 148.24 34.675 ;
    RECT 144.25 33.885 144.46 33.955 ;
    RECT 144.25 34.245 144.46 34.315 ;
    RECT 144.25 34.605 144.46 34.675 ;
    RECT 144.71 33.885 144.92 33.955 ;
    RECT 144.71 34.245 144.92 34.315 ;
    RECT 144.71 34.605 144.92 34.675 ;
    RECT 140.93 33.885 141.14 33.955 ;
    RECT 140.93 34.245 141.14 34.315 ;
    RECT 140.93 34.605 141.14 34.675 ;
    RECT 141.39 33.885 141.6 33.955 ;
    RECT 141.39 34.245 141.6 34.315 ;
    RECT 141.39 34.605 141.6 34.675 ;
    RECT 137.61 33.885 137.82 33.955 ;
    RECT 137.61 34.245 137.82 34.315 ;
    RECT 137.61 34.605 137.82 34.675 ;
    RECT 138.07 33.885 138.28 33.955 ;
    RECT 138.07 34.245 138.28 34.315 ;
    RECT 138.07 34.605 138.28 34.675 ;
    RECT 134.29 33.885 134.5 33.955 ;
    RECT 134.29 34.245 134.5 34.315 ;
    RECT 134.29 34.605 134.5 34.675 ;
    RECT 134.75 33.885 134.96 33.955 ;
    RECT 134.75 34.245 134.96 34.315 ;
    RECT 134.75 34.605 134.96 34.675 ;
    RECT 64.57 33.885 64.78 33.955 ;
    RECT 64.57 34.245 64.78 34.315 ;
    RECT 64.57 34.605 64.78 34.675 ;
    RECT 65.03 33.885 65.24 33.955 ;
    RECT 65.03 34.245 65.24 34.315 ;
    RECT 65.03 34.605 65.24 34.675 ;
    RECT 61.25 34.605 61.46 34.675 ;
    RECT 61.25 34.965 61.46 35.035 ;
    RECT 61.25 35.325 61.46 35.395 ;
    RECT 61.71 34.605 61.92 34.675 ;
    RECT 61.71 34.965 61.92 35.035 ;
    RECT 61.71 35.325 61.92 35.395 ;
    RECT 57.93 34.605 58.14 34.675 ;
    RECT 57.93 34.965 58.14 35.035 ;
    RECT 57.93 35.325 58.14 35.395 ;
    RECT 58.39 34.605 58.6 34.675 ;
    RECT 58.39 34.965 58.6 35.035 ;
    RECT 58.39 35.325 58.6 35.395 ;
    RECT 54.61 34.605 54.82 34.675 ;
    RECT 54.61 34.965 54.82 35.035 ;
    RECT 54.61 35.325 54.82 35.395 ;
    RECT 55.07 34.605 55.28 34.675 ;
    RECT 55.07 34.965 55.28 35.035 ;
    RECT 55.07 35.325 55.28 35.395 ;
    RECT 51.29 34.605 51.5 34.675 ;
    RECT 51.29 34.965 51.5 35.035 ;
    RECT 51.29 35.325 51.5 35.395 ;
    RECT 51.75 34.605 51.96 34.675 ;
    RECT 51.75 34.965 51.96 35.035 ;
    RECT 51.75 35.325 51.96 35.395 ;
    RECT 47.97 34.605 48.18 34.675 ;
    RECT 47.97 34.965 48.18 35.035 ;
    RECT 47.97 35.325 48.18 35.395 ;
    RECT 48.43 34.605 48.64 34.675 ;
    RECT 48.43 34.965 48.64 35.035 ;
    RECT 48.43 35.325 48.64 35.395 ;
    RECT 44.65 34.605 44.86 34.675 ;
    RECT 44.65 34.965 44.86 35.035 ;
    RECT 44.65 35.325 44.86 35.395 ;
    RECT 45.11 34.605 45.32 34.675 ;
    RECT 45.11 34.965 45.32 35.035 ;
    RECT 45.11 35.325 45.32 35.395 ;
    RECT 41.33 34.605 41.54 34.675 ;
    RECT 41.33 34.965 41.54 35.035 ;
    RECT 41.33 35.325 41.54 35.395 ;
    RECT 41.79 34.605 42.0 34.675 ;
    RECT 41.79 34.965 42.0 35.035 ;
    RECT 41.79 35.325 42.0 35.395 ;
    RECT 38.01 34.605 38.22 34.675 ;
    RECT 38.01 34.965 38.22 35.035 ;
    RECT 38.01 35.325 38.22 35.395 ;
    RECT 38.47 34.605 38.68 34.675 ;
    RECT 38.47 34.965 38.68 35.035 ;
    RECT 38.47 35.325 38.68 35.395 ;
    RECT 173.945 34.965 174.015 35.035 ;
    RECT 34.69 34.605 34.9 34.675 ;
    RECT 34.69 34.965 34.9 35.035 ;
    RECT 34.69 35.325 34.9 35.395 ;
    RECT 35.15 34.605 35.36 34.675 ;
    RECT 35.15 34.965 35.36 35.035 ;
    RECT 35.15 35.325 35.36 35.395 ;
    RECT 130.97 34.605 131.18 34.675 ;
    RECT 130.97 34.965 131.18 35.035 ;
    RECT 130.97 35.325 131.18 35.395 ;
    RECT 131.43 34.605 131.64 34.675 ;
    RECT 131.43 34.965 131.64 35.035 ;
    RECT 131.43 35.325 131.64 35.395 ;
    RECT 127.65 34.605 127.86 34.675 ;
    RECT 127.65 34.965 127.86 35.035 ;
    RECT 127.65 35.325 127.86 35.395 ;
    RECT 128.11 34.605 128.32 34.675 ;
    RECT 128.11 34.965 128.32 35.035 ;
    RECT 128.11 35.325 128.32 35.395 ;
    RECT 124.33 34.605 124.54 34.675 ;
    RECT 124.33 34.965 124.54 35.035 ;
    RECT 124.33 35.325 124.54 35.395 ;
    RECT 124.79 34.605 125.0 34.675 ;
    RECT 124.79 34.965 125.0 35.035 ;
    RECT 124.79 35.325 125.0 35.395 ;
    RECT 121.01 34.605 121.22 34.675 ;
    RECT 121.01 34.965 121.22 35.035 ;
    RECT 121.01 35.325 121.22 35.395 ;
    RECT 121.47 34.605 121.68 34.675 ;
    RECT 121.47 34.965 121.68 35.035 ;
    RECT 121.47 35.325 121.68 35.395 ;
    RECT 117.69 34.605 117.9 34.675 ;
    RECT 117.69 34.965 117.9 35.035 ;
    RECT 117.69 35.325 117.9 35.395 ;
    RECT 118.15 34.605 118.36 34.675 ;
    RECT 118.15 34.965 118.36 35.035 ;
    RECT 118.15 35.325 118.36 35.395 ;
    RECT 114.37 34.605 114.58 34.675 ;
    RECT 114.37 34.965 114.58 35.035 ;
    RECT 114.37 35.325 114.58 35.395 ;
    RECT 114.83 34.605 115.04 34.675 ;
    RECT 114.83 34.965 115.04 35.035 ;
    RECT 114.83 35.325 115.04 35.395 ;
    RECT 111.05 34.605 111.26 34.675 ;
    RECT 111.05 34.965 111.26 35.035 ;
    RECT 111.05 35.325 111.26 35.395 ;
    RECT 111.51 34.605 111.72 34.675 ;
    RECT 111.51 34.965 111.72 35.035 ;
    RECT 111.51 35.325 111.72 35.395 ;
    RECT 107.73 34.605 107.94 34.675 ;
    RECT 107.73 34.965 107.94 35.035 ;
    RECT 107.73 35.325 107.94 35.395 ;
    RECT 108.19 34.605 108.4 34.675 ;
    RECT 108.19 34.965 108.4 35.035 ;
    RECT 108.19 35.325 108.4 35.395 ;
    RECT 104.41 34.605 104.62 34.675 ;
    RECT 104.41 34.965 104.62 35.035 ;
    RECT 104.41 35.325 104.62 35.395 ;
    RECT 104.87 34.605 105.08 34.675 ;
    RECT 104.87 34.965 105.08 35.035 ;
    RECT 104.87 35.325 105.08 35.395 ;
    RECT 101.09 34.605 101.3 34.675 ;
    RECT 101.09 34.965 101.3 35.035 ;
    RECT 101.09 35.325 101.3 35.395 ;
    RECT 101.55 34.605 101.76 34.675 ;
    RECT 101.55 34.965 101.76 35.035 ;
    RECT 101.55 35.325 101.76 35.395 ;
    RECT 0.4 34.965 0.47 35.035 ;
    RECT 170.81 34.605 171.02 34.675 ;
    RECT 170.81 34.965 171.02 35.035 ;
    RECT 170.81 35.325 171.02 35.395 ;
    RECT 171.27 34.605 171.48 34.675 ;
    RECT 171.27 34.965 171.48 35.035 ;
    RECT 171.27 35.325 171.48 35.395 ;
    RECT 167.49 34.605 167.7 34.675 ;
    RECT 167.49 34.965 167.7 35.035 ;
    RECT 167.49 35.325 167.7 35.395 ;
    RECT 167.95 34.605 168.16 34.675 ;
    RECT 167.95 34.965 168.16 35.035 ;
    RECT 167.95 35.325 168.16 35.395 ;
    RECT 97.77 34.605 97.98 34.675 ;
    RECT 97.77 34.965 97.98 35.035 ;
    RECT 97.77 35.325 97.98 35.395 ;
    RECT 98.23 34.605 98.44 34.675 ;
    RECT 98.23 34.965 98.44 35.035 ;
    RECT 98.23 35.325 98.44 35.395 ;
    RECT 94.45 34.605 94.66 34.675 ;
    RECT 94.45 34.965 94.66 35.035 ;
    RECT 94.45 35.325 94.66 35.395 ;
    RECT 94.91 34.605 95.12 34.675 ;
    RECT 94.91 34.965 95.12 35.035 ;
    RECT 94.91 35.325 95.12 35.395 ;
    RECT 91.13 34.605 91.34 34.675 ;
    RECT 91.13 34.965 91.34 35.035 ;
    RECT 91.13 35.325 91.34 35.395 ;
    RECT 91.59 34.605 91.8 34.675 ;
    RECT 91.59 34.965 91.8 35.035 ;
    RECT 91.59 35.325 91.8 35.395 ;
    RECT 87.81 34.605 88.02 34.675 ;
    RECT 87.81 34.965 88.02 35.035 ;
    RECT 87.81 35.325 88.02 35.395 ;
    RECT 88.27 34.605 88.48 34.675 ;
    RECT 88.27 34.965 88.48 35.035 ;
    RECT 88.27 35.325 88.48 35.395 ;
    RECT 84.49 34.605 84.7 34.675 ;
    RECT 84.49 34.965 84.7 35.035 ;
    RECT 84.49 35.325 84.7 35.395 ;
    RECT 84.95 34.605 85.16 34.675 ;
    RECT 84.95 34.965 85.16 35.035 ;
    RECT 84.95 35.325 85.16 35.395 ;
    RECT 81.17 34.605 81.38 34.675 ;
    RECT 81.17 34.965 81.38 35.035 ;
    RECT 81.17 35.325 81.38 35.395 ;
    RECT 81.63 34.605 81.84 34.675 ;
    RECT 81.63 34.965 81.84 35.035 ;
    RECT 81.63 35.325 81.84 35.395 ;
    RECT 77.85 34.605 78.06 34.675 ;
    RECT 77.85 34.965 78.06 35.035 ;
    RECT 77.85 35.325 78.06 35.395 ;
    RECT 78.31 34.605 78.52 34.675 ;
    RECT 78.31 34.965 78.52 35.035 ;
    RECT 78.31 35.325 78.52 35.395 ;
    RECT 74.53 34.605 74.74 34.675 ;
    RECT 74.53 34.965 74.74 35.035 ;
    RECT 74.53 35.325 74.74 35.395 ;
    RECT 74.99 34.605 75.2 34.675 ;
    RECT 74.99 34.965 75.2 35.035 ;
    RECT 74.99 35.325 75.2 35.395 ;
    RECT 71.21 34.605 71.42 34.675 ;
    RECT 71.21 34.965 71.42 35.035 ;
    RECT 71.21 35.325 71.42 35.395 ;
    RECT 71.67 34.605 71.88 34.675 ;
    RECT 71.67 34.965 71.88 35.035 ;
    RECT 71.67 35.325 71.88 35.395 ;
    RECT 31.37 34.605 31.58 34.675 ;
    RECT 31.37 34.965 31.58 35.035 ;
    RECT 31.37 35.325 31.58 35.395 ;
    RECT 31.83 34.605 32.04 34.675 ;
    RECT 31.83 34.965 32.04 35.035 ;
    RECT 31.83 35.325 32.04 35.395 ;
    RECT 67.89 34.605 68.1 34.675 ;
    RECT 67.89 34.965 68.1 35.035 ;
    RECT 67.89 35.325 68.1 35.395 ;
    RECT 68.35 34.605 68.56 34.675 ;
    RECT 68.35 34.965 68.56 35.035 ;
    RECT 68.35 35.325 68.56 35.395 ;
    RECT 28.05 34.605 28.26 34.675 ;
    RECT 28.05 34.965 28.26 35.035 ;
    RECT 28.05 35.325 28.26 35.395 ;
    RECT 28.51 34.605 28.72 34.675 ;
    RECT 28.51 34.965 28.72 35.035 ;
    RECT 28.51 35.325 28.72 35.395 ;
    RECT 24.73 34.605 24.94 34.675 ;
    RECT 24.73 34.965 24.94 35.035 ;
    RECT 24.73 35.325 24.94 35.395 ;
    RECT 25.19 34.605 25.4 34.675 ;
    RECT 25.19 34.965 25.4 35.035 ;
    RECT 25.19 35.325 25.4 35.395 ;
    RECT 21.41 34.605 21.62 34.675 ;
    RECT 21.41 34.965 21.62 35.035 ;
    RECT 21.41 35.325 21.62 35.395 ;
    RECT 21.87 34.605 22.08 34.675 ;
    RECT 21.87 34.965 22.08 35.035 ;
    RECT 21.87 35.325 22.08 35.395 ;
    RECT 18.09 34.605 18.3 34.675 ;
    RECT 18.09 34.965 18.3 35.035 ;
    RECT 18.09 35.325 18.3 35.395 ;
    RECT 18.55 34.605 18.76 34.675 ;
    RECT 18.55 34.965 18.76 35.035 ;
    RECT 18.55 35.325 18.76 35.395 ;
    RECT 14.77 34.605 14.98 34.675 ;
    RECT 14.77 34.965 14.98 35.035 ;
    RECT 14.77 35.325 14.98 35.395 ;
    RECT 15.23 34.605 15.44 34.675 ;
    RECT 15.23 34.965 15.44 35.035 ;
    RECT 15.23 35.325 15.44 35.395 ;
    RECT 11.45 34.605 11.66 34.675 ;
    RECT 11.45 34.965 11.66 35.035 ;
    RECT 11.45 35.325 11.66 35.395 ;
    RECT 11.91 34.605 12.12 34.675 ;
    RECT 11.91 34.965 12.12 35.035 ;
    RECT 11.91 35.325 12.12 35.395 ;
    RECT 8.13 34.605 8.34 34.675 ;
    RECT 8.13 34.965 8.34 35.035 ;
    RECT 8.13 35.325 8.34 35.395 ;
    RECT 8.59 34.605 8.8 34.675 ;
    RECT 8.59 34.965 8.8 35.035 ;
    RECT 8.59 35.325 8.8 35.395 ;
    RECT 4.81 34.605 5.02 34.675 ;
    RECT 4.81 34.965 5.02 35.035 ;
    RECT 4.81 35.325 5.02 35.395 ;
    RECT 5.27 34.605 5.48 34.675 ;
    RECT 5.27 34.965 5.48 35.035 ;
    RECT 5.27 35.325 5.48 35.395 ;
    RECT 164.17 34.605 164.38 34.675 ;
    RECT 164.17 34.965 164.38 35.035 ;
    RECT 164.17 35.325 164.38 35.395 ;
    RECT 164.63 34.605 164.84 34.675 ;
    RECT 164.63 34.965 164.84 35.035 ;
    RECT 164.63 35.325 164.84 35.395 ;
    RECT 1.49 34.605 1.7 34.675 ;
    RECT 1.49 34.965 1.7 35.035 ;
    RECT 1.49 35.325 1.7 35.395 ;
    RECT 1.95 34.605 2.16 34.675 ;
    RECT 1.95 34.965 2.16 35.035 ;
    RECT 1.95 35.325 2.16 35.395 ;
    RECT 160.85 34.605 161.06 34.675 ;
    RECT 160.85 34.965 161.06 35.035 ;
    RECT 160.85 35.325 161.06 35.395 ;
    RECT 161.31 34.605 161.52 34.675 ;
    RECT 161.31 34.965 161.52 35.035 ;
    RECT 161.31 35.325 161.52 35.395 ;
    RECT 157.53 34.605 157.74 34.675 ;
    RECT 157.53 34.965 157.74 35.035 ;
    RECT 157.53 35.325 157.74 35.395 ;
    RECT 157.99 34.605 158.2 34.675 ;
    RECT 157.99 34.965 158.2 35.035 ;
    RECT 157.99 35.325 158.2 35.395 ;
    RECT 154.21 34.605 154.42 34.675 ;
    RECT 154.21 34.965 154.42 35.035 ;
    RECT 154.21 35.325 154.42 35.395 ;
    RECT 154.67 34.605 154.88 34.675 ;
    RECT 154.67 34.965 154.88 35.035 ;
    RECT 154.67 35.325 154.88 35.395 ;
    RECT 150.89 34.605 151.1 34.675 ;
    RECT 150.89 34.965 151.1 35.035 ;
    RECT 150.89 35.325 151.1 35.395 ;
    RECT 151.35 34.605 151.56 34.675 ;
    RECT 151.35 34.965 151.56 35.035 ;
    RECT 151.35 35.325 151.56 35.395 ;
    RECT 147.57 34.605 147.78 34.675 ;
    RECT 147.57 34.965 147.78 35.035 ;
    RECT 147.57 35.325 147.78 35.395 ;
    RECT 148.03 34.605 148.24 34.675 ;
    RECT 148.03 34.965 148.24 35.035 ;
    RECT 148.03 35.325 148.24 35.395 ;
    RECT 144.25 34.605 144.46 34.675 ;
    RECT 144.25 34.965 144.46 35.035 ;
    RECT 144.25 35.325 144.46 35.395 ;
    RECT 144.71 34.605 144.92 34.675 ;
    RECT 144.71 34.965 144.92 35.035 ;
    RECT 144.71 35.325 144.92 35.395 ;
    RECT 140.93 34.605 141.14 34.675 ;
    RECT 140.93 34.965 141.14 35.035 ;
    RECT 140.93 35.325 141.14 35.395 ;
    RECT 141.39 34.605 141.6 34.675 ;
    RECT 141.39 34.965 141.6 35.035 ;
    RECT 141.39 35.325 141.6 35.395 ;
    RECT 137.61 34.605 137.82 34.675 ;
    RECT 137.61 34.965 137.82 35.035 ;
    RECT 137.61 35.325 137.82 35.395 ;
    RECT 138.07 34.605 138.28 34.675 ;
    RECT 138.07 34.965 138.28 35.035 ;
    RECT 138.07 35.325 138.28 35.395 ;
    RECT 134.29 34.605 134.5 34.675 ;
    RECT 134.29 34.965 134.5 35.035 ;
    RECT 134.29 35.325 134.5 35.395 ;
    RECT 134.75 34.605 134.96 34.675 ;
    RECT 134.75 34.965 134.96 35.035 ;
    RECT 134.75 35.325 134.96 35.395 ;
    RECT 64.57 34.605 64.78 34.675 ;
    RECT 64.57 34.965 64.78 35.035 ;
    RECT 64.57 35.325 64.78 35.395 ;
    RECT 65.03 34.605 65.24 34.675 ;
    RECT 65.03 34.965 65.24 35.035 ;
    RECT 65.03 35.325 65.24 35.395 ;
    RECT 61.25 54.045 61.46 54.115 ;
    RECT 61.25 54.405 61.46 54.475 ;
    RECT 61.25 54.765 61.46 54.835 ;
    RECT 61.71 54.045 61.92 54.115 ;
    RECT 61.71 54.405 61.92 54.475 ;
    RECT 61.71 54.765 61.92 54.835 ;
    RECT 57.93 54.045 58.14 54.115 ;
    RECT 57.93 54.405 58.14 54.475 ;
    RECT 57.93 54.765 58.14 54.835 ;
    RECT 58.39 54.045 58.6 54.115 ;
    RECT 58.39 54.405 58.6 54.475 ;
    RECT 58.39 54.765 58.6 54.835 ;
    RECT 54.61 54.045 54.82 54.115 ;
    RECT 54.61 54.405 54.82 54.475 ;
    RECT 54.61 54.765 54.82 54.835 ;
    RECT 55.07 54.045 55.28 54.115 ;
    RECT 55.07 54.405 55.28 54.475 ;
    RECT 55.07 54.765 55.28 54.835 ;
    RECT 51.29 54.045 51.5 54.115 ;
    RECT 51.29 54.405 51.5 54.475 ;
    RECT 51.29 54.765 51.5 54.835 ;
    RECT 51.75 54.045 51.96 54.115 ;
    RECT 51.75 54.405 51.96 54.475 ;
    RECT 51.75 54.765 51.96 54.835 ;
    RECT 47.97 54.045 48.18 54.115 ;
    RECT 47.97 54.405 48.18 54.475 ;
    RECT 47.97 54.765 48.18 54.835 ;
    RECT 48.43 54.045 48.64 54.115 ;
    RECT 48.43 54.405 48.64 54.475 ;
    RECT 48.43 54.765 48.64 54.835 ;
    RECT 44.65 54.045 44.86 54.115 ;
    RECT 44.65 54.405 44.86 54.475 ;
    RECT 44.65 54.765 44.86 54.835 ;
    RECT 45.11 54.045 45.32 54.115 ;
    RECT 45.11 54.405 45.32 54.475 ;
    RECT 45.11 54.765 45.32 54.835 ;
    RECT 41.33 54.045 41.54 54.115 ;
    RECT 41.33 54.405 41.54 54.475 ;
    RECT 41.33 54.765 41.54 54.835 ;
    RECT 41.79 54.045 42.0 54.115 ;
    RECT 41.79 54.405 42.0 54.475 ;
    RECT 41.79 54.765 42.0 54.835 ;
    RECT 38.01 54.045 38.22 54.115 ;
    RECT 38.01 54.405 38.22 54.475 ;
    RECT 38.01 54.765 38.22 54.835 ;
    RECT 38.47 54.045 38.68 54.115 ;
    RECT 38.47 54.405 38.68 54.475 ;
    RECT 38.47 54.765 38.68 54.835 ;
    RECT 34.69 54.045 34.9 54.115 ;
    RECT 34.69 54.405 34.9 54.475 ;
    RECT 34.69 54.765 34.9 54.835 ;
    RECT 35.15 54.045 35.36 54.115 ;
    RECT 35.15 54.405 35.36 54.475 ;
    RECT 35.15 54.765 35.36 54.835 ;
    RECT 173.945 54.405 174.015 54.475 ;
    RECT 130.97 54.045 131.18 54.115 ;
    RECT 130.97 54.405 131.18 54.475 ;
    RECT 130.97 54.765 131.18 54.835 ;
    RECT 131.43 54.045 131.64 54.115 ;
    RECT 131.43 54.405 131.64 54.475 ;
    RECT 131.43 54.765 131.64 54.835 ;
    RECT 127.65 54.045 127.86 54.115 ;
    RECT 127.65 54.405 127.86 54.475 ;
    RECT 127.65 54.765 127.86 54.835 ;
    RECT 128.11 54.045 128.32 54.115 ;
    RECT 128.11 54.405 128.32 54.475 ;
    RECT 128.11 54.765 128.32 54.835 ;
    RECT 124.33 54.045 124.54 54.115 ;
    RECT 124.33 54.405 124.54 54.475 ;
    RECT 124.33 54.765 124.54 54.835 ;
    RECT 124.79 54.045 125.0 54.115 ;
    RECT 124.79 54.405 125.0 54.475 ;
    RECT 124.79 54.765 125.0 54.835 ;
    RECT 121.01 54.045 121.22 54.115 ;
    RECT 121.01 54.405 121.22 54.475 ;
    RECT 121.01 54.765 121.22 54.835 ;
    RECT 121.47 54.045 121.68 54.115 ;
    RECT 121.47 54.405 121.68 54.475 ;
    RECT 121.47 54.765 121.68 54.835 ;
    RECT 117.69 54.045 117.9 54.115 ;
    RECT 117.69 54.405 117.9 54.475 ;
    RECT 117.69 54.765 117.9 54.835 ;
    RECT 118.15 54.045 118.36 54.115 ;
    RECT 118.15 54.405 118.36 54.475 ;
    RECT 118.15 54.765 118.36 54.835 ;
    RECT 114.37 54.045 114.58 54.115 ;
    RECT 114.37 54.405 114.58 54.475 ;
    RECT 114.37 54.765 114.58 54.835 ;
    RECT 114.83 54.045 115.04 54.115 ;
    RECT 114.83 54.405 115.04 54.475 ;
    RECT 114.83 54.765 115.04 54.835 ;
    RECT 111.05 54.045 111.26 54.115 ;
    RECT 111.05 54.405 111.26 54.475 ;
    RECT 111.05 54.765 111.26 54.835 ;
    RECT 111.51 54.045 111.72 54.115 ;
    RECT 111.51 54.405 111.72 54.475 ;
    RECT 111.51 54.765 111.72 54.835 ;
    RECT 107.73 54.045 107.94 54.115 ;
    RECT 107.73 54.405 107.94 54.475 ;
    RECT 107.73 54.765 107.94 54.835 ;
    RECT 108.19 54.045 108.4 54.115 ;
    RECT 108.19 54.405 108.4 54.475 ;
    RECT 108.19 54.765 108.4 54.835 ;
    RECT 104.41 54.045 104.62 54.115 ;
    RECT 104.41 54.405 104.62 54.475 ;
    RECT 104.41 54.765 104.62 54.835 ;
    RECT 104.87 54.045 105.08 54.115 ;
    RECT 104.87 54.405 105.08 54.475 ;
    RECT 104.87 54.765 105.08 54.835 ;
    RECT 101.09 54.045 101.3 54.115 ;
    RECT 101.09 54.405 101.3 54.475 ;
    RECT 101.09 54.765 101.3 54.835 ;
    RECT 101.55 54.045 101.76 54.115 ;
    RECT 101.55 54.405 101.76 54.475 ;
    RECT 101.55 54.765 101.76 54.835 ;
    RECT 0.4 54.405 0.47 54.475 ;
    RECT 170.81 54.045 171.02 54.115 ;
    RECT 170.81 54.405 171.02 54.475 ;
    RECT 170.81 54.765 171.02 54.835 ;
    RECT 171.27 54.045 171.48 54.115 ;
    RECT 171.27 54.405 171.48 54.475 ;
    RECT 171.27 54.765 171.48 54.835 ;
    RECT 167.49 54.045 167.7 54.115 ;
    RECT 167.49 54.405 167.7 54.475 ;
    RECT 167.49 54.765 167.7 54.835 ;
    RECT 167.95 54.045 168.16 54.115 ;
    RECT 167.95 54.405 168.16 54.475 ;
    RECT 167.95 54.765 168.16 54.835 ;
    RECT 97.77 54.045 97.98 54.115 ;
    RECT 97.77 54.405 97.98 54.475 ;
    RECT 97.77 54.765 97.98 54.835 ;
    RECT 98.23 54.045 98.44 54.115 ;
    RECT 98.23 54.405 98.44 54.475 ;
    RECT 98.23 54.765 98.44 54.835 ;
    RECT 94.45 54.045 94.66 54.115 ;
    RECT 94.45 54.405 94.66 54.475 ;
    RECT 94.45 54.765 94.66 54.835 ;
    RECT 94.91 54.045 95.12 54.115 ;
    RECT 94.91 54.405 95.12 54.475 ;
    RECT 94.91 54.765 95.12 54.835 ;
    RECT 91.13 54.045 91.34 54.115 ;
    RECT 91.13 54.405 91.34 54.475 ;
    RECT 91.13 54.765 91.34 54.835 ;
    RECT 91.59 54.045 91.8 54.115 ;
    RECT 91.59 54.405 91.8 54.475 ;
    RECT 91.59 54.765 91.8 54.835 ;
    RECT 87.81 54.045 88.02 54.115 ;
    RECT 87.81 54.405 88.02 54.475 ;
    RECT 87.81 54.765 88.02 54.835 ;
    RECT 88.27 54.045 88.48 54.115 ;
    RECT 88.27 54.405 88.48 54.475 ;
    RECT 88.27 54.765 88.48 54.835 ;
    RECT 84.49 54.045 84.7 54.115 ;
    RECT 84.49 54.405 84.7 54.475 ;
    RECT 84.49 54.765 84.7 54.835 ;
    RECT 84.95 54.045 85.16 54.115 ;
    RECT 84.95 54.405 85.16 54.475 ;
    RECT 84.95 54.765 85.16 54.835 ;
    RECT 81.17 54.045 81.38 54.115 ;
    RECT 81.17 54.405 81.38 54.475 ;
    RECT 81.17 54.765 81.38 54.835 ;
    RECT 81.63 54.045 81.84 54.115 ;
    RECT 81.63 54.405 81.84 54.475 ;
    RECT 81.63 54.765 81.84 54.835 ;
    RECT 77.85 54.045 78.06 54.115 ;
    RECT 77.85 54.405 78.06 54.475 ;
    RECT 77.85 54.765 78.06 54.835 ;
    RECT 78.31 54.045 78.52 54.115 ;
    RECT 78.31 54.405 78.52 54.475 ;
    RECT 78.31 54.765 78.52 54.835 ;
    RECT 74.53 54.045 74.74 54.115 ;
    RECT 74.53 54.405 74.74 54.475 ;
    RECT 74.53 54.765 74.74 54.835 ;
    RECT 74.99 54.045 75.2 54.115 ;
    RECT 74.99 54.405 75.2 54.475 ;
    RECT 74.99 54.765 75.2 54.835 ;
    RECT 71.21 54.045 71.42 54.115 ;
    RECT 71.21 54.405 71.42 54.475 ;
    RECT 71.21 54.765 71.42 54.835 ;
    RECT 71.67 54.045 71.88 54.115 ;
    RECT 71.67 54.405 71.88 54.475 ;
    RECT 71.67 54.765 71.88 54.835 ;
    RECT 31.37 54.045 31.58 54.115 ;
    RECT 31.37 54.405 31.58 54.475 ;
    RECT 31.37 54.765 31.58 54.835 ;
    RECT 31.83 54.045 32.04 54.115 ;
    RECT 31.83 54.405 32.04 54.475 ;
    RECT 31.83 54.765 32.04 54.835 ;
    RECT 67.89 54.045 68.1 54.115 ;
    RECT 67.89 54.405 68.1 54.475 ;
    RECT 67.89 54.765 68.1 54.835 ;
    RECT 68.35 54.045 68.56 54.115 ;
    RECT 68.35 54.405 68.56 54.475 ;
    RECT 68.35 54.765 68.56 54.835 ;
    RECT 28.05 54.045 28.26 54.115 ;
    RECT 28.05 54.405 28.26 54.475 ;
    RECT 28.05 54.765 28.26 54.835 ;
    RECT 28.51 54.045 28.72 54.115 ;
    RECT 28.51 54.405 28.72 54.475 ;
    RECT 28.51 54.765 28.72 54.835 ;
    RECT 24.73 54.045 24.94 54.115 ;
    RECT 24.73 54.405 24.94 54.475 ;
    RECT 24.73 54.765 24.94 54.835 ;
    RECT 25.19 54.045 25.4 54.115 ;
    RECT 25.19 54.405 25.4 54.475 ;
    RECT 25.19 54.765 25.4 54.835 ;
    RECT 21.41 54.045 21.62 54.115 ;
    RECT 21.41 54.405 21.62 54.475 ;
    RECT 21.41 54.765 21.62 54.835 ;
    RECT 21.87 54.045 22.08 54.115 ;
    RECT 21.87 54.405 22.08 54.475 ;
    RECT 21.87 54.765 22.08 54.835 ;
    RECT 18.09 54.045 18.3 54.115 ;
    RECT 18.09 54.405 18.3 54.475 ;
    RECT 18.09 54.765 18.3 54.835 ;
    RECT 18.55 54.045 18.76 54.115 ;
    RECT 18.55 54.405 18.76 54.475 ;
    RECT 18.55 54.765 18.76 54.835 ;
    RECT 14.77 54.045 14.98 54.115 ;
    RECT 14.77 54.405 14.98 54.475 ;
    RECT 14.77 54.765 14.98 54.835 ;
    RECT 15.23 54.045 15.44 54.115 ;
    RECT 15.23 54.405 15.44 54.475 ;
    RECT 15.23 54.765 15.44 54.835 ;
    RECT 11.45 54.045 11.66 54.115 ;
    RECT 11.45 54.405 11.66 54.475 ;
    RECT 11.45 54.765 11.66 54.835 ;
    RECT 11.91 54.045 12.12 54.115 ;
    RECT 11.91 54.405 12.12 54.475 ;
    RECT 11.91 54.765 12.12 54.835 ;
    RECT 8.13 54.045 8.34 54.115 ;
    RECT 8.13 54.405 8.34 54.475 ;
    RECT 8.13 54.765 8.34 54.835 ;
    RECT 8.59 54.045 8.8 54.115 ;
    RECT 8.59 54.405 8.8 54.475 ;
    RECT 8.59 54.765 8.8 54.835 ;
    RECT 4.81 54.045 5.02 54.115 ;
    RECT 4.81 54.405 5.02 54.475 ;
    RECT 4.81 54.765 5.02 54.835 ;
    RECT 5.27 54.045 5.48 54.115 ;
    RECT 5.27 54.405 5.48 54.475 ;
    RECT 5.27 54.765 5.48 54.835 ;
    RECT 164.17 54.045 164.38 54.115 ;
    RECT 164.17 54.405 164.38 54.475 ;
    RECT 164.17 54.765 164.38 54.835 ;
    RECT 164.63 54.045 164.84 54.115 ;
    RECT 164.63 54.405 164.84 54.475 ;
    RECT 164.63 54.765 164.84 54.835 ;
    RECT 1.49 54.045 1.7 54.115 ;
    RECT 1.49 54.405 1.7 54.475 ;
    RECT 1.49 54.765 1.7 54.835 ;
    RECT 1.95 54.045 2.16 54.115 ;
    RECT 1.95 54.405 2.16 54.475 ;
    RECT 1.95 54.765 2.16 54.835 ;
    RECT 160.85 54.045 161.06 54.115 ;
    RECT 160.85 54.405 161.06 54.475 ;
    RECT 160.85 54.765 161.06 54.835 ;
    RECT 161.31 54.045 161.52 54.115 ;
    RECT 161.31 54.405 161.52 54.475 ;
    RECT 161.31 54.765 161.52 54.835 ;
    RECT 157.53 54.045 157.74 54.115 ;
    RECT 157.53 54.405 157.74 54.475 ;
    RECT 157.53 54.765 157.74 54.835 ;
    RECT 157.99 54.045 158.2 54.115 ;
    RECT 157.99 54.405 158.2 54.475 ;
    RECT 157.99 54.765 158.2 54.835 ;
    RECT 154.21 54.045 154.42 54.115 ;
    RECT 154.21 54.405 154.42 54.475 ;
    RECT 154.21 54.765 154.42 54.835 ;
    RECT 154.67 54.045 154.88 54.115 ;
    RECT 154.67 54.405 154.88 54.475 ;
    RECT 154.67 54.765 154.88 54.835 ;
    RECT 150.89 54.045 151.1 54.115 ;
    RECT 150.89 54.405 151.1 54.475 ;
    RECT 150.89 54.765 151.1 54.835 ;
    RECT 151.35 54.045 151.56 54.115 ;
    RECT 151.35 54.405 151.56 54.475 ;
    RECT 151.35 54.765 151.56 54.835 ;
    RECT 147.57 54.045 147.78 54.115 ;
    RECT 147.57 54.405 147.78 54.475 ;
    RECT 147.57 54.765 147.78 54.835 ;
    RECT 148.03 54.045 148.24 54.115 ;
    RECT 148.03 54.405 148.24 54.475 ;
    RECT 148.03 54.765 148.24 54.835 ;
    RECT 144.25 54.045 144.46 54.115 ;
    RECT 144.25 54.405 144.46 54.475 ;
    RECT 144.25 54.765 144.46 54.835 ;
    RECT 144.71 54.045 144.92 54.115 ;
    RECT 144.71 54.405 144.92 54.475 ;
    RECT 144.71 54.765 144.92 54.835 ;
    RECT 140.93 54.045 141.14 54.115 ;
    RECT 140.93 54.405 141.14 54.475 ;
    RECT 140.93 54.765 141.14 54.835 ;
    RECT 141.39 54.045 141.6 54.115 ;
    RECT 141.39 54.405 141.6 54.475 ;
    RECT 141.39 54.765 141.6 54.835 ;
    RECT 137.61 54.045 137.82 54.115 ;
    RECT 137.61 54.405 137.82 54.475 ;
    RECT 137.61 54.765 137.82 54.835 ;
    RECT 138.07 54.045 138.28 54.115 ;
    RECT 138.07 54.405 138.28 54.475 ;
    RECT 138.07 54.765 138.28 54.835 ;
    RECT 134.29 54.045 134.5 54.115 ;
    RECT 134.29 54.405 134.5 54.475 ;
    RECT 134.29 54.765 134.5 54.835 ;
    RECT 134.75 54.045 134.96 54.115 ;
    RECT 134.75 54.405 134.96 54.475 ;
    RECT 134.75 54.765 134.96 54.835 ;
    RECT 64.57 54.045 64.78 54.115 ;
    RECT 64.57 54.405 64.78 54.475 ;
    RECT 64.57 54.765 64.78 54.835 ;
    RECT 65.03 54.045 65.24 54.115 ;
    RECT 65.03 54.405 65.24 54.475 ;
    RECT 65.03 54.765 65.24 54.835 ;
    RECT 61.25 53.325 61.46 53.395 ;
    RECT 61.25 53.685 61.46 53.755 ;
    RECT 61.25 54.045 61.46 54.115 ;
    RECT 61.71 53.325 61.92 53.395 ;
    RECT 61.71 53.685 61.92 53.755 ;
    RECT 61.71 54.045 61.92 54.115 ;
    RECT 57.93 53.325 58.14 53.395 ;
    RECT 57.93 53.685 58.14 53.755 ;
    RECT 57.93 54.045 58.14 54.115 ;
    RECT 58.39 53.325 58.6 53.395 ;
    RECT 58.39 53.685 58.6 53.755 ;
    RECT 58.39 54.045 58.6 54.115 ;
    RECT 54.61 53.325 54.82 53.395 ;
    RECT 54.61 53.685 54.82 53.755 ;
    RECT 54.61 54.045 54.82 54.115 ;
    RECT 55.07 53.325 55.28 53.395 ;
    RECT 55.07 53.685 55.28 53.755 ;
    RECT 55.07 54.045 55.28 54.115 ;
    RECT 51.29 53.325 51.5 53.395 ;
    RECT 51.29 53.685 51.5 53.755 ;
    RECT 51.29 54.045 51.5 54.115 ;
    RECT 51.75 53.325 51.96 53.395 ;
    RECT 51.75 53.685 51.96 53.755 ;
    RECT 51.75 54.045 51.96 54.115 ;
    RECT 47.97 53.325 48.18 53.395 ;
    RECT 47.97 53.685 48.18 53.755 ;
    RECT 47.97 54.045 48.18 54.115 ;
    RECT 48.43 53.325 48.64 53.395 ;
    RECT 48.43 53.685 48.64 53.755 ;
    RECT 48.43 54.045 48.64 54.115 ;
    RECT 44.65 53.325 44.86 53.395 ;
    RECT 44.65 53.685 44.86 53.755 ;
    RECT 44.65 54.045 44.86 54.115 ;
    RECT 45.11 53.325 45.32 53.395 ;
    RECT 45.11 53.685 45.32 53.755 ;
    RECT 45.11 54.045 45.32 54.115 ;
    RECT 41.33 53.325 41.54 53.395 ;
    RECT 41.33 53.685 41.54 53.755 ;
    RECT 41.33 54.045 41.54 54.115 ;
    RECT 41.79 53.325 42.0 53.395 ;
    RECT 41.79 53.685 42.0 53.755 ;
    RECT 41.79 54.045 42.0 54.115 ;
    RECT 38.01 53.325 38.22 53.395 ;
    RECT 38.01 53.685 38.22 53.755 ;
    RECT 38.01 54.045 38.22 54.115 ;
    RECT 38.47 53.325 38.68 53.395 ;
    RECT 38.47 53.685 38.68 53.755 ;
    RECT 38.47 54.045 38.68 54.115 ;
    RECT 34.69 53.325 34.9 53.395 ;
    RECT 34.69 53.685 34.9 53.755 ;
    RECT 34.69 54.045 34.9 54.115 ;
    RECT 35.15 53.325 35.36 53.395 ;
    RECT 35.15 53.685 35.36 53.755 ;
    RECT 35.15 54.045 35.36 54.115 ;
    RECT 173.945 53.685 174.015 53.755 ;
    RECT 130.97 53.325 131.18 53.395 ;
    RECT 130.97 53.685 131.18 53.755 ;
    RECT 130.97 54.045 131.18 54.115 ;
    RECT 131.43 53.325 131.64 53.395 ;
    RECT 131.43 53.685 131.64 53.755 ;
    RECT 131.43 54.045 131.64 54.115 ;
    RECT 127.65 53.325 127.86 53.395 ;
    RECT 127.65 53.685 127.86 53.755 ;
    RECT 127.65 54.045 127.86 54.115 ;
    RECT 128.11 53.325 128.32 53.395 ;
    RECT 128.11 53.685 128.32 53.755 ;
    RECT 128.11 54.045 128.32 54.115 ;
    RECT 124.33 53.325 124.54 53.395 ;
    RECT 124.33 53.685 124.54 53.755 ;
    RECT 124.33 54.045 124.54 54.115 ;
    RECT 124.79 53.325 125.0 53.395 ;
    RECT 124.79 53.685 125.0 53.755 ;
    RECT 124.79 54.045 125.0 54.115 ;
    RECT 121.01 53.325 121.22 53.395 ;
    RECT 121.01 53.685 121.22 53.755 ;
    RECT 121.01 54.045 121.22 54.115 ;
    RECT 121.47 53.325 121.68 53.395 ;
    RECT 121.47 53.685 121.68 53.755 ;
    RECT 121.47 54.045 121.68 54.115 ;
    RECT 117.69 53.325 117.9 53.395 ;
    RECT 117.69 53.685 117.9 53.755 ;
    RECT 117.69 54.045 117.9 54.115 ;
    RECT 118.15 53.325 118.36 53.395 ;
    RECT 118.15 53.685 118.36 53.755 ;
    RECT 118.15 54.045 118.36 54.115 ;
    RECT 114.37 53.325 114.58 53.395 ;
    RECT 114.37 53.685 114.58 53.755 ;
    RECT 114.37 54.045 114.58 54.115 ;
    RECT 114.83 53.325 115.04 53.395 ;
    RECT 114.83 53.685 115.04 53.755 ;
    RECT 114.83 54.045 115.04 54.115 ;
    RECT 111.05 53.325 111.26 53.395 ;
    RECT 111.05 53.685 111.26 53.755 ;
    RECT 111.05 54.045 111.26 54.115 ;
    RECT 111.51 53.325 111.72 53.395 ;
    RECT 111.51 53.685 111.72 53.755 ;
    RECT 111.51 54.045 111.72 54.115 ;
    RECT 107.73 53.325 107.94 53.395 ;
    RECT 107.73 53.685 107.94 53.755 ;
    RECT 107.73 54.045 107.94 54.115 ;
    RECT 108.19 53.325 108.4 53.395 ;
    RECT 108.19 53.685 108.4 53.755 ;
    RECT 108.19 54.045 108.4 54.115 ;
    RECT 104.41 53.325 104.62 53.395 ;
    RECT 104.41 53.685 104.62 53.755 ;
    RECT 104.41 54.045 104.62 54.115 ;
    RECT 104.87 53.325 105.08 53.395 ;
    RECT 104.87 53.685 105.08 53.755 ;
    RECT 104.87 54.045 105.08 54.115 ;
    RECT 101.09 53.325 101.3 53.395 ;
    RECT 101.09 53.685 101.3 53.755 ;
    RECT 101.09 54.045 101.3 54.115 ;
    RECT 101.55 53.325 101.76 53.395 ;
    RECT 101.55 53.685 101.76 53.755 ;
    RECT 101.55 54.045 101.76 54.115 ;
    RECT 0.4 53.685 0.47 53.755 ;
    RECT 170.81 53.325 171.02 53.395 ;
    RECT 170.81 53.685 171.02 53.755 ;
    RECT 170.81 54.045 171.02 54.115 ;
    RECT 171.27 53.325 171.48 53.395 ;
    RECT 171.27 53.685 171.48 53.755 ;
    RECT 171.27 54.045 171.48 54.115 ;
    RECT 167.49 53.325 167.7 53.395 ;
    RECT 167.49 53.685 167.7 53.755 ;
    RECT 167.49 54.045 167.7 54.115 ;
    RECT 167.95 53.325 168.16 53.395 ;
    RECT 167.95 53.685 168.16 53.755 ;
    RECT 167.95 54.045 168.16 54.115 ;
    RECT 97.77 53.325 97.98 53.395 ;
    RECT 97.77 53.685 97.98 53.755 ;
    RECT 97.77 54.045 97.98 54.115 ;
    RECT 98.23 53.325 98.44 53.395 ;
    RECT 98.23 53.685 98.44 53.755 ;
    RECT 98.23 54.045 98.44 54.115 ;
    RECT 94.45 53.325 94.66 53.395 ;
    RECT 94.45 53.685 94.66 53.755 ;
    RECT 94.45 54.045 94.66 54.115 ;
    RECT 94.91 53.325 95.12 53.395 ;
    RECT 94.91 53.685 95.12 53.755 ;
    RECT 94.91 54.045 95.12 54.115 ;
    RECT 91.13 53.325 91.34 53.395 ;
    RECT 91.13 53.685 91.34 53.755 ;
    RECT 91.13 54.045 91.34 54.115 ;
    RECT 91.59 53.325 91.8 53.395 ;
    RECT 91.59 53.685 91.8 53.755 ;
    RECT 91.59 54.045 91.8 54.115 ;
    RECT 87.81 53.325 88.02 53.395 ;
    RECT 87.81 53.685 88.02 53.755 ;
    RECT 87.81 54.045 88.02 54.115 ;
    RECT 88.27 53.325 88.48 53.395 ;
    RECT 88.27 53.685 88.48 53.755 ;
    RECT 88.27 54.045 88.48 54.115 ;
    RECT 84.49 53.325 84.7 53.395 ;
    RECT 84.49 53.685 84.7 53.755 ;
    RECT 84.49 54.045 84.7 54.115 ;
    RECT 84.95 53.325 85.16 53.395 ;
    RECT 84.95 53.685 85.16 53.755 ;
    RECT 84.95 54.045 85.16 54.115 ;
    RECT 81.17 53.325 81.38 53.395 ;
    RECT 81.17 53.685 81.38 53.755 ;
    RECT 81.17 54.045 81.38 54.115 ;
    RECT 81.63 53.325 81.84 53.395 ;
    RECT 81.63 53.685 81.84 53.755 ;
    RECT 81.63 54.045 81.84 54.115 ;
    RECT 77.85 53.325 78.06 53.395 ;
    RECT 77.85 53.685 78.06 53.755 ;
    RECT 77.85 54.045 78.06 54.115 ;
    RECT 78.31 53.325 78.52 53.395 ;
    RECT 78.31 53.685 78.52 53.755 ;
    RECT 78.31 54.045 78.52 54.115 ;
    RECT 74.53 53.325 74.74 53.395 ;
    RECT 74.53 53.685 74.74 53.755 ;
    RECT 74.53 54.045 74.74 54.115 ;
    RECT 74.99 53.325 75.2 53.395 ;
    RECT 74.99 53.685 75.2 53.755 ;
    RECT 74.99 54.045 75.2 54.115 ;
    RECT 71.21 53.325 71.42 53.395 ;
    RECT 71.21 53.685 71.42 53.755 ;
    RECT 71.21 54.045 71.42 54.115 ;
    RECT 71.67 53.325 71.88 53.395 ;
    RECT 71.67 53.685 71.88 53.755 ;
    RECT 71.67 54.045 71.88 54.115 ;
    RECT 31.37 53.325 31.58 53.395 ;
    RECT 31.37 53.685 31.58 53.755 ;
    RECT 31.37 54.045 31.58 54.115 ;
    RECT 31.83 53.325 32.04 53.395 ;
    RECT 31.83 53.685 32.04 53.755 ;
    RECT 31.83 54.045 32.04 54.115 ;
    RECT 67.89 53.325 68.1 53.395 ;
    RECT 67.89 53.685 68.1 53.755 ;
    RECT 67.89 54.045 68.1 54.115 ;
    RECT 68.35 53.325 68.56 53.395 ;
    RECT 68.35 53.685 68.56 53.755 ;
    RECT 68.35 54.045 68.56 54.115 ;
    RECT 28.05 53.325 28.26 53.395 ;
    RECT 28.05 53.685 28.26 53.755 ;
    RECT 28.05 54.045 28.26 54.115 ;
    RECT 28.51 53.325 28.72 53.395 ;
    RECT 28.51 53.685 28.72 53.755 ;
    RECT 28.51 54.045 28.72 54.115 ;
    RECT 24.73 53.325 24.94 53.395 ;
    RECT 24.73 53.685 24.94 53.755 ;
    RECT 24.73 54.045 24.94 54.115 ;
    RECT 25.19 53.325 25.4 53.395 ;
    RECT 25.19 53.685 25.4 53.755 ;
    RECT 25.19 54.045 25.4 54.115 ;
    RECT 21.41 53.325 21.62 53.395 ;
    RECT 21.41 53.685 21.62 53.755 ;
    RECT 21.41 54.045 21.62 54.115 ;
    RECT 21.87 53.325 22.08 53.395 ;
    RECT 21.87 53.685 22.08 53.755 ;
    RECT 21.87 54.045 22.08 54.115 ;
    RECT 18.09 53.325 18.3 53.395 ;
    RECT 18.09 53.685 18.3 53.755 ;
    RECT 18.09 54.045 18.3 54.115 ;
    RECT 18.55 53.325 18.76 53.395 ;
    RECT 18.55 53.685 18.76 53.755 ;
    RECT 18.55 54.045 18.76 54.115 ;
    RECT 14.77 53.325 14.98 53.395 ;
    RECT 14.77 53.685 14.98 53.755 ;
    RECT 14.77 54.045 14.98 54.115 ;
    RECT 15.23 53.325 15.44 53.395 ;
    RECT 15.23 53.685 15.44 53.755 ;
    RECT 15.23 54.045 15.44 54.115 ;
    RECT 11.45 53.325 11.66 53.395 ;
    RECT 11.45 53.685 11.66 53.755 ;
    RECT 11.45 54.045 11.66 54.115 ;
    RECT 11.91 53.325 12.12 53.395 ;
    RECT 11.91 53.685 12.12 53.755 ;
    RECT 11.91 54.045 12.12 54.115 ;
    RECT 8.13 53.325 8.34 53.395 ;
    RECT 8.13 53.685 8.34 53.755 ;
    RECT 8.13 54.045 8.34 54.115 ;
    RECT 8.59 53.325 8.8 53.395 ;
    RECT 8.59 53.685 8.8 53.755 ;
    RECT 8.59 54.045 8.8 54.115 ;
    RECT 4.81 53.325 5.02 53.395 ;
    RECT 4.81 53.685 5.02 53.755 ;
    RECT 4.81 54.045 5.02 54.115 ;
    RECT 5.27 53.325 5.48 53.395 ;
    RECT 5.27 53.685 5.48 53.755 ;
    RECT 5.27 54.045 5.48 54.115 ;
    RECT 164.17 53.325 164.38 53.395 ;
    RECT 164.17 53.685 164.38 53.755 ;
    RECT 164.17 54.045 164.38 54.115 ;
    RECT 164.63 53.325 164.84 53.395 ;
    RECT 164.63 53.685 164.84 53.755 ;
    RECT 164.63 54.045 164.84 54.115 ;
    RECT 1.49 53.325 1.7 53.395 ;
    RECT 1.49 53.685 1.7 53.755 ;
    RECT 1.49 54.045 1.7 54.115 ;
    RECT 1.95 53.325 2.16 53.395 ;
    RECT 1.95 53.685 2.16 53.755 ;
    RECT 1.95 54.045 2.16 54.115 ;
    RECT 160.85 53.325 161.06 53.395 ;
    RECT 160.85 53.685 161.06 53.755 ;
    RECT 160.85 54.045 161.06 54.115 ;
    RECT 161.31 53.325 161.52 53.395 ;
    RECT 161.31 53.685 161.52 53.755 ;
    RECT 161.31 54.045 161.52 54.115 ;
    RECT 157.53 53.325 157.74 53.395 ;
    RECT 157.53 53.685 157.74 53.755 ;
    RECT 157.53 54.045 157.74 54.115 ;
    RECT 157.99 53.325 158.2 53.395 ;
    RECT 157.99 53.685 158.2 53.755 ;
    RECT 157.99 54.045 158.2 54.115 ;
    RECT 154.21 53.325 154.42 53.395 ;
    RECT 154.21 53.685 154.42 53.755 ;
    RECT 154.21 54.045 154.42 54.115 ;
    RECT 154.67 53.325 154.88 53.395 ;
    RECT 154.67 53.685 154.88 53.755 ;
    RECT 154.67 54.045 154.88 54.115 ;
    RECT 150.89 53.325 151.1 53.395 ;
    RECT 150.89 53.685 151.1 53.755 ;
    RECT 150.89 54.045 151.1 54.115 ;
    RECT 151.35 53.325 151.56 53.395 ;
    RECT 151.35 53.685 151.56 53.755 ;
    RECT 151.35 54.045 151.56 54.115 ;
    RECT 147.57 53.325 147.78 53.395 ;
    RECT 147.57 53.685 147.78 53.755 ;
    RECT 147.57 54.045 147.78 54.115 ;
    RECT 148.03 53.325 148.24 53.395 ;
    RECT 148.03 53.685 148.24 53.755 ;
    RECT 148.03 54.045 148.24 54.115 ;
    RECT 144.25 53.325 144.46 53.395 ;
    RECT 144.25 53.685 144.46 53.755 ;
    RECT 144.25 54.045 144.46 54.115 ;
    RECT 144.71 53.325 144.92 53.395 ;
    RECT 144.71 53.685 144.92 53.755 ;
    RECT 144.71 54.045 144.92 54.115 ;
    RECT 140.93 53.325 141.14 53.395 ;
    RECT 140.93 53.685 141.14 53.755 ;
    RECT 140.93 54.045 141.14 54.115 ;
    RECT 141.39 53.325 141.6 53.395 ;
    RECT 141.39 53.685 141.6 53.755 ;
    RECT 141.39 54.045 141.6 54.115 ;
    RECT 137.61 53.325 137.82 53.395 ;
    RECT 137.61 53.685 137.82 53.755 ;
    RECT 137.61 54.045 137.82 54.115 ;
    RECT 138.07 53.325 138.28 53.395 ;
    RECT 138.07 53.685 138.28 53.755 ;
    RECT 138.07 54.045 138.28 54.115 ;
    RECT 134.29 53.325 134.5 53.395 ;
    RECT 134.29 53.685 134.5 53.755 ;
    RECT 134.29 54.045 134.5 54.115 ;
    RECT 134.75 53.325 134.96 53.395 ;
    RECT 134.75 53.685 134.96 53.755 ;
    RECT 134.75 54.045 134.96 54.115 ;
    RECT 64.57 53.325 64.78 53.395 ;
    RECT 64.57 53.685 64.78 53.755 ;
    RECT 64.57 54.045 64.78 54.115 ;
    RECT 65.03 53.325 65.24 53.395 ;
    RECT 65.03 53.685 65.24 53.755 ;
    RECT 65.03 54.045 65.24 54.115 ;
    RECT 61.25 52.605 61.46 52.675 ;
    RECT 61.25 52.965 61.46 53.035 ;
    RECT 61.25 53.325 61.46 53.395 ;
    RECT 61.71 52.605 61.92 52.675 ;
    RECT 61.71 52.965 61.92 53.035 ;
    RECT 61.71 53.325 61.92 53.395 ;
    RECT 57.93 52.605 58.14 52.675 ;
    RECT 57.93 52.965 58.14 53.035 ;
    RECT 57.93 53.325 58.14 53.395 ;
    RECT 58.39 52.605 58.6 52.675 ;
    RECT 58.39 52.965 58.6 53.035 ;
    RECT 58.39 53.325 58.6 53.395 ;
    RECT 54.61 52.605 54.82 52.675 ;
    RECT 54.61 52.965 54.82 53.035 ;
    RECT 54.61 53.325 54.82 53.395 ;
    RECT 55.07 52.605 55.28 52.675 ;
    RECT 55.07 52.965 55.28 53.035 ;
    RECT 55.07 53.325 55.28 53.395 ;
    RECT 51.29 52.605 51.5 52.675 ;
    RECT 51.29 52.965 51.5 53.035 ;
    RECT 51.29 53.325 51.5 53.395 ;
    RECT 51.75 52.605 51.96 52.675 ;
    RECT 51.75 52.965 51.96 53.035 ;
    RECT 51.75 53.325 51.96 53.395 ;
    RECT 47.97 52.605 48.18 52.675 ;
    RECT 47.97 52.965 48.18 53.035 ;
    RECT 47.97 53.325 48.18 53.395 ;
    RECT 48.43 52.605 48.64 52.675 ;
    RECT 48.43 52.965 48.64 53.035 ;
    RECT 48.43 53.325 48.64 53.395 ;
    RECT 44.65 52.605 44.86 52.675 ;
    RECT 44.65 52.965 44.86 53.035 ;
    RECT 44.65 53.325 44.86 53.395 ;
    RECT 45.11 52.605 45.32 52.675 ;
    RECT 45.11 52.965 45.32 53.035 ;
    RECT 45.11 53.325 45.32 53.395 ;
    RECT 41.33 52.605 41.54 52.675 ;
    RECT 41.33 52.965 41.54 53.035 ;
    RECT 41.33 53.325 41.54 53.395 ;
    RECT 41.79 52.605 42.0 52.675 ;
    RECT 41.79 52.965 42.0 53.035 ;
    RECT 41.79 53.325 42.0 53.395 ;
    RECT 38.01 52.605 38.22 52.675 ;
    RECT 38.01 52.965 38.22 53.035 ;
    RECT 38.01 53.325 38.22 53.395 ;
    RECT 38.47 52.605 38.68 52.675 ;
    RECT 38.47 52.965 38.68 53.035 ;
    RECT 38.47 53.325 38.68 53.395 ;
    RECT 34.69 52.605 34.9 52.675 ;
    RECT 34.69 52.965 34.9 53.035 ;
    RECT 34.69 53.325 34.9 53.395 ;
    RECT 35.15 52.605 35.36 52.675 ;
    RECT 35.15 52.965 35.36 53.035 ;
    RECT 35.15 53.325 35.36 53.395 ;
    RECT 173.945 52.965 174.015 53.035 ;
    RECT 130.97 52.605 131.18 52.675 ;
    RECT 130.97 52.965 131.18 53.035 ;
    RECT 130.97 53.325 131.18 53.395 ;
    RECT 131.43 52.605 131.64 52.675 ;
    RECT 131.43 52.965 131.64 53.035 ;
    RECT 131.43 53.325 131.64 53.395 ;
    RECT 127.65 52.605 127.86 52.675 ;
    RECT 127.65 52.965 127.86 53.035 ;
    RECT 127.65 53.325 127.86 53.395 ;
    RECT 128.11 52.605 128.32 52.675 ;
    RECT 128.11 52.965 128.32 53.035 ;
    RECT 128.11 53.325 128.32 53.395 ;
    RECT 124.33 52.605 124.54 52.675 ;
    RECT 124.33 52.965 124.54 53.035 ;
    RECT 124.33 53.325 124.54 53.395 ;
    RECT 124.79 52.605 125.0 52.675 ;
    RECT 124.79 52.965 125.0 53.035 ;
    RECT 124.79 53.325 125.0 53.395 ;
    RECT 121.01 52.605 121.22 52.675 ;
    RECT 121.01 52.965 121.22 53.035 ;
    RECT 121.01 53.325 121.22 53.395 ;
    RECT 121.47 52.605 121.68 52.675 ;
    RECT 121.47 52.965 121.68 53.035 ;
    RECT 121.47 53.325 121.68 53.395 ;
    RECT 117.69 52.605 117.9 52.675 ;
    RECT 117.69 52.965 117.9 53.035 ;
    RECT 117.69 53.325 117.9 53.395 ;
    RECT 118.15 52.605 118.36 52.675 ;
    RECT 118.15 52.965 118.36 53.035 ;
    RECT 118.15 53.325 118.36 53.395 ;
    RECT 114.37 52.605 114.58 52.675 ;
    RECT 114.37 52.965 114.58 53.035 ;
    RECT 114.37 53.325 114.58 53.395 ;
    RECT 114.83 52.605 115.04 52.675 ;
    RECT 114.83 52.965 115.04 53.035 ;
    RECT 114.83 53.325 115.04 53.395 ;
    RECT 111.05 52.605 111.26 52.675 ;
    RECT 111.05 52.965 111.26 53.035 ;
    RECT 111.05 53.325 111.26 53.395 ;
    RECT 111.51 52.605 111.72 52.675 ;
    RECT 111.51 52.965 111.72 53.035 ;
    RECT 111.51 53.325 111.72 53.395 ;
    RECT 107.73 52.605 107.94 52.675 ;
    RECT 107.73 52.965 107.94 53.035 ;
    RECT 107.73 53.325 107.94 53.395 ;
    RECT 108.19 52.605 108.4 52.675 ;
    RECT 108.19 52.965 108.4 53.035 ;
    RECT 108.19 53.325 108.4 53.395 ;
    RECT 104.41 52.605 104.62 52.675 ;
    RECT 104.41 52.965 104.62 53.035 ;
    RECT 104.41 53.325 104.62 53.395 ;
    RECT 104.87 52.605 105.08 52.675 ;
    RECT 104.87 52.965 105.08 53.035 ;
    RECT 104.87 53.325 105.08 53.395 ;
    RECT 101.09 52.605 101.3 52.675 ;
    RECT 101.09 52.965 101.3 53.035 ;
    RECT 101.09 53.325 101.3 53.395 ;
    RECT 101.55 52.605 101.76 52.675 ;
    RECT 101.55 52.965 101.76 53.035 ;
    RECT 101.55 53.325 101.76 53.395 ;
    RECT 0.4 52.965 0.47 53.035 ;
    RECT 170.81 52.605 171.02 52.675 ;
    RECT 170.81 52.965 171.02 53.035 ;
    RECT 170.81 53.325 171.02 53.395 ;
    RECT 171.27 52.605 171.48 52.675 ;
    RECT 171.27 52.965 171.48 53.035 ;
    RECT 171.27 53.325 171.48 53.395 ;
    RECT 167.49 52.605 167.7 52.675 ;
    RECT 167.49 52.965 167.7 53.035 ;
    RECT 167.49 53.325 167.7 53.395 ;
    RECT 167.95 52.605 168.16 52.675 ;
    RECT 167.95 52.965 168.16 53.035 ;
    RECT 167.95 53.325 168.16 53.395 ;
    RECT 97.77 52.605 97.98 52.675 ;
    RECT 97.77 52.965 97.98 53.035 ;
    RECT 97.77 53.325 97.98 53.395 ;
    RECT 98.23 52.605 98.44 52.675 ;
    RECT 98.23 52.965 98.44 53.035 ;
    RECT 98.23 53.325 98.44 53.395 ;
    RECT 94.45 52.605 94.66 52.675 ;
    RECT 94.45 52.965 94.66 53.035 ;
    RECT 94.45 53.325 94.66 53.395 ;
    RECT 94.91 52.605 95.12 52.675 ;
    RECT 94.91 52.965 95.12 53.035 ;
    RECT 94.91 53.325 95.12 53.395 ;
    RECT 91.13 52.605 91.34 52.675 ;
    RECT 91.13 52.965 91.34 53.035 ;
    RECT 91.13 53.325 91.34 53.395 ;
    RECT 91.59 52.605 91.8 52.675 ;
    RECT 91.59 52.965 91.8 53.035 ;
    RECT 91.59 53.325 91.8 53.395 ;
    RECT 87.81 52.605 88.02 52.675 ;
    RECT 87.81 52.965 88.02 53.035 ;
    RECT 87.81 53.325 88.02 53.395 ;
    RECT 88.27 52.605 88.48 52.675 ;
    RECT 88.27 52.965 88.48 53.035 ;
    RECT 88.27 53.325 88.48 53.395 ;
    RECT 84.49 52.605 84.7 52.675 ;
    RECT 84.49 52.965 84.7 53.035 ;
    RECT 84.49 53.325 84.7 53.395 ;
    RECT 84.95 52.605 85.16 52.675 ;
    RECT 84.95 52.965 85.16 53.035 ;
    RECT 84.95 53.325 85.16 53.395 ;
    RECT 81.17 52.605 81.38 52.675 ;
    RECT 81.17 52.965 81.38 53.035 ;
    RECT 81.17 53.325 81.38 53.395 ;
    RECT 81.63 52.605 81.84 52.675 ;
    RECT 81.63 52.965 81.84 53.035 ;
    RECT 81.63 53.325 81.84 53.395 ;
    RECT 77.85 52.605 78.06 52.675 ;
    RECT 77.85 52.965 78.06 53.035 ;
    RECT 77.85 53.325 78.06 53.395 ;
    RECT 78.31 52.605 78.52 52.675 ;
    RECT 78.31 52.965 78.52 53.035 ;
    RECT 78.31 53.325 78.52 53.395 ;
    RECT 74.53 52.605 74.74 52.675 ;
    RECT 74.53 52.965 74.74 53.035 ;
    RECT 74.53 53.325 74.74 53.395 ;
    RECT 74.99 52.605 75.2 52.675 ;
    RECT 74.99 52.965 75.2 53.035 ;
    RECT 74.99 53.325 75.2 53.395 ;
    RECT 71.21 52.605 71.42 52.675 ;
    RECT 71.21 52.965 71.42 53.035 ;
    RECT 71.21 53.325 71.42 53.395 ;
    RECT 71.67 52.605 71.88 52.675 ;
    RECT 71.67 52.965 71.88 53.035 ;
    RECT 71.67 53.325 71.88 53.395 ;
    RECT 31.37 52.605 31.58 52.675 ;
    RECT 31.37 52.965 31.58 53.035 ;
    RECT 31.37 53.325 31.58 53.395 ;
    RECT 31.83 52.605 32.04 52.675 ;
    RECT 31.83 52.965 32.04 53.035 ;
    RECT 31.83 53.325 32.04 53.395 ;
    RECT 67.89 52.605 68.1 52.675 ;
    RECT 67.89 52.965 68.1 53.035 ;
    RECT 67.89 53.325 68.1 53.395 ;
    RECT 68.35 52.605 68.56 52.675 ;
    RECT 68.35 52.965 68.56 53.035 ;
    RECT 68.35 53.325 68.56 53.395 ;
    RECT 28.05 52.605 28.26 52.675 ;
    RECT 28.05 52.965 28.26 53.035 ;
    RECT 28.05 53.325 28.26 53.395 ;
    RECT 28.51 52.605 28.72 52.675 ;
    RECT 28.51 52.965 28.72 53.035 ;
    RECT 28.51 53.325 28.72 53.395 ;
    RECT 24.73 52.605 24.94 52.675 ;
    RECT 24.73 52.965 24.94 53.035 ;
    RECT 24.73 53.325 24.94 53.395 ;
    RECT 25.19 52.605 25.4 52.675 ;
    RECT 25.19 52.965 25.4 53.035 ;
    RECT 25.19 53.325 25.4 53.395 ;
    RECT 21.41 52.605 21.62 52.675 ;
    RECT 21.41 52.965 21.62 53.035 ;
    RECT 21.41 53.325 21.62 53.395 ;
    RECT 21.87 52.605 22.08 52.675 ;
    RECT 21.87 52.965 22.08 53.035 ;
    RECT 21.87 53.325 22.08 53.395 ;
    RECT 18.09 52.605 18.3 52.675 ;
    RECT 18.09 52.965 18.3 53.035 ;
    RECT 18.09 53.325 18.3 53.395 ;
    RECT 18.55 52.605 18.76 52.675 ;
    RECT 18.55 52.965 18.76 53.035 ;
    RECT 18.55 53.325 18.76 53.395 ;
    RECT 14.77 52.605 14.98 52.675 ;
    RECT 14.77 52.965 14.98 53.035 ;
    RECT 14.77 53.325 14.98 53.395 ;
    RECT 15.23 52.605 15.44 52.675 ;
    RECT 15.23 52.965 15.44 53.035 ;
    RECT 15.23 53.325 15.44 53.395 ;
    RECT 11.45 52.605 11.66 52.675 ;
    RECT 11.45 52.965 11.66 53.035 ;
    RECT 11.45 53.325 11.66 53.395 ;
    RECT 11.91 52.605 12.12 52.675 ;
    RECT 11.91 52.965 12.12 53.035 ;
    RECT 11.91 53.325 12.12 53.395 ;
    RECT 8.13 52.605 8.34 52.675 ;
    RECT 8.13 52.965 8.34 53.035 ;
    RECT 8.13 53.325 8.34 53.395 ;
    RECT 8.59 52.605 8.8 52.675 ;
    RECT 8.59 52.965 8.8 53.035 ;
    RECT 8.59 53.325 8.8 53.395 ;
    RECT 4.81 52.605 5.02 52.675 ;
    RECT 4.81 52.965 5.02 53.035 ;
    RECT 4.81 53.325 5.02 53.395 ;
    RECT 5.27 52.605 5.48 52.675 ;
    RECT 5.27 52.965 5.48 53.035 ;
    RECT 5.27 53.325 5.48 53.395 ;
    RECT 164.17 52.605 164.38 52.675 ;
    RECT 164.17 52.965 164.38 53.035 ;
    RECT 164.17 53.325 164.38 53.395 ;
    RECT 164.63 52.605 164.84 52.675 ;
    RECT 164.63 52.965 164.84 53.035 ;
    RECT 164.63 53.325 164.84 53.395 ;
    RECT 1.49 52.605 1.7 52.675 ;
    RECT 1.49 52.965 1.7 53.035 ;
    RECT 1.49 53.325 1.7 53.395 ;
    RECT 1.95 52.605 2.16 52.675 ;
    RECT 1.95 52.965 2.16 53.035 ;
    RECT 1.95 53.325 2.16 53.395 ;
    RECT 160.85 52.605 161.06 52.675 ;
    RECT 160.85 52.965 161.06 53.035 ;
    RECT 160.85 53.325 161.06 53.395 ;
    RECT 161.31 52.605 161.52 52.675 ;
    RECT 161.31 52.965 161.52 53.035 ;
    RECT 161.31 53.325 161.52 53.395 ;
    RECT 157.53 52.605 157.74 52.675 ;
    RECT 157.53 52.965 157.74 53.035 ;
    RECT 157.53 53.325 157.74 53.395 ;
    RECT 157.99 52.605 158.2 52.675 ;
    RECT 157.99 52.965 158.2 53.035 ;
    RECT 157.99 53.325 158.2 53.395 ;
    RECT 154.21 52.605 154.42 52.675 ;
    RECT 154.21 52.965 154.42 53.035 ;
    RECT 154.21 53.325 154.42 53.395 ;
    RECT 154.67 52.605 154.88 52.675 ;
    RECT 154.67 52.965 154.88 53.035 ;
    RECT 154.67 53.325 154.88 53.395 ;
    RECT 150.89 52.605 151.1 52.675 ;
    RECT 150.89 52.965 151.1 53.035 ;
    RECT 150.89 53.325 151.1 53.395 ;
    RECT 151.35 52.605 151.56 52.675 ;
    RECT 151.35 52.965 151.56 53.035 ;
    RECT 151.35 53.325 151.56 53.395 ;
    RECT 147.57 52.605 147.78 52.675 ;
    RECT 147.57 52.965 147.78 53.035 ;
    RECT 147.57 53.325 147.78 53.395 ;
    RECT 148.03 52.605 148.24 52.675 ;
    RECT 148.03 52.965 148.24 53.035 ;
    RECT 148.03 53.325 148.24 53.395 ;
    RECT 144.25 52.605 144.46 52.675 ;
    RECT 144.25 52.965 144.46 53.035 ;
    RECT 144.25 53.325 144.46 53.395 ;
    RECT 144.71 52.605 144.92 52.675 ;
    RECT 144.71 52.965 144.92 53.035 ;
    RECT 144.71 53.325 144.92 53.395 ;
    RECT 140.93 52.605 141.14 52.675 ;
    RECT 140.93 52.965 141.14 53.035 ;
    RECT 140.93 53.325 141.14 53.395 ;
    RECT 141.39 52.605 141.6 52.675 ;
    RECT 141.39 52.965 141.6 53.035 ;
    RECT 141.39 53.325 141.6 53.395 ;
    RECT 137.61 52.605 137.82 52.675 ;
    RECT 137.61 52.965 137.82 53.035 ;
    RECT 137.61 53.325 137.82 53.395 ;
    RECT 138.07 52.605 138.28 52.675 ;
    RECT 138.07 52.965 138.28 53.035 ;
    RECT 138.07 53.325 138.28 53.395 ;
    RECT 134.29 52.605 134.5 52.675 ;
    RECT 134.29 52.965 134.5 53.035 ;
    RECT 134.29 53.325 134.5 53.395 ;
    RECT 134.75 52.605 134.96 52.675 ;
    RECT 134.75 52.965 134.96 53.035 ;
    RECT 134.75 53.325 134.96 53.395 ;
    RECT 64.57 52.605 64.78 52.675 ;
    RECT 64.57 52.965 64.78 53.035 ;
    RECT 64.57 53.325 64.78 53.395 ;
    RECT 65.03 52.605 65.24 52.675 ;
    RECT 65.03 52.965 65.24 53.035 ;
    RECT 65.03 53.325 65.24 53.395 ;
    RECT 61.25 51.885 61.46 51.955 ;
    RECT 61.25 52.245 61.46 52.315 ;
    RECT 61.25 52.605 61.46 52.675 ;
    RECT 61.71 51.885 61.92 51.955 ;
    RECT 61.71 52.245 61.92 52.315 ;
    RECT 61.71 52.605 61.92 52.675 ;
    RECT 57.93 51.885 58.14 51.955 ;
    RECT 57.93 52.245 58.14 52.315 ;
    RECT 57.93 52.605 58.14 52.675 ;
    RECT 58.39 51.885 58.6 51.955 ;
    RECT 58.39 52.245 58.6 52.315 ;
    RECT 58.39 52.605 58.6 52.675 ;
    RECT 54.61 51.885 54.82 51.955 ;
    RECT 54.61 52.245 54.82 52.315 ;
    RECT 54.61 52.605 54.82 52.675 ;
    RECT 55.07 51.885 55.28 51.955 ;
    RECT 55.07 52.245 55.28 52.315 ;
    RECT 55.07 52.605 55.28 52.675 ;
    RECT 51.29 51.885 51.5 51.955 ;
    RECT 51.29 52.245 51.5 52.315 ;
    RECT 51.29 52.605 51.5 52.675 ;
    RECT 51.75 51.885 51.96 51.955 ;
    RECT 51.75 52.245 51.96 52.315 ;
    RECT 51.75 52.605 51.96 52.675 ;
    RECT 47.97 51.885 48.18 51.955 ;
    RECT 47.97 52.245 48.18 52.315 ;
    RECT 47.97 52.605 48.18 52.675 ;
    RECT 48.43 51.885 48.64 51.955 ;
    RECT 48.43 52.245 48.64 52.315 ;
    RECT 48.43 52.605 48.64 52.675 ;
    RECT 44.65 51.885 44.86 51.955 ;
    RECT 44.65 52.245 44.86 52.315 ;
    RECT 44.65 52.605 44.86 52.675 ;
    RECT 45.11 51.885 45.32 51.955 ;
    RECT 45.11 52.245 45.32 52.315 ;
    RECT 45.11 52.605 45.32 52.675 ;
    RECT 41.33 51.885 41.54 51.955 ;
    RECT 41.33 52.245 41.54 52.315 ;
    RECT 41.33 52.605 41.54 52.675 ;
    RECT 41.79 51.885 42.0 51.955 ;
    RECT 41.79 52.245 42.0 52.315 ;
    RECT 41.79 52.605 42.0 52.675 ;
    RECT 38.01 51.885 38.22 51.955 ;
    RECT 38.01 52.245 38.22 52.315 ;
    RECT 38.01 52.605 38.22 52.675 ;
    RECT 38.47 51.885 38.68 51.955 ;
    RECT 38.47 52.245 38.68 52.315 ;
    RECT 38.47 52.605 38.68 52.675 ;
    RECT 34.69 51.885 34.9 51.955 ;
    RECT 34.69 52.245 34.9 52.315 ;
    RECT 34.69 52.605 34.9 52.675 ;
    RECT 35.15 51.885 35.36 51.955 ;
    RECT 35.15 52.245 35.36 52.315 ;
    RECT 35.15 52.605 35.36 52.675 ;
    RECT 173.945 52.245 174.015 52.315 ;
    RECT 130.97 51.885 131.18 51.955 ;
    RECT 130.97 52.245 131.18 52.315 ;
    RECT 130.97 52.605 131.18 52.675 ;
    RECT 131.43 51.885 131.64 51.955 ;
    RECT 131.43 52.245 131.64 52.315 ;
    RECT 131.43 52.605 131.64 52.675 ;
    RECT 127.65 51.885 127.86 51.955 ;
    RECT 127.65 52.245 127.86 52.315 ;
    RECT 127.65 52.605 127.86 52.675 ;
    RECT 128.11 51.885 128.32 51.955 ;
    RECT 128.11 52.245 128.32 52.315 ;
    RECT 128.11 52.605 128.32 52.675 ;
    RECT 124.33 51.885 124.54 51.955 ;
    RECT 124.33 52.245 124.54 52.315 ;
    RECT 124.33 52.605 124.54 52.675 ;
    RECT 124.79 51.885 125.0 51.955 ;
    RECT 124.79 52.245 125.0 52.315 ;
    RECT 124.79 52.605 125.0 52.675 ;
    RECT 121.01 51.885 121.22 51.955 ;
    RECT 121.01 52.245 121.22 52.315 ;
    RECT 121.01 52.605 121.22 52.675 ;
    RECT 121.47 51.885 121.68 51.955 ;
    RECT 121.47 52.245 121.68 52.315 ;
    RECT 121.47 52.605 121.68 52.675 ;
    RECT 117.69 51.885 117.9 51.955 ;
    RECT 117.69 52.245 117.9 52.315 ;
    RECT 117.69 52.605 117.9 52.675 ;
    RECT 118.15 51.885 118.36 51.955 ;
    RECT 118.15 52.245 118.36 52.315 ;
    RECT 118.15 52.605 118.36 52.675 ;
    RECT 114.37 51.885 114.58 51.955 ;
    RECT 114.37 52.245 114.58 52.315 ;
    RECT 114.37 52.605 114.58 52.675 ;
    RECT 114.83 51.885 115.04 51.955 ;
    RECT 114.83 52.245 115.04 52.315 ;
    RECT 114.83 52.605 115.04 52.675 ;
    RECT 111.05 51.885 111.26 51.955 ;
    RECT 111.05 52.245 111.26 52.315 ;
    RECT 111.05 52.605 111.26 52.675 ;
    RECT 111.51 51.885 111.72 51.955 ;
    RECT 111.51 52.245 111.72 52.315 ;
    RECT 111.51 52.605 111.72 52.675 ;
    RECT 107.73 51.885 107.94 51.955 ;
    RECT 107.73 52.245 107.94 52.315 ;
    RECT 107.73 52.605 107.94 52.675 ;
    RECT 108.19 51.885 108.4 51.955 ;
    RECT 108.19 52.245 108.4 52.315 ;
    RECT 108.19 52.605 108.4 52.675 ;
    RECT 104.41 51.885 104.62 51.955 ;
    RECT 104.41 52.245 104.62 52.315 ;
    RECT 104.41 52.605 104.62 52.675 ;
    RECT 104.87 51.885 105.08 51.955 ;
    RECT 104.87 52.245 105.08 52.315 ;
    RECT 104.87 52.605 105.08 52.675 ;
    RECT 101.09 51.885 101.3 51.955 ;
    RECT 101.09 52.245 101.3 52.315 ;
    RECT 101.09 52.605 101.3 52.675 ;
    RECT 101.55 51.885 101.76 51.955 ;
    RECT 101.55 52.245 101.76 52.315 ;
    RECT 101.55 52.605 101.76 52.675 ;
    RECT 0.4 52.245 0.47 52.315 ;
    RECT 170.81 51.885 171.02 51.955 ;
    RECT 170.81 52.245 171.02 52.315 ;
    RECT 170.81 52.605 171.02 52.675 ;
    RECT 171.27 51.885 171.48 51.955 ;
    RECT 171.27 52.245 171.48 52.315 ;
    RECT 171.27 52.605 171.48 52.675 ;
    RECT 167.49 51.885 167.7 51.955 ;
    RECT 167.49 52.245 167.7 52.315 ;
    RECT 167.49 52.605 167.7 52.675 ;
    RECT 167.95 51.885 168.16 51.955 ;
    RECT 167.95 52.245 168.16 52.315 ;
    RECT 167.95 52.605 168.16 52.675 ;
    RECT 97.77 51.885 97.98 51.955 ;
    RECT 97.77 52.245 97.98 52.315 ;
    RECT 97.77 52.605 97.98 52.675 ;
    RECT 98.23 51.885 98.44 51.955 ;
    RECT 98.23 52.245 98.44 52.315 ;
    RECT 98.23 52.605 98.44 52.675 ;
    RECT 94.45 51.885 94.66 51.955 ;
    RECT 94.45 52.245 94.66 52.315 ;
    RECT 94.45 52.605 94.66 52.675 ;
    RECT 94.91 51.885 95.12 51.955 ;
    RECT 94.91 52.245 95.12 52.315 ;
    RECT 94.91 52.605 95.12 52.675 ;
    RECT 91.13 51.885 91.34 51.955 ;
    RECT 91.13 52.245 91.34 52.315 ;
    RECT 91.13 52.605 91.34 52.675 ;
    RECT 91.59 51.885 91.8 51.955 ;
    RECT 91.59 52.245 91.8 52.315 ;
    RECT 91.59 52.605 91.8 52.675 ;
    RECT 87.81 51.885 88.02 51.955 ;
    RECT 87.81 52.245 88.02 52.315 ;
    RECT 87.81 52.605 88.02 52.675 ;
    RECT 88.27 51.885 88.48 51.955 ;
    RECT 88.27 52.245 88.48 52.315 ;
    RECT 88.27 52.605 88.48 52.675 ;
    RECT 84.49 51.885 84.7 51.955 ;
    RECT 84.49 52.245 84.7 52.315 ;
    RECT 84.49 52.605 84.7 52.675 ;
    RECT 84.95 51.885 85.16 51.955 ;
    RECT 84.95 52.245 85.16 52.315 ;
    RECT 84.95 52.605 85.16 52.675 ;
    RECT 81.17 51.885 81.38 51.955 ;
    RECT 81.17 52.245 81.38 52.315 ;
    RECT 81.17 52.605 81.38 52.675 ;
    RECT 81.63 51.885 81.84 51.955 ;
    RECT 81.63 52.245 81.84 52.315 ;
    RECT 81.63 52.605 81.84 52.675 ;
    RECT 77.85 51.885 78.06 51.955 ;
    RECT 77.85 52.245 78.06 52.315 ;
    RECT 77.85 52.605 78.06 52.675 ;
    RECT 78.31 51.885 78.52 51.955 ;
    RECT 78.31 52.245 78.52 52.315 ;
    RECT 78.31 52.605 78.52 52.675 ;
    RECT 74.53 51.885 74.74 51.955 ;
    RECT 74.53 52.245 74.74 52.315 ;
    RECT 74.53 52.605 74.74 52.675 ;
    RECT 74.99 51.885 75.2 51.955 ;
    RECT 74.99 52.245 75.2 52.315 ;
    RECT 74.99 52.605 75.2 52.675 ;
    RECT 71.21 51.885 71.42 51.955 ;
    RECT 71.21 52.245 71.42 52.315 ;
    RECT 71.21 52.605 71.42 52.675 ;
    RECT 71.67 51.885 71.88 51.955 ;
    RECT 71.67 52.245 71.88 52.315 ;
    RECT 71.67 52.605 71.88 52.675 ;
    RECT 31.37 51.885 31.58 51.955 ;
    RECT 31.37 52.245 31.58 52.315 ;
    RECT 31.37 52.605 31.58 52.675 ;
    RECT 31.83 51.885 32.04 51.955 ;
    RECT 31.83 52.245 32.04 52.315 ;
    RECT 31.83 52.605 32.04 52.675 ;
    RECT 67.89 51.885 68.1 51.955 ;
    RECT 67.89 52.245 68.1 52.315 ;
    RECT 67.89 52.605 68.1 52.675 ;
    RECT 68.35 51.885 68.56 51.955 ;
    RECT 68.35 52.245 68.56 52.315 ;
    RECT 68.35 52.605 68.56 52.675 ;
    RECT 28.05 51.885 28.26 51.955 ;
    RECT 28.05 52.245 28.26 52.315 ;
    RECT 28.05 52.605 28.26 52.675 ;
    RECT 28.51 51.885 28.72 51.955 ;
    RECT 28.51 52.245 28.72 52.315 ;
    RECT 28.51 52.605 28.72 52.675 ;
    RECT 24.73 51.885 24.94 51.955 ;
    RECT 24.73 52.245 24.94 52.315 ;
    RECT 24.73 52.605 24.94 52.675 ;
    RECT 25.19 51.885 25.4 51.955 ;
    RECT 25.19 52.245 25.4 52.315 ;
    RECT 25.19 52.605 25.4 52.675 ;
    RECT 21.41 51.885 21.62 51.955 ;
    RECT 21.41 52.245 21.62 52.315 ;
    RECT 21.41 52.605 21.62 52.675 ;
    RECT 21.87 51.885 22.08 51.955 ;
    RECT 21.87 52.245 22.08 52.315 ;
    RECT 21.87 52.605 22.08 52.675 ;
    RECT 18.09 51.885 18.3 51.955 ;
    RECT 18.09 52.245 18.3 52.315 ;
    RECT 18.09 52.605 18.3 52.675 ;
    RECT 18.55 51.885 18.76 51.955 ;
    RECT 18.55 52.245 18.76 52.315 ;
    RECT 18.55 52.605 18.76 52.675 ;
    RECT 14.77 51.885 14.98 51.955 ;
    RECT 14.77 52.245 14.98 52.315 ;
    RECT 14.77 52.605 14.98 52.675 ;
    RECT 15.23 51.885 15.44 51.955 ;
    RECT 15.23 52.245 15.44 52.315 ;
    RECT 15.23 52.605 15.44 52.675 ;
    RECT 11.45 51.885 11.66 51.955 ;
    RECT 11.45 52.245 11.66 52.315 ;
    RECT 11.45 52.605 11.66 52.675 ;
    RECT 11.91 51.885 12.12 51.955 ;
    RECT 11.91 52.245 12.12 52.315 ;
    RECT 11.91 52.605 12.12 52.675 ;
    RECT 8.13 51.885 8.34 51.955 ;
    RECT 8.13 52.245 8.34 52.315 ;
    RECT 8.13 52.605 8.34 52.675 ;
    RECT 8.59 51.885 8.8 51.955 ;
    RECT 8.59 52.245 8.8 52.315 ;
    RECT 8.59 52.605 8.8 52.675 ;
    RECT 4.81 51.885 5.02 51.955 ;
    RECT 4.81 52.245 5.02 52.315 ;
    RECT 4.81 52.605 5.02 52.675 ;
    RECT 5.27 51.885 5.48 51.955 ;
    RECT 5.27 52.245 5.48 52.315 ;
    RECT 5.27 52.605 5.48 52.675 ;
    RECT 164.17 51.885 164.38 51.955 ;
    RECT 164.17 52.245 164.38 52.315 ;
    RECT 164.17 52.605 164.38 52.675 ;
    RECT 164.63 51.885 164.84 51.955 ;
    RECT 164.63 52.245 164.84 52.315 ;
    RECT 164.63 52.605 164.84 52.675 ;
    RECT 1.49 51.885 1.7 51.955 ;
    RECT 1.49 52.245 1.7 52.315 ;
    RECT 1.49 52.605 1.7 52.675 ;
    RECT 1.95 51.885 2.16 51.955 ;
    RECT 1.95 52.245 2.16 52.315 ;
    RECT 1.95 52.605 2.16 52.675 ;
    RECT 160.85 51.885 161.06 51.955 ;
    RECT 160.85 52.245 161.06 52.315 ;
    RECT 160.85 52.605 161.06 52.675 ;
    RECT 161.31 51.885 161.52 51.955 ;
    RECT 161.31 52.245 161.52 52.315 ;
    RECT 161.31 52.605 161.52 52.675 ;
    RECT 157.53 51.885 157.74 51.955 ;
    RECT 157.53 52.245 157.74 52.315 ;
    RECT 157.53 52.605 157.74 52.675 ;
    RECT 157.99 51.885 158.2 51.955 ;
    RECT 157.99 52.245 158.2 52.315 ;
    RECT 157.99 52.605 158.2 52.675 ;
    RECT 154.21 51.885 154.42 51.955 ;
    RECT 154.21 52.245 154.42 52.315 ;
    RECT 154.21 52.605 154.42 52.675 ;
    RECT 154.67 51.885 154.88 51.955 ;
    RECT 154.67 52.245 154.88 52.315 ;
    RECT 154.67 52.605 154.88 52.675 ;
    RECT 150.89 51.885 151.1 51.955 ;
    RECT 150.89 52.245 151.1 52.315 ;
    RECT 150.89 52.605 151.1 52.675 ;
    RECT 151.35 51.885 151.56 51.955 ;
    RECT 151.35 52.245 151.56 52.315 ;
    RECT 151.35 52.605 151.56 52.675 ;
    RECT 147.57 51.885 147.78 51.955 ;
    RECT 147.57 52.245 147.78 52.315 ;
    RECT 147.57 52.605 147.78 52.675 ;
    RECT 148.03 51.885 148.24 51.955 ;
    RECT 148.03 52.245 148.24 52.315 ;
    RECT 148.03 52.605 148.24 52.675 ;
    RECT 144.25 51.885 144.46 51.955 ;
    RECT 144.25 52.245 144.46 52.315 ;
    RECT 144.25 52.605 144.46 52.675 ;
    RECT 144.71 51.885 144.92 51.955 ;
    RECT 144.71 52.245 144.92 52.315 ;
    RECT 144.71 52.605 144.92 52.675 ;
    RECT 140.93 51.885 141.14 51.955 ;
    RECT 140.93 52.245 141.14 52.315 ;
    RECT 140.93 52.605 141.14 52.675 ;
    RECT 141.39 51.885 141.6 51.955 ;
    RECT 141.39 52.245 141.6 52.315 ;
    RECT 141.39 52.605 141.6 52.675 ;
    RECT 137.61 51.885 137.82 51.955 ;
    RECT 137.61 52.245 137.82 52.315 ;
    RECT 137.61 52.605 137.82 52.675 ;
    RECT 138.07 51.885 138.28 51.955 ;
    RECT 138.07 52.245 138.28 52.315 ;
    RECT 138.07 52.605 138.28 52.675 ;
    RECT 134.29 51.885 134.5 51.955 ;
    RECT 134.29 52.245 134.5 52.315 ;
    RECT 134.29 52.605 134.5 52.675 ;
    RECT 134.75 51.885 134.96 51.955 ;
    RECT 134.75 52.245 134.96 52.315 ;
    RECT 134.75 52.605 134.96 52.675 ;
    RECT 64.57 51.885 64.78 51.955 ;
    RECT 64.57 52.245 64.78 52.315 ;
    RECT 64.57 52.605 64.78 52.675 ;
    RECT 65.03 51.885 65.24 51.955 ;
    RECT 65.03 52.245 65.24 52.315 ;
    RECT 65.03 52.605 65.24 52.675 ;
    RECT 61.25 51.165 61.46 51.235 ;
    RECT 61.25 51.525 61.46 51.595 ;
    RECT 61.25 51.885 61.46 51.955 ;
    RECT 61.71 51.165 61.92 51.235 ;
    RECT 61.71 51.525 61.92 51.595 ;
    RECT 61.71 51.885 61.92 51.955 ;
    RECT 57.93 51.165 58.14 51.235 ;
    RECT 57.93 51.525 58.14 51.595 ;
    RECT 57.93 51.885 58.14 51.955 ;
    RECT 58.39 51.165 58.6 51.235 ;
    RECT 58.39 51.525 58.6 51.595 ;
    RECT 58.39 51.885 58.6 51.955 ;
    RECT 54.61 51.165 54.82 51.235 ;
    RECT 54.61 51.525 54.82 51.595 ;
    RECT 54.61 51.885 54.82 51.955 ;
    RECT 55.07 51.165 55.28 51.235 ;
    RECT 55.07 51.525 55.28 51.595 ;
    RECT 55.07 51.885 55.28 51.955 ;
    RECT 51.29 51.165 51.5 51.235 ;
    RECT 51.29 51.525 51.5 51.595 ;
    RECT 51.29 51.885 51.5 51.955 ;
    RECT 51.75 51.165 51.96 51.235 ;
    RECT 51.75 51.525 51.96 51.595 ;
    RECT 51.75 51.885 51.96 51.955 ;
    RECT 47.97 51.165 48.18 51.235 ;
    RECT 47.97 51.525 48.18 51.595 ;
    RECT 47.97 51.885 48.18 51.955 ;
    RECT 48.43 51.165 48.64 51.235 ;
    RECT 48.43 51.525 48.64 51.595 ;
    RECT 48.43 51.885 48.64 51.955 ;
    RECT 44.65 51.165 44.86 51.235 ;
    RECT 44.65 51.525 44.86 51.595 ;
    RECT 44.65 51.885 44.86 51.955 ;
    RECT 45.11 51.165 45.32 51.235 ;
    RECT 45.11 51.525 45.32 51.595 ;
    RECT 45.11 51.885 45.32 51.955 ;
    RECT 41.33 51.165 41.54 51.235 ;
    RECT 41.33 51.525 41.54 51.595 ;
    RECT 41.33 51.885 41.54 51.955 ;
    RECT 41.79 51.165 42.0 51.235 ;
    RECT 41.79 51.525 42.0 51.595 ;
    RECT 41.79 51.885 42.0 51.955 ;
    RECT 38.01 51.165 38.22 51.235 ;
    RECT 38.01 51.525 38.22 51.595 ;
    RECT 38.01 51.885 38.22 51.955 ;
    RECT 38.47 51.165 38.68 51.235 ;
    RECT 38.47 51.525 38.68 51.595 ;
    RECT 38.47 51.885 38.68 51.955 ;
    RECT 34.69 51.165 34.9 51.235 ;
    RECT 34.69 51.525 34.9 51.595 ;
    RECT 34.69 51.885 34.9 51.955 ;
    RECT 35.15 51.165 35.36 51.235 ;
    RECT 35.15 51.525 35.36 51.595 ;
    RECT 35.15 51.885 35.36 51.955 ;
    RECT 173.945 51.525 174.015 51.595 ;
    RECT 130.97 51.165 131.18 51.235 ;
    RECT 130.97 51.525 131.18 51.595 ;
    RECT 130.97 51.885 131.18 51.955 ;
    RECT 131.43 51.165 131.64 51.235 ;
    RECT 131.43 51.525 131.64 51.595 ;
    RECT 131.43 51.885 131.64 51.955 ;
    RECT 127.65 51.165 127.86 51.235 ;
    RECT 127.65 51.525 127.86 51.595 ;
    RECT 127.65 51.885 127.86 51.955 ;
    RECT 128.11 51.165 128.32 51.235 ;
    RECT 128.11 51.525 128.32 51.595 ;
    RECT 128.11 51.885 128.32 51.955 ;
    RECT 124.33 51.165 124.54 51.235 ;
    RECT 124.33 51.525 124.54 51.595 ;
    RECT 124.33 51.885 124.54 51.955 ;
    RECT 124.79 51.165 125.0 51.235 ;
    RECT 124.79 51.525 125.0 51.595 ;
    RECT 124.79 51.885 125.0 51.955 ;
    RECT 121.01 51.165 121.22 51.235 ;
    RECT 121.01 51.525 121.22 51.595 ;
    RECT 121.01 51.885 121.22 51.955 ;
    RECT 121.47 51.165 121.68 51.235 ;
    RECT 121.47 51.525 121.68 51.595 ;
    RECT 121.47 51.885 121.68 51.955 ;
    RECT 117.69 51.165 117.9 51.235 ;
    RECT 117.69 51.525 117.9 51.595 ;
    RECT 117.69 51.885 117.9 51.955 ;
    RECT 118.15 51.165 118.36 51.235 ;
    RECT 118.15 51.525 118.36 51.595 ;
    RECT 118.15 51.885 118.36 51.955 ;
    RECT 114.37 51.165 114.58 51.235 ;
    RECT 114.37 51.525 114.58 51.595 ;
    RECT 114.37 51.885 114.58 51.955 ;
    RECT 114.83 51.165 115.04 51.235 ;
    RECT 114.83 51.525 115.04 51.595 ;
    RECT 114.83 51.885 115.04 51.955 ;
    RECT 111.05 51.165 111.26 51.235 ;
    RECT 111.05 51.525 111.26 51.595 ;
    RECT 111.05 51.885 111.26 51.955 ;
    RECT 111.51 51.165 111.72 51.235 ;
    RECT 111.51 51.525 111.72 51.595 ;
    RECT 111.51 51.885 111.72 51.955 ;
    RECT 107.73 51.165 107.94 51.235 ;
    RECT 107.73 51.525 107.94 51.595 ;
    RECT 107.73 51.885 107.94 51.955 ;
    RECT 108.19 51.165 108.4 51.235 ;
    RECT 108.19 51.525 108.4 51.595 ;
    RECT 108.19 51.885 108.4 51.955 ;
    RECT 104.41 51.165 104.62 51.235 ;
    RECT 104.41 51.525 104.62 51.595 ;
    RECT 104.41 51.885 104.62 51.955 ;
    RECT 104.87 51.165 105.08 51.235 ;
    RECT 104.87 51.525 105.08 51.595 ;
    RECT 104.87 51.885 105.08 51.955 ;
    RECT 101.09 51.165 101.3 51.235 ;
    RECT 101.09 51.525 101.3 51.595 ;
    RECT 101.09 51.885 101.3 51.955 ;
    RECT 101.55 51.165 101.76 51.235 ;
    RECT 101.55 51.525 101.76 51.595 ;
    RECT 101.55 51.885 101.76 51.955 ;
    RECT 0.4 51.525 0.47 51.595 ;
    RECT 170.81 51.165 171.02 51.235 ;
    RECT 170.81 51.525 171.02 51.595 ;
    RECT 170.81 51.885 171.02 51.955 ;
    RECT 171.27 51.165 171.48 51.235 ;
    RECT 171.27 51.525 171.48 51.595 ;
    RECT 171.27 51.885 171.48 51.955 ;
    RECT 167.49 51.165 167.7 51.235 ;
    RECT 167.49 51.525 167.7 51.595 ;
    RECT 167.49 51.885 167.7 51.955 ;
    RECT 167.95 51.165 168.16 51.235 ;
    RECT 167.95 51.525 168.16 51.595 ;
    RECT 167.95 51.885 168.16 51.955 ;
    RECT 97.77 51.165 97.98 51.235 ;
    RECT 97.77 51.525 97.98 51.595 ;
    RECT 97.77 51.885 97.98 51.955 ;
    RECT 98.23 51.165 98.44 51.235 ;
    RECT 98.23 51.525 98.44 51.595 ;
    RECT 98.23 51.885 98.44 51.955 ;
    RECT 94.45 51.165 94.66 51.235 ;
    RECT 94.45 51.525 94.66 51.595 ;
    RECT 94.45 51.885 94.66 51.955 ;
    RECT 94.91 51.165 95.12 51.235 ;
    RECT 94.91 51.525 95.12 51.595 ;
    RECT 94.91 51.885 95.12 51.955 ;
    RECT 91.13 51.165 91.34 51.235 ;
    RECT 91.13 51.525 91.34 51.595 ;
    RECT 91.13 51.885 91.34 51.955 ;
    RECT 91.59 51.165 91.8 51.235 ;
    RECT 91.59 51.525 91.8 51.595 ;
    RECT 91.59 51.885 91.8 51.955 ;
    RECT 87.81 51.165 88.02 51.235 ;
    RECT 87.81 51.525 88.02 51.595 ;
    RECT 87.81 51.885 88.02 51.955 ;
    RECT 88.27 51.165 88.48 51.235 ;
    RECT 88.27 51.525 88.48 51.595 ;
    RECT 88.27 51.885 88.48 51.955 ;
    RECT 84.49 51.165 84.7 51.235 ;
    RECT 84.49 51.525 84.7 51.595 ;
    RECT 84.49 51.885 84.7 51.955 ;
    RECT 84.95 51.165 85.16 51.235 ;
    RECT 84.95 51.525 85.16 51.595 ;
    RECT 84.95 51.885 85.16 51.955 ;
    RECT 81.17 51.165 81.38 51.235 ;
    RECT 81.17 51.525 81.38 51.595 ;
    RECT 81.17 51.885 81.38 51.955 ;
    RECT 81.63 51.165 81.84 51.235 ;
    RECT 81.63 51.525 81.84 51.595 ;
    RECT 81.63 51.885 81.84 51.955 ;
    RECT 77.85 51.165 78.06 51.235 ;
    RECT 77.85 51.525 78.06 51.595 ;
    RECT 77.85 51.885 78.06 51.955 ;
    RECT 78.31 51.165 78.52 51.235 ;
    RECT 78.31 51.525 78.52 51.595 ;
    RECT 78.31 51.885 78.52 51.955 ;
    RECT 74.53 51.165 74.74 51.235 ;
    RECT 74.53 51.525 74.74 51.595 ;
    RECT 74.53 51.885 74.74 51.955 ;
    RECT 74.99 51.165 75.2 51.235 ;
    RECT 74.99 51.525 75.2 51.595 ;
    RECT 74.99 51.885 75.2 51.955 ;
    RECT 71.21 51.165 71.42 51.235 ;
    RECT 71.21 51.525 71.42 51.595 ;
    RECT 71.21 51.885 71.42 51.955 ;
    RECT 71.67 51.165 71.88 51.235 ;
    RECT 71.67 51.525 71.88 51.595 ;
    RECT 71.67 51.885 71.88 51.955 ;
    RECT 31.37 51.165 31.58 51.235 ;
    RECT 31.37 51.525 31.58 51.595 ;
    RECT 31.37 51.885 31.58 51.955 ;
    RECT 31.83 51.165 32.04 51.235 ;
    RECT 31.83 51.525 32.04 51.595 ;
    RECT 31.83 51.885 32.04 51.955 ;
    RECT 67.89 51.165 68.1 51.235 ;
    RECT 67.89 51.525 68.1 51.595 ;
    RECT 67.89 51.885 68.1 51.955 ;
    RECT 68.35 51.165 68.56 51.235 ;
    RECT 68.35 51.525 68.56 51.595 ;
    RECT 68.35 51.885 68.56 51.955 ;
    RECT 28.05 51.165 28.26 51.235 ;
    RECT 28.05 51.525 28.26 51.595 ;
    RECT 28.05 51.885 28.26 51.955 ;
    RECT 28.51 51.165 28.72 51.235 ;
    RECT 28.51 51.525 28.72 51.595 ;
    RECT 28.51 51.885 28.72 51.955 ;
    RECT 24.73 51.165 24.94 51.235 ;
    RECT 24.73 51.525 24.94 51.595 ;
    RECT 24.73 51.885 24.94 51.955 ;
    RECT 25.19 51.165 25.4 51.235 ;
    RECT 25.19 51.525 25.4 51.595 ;
    RECT 25.19 51.885 25.4 51.955 ;
    RECT 21.41 51.165 21.62 51.235 ;
    RECT 21.41 51.525 21.62 51.595 ;
    RECT 21.41 51.885 21.62 51.955 ;
    RECT 21.87 51.165 22.08 51.235 ;
    RECT 21.87 51.525 22.08 51.595 ;
    RECT 21.87 51.885 22.08 51.955 ;
    RECT 18.09 51.165 18.3 51.235 ;
    RECT 18.09 51.525 18.3 51.595 ;
    RECT 18.09 51.885 18.3 51.955 ;
    RECT 18.55 51.165 18.76 51.235 ;
    RECT 18.55 51.525 18.76 51.595 ;
    RECT 18.55 51.885 18.76 51.955 ;
    RECT 14.77 51.165 14.98 51.235 ;
    RECT 14.77 51.525 14.98 51.595 ;
    RECT 14.77 51.885 14.98 51.955 ;
    RECT 15.23 51.165 15.44 51.235 ;
    RECT 15.23 51.525 15.44 51.595 ;
    RECT 15.23 51.885 15.44 51.955 ;
    RECT 11.45 51.165 11.66 51.235 ;
    RECT 11.45 51.525 11.66 51.595 ;
    RECT 11.45 51.885 11.66 51.955 ;
    RECT 11.91 51.165 12.12 51.235 ;
    RECT 11.91 51.525 12.12 51.595 ;
    RECT 11.91 51.885 12.12 51.955 ;
    RECT 8.13 51.165 8.34 51.235 ;
    RECT 8.13 51.525 8.34 51.595 ;
    RECT 8.13 51.885 8.34 51.955 ;
    RECT 8.59 51.165 8.8 51.235 ;
    RECT 8.59 51.525 8.8 51.595 ;
    RECT 8.59 51.885 8.8 51.955 ;
    RECT 4.81 51.165 5.02 51.235 ;
    RECT 4.81 51.525 5.02 51.595 ;
    RECT 4.81 51.885 5.02 51.955 ;
    RECT 5.27 51.165 5.48 51.235 ;
    RECT 5.27 51.525 5.48 51.595 ;
    RECT 5.27 51.885 5.48 51.955 ;
    RECT 164.17 51.165 164.38 51.235 ;
    RECT 164.17 51.525 164.38 51.595 ;
    RECT 164.17 51.885 164.38 51.955 ;
    RECT 164.63 51.165 164.84 51.235 ;
    RECT 164.63 51.525 164.84 51.595 ;
    RECT 164.63 51.885 164.84 51.955 ;
    RECT 1.49 51.165 1.7 51.235 ;
    RECT 1.49 51.525 1.7 51.595 ;
    RECT 1.49 51.885 1.7 51.955 ;
    RECT 1.95 51.165 2.16 51.235 ;
    RECT 1.95 51.525 2.16 51.595 ;
    RECT 1.95 51.885 2.16 51.955 ;
    RECT 160.85 51.165 161.06 51.235 ;
    RECT 160.85 51.525 161.06 51.595 ;
    RECT 160.85 51.885 161.06 51.955 ;
    RECT 161.31 51.165 161.52 51.235 ;
    RECT 161.31 51.525 161.52 51.595 ;
    RECT 161.31 51.885 161.52 51.955 ;
    RECT 157.53 51.165 157.74 51.235 ;
    RECT 157.53 51.525 157.74 51.595 ;
    RECT 157.53 51.885 157.74 51.955 ;
    RECT 157.99 51.165 158.2 51.235 ;
    RECT 157.99 51.525 158.2 51.595 ;
    RECT 157.99 51.885 158.2 51.955 ;
    RECT 154.21 51.165 154.42 51.235 ;
    RECT 154.21 51.525 154.42 51.595 ;
    RECT 154.21 51.885 154.42 51.955 ;
    RECT 154.67 51.165 154.88 51.235 ;
    RECT 154.67 51.525 154.88 51.595 ;
    RECT 154.67 51.885 154.88 51.955 ;
    RECT 150.89 51.165 151.1 51.235 ;
    RECT 150.89 51.525 151.1 51.595 ;
    RECT 150.89 51.885 151.1 51.955 ;
    RECT 151.35 51.165 151.56 51.235 ;
    RECT 151.35 51.525 151.56 51.595 ;
    RECT 151.35 51.885 151.56 51.955 ;
    RECT 147.57 51.165 147.78 51.235 ;
    RECT 147.57 51.525 147.78 51.595 ;
    RECT 147.57 51.885 147.78 51.955 ;
    RECT 148.03 51.165 148.24 51.235 ;
    RECT 148.03 51.525 148.24 51.595 ;
    RECT 148.03 51.885 148.24 51.955 ;
    RECT 144.25 51.165 144.46 51.235 ;
    RECT 144.25 51.525 144.46 51.595 ;
    RECT 144.25 51.885 144.46 51.955 ;
    RECT 144.71 51.165 144.92 51.235 ;
    RECT 144.71 51.525 144.92 51.595 ;
    RECT 144.71 51.885 144.92 51.955 ;
    RECT 140.93 51.165 141.14 51.235 ;
    RECT 140.93 51.525 141.14 51.595 ;
    RECT 140.93 51.885 141.14 51.955 ;
    RECT 141.39 51.165 141.6 51.235 ;
    RECT 141.39 51.525 141.6 51.595 ;
    RECT 141.39 51.885 141.6 51.955 ;
    RECT 137.61 51.165 137.82 51.235 ;
    RECT 137.61 51.525 137.82 51.595 ;
    RECT 137.61 51.885 137.82 51.955 ;
    RECT 138.07 51.165 138.28 51.235 ;
    RECT 138.07 51.525 138.28 51.595 ;
    RECT 138.07 51.885 138.28 51.955 ;
    RECT 134.29 51.165 134.5 51.235 ;
    RECT 134.29 51.525 134.5 51.595 ;
    RECT 134.29 51.885 134.5 51.955 ;
    RECT 134.75 51.165 134.96 51.235 ;
    RECT 134.75 51.525 134.96 51.595 ;
    RECT 134.75 51.885 134.96 51.955 ;
    RECT 64.57 51.165 64.78 51.235 ;
    RECT 64.57 51.525 64.78 51.595 ;
    RECT 64.57 51.885 64.78 51.955 ;
    RECT 65.03 51.165 65.24 51.235 ;
    RECT 65.03 51.525 65.24 51.595 ;
    RECT 65.03 51.885 65.24 51.955 ;
    RECT 61.25 50.445 61.46 50.515 ;
    RECT 61.25 50.805 61.46 50.875 ;
    RECT 61.25 51.165 61.46 51.235 ;
    RECT 61.71 50.445 61.92 50.515 ;
    RECT 61.71 50.805 61.92 50.875 ;
    RECT 61.71 51.165 61.92 51.235 ;
    RECT 57.93 50.445 58.14 50.515 ;
    RECT 57.93 50.805 58.14 50.875 ;
    RECT 57.93 51.165 58.14 51.235 ;
    RECT 58.39 50.445 58.6 50.515 ;
    RECT 58.39 50.805 58.6 50.875 ;
    RECT 58.39 51.165 58.6 51.235 ;
    RECT 54.61 50.445 54.82 50.515 ;
    RECT 54.61 50.805 54.82 50.875 ;
    RECT 54.61 51.165 54.82 51.235 ;
    RECT 55.07 50.445 55.28 50.515 ;
    RECT 55.07 50.805 55.28 50.875 ;
    RECT 55.07 51.165 55.28 51.235 ;
    RECT 51.29 50.445 51.5 50.515 ;
    RECT 51.29 50.805 51.5 50.875 ;
    RECT 51.29 51.165 51.5 51.235 ;
    RECT 51.75 50.445 51.96 50.515 ;
    RECT 51.75 50.805 51.96 50.875 ;
    RECT 51.75 51.165 51.96 51.235 ;
    RECT 47.97 50.445 48.18 50.515 ;
    RECT 47.97 50.805 48.18 50.875 ;
    RECT 47.97 51.165 48.18 51.235 ;
    RECT 48.43 50.445 48.64 50.515 ;
    RECT 48.43 50.805 48.64 50.875 ;
    RECT 48.43 51.165 48.64 51.235 ;
    RECT 44.65 50.445 44.86 50.515 ;
    RECT 44.65 50.805 44.86 50.875 ;
    RECT 44.65 51.165 44.86 51.235 ;
    RECT 45.11 50.445 45.32 50.515 ;
    RECT 45.11 50.805 45.32 50.875 ;
    RECT 45.11 51.165 45.32 51.235 ;
    RECT 41.33 50.445 41.54 50.515 ;
    RECT 41.33 50.805 41.54 50.875 ;
    RECT 41.33 51.165 41.54 51.235 ;
    RECT 41.79 50.445 42.0 50.515 ;
    RECT 41.79 50.805 42.0 50.875 ;
    RECT 41.79 51.165 42.0 51.235 ;
    RECT 38.01 50.445 38.22 50.515 ;
    RECT 38.01 50.805 38.22 50.875 ;
    RECT 38.01 51.165 38.22 51.235 ;
    RECT 38.47 50.445 38.68 50.515 ;
    RECT 38.47 50.805 38.68 50.875 ;
    RECT 38.47 51.165 38.68 51.235 ;
    RECT 34.69 50.445 34.9 50.515 ;
    RECT 34.69 50.805 34.9 50.875 ;
    RECT 34.69 51.165 34.9 51.235 ;
    RECT 35.15 50.445 35.36 50.515 ;
    RECT 35.15 50.805 35.36 50.875 ;
    RECT 35.15 51.165 35.36 51.235 ;
    RECT 173.945 50.805 174.015 50.875 ;
    RECT 130.97 50.445 131.18 50.515 ;
    RECT 130.97 50.805 131.18 50.875 ;
    RECT 130.97 51.165 131.18 51.235 ;
    RECT 131.43 50.445 131.64 50.515 ;
    RECT 131.43 50.805 131.64 50.875 ;
    RECT 131.43 51.165 131.64 51.235 ;
    RECT 127.65 50.445 127.86 50.515 ;
    RECT 127.65 50.805 127.86 50.875 ;
    RECT 127.65 51.165 127.86 51.235 ;
    RECT 128.11 50.445 128.32 50.515 ;
    RECT 128.11 50.805 128.32 50.875 ;
    RECT 128.11 51.165 128.32 51.235 ;
    RECT 124.33 50.445 124.54 50.515 ;
    RECT 124.33 50.805 124.54 50.875 ;
    RECT 124.33 51.165 124.54 51.235 ;
    RECT 124.79 50.445 125.0 50.515 ;
    RECT 124.79 50.805 125.0 50.875 ;
    RECT 124.79 51.165 125.0 51.235 ;
    RECT 121.01 50.445 121.22 50.515 ;
    RECT 121.01 50.805 121.22 50.875 ;
    RECT 121.01 51.165 121.22 51.235 ;
    RECT 121.47 50.445 121.68 50.515 ;
    RECT 121.47 50.805 121.68 50.875 ;
    RECT 121.47 51.165 121.68 51.235 ;
    RECT 117.69 50.445 117.9 50.515 ;
    RECT 117.69 50.805 117.9 50.875 ;
    RECT 117.69 51.165 117.9 51.235 ;
    RECT 118.15 50.445 118.36 50.515 ;
    RECT 118.15 50.805 118.36 50.875 ;
    RECT 118.15 51.165 118.36 51.235 ;
    RECT 114.37 50.445 114.58 50.515 ;
    RECT 114.37 50.805 114.58 50.875 ;
    RECT 114.37 51.165 114.58 51.235 ;
    RECT 114.83 50.445 115.04 50.515 ;
    RECT 114.83 50.805 115.04 50.875 ;
    RECT 114.83 51.165 115.04 51.235 ;
    RECT 111.05 50.445 111.26 50.515 ;
    RECT 111.05 50.805 111.26 50.875 ;
    RECT 111.05 51.165 111.26 51.235 ;
    RECT 111.51 50.445 111.72 50.515 ;
    RECT 111.51 50.805 111.72 50.875 ;
    RECT 111.51 51.165 111.72 51.235 ;
    RECT 107.73 50.445 107.94 50.515 ;
    RECT 107.73 50.805 107.94 50.875 ;
    RECT 107.73 51.165 107.94 51.235 ;
    RECT 108.19 50.445 108.4 50.515 ;
    RECT 108.19 50.805 108.4 50.875 ;
    RECT 108.19 51.165 108.4 51.235 ;
    RECT 104.41 50.445 104.62 50.515 ;
    RECT 104.41 50.805 104.62 50.875 ;
    RECT 104.41 51.165 104.62 51.235 ;
    RECT 104.87 50.445 105.08 50.515 ;
    RECT 104.87 50.805 105.08 50.875 ;
    RECT 104.87 51.165 105.08 51.235 ;
    RECT 101.09 50.445 101.3 50.515 ;
    RECT 101.09 50.805 101.3 50.875 ;
    RECT 101.09 51.165 101.3 51.235 ;
    RECT 101.55 50.445 101.76 50.515 ;
    RECT 101.55 50.805 101.76 50.875 ;
    RECT 101.55 51.165 101.76 51.235 ;
    RECT 0.4 50.805 0.47 50.875 ;
    RECT 170.81 50.445 171.02 50.515 ;
    RECT 170.81 50.805 171.02 50.875 ;
    RECT 170.81 51.165 171.02 51.235 ;
    RECT 171.27 50.445 171.48 50.515 ;
    RECT 171.27 50.805 171.48 50.875 ;
    RECT 171.27 51.165 171.48 51.235 ;
    RECT 167.49 50.445 167.7 50.515 ;
    RECT 167.49 50.805 167.7 50.875 ;
    RECT 167.49 51.165 167.7 51.235 ;
    RECT 167.95 50.445 168.16 50.515 ;
    RECT 167.95 50.805 168.16 50.875 ;
    RECT 167.95 51.165 168.16 51.235 ;
    RECT 97.77 50.445 97.98 50.515 ;
    RECT 97.77 50.805 97.98 50.875 ;
    RECT 97.77 51.165 97.98 51.235 ;
    RECT 98.23 50.445 98.44 50.515 ;
    RECT 98.23 50.805 98.44 50.875 ;
    RECT 98.23 51.165 98.44 51.235 ;
    RECT 94.45 50.445 94.66 50.515 ;
    RECT 94.45 50.805 94.66 50.875 ;
    RECT 94.45 51.165 94.66 51.235 ;
    RECT 94.91 50.445 95.12 50.515 ;
    RECT 94.91 50.805 95.12 50.875 ;
    RECT 94.91 51.165 95.12 51.235 ;
    RECT 91.13 50.445 91.34 50.515 ;
    RECT 91.13 50.805 91.34 50.875 ;
    RECT 91.13 51.165 91.34 51.235 ;
    RECT 91.59 50.445 91.8 50.515 ;
    RECT 91.59 50.805 91.8 50.875 ;
    RECT 91.59 51.165 91.8 51.235 ;
    RECT 87.81 50.445 88.02 50.515 ;
    RECT 87.81 50.805 88.02 50.875 ;
    RECT 87.81 51.165 88.02 51.235 ;
    RECT 88.27 50.445 88.48 50.515 ;
    RECT 88.27 50.805 88.48 50.875 ;
    RECT 88.27 51.165 88.48 51.235 ;
    RECT 84.49 50.445 84.7 50.515 ;
    RECT 84.49 50.805 84.7 50.875 ;
    RECT 84.49 51.165 84.7 51.235 ;
    RECT 84.95 50.445 85.16 50.515 ;
    RECT 84.95 50.805 85.16 50.875 ;
    RECT 84.95 51.165 85.16 51.235 ;
    RECT 81.17 50.445 81.38 50.515 ;
    RECT 81.17 50.805 81.38 50.875 ;
    RECT 81.17 51.165 81.38 51.235 ;
    RECT 81.63 50.445 81.84 50.515 ;
    RECT 81.63 50.805 81.84 50.875 ;
    RECT 81.63 51.165 81.84 51.235 ;
    RECT 77.85 50.445 78.06 50.515 ;
    RECT 77.85 50.805 78.06 50.875 ;
    RECT 77.85 51.165 78.06 51.235 ;
    RECT 78.31 50.445 78.52 50.515 ;
    RECT 78.31 50.805 78.52 50.875 ;
    RECT 78.31 51.165 78.52 51.235 ;
    RECT 74.53 50.445 74.74 50.515 ;
    RECT 74.53 50.805 74.74 50.875 ;
    RECT 74.53 51.165 74.74 51.235 ;
    RECT 74.99 50.445 75.2 50.515 ;
    RECT 74.99 50.805 75.2 50.875 ;
    RECT 74.99 51.165 75.2 51.235 ;
    RECT 71.21 50.445 71.42 50.515 ;
    RECT 71.21 50.805 71.42 50.875 ;
    RECT 71.21 51.165 71.42 51.235 ;
    RECT 71.67 50.445 71.88 50.515 ;
    RECT 71.67 50.805 71.88 50.875 ;
    RECT 71.67 51.165 71.88 51.235 ;
    RECT 31.37 50.445 31.58 50.515 ;
    RECT 31.37 50.805 31.58 50.875 ;
    RECT 31.37 51.165 31.58 51.235 ;
    RECT 31.83 50.445 32.04 50.515 ;
    RECT 31.83 50.805 32.04 50.875 ;
    RECT 31.83 51.165 32.04 51.235 ;
    RECT 67.89 50.445 68.1 50.515 ;
    RECT 67.89 50.805 68.1 50.875 ;
    RECT 67.89 51.165 68.1 51.235 ;
    RECT 68.35 50.445 68.56 50.515 ;
    RECT 68.35 50.805 68.56 50.875 ;
    RECT 68.35 51.165 68.56 51.235 ;
    RECT 28.05 50.445 28.26 50.515 ;
    RECT 28.05 50.805 28.26 50.875 ;
    RECT 28.05 51.165 28.26 51.235 ;
    RECT 28.51 50.445 28.72 50.515 ;
    RECT 28.51 50.805 28.72 50.875 ;
    RECT 28.51 51.165 28.72 51.235 ;
    RECT 24.73 50.445 24.94 50.515 ;
    RECT 24.73 50.805 24.94 50.875 ;
    RECT 24.73 51.165 24.94 51.235 ;
    RECT 25.19 50.445 25.4 50.515 ;
    RECT 25.19 50.805 25.4 50.875 ;
    RECT 25.19 51.165 25.4 51.235 ;
    RECT 21.41 50.445 21.62 50.515 ;
    RECT 21.41 50.805 21.62 50.875 ;
    RECT 21.41 51.165 21.62 51.235 ;
    RECT 21.87 50.445 22.08 50.515 ;
    RECT 21.87 50.805 22.08 50.875 ;
    RECT 21.87 51.165 22.08 51.235 ;
    RECT 18.09 50.445 18.3 50.515 ;
    RECT 18.09 50.805 18.3 50.875 ;
    RECT 18.09 51.165 18.3 51.235 ;
    RECT 18.55 50.445 18.76 50.515 ;
    RECT 18.55 50.805 18.76 50.875 ;
    RECT 18.55 51.165 18.76 51.235 ;
    RECT 14.77 50.445 14.98 50.515 ;
    RECT 14.77 50.805 14.98 50.875 ;
    RECT 14.77 51.165 14.98 51.235 ;
    RECT 15.23 50.445 15.44 50.515 ;
    RECT 15.23 50.805 15.44 50.875 ;
    RECT 15.23 51.165 15.44 51.235 ;
    RECT 11.45 50.445 11.66 50.515 ;
    RECT 11.45 50.805 11.66 50.875 ;
    RECT 11.45 51.165 11.66 51.235 ;
    RECT 11.91 50.445 12.12 50.515 ;
    RECT 11.91 50.805 12.12 50.875 ;
    RECT 11.91 51.165 12.12 51.235 ;
    RECT 8.13 50.445 8.34 50.515 ;
    RECT 8.13 50.805 8.34 50.875 ;
    RECT 8.13 51.165 8.34 51.235 ;
    RECT 8.59 50.445 8.8 50.515 ;
    RECT 8.59 50.805 8.8 50.875 ;
    RECT 8.59 51.165 8.8 51.235 ;
    RECT 4.81 50.445 5.02 50.515 ;
    RECT 4.81 50.805 5.02 50.875 ;
    RECT 4.81 51.165 5.02 51.235 ;
    RECT 5.27 50.445 5.48 50.515 ;
    RECT 5.27 50.805 5.48 50.875 ;
    RECT 5.27 51.165 5.48 51.235 ;
    RECT 164.17 50.445 164.38 50.515 ;
    RECT 164.17 50.805 164.38 50.875 ;
    RECT 164.17 51.165 164.38 51.235 ;
    RECT 164.63 50.445 164.84 50.515 ;
    RECT 164.63 50.805 164.84 50.875 ;
    RECT 164.63 51.165 164.84 51.235 ;
    RECT 1.49 50.445 1.7 50.515 ;
    RECT 1.49 50.805 1.7 50.875 ;
    RECT 1.49 51.165 1.7 51.235 ;
    RECT 1.95 50.445 2.16 50.515 ;
    RECT 1.95 50.805 2.16 50.875 ;
    RECT 1.95 51.165 2.16 51.235 ;
    RECT 160.85 50.445 161.06 50.515 ;
    RECT 160.85 50.805 161.06 50.875 ;
    RECT 160.85 51.165 161.06 51.235 ;
    RECT 161.31 50.445 161.52 50.515 ;
    RECT 161.31 50.805 161.52 50.875 ;
    RECT 161.31 51.165 161.52 51.235 ;
    RECT 157.53 50.445 157.74 50.515 ;
    RECT 157.53 50.805 157.74 50.875 ;
    RECT 157.53 51.165 157.74 51.235 ;
    RECT 157.99 50.445 158.2 50.515 ;
    RECT 157.99 50.805 158.2 50.875 ;
    RECT 157.99 51.165 158.2 51.235 ;
    RECT 154.21 50.445 154.42 50.515 ;
    RECT 154.21 50.805 154.42 50.875 ;
    RECT 154.21 51.165 154.42 51.235 ;
    RECT 154.67 50.445 154.88 50.515 ;
    RECT 154.67 50.805 154.88 50.875 ;
    RECT 154.67 51.165 154.88 51.235 ;
    RECT 150.89 50.445 151.1 50.515 ;
    RECT 150.89 50.805 151.1 50.875 ;
    RECT 150.89 51.165 151.1 51.235 ;
    RECT 151.35 50.445 151.56 50.515 ;
    RECT 151.35 50.805 151.56 50.875 ;
    RECT 151.35 51.165 151.56 51.235 ;
    RECT 147.57 50.445 147.78 50.515 ;
    RECT 147.57 50.805 147.78 50.875 ;
    RECT 147.57 51.165 147.78 51.235 ;
    RECT 148.03 50.445 148.24 50.515 ;
    RECT 148.03 50.805 148.24 50.875 ;
    RECT 148.03 51.165 148.24 51.235 ;
    RECT 144.25 50.445 144.46 50.515 ;
    RECT 144.25 50.805 144.46 50.875 ;
    RECT 144.25 51.165 144.46 51.235 ;
    RECT 144.71 50.445 144.92 50.515 ;
    RECT 144.71 50.805 144.92 50.875 ;
    RECT 144.71 51.165 144.92 51.235 ;
    RECT 140.93 50.445 141.14 50.515 ;
    RECT 140.93 50.805 141.14 50.875 ;
    RECT 140.93 51.165 141.14 51.235 ;
    RECT 141.39 50.445 141.6 50.515 ;
    RECT 141.39 50.805 141.6 50.875 ;
    RECT 141.39 51.165 141.6 51.235 ;
    RECT 137.61 50.445 137.82 50.515 ;
    RECT 137.61 50.805 137.82 50.875 ;
    RECT 137.61 51.165 137.82 51.235 ;
    RECT 138.07 50.445 138.28 50.515 ;
    RECT 138.07 50.805 138.28 50.875 ;
    RECT 138.07 51.165 138.28 51.235 ;
    RECT 134.29 50.445 134.5 50.515 ;
    RECT 134.29 50.805 134.5 50.875 ;
    RECT 134.29 51.165 134.5 51.235 ;
    RECT 134.75 50.445 134.96 50.515 ;
    RECT 134.75 50.805 134.96 50.875 ;
    RECT 134.75 51.165 134.96 51.235 ;
    RECT 64.57 50.445 64.78 50.515 ;
    RECT 64.57 50.805 64.78 50.875 ;
    RECT 64.57 51.165 64.78 51.235 ;
    RECT 65.03 50.445 65.24 50.515 ;
    RECT 65.03 50.805 65.24 50.875 ;
    RECT 65.03 51.165 65.24 51.235 ;
    RECT 175.75 51.525 175.96 51.595 ;
    RECT 186.51 35.592 186.58 35.662 ;
    RECT 174.56 56.925 174.63 57.715 ;
    RECT 175.16 56.925 175.37 56.995 ;
    RECT 175.16 57.28 175.37 57.35 ;
    RECT 175.16 57.645 175.37 57.715 ;
    RECT 176.325 57.37 177.125 57.44 ;
    RECT 178.79 57.195 179.025 57.265 ;
    RECT 179.85 57.195 180.11 57.265 ;
    RECT 181.825 57.195 182.055 57.265 ;
    RECT 182.54 57.195 182.8 57.265 ;
    RECT 183.71 57.195 183.78 57.265 ;
    RECT 187.045 57.195 187.255 57.265 ;
    RECT 187.43 57.195 187.7 57.265 ;
    RECT 191.485 57.195 191.555 57.265 ;
    RECT 191.815 57.195 192.08 57.265 ;
    RECT 193.57 57.195 193.83 57.265 ;
    RECT 194.015 57.195 194.085 57.265 ;
    RECT 194.505 57.195 194.765 57.265 ;
    RECT 195.63 57.195 195.84 57.265 ;
    RECT 197.44 57.37 198.255 57.44 ;
    RECT 199.245 56.925 199.515 56.995 ;
    RECT 199.245 57.28 199.515 57.35 ;
    RECT 199.245 57.645 199.515 57.715 ;
    RECT 174.56 56.205 174.63 56.995 ;
    RECT 175.16 56.205 175.37 56.275 ;
    RECT 175.16 56.56 175.37 56.63 ;
    RECT 175.16 56.925 175.37 56.995 ;
    RECT 176.325 56.65 177.125 56.72 ;
    RECT 178.79 56.475 179.025 56.545 ;
    RECT 179.85 56.475 180.11 56.545 ;
    RECT 181.825 56.475 182.055 56.545 ;
    RECT 182.54 56.475 182.8 56.545 ;
    RECT 183.71 56.475 183.78 56.545 ;
    RECT 187.045 56.475 187.255 56.545 ;
    RECT 187.43 56.475 187.7 56.545 ;
    RECT 191.485 56.475 191.555 56.545 ;
    RECT 191.815 56.475 192.08 56.545 ;
    RECT 193.57 56.475 193.83 56.545 ;
    RECT 194.015 56.475 194.085 56.545 ;
    RECT 194.505 56.475 194.765 56.545 ;
    RECT 195.63 56.475 195.84 56.545 ;
    RECT 197.44 56.65 198.255 56.72 ;
    RECT 199.245 56.205 199.515 56.275 ;
    RECT 199.245 56.56 199.515 56.63 ;
    RECT 199.245 56.925 199.515 56.995 ;
    RECT 188.225 41.352 188.295 41.422 ;
    RECT 198.605 50.805 198.815 50.875 ;
    RECT 192.85 50.715 193.06 50.785 ;
    RECT 175.75 26.325 175.96 26.395 ;
    RECT 175.75 25.605 175.96 25.675 ;
    RECT 175.75 24.885 175.96 24.955 ;
    RECT 175.75 24.165 175.96 24.235 ;
    RECT 174.56 55.485 174.63 56.275 ;
    RECT 175.16 55.485 175.37 55.555 ;
    RECT 175.16 55.84 175.37 55.91 ;
    RECT 175.16 56.205 175.37 56.275 ;
    RECT 176.325 55.93 177.125 56.0 ;
    RECT 178.79 55.755 179.025 55.825 ;
    RECT 179.85 55.755 180.11 55.825 ;
    RECT 181.825 55.755 182.055 55.825 ;
    RECT 182.54 55.755 182.8 55.825 ;
    RECT 183.71 55.755 183.78 55.825 ;
    RECT 187.045 55.755 187.255 55.825 ;
    RECT 187.43 55.755 187.7 55.825 ;
    RECT 191.485 55.755 191.555 55.825 ;
    RECT 191.815 55.755 192.08 55.825 ;
    RECT 193.57 55.755 193.83 55.825 ;
    RECT 194.015 55.755 194.085 55.825 ;
    RECT 194.505 55.755 194.765 55.825 ;
    RECT 195.63 55.755 195.84 55.825 ;
    RECT 197.44 55.93 198.255 56.0 ;
    RECT 199.245 55.485 199.515 55.555 ;
    RECT 199.245 55.84 199.515 55.91 ;
    RECT 199.245 56.205 199.515 56.275 ;
    RECT 174.56 54.765 174.63 55.555 ;
    RECT 175.16 54.765 175.37 54.835 ;
    RECT 175.16 55.12 175.37 55.19 ;
    RECT 175.16 55.485 175.37 55.555 ;
    RECT 176.325 55.21 177.125 55.28 ;
    RECT 178.79 55.035 179.025 55.105 ;
    RECT 179.85 55.035 180.11 55.105 ;
    RECT 181.825 55.035 182.055 55.105 ;
    RECT 182.54 55.035 182.8 55.105 ;
    RECT 183.71 55.035 183.78 55.105 ;
    RECT 187.045 55.035 187.255 55.105 ;
    RECT 187.43 55.035 187.7 55.105 ;
    RECT 191.485 55.035 191.555 55.105 ;
    RECT 191.815 55.035 192.08 55.105 ;
    RECT 193.57 55.035 193.83 55.105 ;
    RECT 194.015 55.035 194.085 55.105 ;
    RECT 194.505 55.035 194.765 55.105 ;
    RECT 195.63 55.035 195.84 55.105 ;
    RECT 197.44 55.21 198.255 55.28 ;
    RECT 199.245 54.765 199.515 54.835 ;
    RECT 199.245 55.12 199.515 55.19 ;
    RECT 199.245 55.485 199.515 55.555 ;
    RECT 174.56 54.045 174.63 54.835 ;
    RECT 175.16 54.045 175.37 54.115 ;
    RECT 175.16 54.4 175.37 54.47 ;
    RECT 175.16 54.765 175.37 54.835 ;
    RECT 176.325 54.49 177.125 54.56 ;
    RECT 178.79 54.315 179.025 54.385 ;
    RECT 179.85 54.315 180.11 54.385 ;
    RECT 181.825 54.315 182.055 54.385 ;
    RECT 182.54 54.315 182.8 54.385 ;
    RECT 183.71 54.315 183.78 54.385 ;
    RECT 187.045 54.315 187.255 54.385 ;
    RECT 187.43 54.315 187.7 54.385 ;
    RECT 191.485 54.315 191.555 54.385 ;
    RECT 191.815 54.315 192.08 54.385 ;
    RECT 193.57 54.315 193.83 54.385 ;
    RECT 194.015 54.315 194.085 54.385 ;
    RECT 194.505 54.315 194.765 54.385 ;
    RECT 195.63 54.315 195.84 54.385 ;
    RECT 197.44 54.49 198.255 54.56 ;
    RECT 199.245 54.045 199.515 54.115 ;
    RECT 199.245 54.4 199.515 54.47 ;
    RECT 199.245 54.765 199.515 54.835 ;
    RECT 198.605 48.645 198.815 48.715 ;
    RECT 174.56 53.325 174.63 54.115 ;
    RECT 175.16 53.325 175.37 53.395 ;
    RECT 175.16 53.68 175.37 53.75 ;
    RECT 175.16 54.045 175.37 54.115 ;
    RECT 176.325 53.77 177.125 53.84 ;
    RECT 178.79 53.595 179.025 53.665 ;
    RECT 179.85 53.595 180.11 53.665 ;
    RECT 181.825 53.595 182.055 53.665 ;
    RECT 182.54 53.595 182.8 53.665 ;
    RECT 183.71 53.595 183.78 53.665 ;
    RECT 187.045 53.595 187.255 53.665 ;
    RECT 187.43 53.595 187.7 53.665 ;
    RECT 191.485 53.595 191.555 53.665 ;
    RECT 191.815 53.595 192.08 53.665 ;
    RECT 193.57 53.595 193.83 53.665 ;
    RECT 194.015 53.595 194.085 53.665 ;
    RECT 194.505 53.595 194.765 53.665 ;
    RECT 195.63 53.595 195.84 53.665 ;
    RECT 197.44 53.77 198.255 53.84 ;
    RECT 199.245 53.325 199.515 53.395 ;
    RECT 199.245 53.68 199.515 53.75 ;
    RECT 199.245 54.045 199.515 54.115 ;
    RECT 174.56 52.605 174.63 53.395 ;
    RECT 175.16 52.605 175.37 52.675 ;
    RECT 175.16 52.96 175.37 53.03 ;
    RECT 175.16 53.325 175.37 53.395 ;
    RECT 176.325 53.05 177.125 53.12 ;
    RECT 178.79 52.875 179.025 52.945 ;
    RECT 179.85 52.875 180.11 52.945 ;
    RECT 181.825 52.875 182.055 52.945 ;
    RECT 182.54 52.875 182.8 52.945 ;
    RECT 183.71 52.875 183.78 52.945 ;
    RECT 187.045 52.875 187.255 52.945 ;
    RECT 187.43 52.875 187.7 52.945 ;
    RECT 191.485 52.875 191.555 52.945 ;
    RECT 191.815 52.875 192.08 52.945 ;
    RECT 193.57 52.875 193.83 52.945 ;
    RECT 194.015 52.875 194.085 52.945 ;
    RECT 194.505 52.875 194.765 52.945 ;
    RECT 195.63 52.875 195.84 52.945 ;
    RECT 197.44 53.05 198.255 53.12 ;
    RECT 199.245 52.605 199.515 52.675 ;
    RECT 199.245 52.96 199.515 53.03 ;
    RECT 199.245 53.325 199.515 53.395 ;
    RECT 174.56 51.885 174.63 52.675 ;
    RECT 175.16 51.885 175.37 51.955 ;
    RECT 175.16 52.24 175.37 52.31 ;
    RECT 175.16 52.605 175.37 52.675 ;
    RECT 176.325 52.33 177.125 52.4 ;
    RECT 178.79 52.155 179.025 52.225 ;
    RECT 179.85 52.155 180.11 52.225 ;
    RECT 181.825 52.155 182.055 52.225 ;
    RECT 182.54 52.155 182.8 52.225 ;
    RECT 183.71 52.155 183.78 52.225 ;
    RECT 187.045 52.155 187.255 52.225 ;
    RECT 187.43 52.155 187.7 52.225 ;
    RECT 191.485 52.155 191.555 52.225 ;
    RECT 191.815 52.155 192.08 52.225 ;
    RECT 193.57 52.155 193.83 52.225 ;
    RECT 194.015 52.155 194.085 52.225 ;
    RECT 194.505 52.155 194.765 52.225 ;
    RECT 195.63 52.155 195.84 52.225 ;
    RECT 197.44 52.33 198.255 52.4 ;
    RECT 199.245 51.885 199.515 51.955 ;
    RECT 199.245 52.24 199.515 52.31 ;
    RECT 199.245 52.605 199.515 52.675 ;
    RECT 174.56 51.165 174.63 51.955 ;
    RECT 175.16 51.165 175.37 51.235 ;
    RECT 175.16 51.52 175.37 51.59 ;
    RECT 175.16 51.885 175.37 51.955 ;
    RECT 176.325 51.61 177.125 51.68 ;
    RECT 178.79 51.435 179.025 51.505 ;
    RECT 179.85 51.435 180.11 51.505 ;
    RECT 181.825 51.435 182.055 51.505 ;
    RECT 182.54 51.435 182.8 51.505 ;
    RECT 183.71 51.435 183.78 51.505 ;
    RECT 187.045 51.435 187.255 51.505 ;
    RECT 187.43 51.435 187.7 51.505 ;
    RECT 191.485 51.435 191.555 51.505 ;
    RECT 191.815 51.435 192.08 51.505 ;
    RECT 193.57 51.435 193.83 51.505 ;
    RECT 194.015 51.435 194.085 51.505 ;
    RECT 194.505 51.435 194.765 51.505 ;
    RECT 195.63 51.435 195.84 51.505 ;
    RECT 197.44 51.61 198.255 51.68 ;
    RECT 199.245 51.165 199.515 51.235 ;
    RECT 199.245 51.52 199.515 51.59 ;
    RECT 199.245 51.885 199.515 51.955 ;
    RECT 174.56 50.445 174.63 51.235 ;
    RECT 175.16 50.445 175.37 50.515 ;
    RECT 175.16 50.8 175.37 50.87 ;
    RECT 175.16 51.165 175.37 51.235 ;
    RECT 176.325 50.89 177.125 50.96 ;
    RECT 178.79 50.715 179.025 50.785 ;
    RECT 179.85 50.715 180.11 50.785 ;
    RECT 181.825 50.715 182.055 50.785 ;
    RECT 182.54 50.715 182.8 50.785 ;
    RECT 183.71 50.715 183.78 50.785 ;
    RECT 187.045 50.715 187.255 50.785 ;
    RECT 187.43 50.715 187.7 50.785 ;
    RECT 191.485 50.715 191.555 50.785 ;
    RECT 191.815 50.715 192.08 50.785 ;
    RECT 193.57 50.715 193.83 50.785 ;
    RECT 194.015 50.715 194.085 50.785 ;
    RECT 194.505 50.715 194.765 50.785 ;
    RECT 195.63 50.715 195.84 50.785 ;
    RECT 197.44 50.89 198.255 50.96 ;
    RECT 199.245 50.445 199.515 50.515 ;
    RECT 199.245 50.8 199.515 50.87 ;
    RECT 199.245 51.165 199.515 51.235 ;
    RECT 174.56 49.725 174.63 50.515 ;
    RECT 175.16 49.725 175.37 49.795 ;
    RECT 175.16 50.08 175.37 50.15 ;
    RECT 175.16 50.445 175.37 50.515 ;
    RECT 176.325 50.17 177.125 50.24 ;
    RECT 178.79 49.995 179.025 50.065 ;
    RECT 179.85 49.995 180.11 50.065 ;
    RECT 181.825 49.995 182.055 50.065 ;
    RECT 182.54 49.995 182.8 50.065 ;
    RECT 183.71 49.995 183.78 50.065 ;
    RECT 187.045 49.995 187.255 50.065 ;
    RECT 187.43 49.995 187.7 50.065 ;
    RECT 191.485 49.995 191.555 50.065 ;
    RECT 191.815 49.995 192.08 50.065 ;
    RECT 193.57 49.995 193.83 50.065 ;
    RECT 194.015 49.995 194.085 50.065 ;
    RECT 194.505 49.995 194.765 50.065 ;
    RECT 195.63 49.995 195.84 50.065 ;
    RECT 197.44 50.17 198.255 50.24 ;
    RECT 199.245 49.725 199.515 49.795 ;
    RECT 199.245 50.08 199.515 50.15 ;
    RECT 199.245 50.445 199.515 50.515 ;
    RECT 174.56 49.005 174.63 49.795 ;
    RECT 175.16 49.005 175.37 49.075 ;
    RECT 175.16 49.36 175.37 49.43 ;
    RECT 175.16 49.725 175.37 49.795 ;
    RECT 176.325 49.45 177.125 49.52 ;
    RECT 178.79 49.275 179.025 49.345 ;
    RECT 179.85 49.275 180.11 49.345 ;
    RECT 181.825 49.275 182.055 49.345 ;
    RECT 182.54 49.275 182.8 49.345 ;
    RECT 183.71 49.275 183.78 49.345 ;
    RECT 187.045 49.275 187.255 49.345 ;
    RECT 187.43 49.275 187.7 49.345 ;
    RECT 191.485 49.275 191.555 49.345 ;
    RECT 191.815 49.275 192.08 49.345 ;
    RECT 193.57 49.275 193.83 49.345 ;
    RECT 194.015 49.275 194.085 49.345 ;
    RECT 194.505 49.275 194.765 49.345 ;
    RECT 195.63 49.275 195.84 49.345 ;
    RECT 197.44 49.45 198.255 49.52 ;
    RECT 199.245 49.005 199.515 49.075 ;
    RECT 199.245 49.36 199.515 49.43 ;
    RECT 199.245 49.725 199.515 49.795 ;
    RECT 186.51 34.872 186.58 34.942 ;
    RECT 180.81 50.712 181.02 50.782 ;
    RECT 174.56 58.385 174.63 59.175 ;
    RECT 175.16 58.385 175.37 58.455 ;
    RECT 175.16 58.74 175.37 58.81 ;
    RECT 175.16 59.105 175.37 59.175 ;
    RECT 176.325 58.83 177.125 58.9 ;
    RECT 178.79 58.655 179.025 58.725 ;
    RECT 179.85 58.655 180.11 58.725 ;
    RECT 181.825 58.655 182.055 58.725 ;
    RECT 182.54 58.655 182.8 58.725 ;
    RECT 183.71 58.655 183.78 58.725 ;
    RECT 187.045 58.655 187.255 58.725 ;
    RECT 187.43 58.655 187.7 58.725 ;
    RECT 191.485 58.655 191.555 58.725 ;
    RECT 191.815 58.655 192.08 58.725 ;
    RECT 193.57 58.655 193.83 58.725 ;
    RECT 194.015 58.655 194.085 58.725 ;
    RECT 194.505 58.655 194.765 58.725 ;
    RECT 195.63 58.655 195.84 58.725 ;
    RECT 197.44 58.83 198.255 58.9 ;
    RECT 199.245 58.385 199.515 58.455 ;
    RECT 199.245 58.74 199.515 58.81 ;
    RECT 199.245 59.105 199.515 59.175 ;
    RECT 175.75 50.805 175.96 50.875 ;
    RECT 175.75 23.445 175.96 23.515 ;
    RECT 188.225 40.632 188.295 40.702 ;
    RECT 175.75 22.725 175.96 22.795 ;
    RECT 192.85 48.555 193.06 48.625 ;
    RECT 175.75 22.005 175.96 22.075 ;
    RECT 180.81 48.552 181.02 48.622 ;
    RECT 174.56 48.285 174.63 49.075 ;
    RECT 175.16 48.285 175.37 48.355 ;
    RECT 175.16 48.64 175.37 48.71 ;
    RECT 175.16 49.005 175.37 49.075 ;
    RECT 176.325 48.73 177.125 48.8 ;
    RECT 178.79 48.555 179.025 48.625 ;
    RECT 179.85 48.555 180.11 48.625 ;
    RECT 181.825 48.555 182.055 48.625 ;
    RECT 182.54 48.555 182.8 48.625 ;
    RECT 183.71 48.555 183.78 48.625 ;
    RECT 187.045 48.555 187.255 48.625 ;
    RECT 187.43 48.555 187.7 48.625 ;
    RECT 191.485 48.555 191.555 48.625 ;
    RECT 191.815 48.555 192.08 48.625 ;
    RECT 193.57 48.555 193.83 48.625 ;
    RECT 194.015 48.555 194.085 48.625 ;
    RECT 194.505 48.555 194.765 48.625 ;
    RECT 195.63 48.555 195.84 48.625 ;
    RECT 197.44 48.73 198.255 48.8 ;
    RECT 199.245 48.285 199.515 48.355 ;
    RECT 199.245 48.64 199.515 48.71 ;
    RECT 199.245 49.005 199.515 49.075 ;
    RECT 174.56 47.565 174.63 48.355 ;
    RECT 175.16 47.565 175.37 47.635 ;
    RECT 175.16 47.92 175.37 47.99 ;
    RECT 175.16 48.285 175.37 48.355 ;
    RECT 176.325 48.01 177.125 48.08 ;
    RECT 178.79 47.835 179.025 47.905 ;
    RECT 179.85 47.835 180.11 47.905 ;
    RECT 181.825 47.835 182.055 47.905 ;
    RECT 182.54 47.835 182.8 47.905 ;
    RECT 183.71 47.835 183.78 47.905 ;
    RECT 187.045 47.835 187.255 47.905 ;
    RECT 187.43 47.835 187.7 47.905 ;
    RECT 191.485 47.835 191.555 47.905 ;
    RECT 191.815 47.835 192.08 47.905 ;
    RECT 193.57 47.835 193.83 47.905 ;
    RECT 194.015 47.835 194.085 47.905 ;
    RECT 194.505 47.835 194.765 47.905 ;
    RECT 195.63 47.835 195.84 47.905 ;
    RECT 197.44 48.01 198.255 48.08 ;
    RECT 199.245 47.565 199.515 47.635 ;
    RECT 199.245 47.92 199.515 47.99 ;
    RECT 199.245 48.285 199.515 48.355 ;
    RECT 174.56 46.845 174.63 47.635 ;
    RECT 175.16 46.845 175.37 46.915 ;
    RECT 175.16 47.2 175.37 47.27 ;
    RECT 175.16 47.565 175.37 47.635 ;
    RECT 176.325 47.29 177.125 47.36 ;
    RECT 178.79 47.115 179.025 47.185 ;
    RECT 179.85 47.115 180.11 47.185 ;
    RECT 181.825 47.115 182.055 47.185 ;
    RECT 182.54 47.115 182.8 47.185 ;
    RECT 183.71 47.115 183.78 47.185 ;
    RECT 187.045 47.115 187.255 47.185 ;
    RECT 187.43 47.115 187.7 47.185 ;
    RECT 191.485 47.115 191.555 47.185 ;
    RECT 191.815 47.115 192.08 47.185 ;
    RECT 193.57 47.115 193.83 47.185 ;
    RECT 194.015 47.115 194.085 47.185 ;
    RECT 194.505 47.115 194.765 47.185 ;
    RECT 195.63 47.115 195.84 47.185 ;
    RECT 197.44 47.29 198.255 47.36 ;
    RECT 199.245 46.845 199.515 46.915 ;
    RECT 199.245 47.2 199.515 47.27 ;
    RECT 199.245 47.565 199.515 47.635 ;
    RECT 175.75 48.645 175.96 48.715 ;
    RECT 174.56 46.125 174.63 46.915 ;
    RECT 175.16 46.125 175.37 46.195 ;
    RECT 175.16 46.48 175.37 46.55 ;
    RECT 175.16 46.845 175.37 46.915 ;
    RECT 176.325 46.57 177.125 46.64 ;
    RECT 178.79 46.395 179.025 46.465 ;
    RECT 179.85 46.395 180.11 46.465 ;
    RECT 181.825 46.395 182.055 46.465 ;
    RECT 182.54 46.395 182.8 46.465 ;
    RECT 183.71 46.395 183.78 46.465 ;
    RECT 187.045 46.395 187.255 46.465 ;
    RECT 187.43 46.395 187.7 46.465 ;
    RECT 191.485 46.395 191.555 46.465 ;
    RECT 191.815 46.395 192.08 46.465 ;
    RECT 193.57 46.395 193.83 46.465 ;
    RECT 194.015 46.395 194.085 46.465 ;
    RECT 194.505 46.395 194.765 46.465 ;
    RECT 195.63 46.395 195.84 46.465 ;
    RECT 197.44 46.57 198.255 46.64 ;
    RECT 199.245 46.125 199.515 46.195 ;
    RECT 199.245 46.48 199.515 46.55 ;
    RECT 199.245 46.845 199.515 46.915 ;
    RECT 198.605 50.085 198.815 50.155 ;
    RECT 174.56 45.405 174.63 46.195 ;
    RECT 175.16 45.405 175.37 45.475 ;
    RECT 175.16 45.76 175.37 45.83 ;
    RECT 175.16 46.125 175.37 46.195 ;
    RECT 176.325 45.85 177.125 45.92 ;
    RECT 178.79 45.675 179.025 45.745 ;
    RECT 179.85 45.675 180.11 45.745 ;
    RECT 181.825 45.675 182.055 45.745 ;
    RECT 182.54 45.675 182.8 45.745 ;
    RECT 183.71 45.675 183.78 45.745 ;
    RECT 187.045 45.675 187.255 45.745 ;
    RECT 187.43 45.675 187.7 45.745 ;
    RECT 191.485 45.675 191.555 45.745 ;
    RECT 191.815 45.675 192.08 45.745 ;
    RECT 193.57 45.675 193.83 45.745 ;
    RECT 194.015 45.675 194.085 45.745 ;
    RECT 194.505 45.675 194.765 45.745 ;
    RECT 195.63 45.675 195.84 45.745 ;
    RECT 197.44 45.85 198.255 45.92 ;
    RECT 199.245 45.405 199.515 45.475 ;
    RECT 199.245 45.76 199.515 45.83 ;
    RECT 199.245 46.125 199.515 46.195 ;
    RECT 174.56 44.685 174.63 45.475 ;
    RECT 175.16 44.685 175.37 44.755 ;
    RECT 175.16 45.04 175.37 45.11 ;
    RECT 175.16 45.405 175.37 45.475 ;
    RECT 176.325 45.13 177.125 45.2 ;
    RECT 178.79 44.955 179.025 45.025 ;
    RECT 179.85 44.955 180.11 45.025 ;
    RECT 181.825 44.955 182.055 45.025 ;
    RECT 182.54 44.955 182.8 45.025 ;
    RECT 183.71 44.955 183.78 45.025 ;
    RECT 187.045 44.955 187.255 45.025 ;
    RECT 187.43 44.955 187.7 45.025 ;
    RECT 191.485 44.955 191.555 45.025 ;
    RECT 191.815 44.955 192.08 45.025 ;
    RECT 193.57 44.955 193.83 45.025 ;
    RECT 194.015 44.955 194.085 45.025 ;
    RECT 194.505 44.955 194.765 45.025 ;
    RECT 195.63 44.955 195.84 45.025 ;
    RECT 197.44 45.13 198.255 45.2 ;
    RECT 199.245 44.685 199.515 44.755 ;
    RECT 199.245 45.04 199.515 45.11 ;
    RECT 199.245 45.405 199.515 45.475 ;
    RECT 192.85 49.995 193.06 50.065 ;
    RECT 174.56 43.965 174.63 44.755 ;
    RECT 175.16 43.965 175.37 44.035 ;
    RECT 175.16 44.32 175.37 44.39 ;
    RECT 175.16 44.685 175.37 44.755 ;
    RECT 176.325 44.41 177.125 44.48 ;
    RECT 178.79 44.235 179.025 44.305 ;
    RECT 179.85 44.235 180.11 44.305 ;
    RECT 181.825 44.235 182.055 44.305 ;
    RECT 182.54 44.235 182.8 44.305 ;
    RECT 183.71 44.235 183.78 44.305 ;
    RECT 187.045 44.235 187.255 44.305 ;
    RECT 187.43 44.235 187.7 44.305 ;
    RECT 191.485 44.235 191.555 44.305 ;
    RECT 191.815 44.235 192.08 44.305 ;
    RECT 193.57 44.235 193.83 44.305 ;
    RECT 194.015 44.235 194.085 44.305 ;
    RECT 194.505 44.235 194.765 44.305 ;
    RECT 195.63 44.235 195.84 44.305 ;
    RECT 197.44 44.41 198.255 44.48 ;
    RECT 199.245 43.965 199.515 44.035 ;
    RECT 199.245 44.32 199.515 44.39 ;
    RECT 199.245 44.685 199.515 44.755 ;
    RECT 174.56 43.245 174.63 44.035 ;
    RECT 175.16 43.245 175.37 43.315 ;
    RECT 175.16 43.6 175.37 43.67 ;
    RECT 175.16 43.965 175.37 44.035 ;
    RECT 176.325 43.69 177.125 43.76 ;
    RECT 178.79 43.515 179.025 43.585 ;
    RECT 179.85 43.515 180.11 43.585 ;
    RECT 181.825 43.515 182.055 43.585 ;
    RECT 182.54 43.515 182.8 43.585 ;
    RECT 183.71 43.515 183.78 43.585 ;
    RECT 187.045 43.515 187.255 43.585 ;
    RECT 187.43 43.515 187.7 43.585 ;
    RECT 191.485 43.515 191.555 43.585 ;
    RECT 191.815 43.515 192.08 43.585 ;
    RECT 193.57 43.515 193.83 43.585 ;
    RECT 194.015 43.515 194.085 43.585 ;
    RECT 194.505 43.515 194.765 43.585 ;
    RECT 195.63 43.515 195.84 43.585 ;
    RECT 197.44 43.69 198.255 43.76 ;
    RECT 199.245 43.245 199.515 43.315 ;
    RECT 199.245 43.6 199.515 43.67 ;
    RECT 199.245 43.965 199.515 44.035 ;
    RECT 174.56 42.525 174.63 43.315 ;
    RECT 175.16 42.525 175.37 42.595 ;
    RECT 175.16 42.88 175.37 42.95 ;
    RECT 175.16 43.245 175.37 43.315 ;
    RECT 176.325 42.97 177.125 43.04 ;
    RECT 178.79 42.795 179.025 42.865 ;
    RECT 179.85 42.795 180.11 42.865 ;
    RECT 181.825 42.795 182.055 42.865 ;
    RECT 182.54 42.795 182.8 42.865 ;
    RECT 183.71 42.795 183.78 42.865 ;
    RECT 187.045 42.795 187.255 42.865 ;
    RECT 187.43 42.795 187.7 42.865 ;
    RECT 191.485 42.795 191.555 42.865 ;
    RECT 191.815 42.795 192.08 42.865 ;
    RECT 193.57 42.795 193.83 42.865 ;
    RECT 194.015 42.795 194.085 42.865 ;
    RECT 194.505 42.795 194.765 42.865 ;
    RECT 195.63 42.795 195.84 42.865 ;
    RECT 197.44 42.97 198.255 43.04 ;
    RECT 199.245 42.525 199.515 42.595 ;
    RECT 199.245 42.88 199.515 42.95 ;
    RECT 199.245 43.245 199.515 43.315 ;
    RECT 174.56 41.805 174.63 42.595 ;
    RECT 175.16 41.805 175.37 41.875 ;
    RECT 175.16 42.16 175.37 42.23 ;
    RECT 175.16 42.525 175.37 42.595 ;
    RECT 176.325 42.25 177.125 42.32 ;
    RECT 178.79 42.075 179.025 42.145 ;
    RECT 179.85 42.075 180.11 42.145 ;
    RECT 181.825 42.075 182.055 42.145 ;
    RECT 182.54 42.075 182.8 42.145 ;
    RECT 183.71 42.075 183.78 42.145 ;
    RECT 187.045 42.075 187.255 42.145 ;
    RECT 187.43 42.075 187.7 42.145 ;
    RECT 191.485 42.075 191.555 42.145 ;
    RECT 191.815 42.075 192.08 42.145 ;
    RECT 193.57 42.075 193.83 42.145 ;
    RECT 194.015 42.075 194.085 42.145 ;
    RECT 194.505 42.075 194.765 42.145 ;
    RECT 195.63 42.075 195.84 42.145 ;
    RECT 197.44 42.25 198.255 42.32 ;
    RECT 199.245 41.805 199.515 41.875 ;
    RECT 199.245 42.16 199.515 42.23 ;
    RECT 199.245 42.525 199.515 42.595 ;
    RECT 188.225 39.912 188.295 39.982 ;
    RECT 198.605 47.925 198.815 47.995 ;
    RECT 175.75 21.285 175.96 21.355 ;
    RECT 175.75 20.565 175.96 20.635 ;
    RECT 180.81 49.992 181.02 50.062 ;
    RECT 175.75 50.085 175.96 50.155 ;
    RECT 185.115 57.192 185.185 57.262 ;
    RECT 198.605 49.365 198.815 49.435 ;
    RECT 185.315 54.312 185.385 54.382 ;
    RECT 192.85 49.275 193.06 49.345 ;
    RECT 188.225 39.192 188.295 39.262 ;
    RECT 193.595 13.27 193.805 13.34 ;
    RECT 185.115 56.472 185.185 56.542 ;
    RECT 180.81 49.272 181.02 49.342 ;
    RECT 175.75 49.365 175.96 49.435 ;
    RECT 185.315 53.592 185.385 53.662 ;
    RECT 192.85 26.945 193.06 27.015 ;
    RECT 192.85 26.225 193.06 26.295 ;
    RECT 188.225 38.472 188.295 38.542 ;
    RECT 192.85 24.065 193.06 24.135 ;
    RECT 191.02 19.752 191.23 19.822 ;
    RECT 191.02 18.312 191.23 18.382 ;
    RECT 191.02 16.872 191.23 16.942 ;
    RECT 191.02 11.84 191.23 11.91 ;
    RECT 185.315 52.872 185.385 52.942 ;
    RECT 188.225 37.752 188.295 37.822 ;
    RECT 185.715 46.392 185.785 46.462 ;
    RECT 188.225 37.032 188.295 37.102 ;
    RECT 185.315 52.152 185.385 52.222 ;
    RECT 185.91 45.672 185.98 45.742 ;
    RECT 185.515 51.432 185.585 51.502 ;
    RECT 188.225 36.312 188.295 36.382 ;
    RECT 185.91 44.952 185.98 45.022 ;
    RECT 190.122 24.792 190.192 24.862 ;
    RECT 190.04 26.945 190.25 27.015 ;
    RECT 190.04 26.225 190.25 26.295 ;
    RECT 190.04 25.512 190.25 25.582 ;
    RECT 190.04 24.065 190.25 24.135 ;
    RECT 188.225 35.592 188.295 35.662 ;
    RECT 198.605 55.845 198.815 55.915 ;
    RECT 185.515 50.712 185.585 50.782 ;
    RECT 187.46 26.945 187.67 27.015 ;
    RECT 199.28 58.145 199.49 58.215 ;
    RECT 187.46 26.225 187.67 26.295 ;
    RECT 187.46 24.065 187.67 24.135 ;
    RECT 184.915 26.945 184.985 27.015 ;
    RECT 184.915 26.225 184.985 26.295 ;
    RECT 185.91 44.232 185.98 44.302 ;
    RECT 184.915 24.065 184.985 24.135 ;
    RECT 192.85 55.755 193.06 55.825 ;
    RECT 180.81 55.752 181.02 55.822 ;
    RECT 175.75 55.845 175.96 55.915 ;
    RECT 174.56 57.645 174.63 57.715 ;
    RECT 174.56 58.385 174.63 58.455 ;
    RECT 175.16 57.645 175.37 57.715 ;
    RECT 175.16 58.385 175.37 58.455 ;
    RECT 177.345 57.905 177.615 57.975 ;
    RECT 178.31 57.905 178.38 57.975 ;
    RECT 178.765 57.725 179.025 57.795 ;
    RECT 179.85 57.905 180.115 57.975 ;
    RECT 183.71 58.27 183.78 58.34 ;
    RECT 187.425 57.905 187.685 57.975 ;
    RECT 190.04 57.91 190.25 57.98 ;
    RECT 192.82 57.905 193.09 57.975 ;
    RECT 194.015 58.27 194.085 58.34 ;
    RECT 194.505 57.905 194.755 57.975 ;
    RECT 195.63 57.725 195.84 57.795 ;
    RECT 196.185 57.905 196.255 57.975 ;
    RECT 196.78 57.905 197.05 57.975 ;
    RECT 199.245 57.645 199.515 57.715 ;
    RECT 199.245 58.385 199.515 58.455 ;
    RECT 196.81 58.272 197.02 58.342 ;
    RECT 196.185 58.272 196.255 58.342 ;
    RECT 194.535 58.272 194.745 58.342 ;
    RECT 194.015 57.907 194.085 57.977 ;
    RECT 184.12 34.152 184.33 34.222 ;
    RECT 184.12 14.697 184.33 14.767 ;
    RECT 192.85 58.272 193.06 58.342 ;
    RECT 190.04 58.272 190.25 58.342 ;
    RECT 183.085 34.152 183.295 34.222 ;
    RECT 198.605 55.125 198.815 55.195 ;
    RECT 183.085 14.697 183.295 14.767 ;
    RECT 181.455 26.945 181.665 27.015 ;
    RECT 181.455 26.225 181.665 26.295 ;
    RECT 181.455 24.065 181.665 24.135 ;
    RECT 185.515 49.992 185.585 50.062 ;
    RECT 174.56 41.085 174.63 41.875 ;
    RECT 175.16 41.085 175.37 41.155 ;
    RECT 175.16 41.44 175.37 41.51 ;
    RECT 175.16 41.805 175.37 41.875 ;
    RECT 176.325 41.53 177.125 41.6 ;
    RECT 178.79 41.355 179.025 41.425 ;
    RECT 179.85 41.355 180.11 41.425 ;
    RECT 181.825 41.355 182.055 41.425 ;
    RECT 182.54 41.355 182.8 41.425 ;
    RECT 183.71 41.355 183.78 41.425 ;
    RECT 187.045 41.355 187.255 41.425 ;
    RECT 187.43 41.355 187.7 41.425 ;
    RECT 191.485 41.355 191.555 41.425 ;
    RECT 191.815 41.355 192.08 41.425 ;
    RECT 193.57 41.355 193.83 41.425 ;
    RECT 194.015 41.355 194.085 41.425 ;
    RECT 194.505 41.355 194.765 41.425 ;
    RECT 195.63 41.355 195.84 41.425 ;
    RECT 197.44 41.53 198.255 41.6 ;
    RECT 199.245 41.085 199.515 41.155 ;
    RECT 199.245 41.44 199.515 41.51 ;
    RECT 199.245 41.805 199.515 41.875 ;
    RECT 174.56 40.365 174.63 41.155 ;
    RECT 175.16 40.365 175.37 40.435 ;
    RECT 175.16 40.72 175.37 40.79 ;
    RECT 175.16 41.085 175.37 41.155 ;
    RECT 176.325 40.81 177.125 40.88 ;
    RECT 178.79 40.635 179.025 40.705 ;
    RECT 179.85 40.635 180.11 40.705 ;
    RECT 181.825 40.635 182.055 40.705 ;
    RECT 182.54 40.635 182.8 40.705 ;
    RECT 183.71 40.635 183.78 40.705 ;
    RECT 187.045 40.635 187.255 40.705 ;
    RECT 187.43 40.635 187.7 40.705 ;
    RECT 191.485 40.635 191.555 40.705 ;
    RECT 191.815 40.635 192.08 40.705 ;
    RECT 193.57 40.635 193.83 40.705 ;
    RECT 194.015 40.635 194.085 40.705 ;
    RECT 194.505 40.635 194.765 40.705 ;
    RECT 195.63 40.635 195.84 40.705 ;
    RECT 197.44 40.81 198.255 40.88 ;
    RECT 199.245 40.365 199.515 40.435 ;
    RECT 199.245 40.72 199.515 40.79 ;
    RECT 199.245 41.085 199.515 41.155 ;
    RECT 174.56 39.645 174.63 40.435 ;
    RECT 175.16 39.645 175.37 39.715 ;
    RECT 175.16 40.0 175.37 40.07 ;
    RECT 175.16 40.365 175.37 40.435 ;
    RECT 176.325 40.09 177.125 40.16 ;
    RECT 178.79 39.915 179.025 39.985 ;
    RECT 179.85 39.915 180.11 39.985 ;
    RECT 181.825 39.915 182.055 39.985 ;
    RECT 182.54 39.915 182.8 39.985 ;
    RECT 183.71 39.915 183.78 39.985 ;
    RECT 187.045 39.915 187.255 39.985 ;
    RECT 187.43 39.915 187.7 39.985 ;
    RECT 191.485 39.915 191.555 39.985 ;
    RECT 191.815 39.915 192.08 39.985 ;
    RECT 193.57 39.915 193.83 39.985 ;
    RECT 194.015 39.915 194.085 39.985 ;
    RECT 194.505 39.915 194.765 39.985 ;
    RECT 195.63 39.915 195.84 39.985 ;
    RECT 197.44 40.09 198.255 40.16 ;
    RECT 199.245 39.645 199.515 39.715 ;
    RECT 199.245 40.0 199.515 40.07 ;
    RECT 199.245 40.365 199.515 40.435 ;
    RECT 174.56 38.925 174.63 39.715 ;
    RECT 175.16 38.925 175.37 38.995 ;
    RECT 175.16 39.28 175.37 39.35 ;
    RECT 175.16 39.645 175.37 39.715 ;
    RECT 176.325 39.37 177.125 39.44 ;
    RECT 178.79 39.195 179.025 39.265 ;
    RECT 179.85 39.195 180.11 39.265 ;
    RECT 181.825 39.195 182.055 39.265 ;
    RECT 182.54 39.195 182.8 39.265 ;
    RECT 183.71 39.195 183.78 39.265 ;
    RECT 187.045 39.195 187.255 39.265 ;
    RECT 187.43 39.195 187.7 39.265 ;
    RECT 191.485 39.195 191.555 39.265 ;
    RECT 191.815 39.195 192.08 39.265 ;
    RECT 193.57 39.195 193.83 39.265 ;
    RECT 194.015 39.195 194.085 39.265 ;
    RECT 194.505 39.195 194.765 39.265 ;
    RECT 195.63 39.195 195.84 39.265 ;
    RECT 197.44 39.37 198.255 39.44 ;
    RECT 199.245 38.925 199.515 38.995 ;
    RECT 199.245 39.28 199.515 39.35 ;
    RECT 199.245 39.645 199.515 39.715 ;
    RECT 174.56 38.205 174.63 38.995 ;
    RECT 175.16 38.205 175.37 38.275 ;
    RECT 175.16 38.56 175.37 38.63 ;
    RECT 175.16 38.925 175.37 38.995 ;
    RECT 176.325 38.65 177.125 38.72 ;
    RECT 178.79 38.475 179.025 38.545 ;
    RECT 179.85 38.475 180.11 38.545 ;
    RECT 181.825 38.475 182.055 38.545 ;
    RECT 182.54 38.475 182.8 38.545 ;
    RECT 183.71 38.475 183.78 38.545 ;
    RECT 187.045 38.475 187.255 38.545 ;
    RECT 187.43 38.475 187.7 38.545 ;
    RECT 191.485 38.475 191.555 38.545 ;
    RECT 191.815 38.475 192.08 38.545 ;
    RECT 193.57 38.475 193.83 38.545 ;
    RECT 194.015 38.475 194.085 38.545 ;
    RECT 194.505 38.475 194.765 38.545 ;
    RECT 195.63 38.475 195.84 38.545 ;
    RECT 197.44 38.65 198.255 38.72 ;
    RECT 199.245 38.205 199.515 38.275 ;
    RECT 199.245 38.56 199.515 38.63 ;
    RECT 199.245 38.925 199.515 38.995 ;
    RECT 174.56 37.485 174.63 38.275 ;
    RECT 175.16 37.485 175.37 37.555 ;
    RECT 175.16 37.84 175.37 37.91 ;
    RECT 175.16 38.205 175.37 38.275 ;
    RECT 176.325 37.93 177.125 38.0 ;
    RECT 178.79 37.755 179.025 37.825 ;
    RECT 179.85 37.755 180.11 37.825 ;
    RECT 181.825 37.755 182.055 37.825 ;
    RECT 182.54 37.755 182.8 37.825 ;
    RECT 183.71 37.755 183.78 37.825 ;
    RECT 187.045 37.755 187.255 37.825 ;
    RECT 187.43 37.755 187.7 37.825 ;
    RECT 191.485 37.755 191.555 37.825 ;
    RECT 191.815 37.755 192.08 37.825 ;
    RECT 193.57 37.755 193.83 37.825 ;
    RECT 194.015 37.755 194.085 37.825 ;
    RECT 194.505 37.755 194.765 37.825 ;
    RECT 195.63 37.755 195.84 37.825 ;
    RECT 197.44 37.93 198.255 38.0 ;
    RECT 199.245 37.485 199.515 37.555 ;
    RECT 199.245 37.84 199.515 37.91 ;
    RECT 199.245 38.205 199.515 38.275 ;
    RECT 185.91 43.512 185.98 43.582 ;
    RECT 174.56 36.765 174.63 37.555 ;
    RECT 175.16 36.765 175.37 36.835 ;
    RECT 175.16 37.12 175.37 37.19 ;
    RECT 175.16 37.485 175.37 37.555 ;
    RECT 176.325 37.21 177.125 37.28 ;
    RECT 178.79 37.035 179.025 37.105 ;
    RECT 179.85 37.035 180.11 37.105 ;
    RECT 181.825 37.035 182.055 37.105 ;
    RECT 182.54 37.035 182.8 37.105 ;
    RECT 183.71 37.035 183.78 37.105 ;
    RECT 187.045 37.035 187.255 37.105 ;
    RECT 187.43 37.035 187.7 37.105 ;
    RECT 191.485 37.035 191.555 37.105 ;
    RECT 191.815 37.035 192.08 37.105 ;
    RECT 193.57 37.035 193.83 37.105 ;
    RECT 194.015 37.035 194.085 37.105 ;
    RECT 194.505 37.035 194.765 37.105 ;
    RECT 195.63 37.035 195.84 37.105 ;
    RECT 197.44 37.21 198.255 37.28 ;
    RECT 199.245 36.765 199.515 36.835 ;
    RECT 199.245 37.12 199.515 37.19 ;
    RECT 199.245 37.485 199.515 37.555 ;
    RECT 174.56 36.045 174.63 36.835 ;
    RECT 175.16 36.045 175.37 36.115 ;
    RECT 175.16 36.4 175.37 36.47 ;
    RECT 175.16 36.765 175.37 36.835 ;
    RECT 176.325 36.49 177.125 36.56 ;
    RECT 178.79 36.315 179.025 36.385 ;
    RECT 179.85 36.315 180.11 36.385 ;
    RECT 181.825 36.315 182.055 36.385 ;
    RECT 182.54 36.315 182.8 36.385 ;
    RECT 183.71 36.315 183.78 36.385 ;
    RECT 187.045 36.315 187.255 36.385 ;
    RECT 187.43 36.315 187.7 36.385 ;
    RECT 191.485 36.315 191.555 36.385 ;
    RECT 191.815 36.315 192.08 36.385 ;
    RECT 193.57 36.315 193.83 36.385 ;
    RECT 194.015 36.315 194.085 36.385 ;
    RECT 194.505 36.315 194.765 36.385 ;
    RECT 195.63 36.315 195.84 36.385 ;
    RECT 197.44 36.49 198.255 36.56 ;
    RECT 199.245 36.045 199.515 36.115 ;
    RECT 199.245 36.4 199.515 36.47 ;
    RECT 199.245 36.765 199.515 36.835 ;
    RECT 174.56 35.325 174.63 36.115 ;
    RECT 175.16 35.325 175.37 35.395 ;
    RECT 175.16 35.68 175.37 35.75 ;
    RECT 175.16 36.045 175.37 36.115 ;
    RECT 176.325 35.77 177.125 35.84 ;
    RECT 178.79 35.595 179.025 35.665 ;
    RECT 179.85 35.595 180.11 35.665 ;
    RECT 181.825 35.595 182.055 35.665 ;
    RECT 182.54 35.595 182.8 35.665 ;
    RECT 183.71 35.595 183.78 35.665 ;
    RECT 187.045 35.595 187.255 35.665 ;
    RECT 187.43 35.595 187.7 35.665 ;
    RECT 191.485 35.595 191.555 35.665 ;
    RECT 191.815 35.595 192.08 35.665 ;
    RECT 193.57 35.595 193.83 35.665 ;
    RECT 194.015 35.595 194.085 35.665 ;
    RECT 194.505 35.595 194.765 35.665 ;
    RECT 195.63 35.595 195.84 35.665 ;
    RECT 197.44 35.77 198.255 35.84 ;
    RECT 199.245 35.325 199.515 35.395 ;
    RECT 199.245 35.68 199.515 35.75 ;
    RECT 199.245 36.045 199.515 36.115 ;
    RECT 174.56 34.605 174.63 35.395 ;
    RECT 175.16 34.605 175.37 34.675 ;
    RECT 175.16 34.96 175.37 35.03 ;
    RECT 175.16 35.325 175.37 35.395 ;
    RECT 176.325 35.05 177.125 35.12 ;
    RECT 178.79 34.875 179.025 34.945 ;
    RECT 179.85 34.875 180.11 34.945 ;
    RECT 181.825 34.875 182.055 34.945 ;
    RECT 182.54 34.875 182.8 34.945 ;
    RECT 183.71 34.875 183.78 34.945 ;
    RECT 187.045 34.875 187.255 34.945 ;
    RECT 187.43 34.875 187.7 34.945 ;
    RECT 191.485 34.875 191.555 34.945 ;
    RECT 191.815 34.875 192.08 34.945 ;
    RECT 193.57 34.875 193.83 34.945 ;
    RECT 194.015 34.875 194.085 34.945 ;
    RECT 194.505 34.875 194.765 34.945 ;
    RECT 195.63 34.875 195.84 34.945 ;
    RECT 197.44 35.05 198.255 35.12 ;
    RECT 199.245 34.605 199.515 34.675 ;
    RECT 199.245 34.96 199.515 35.03 ;
    RECT 199.245 35.325 199.515 35.395 ;
    RECT 192.85 55.035 193.06 55.105 ;
    RECT 187.46 58.272 187.67 58.342 ;
    RECT 183.715 57.907 183.785 57.977 ;
    RECT 180.81 55.032 181.02 55.102 ;
    RECT 185.515 49.272 185.585 49.342 ;
    RECT 179.88 58.272 180.09 58.342 ;
    RECT 178.23 58.272 178.44 58.342 ;
    RECT 177.375 58.272 177.585 58.342 ;
    RECT 175.75 55.125 175.96 55.195 ;
    RECT 186.11 42.792 186.18 42.862 ;
    RECT 174.56 58.145 174.63 58.215 ;
    RECT 186.11 42.072 186.18 42.142 ;
    RECT 180.81 34.872 181.02 34.942 ;
    RECT 175.75 34.965 175.96 35.035 ;
    RECT 198.605 57.722 198.815 57.792 ;
    RECT 193.595 57.907 193.805 57.977 ;
    RECT 191.02 57.907 191.23 57.977 ;
    RECT 184.915 57.907 184.985 57.977 ;
    RECT 184.12 57.907 184.33 57.977 ;
    RECT 183.085 57.907 183.295 57.977 ;
    RECT 180.81 57.907 181.02 57.977 ;
    RECT 188.225 56.472 188.295 56.542 ;
    RECT 185.115 55.752 185.185 55.822 ;
    RECT 175.75 57.722 175.96 57.792 ;
    RECT 198.605 34.245 198.815 34.315 ;
    RECT 198.605 33.525 198.815 33.595 ;
    RECT 198.605 32.805 198.815 32.875 ;
    RECT 198.605 32.085 198.815 32.155 ;
    RECT 198.605 31.365 198.815 31.435 ;
    RECT 198.605 30.645 198.815 30.715 ;
    RECT 198.605 29.925 198.815 29.995 ;
    RECT 198.605 29.205 198.815 29.275 ;
    RECT 198.605 28.485 198.815 28.555 ;
    RECT 198.045 57.722 198.255 57.792 ;
    RECT 198.605 27.765 198.815 27.835 ;
    RECT 185.115 55.032 185.185 55.102 ;
    RECT 198.605 27.045 198.815 27.115 ;
    RECT 198.605 26.325 198.815 26.395 ;
    RECT 198.605 25.605 198.815 25.675 ;
    RECT 198.605 24.885 198.815 24.955 ;
    RECT 198.605 24.165 198.815 24.235 ;
    RECT 198.605 23.445 198.815 23.515 ;
    RECT 198.605 22.725 198.815 22.795 ;
    RECT 198.605 22.005 198.815 22.075 ;
    RECT 188.225 45.672 188.295 45.742 ;
    RECT 198.605 21.285 198.815 21.355 ;
    RECT 198.605 20.565 198.815 20.635 ;
    RECT 198.605 19.845 198.815 19.915 ;
    RECT 188.225 44.952 188.295 45.022 ;
    RECT 192.85 41.355 193.06 41.425 ;
    RECT 198.605 19.125 198.815 19.195 ;
    RECT 180.81 41.352 181.02 41.422 ;
    RECT 198.605 18.405 198.815 18.475 ;
    RECT 198.605 17.685 198.815 17.755 ;
    RECT 198.605 16.965 198.815 17.035 ;
    RECT 198.605 16.245 198.815 16.315 ;
    RECT 175.75 41.445 175.96 41.515 ;
    RECT 198.605 15.525 198.815 15.595 ;
    RECT 198.605 14.805 198.815 14.875 ;
    RECT 198.605 14.085 198.815 14.155 ;
    RECT 198.605 13.365 198.815 13.435 ;
    RECT 198.605 12.645 198.815 12.715 ;
    RECT 188.225 50.712 188.295 50.782 ;
    RECT 186.11 41.352 186.18 41.422 ;
    RECT 188.225 44.232 188.295 44.302 ;
    RECT 198.605 40.725 198.815 40.795 ;
    RECT 198.605 11.925 198.815 11.995 ;
    RECT 186.11 40.632 186.18 40.702 ;
    RECT 192.85 40.635 193.06 40.705 ;
    RECT 180.81 40.632 181.02 40.702 ;
    RECT 188.225 49.992 188.295 50.062 ;
    RECT 175.75 40.725 175.96 40.795 ;
    RECT 188.225 43.512 188.295 43.582 ;
    RECT 186.51 58.652 186.58 58.722 ;
    RECT 186.31 39.912 186.38 39.982 ;
    RECT 188.225 34.872 188.295 34.942 ;
    RECT 176.355 57.722 176.565 57.792 ;
    RECT 198.605 40.005 198.815 40.075 ;
    RECT 174.56 11.565 174.63 34.675 ;
    RECT 175.16 11.565 175.37 11.99 ;
    RECT 175.16 12.285 175.37 12.355 ;
    RECT 175.16 12.645 175.37 12.715 ;
    RECT 175.16 13.005 175.37 13.075 ;
    RECT 175.16 13.365 175.37 13.435 ;
    RECT 175.16 13.725 175.37 13.795 ;
    RECT 175.16 14.085 175.37 14.155 ;
    RECT 175.16 14.445 175.37 14.515 ;
    RECT 175.16 14.805 175.37 14.875 ;
    RECT 175.16 15.165 175.37 15.235 ;
    RECT 175.16 15.525 175.37 15.595 ;
    RECT 175.16 15.885 175.37 15.955 ;
    RECT 175.16 16.245 175.37 16.315 ;
    RECT 175.16 16.605 175.37 16.675 ;
    RECT 175.16 16.965 175.37 17.035 ;
    RECT 175.16 17.325 175.37 17.395 ;
    RECT 175.16 17.685 175.37 17.755 ;
    RECT 175.16 18.045 175.37 18.115 ;
    RECT 175.16 18.405 175.37 18.475 ;
    RECT 175.16 18.765 175.37 18.835 ;
    RECT 175.16 19.125 175.37 19.195 ;
    RECT 175.16 19.485 175.37 19.555 ;
    RECT 175.16 19.845 175.37 19.915 ;
    RECT 175.16 20.205 175.37 20.275 ;
    RECT 175.16 20.565 175.37 20.635 ;
    RECT 175.16 20.925 175.37 20.995 ;
    RECT 175.16 21.285 175.37 21.355 ;
    RECT 175.16 21.645 175.37 21.715 ;
    RECT 175.16 22.005 175.37 22.075 ;
    RECT 175.16 22.365 175.37 22.435 ;
    RECT 175.16 22.725 175.37 22.795 ;
    RECT 175.16 23.085 175.37 23.155 ;
    RECT 175.16 23.445 175.37 23.515 ;
    RECT 175.16 23.805 175.37 23.875 ;
    RECT 175.16 24.165 175.37 24.235 ;
    RECT 175.16 24.525 175.37 24.595 ;
    RECT 175.16 24.885 175.37 24.955 ;
    RECT 175.16 25.245 175.37 25.315 ;
    RECT 175.16 25.605 175.37 25.675 ;
    RECT 175.16 25.965 175.37 26.035 ;
    RECT 175.16 26.325 175.37 26.395 ;
    RECT 175.16 26.685 175.37 26.755 ;
    RECT 175.16 27.045 175.37 27.115 ;
    RECT 175.16 27.405 175.37 27.475 ;
    RECT 175.16 27.765 175.37 27.835 ;
    RECT 175.16 28.125 175.37 28.195 ;
    RECT 175.16 28.485 175.37 28.555 ;
    RECT 175.16 28.845 175.37 28.915 ;
    RECT 175.16 29.205 175.37 29.275 ;
    RECT 175.16 29.565 175.37 29.635 ;
    RECT 175.16 29.925 175.37 29.995 ;
    RECT 175.16 30.285 175.37 30.355 ;
    RECT 175.16 30.645 175.37 30.715 ;
    RECT 175.16 31.005 175.37 31.075 ;
    RECT 175.16 31.365 175.37 31.435 ;
    RECT 175.16 31.725 175.37 31.795 ;
    RECT 175.16 32.085 175.37 32.155 ;
    RECT 175.16 32.445 175.37 32.515 ;
    RECT 175.16 32.805 175.37 32.875 ;
    RECT 175.16 33.165 175.37 33.235 ;
    RECT 175.16 33.525 175.37 33.595 ;
    RECT 175.16 33.885 175.37 33.955 ;
    RECT 175.16 34.245 175.37 34.315 ;
    RECT 175.16 34.605 175.37 34.675 ;
    RECT 176.355 12.01 177.095 12.08 ;
    RECT 176.355 12.73 177.095 12.8 ;
    RECT 176.355 13.445 177.095 13.515 ;
    RECT 176.355 14.17 177.095 14.24 ;
    RECT 176.355 14.89 177.095 14.96 ;
    RECT 176.355 15.61 177.095 15.68 ;
    RECT 176.355 16.325 177.095 16.395 ;
    RECT 176.355 17.05 177.095 17.12 ;
    RECT 176.355 17.77 177.095 17.84 ;
    RECT 176.355 18.485 177.095 18.555 ;
    RECT 176.355 19.21 177.095 19.28 ;
    RECT 176.355 19.93 177.095 20.0 ;
    RECT 176.355 20.65 177.095 20.72 ;
    RECT 176.355 21.37 177.095 21.44 ;
    RECT 176.355 22.09 177.095 22.16 ;
    RECT 176.355 22.81 177.095 22.88 ;
    RECT 176.355 23.53 177.095 23.6 ;
    RECT 176.355 24.25 177.095 24.32 ;
    RECT 176.355 24.97 177.095 25.04 ;
    RECT 176.355 25.69 177.095 25.76 ;
    RECT 176.355 26.41 177.095 26.48 ;
    RECT 176.355 27.13 177.095 27.2 ;
    RECT 176.355 27.845 177.095 27.915 ;
    RECT 176.355 28.565 177.095 28.635 ;
    RECT 176.355 29.29 177.095 29.36 ;
    RECT 176.355 30.01 177.095 30.08 ;
    RECT 176.355 30.73 177.095 30.8 ;
    RECT 176.355 31.45 177.095 31.52 ;
    RECT 176.355 32.17 177.095 32.24 ;
    RECT 176.355 32.885 177.095 32.955 ;
    RECT 176.355 33.605 177.095 33.675 ;
    RECT 176.355 34.33 177.095 34.4 ;
    RECT 178.8 34.15 179.01 34.22 ;
    RECT 178.815 11.835 179.025 11.905 ;
    RECT 178.815 12.55 179.025 12.62 ;
    RECT 178.815 13.265 179.025 13.335 ;
    RECT 178.815 13.98 179.025 14.05 ;
    RECT 178.815 14.695 179.025 14.765 ;
    RECT 178.815 15.435 179.025 15.505 ;
    RECT 178.815 16.15 179.025 16.22 ;
    RECT 178.815 16.87 179.025 16.94 ;
    RECT 178.815 17.59 179.025 17.66 ;
    RECT 178.815 18.31 179.025 18.38 ;
    RECT 178.815 19.03 179.025 19.1 ;
    RECT 178.815 19.75 179.025 19.82 ;
    RECT 178.815 22.63 179.025 22.7 ;
    RECT 178.815 23.35 179.025 23.42 ;
    RECT 178.815 24.79 179.025 24.86 ;
    RECT 178.815 26.235 179.025 26.305 ;
    RECT 178.815 26.955 179.025 27.025 ;
    RECT 178.815 27.675 179.025 27.745 ;
    RECT 178.815 28.39 179.025 28.46 ;
    RECT 178.815 29.11 179.025 29.18 ;
    RECT 178.815 29.83 179.025 29.9 ;
    RECT 178.815 30.55 179.025 30.62 ;
    RECT 178.815 31.275 179.025 31.345 ;
    RECT 178.815 31.995 179.025 32.065 ;
    RECT 178.815 32.715 179.025 32.785 ;
    RECT 178.815 33.43 179.025 33.5 ;
    RECT 179.85 11.835 180.11 11.905 ;
    RECT 179.85 12.55 180.11 12.62 ;
    RECT 179.85 13.265 180.11 13.335 ;
    RECT 179.85 15.435 180.11 15.505 ;
    RECT 179.85 16.15 180.11 16.22 ;
    RECT 179.85 16.87 180.11 16.94 ;
    RECT 179.85 17.59 180.11 17.66 ;
    RECT 179.85 19.75 180.11 19.82 ;
    RECT 179.85 23.35 180.11 23.42 ;
    RECT 179.85 26.235 180.11 26.305 ;
    RECT 179.85 26.955 180.11 27.025 ;
    RECT 179.85 27.675 180.11 27.745 ;
    RECT 179.85 29.83 180.11 29.9 ;
    RECT 179.85 30.55 180.11 30.62 ;
    RECT 179.85 31.275 180.11 31.345 ;
    RECT 179.85 31.995 180.11 32.065 ;
    RECT 179.85 32.715 180.11 32.785 ;
    RECT 179.85 33.43 180.11 33.5 ;
    RECT 179.88 13.985 180.09 14.055 ;
    RECT 179.88 14.7 180.09 14.77 ;
    RECT 179.88 18.315 180.09 18.385 ;
    RECT 179.88 19.03 180.09 19.1 ;
    RECT 179.88 29.12 180.09 29.19 ;
    RECT 179.88 34.155 180.09 34.225 ;
    RECT 180.79 11.835 181.04 11.905 ;
    RECT 180.79 12.55 181.04 12.62 ;
    RECT 180.79 13.265 181.04 13.335 ;
    RECT 180.79 16.15 181.04 16.22 ;
    RECT 180.79 16.87 181.04 16.94 ;
    RECT 180.79 17.59 181.04 17.66 ;
    RECT 180.79 19.75 181.04 19.82 ;
    RECT 180.79 20.47 181.04 20.54 ;
    RECT 180.79 21.915 181.04 21.985 ;
    RECT 180.79 29.83 181.01 29.9 ;
    RECT 180.795 23.35 181.04 23.42 ;
    RECT 180.795 27.675 181.015 27.745 ;
    RECT 180.8 30.55 181.02 30.62 ;
    RECT 180.8 31.275 181.02 31.345 ;
    RECT 180.8 31.995 181.02 32.065 ;
    RECT 180.805 25.51 181.04 25.58 ;
    RECT 180.805 33.43 181.04 33.5 ;
    RECT 180.81 24.065 181.02 24.135 ;
    RECT 180.81 26.225 181.02 26.295 ;
    RECT 180.81 26.945 181.02 27.015 ;
    RECT 180.81 32.715 181.03 32.785 ;
    RECT 181.245 13.265 181.315 13.335 ;
    RECT 181.245 16.87 181.315 16.94 ;
    RECT 181.245 19.75 181.315 19.82 ;
    RECT 181.245 20.47 181.315 20.54 ;
    RECT 181.245 21.915 181.315 21.985 ;
    RECT 181.245 23.35 181.315 23.42 ;
    RECT 181.245 25.51 181.315 25.58 ;
    RECT 181.455 14.7 181.525 14.77 ;
    RECT 181.455 18.315 181.665 18.385 ;
    RECT 181.455 19.03 181.665 19.1 ;
    RECT 181.455 29.12 181.665 29.19 ;
    RECT 181.49 13.985 181.56 14.055 ;
    RECT 181.595 14.7 181.665 14.77 ;
    RECT 181.825 13.265 182.055 13.335 ;
    RECT 181.825 13.98 182.055 14.05 ;
    RECT 181.825 16.87 182.055 16.94 ;
    RECT 181.825 19.75 182.055 19.82 ;
    RECT 181.825 20.47 182.055 20.54 ;
    RECT 181.825 21.915 182.055 21.985 ;
    RECT 181.825 22.63 182.055 22.7 ;
    RECT 181.825 23.35 182.055 23.42 ;
    RECT 181.825 24.79 182.055 24.86 ;
    RECT 181.825 25.51 182.055 25.58 ;
    RECT 182.535 13.98 182.805 14.05 ;
    RECT 182.535 16.87 182.805 16.94 ;
    RECT 182.535 19.75 182.805 19.82 ;
    RECT 182.535 20.47 182.805 20.54 ;
    RECT 182.535 21.915 182.805 21.985 ;
    RECT 182.535 22.63 182.805 22.7 ;
    RECT 182.535 23.35 182.805 23.42 ;
    RECT 182.535 24.79 182.805 24.86 ;
    RECT 182.535 25.51 182.805 25.58 ;
    RECT 182.54 13.265 182.8 13.335 ;
    RECT 182.54 27.675 182.8 27.745 ;
    RECT 183.06 13.265 183.32 13.335 ;
    RECT 183.085 24.065 183.295 24.135 ;
    RECT 183.085 26.225 183.295 26.295 ;
    RECT 183.085 26.945 183.295 27.015 ;
    RECT 183.71 15.43 183.78 15.5 ;
    RECT 184.105 13.265 184.345 13.335 ;
    RECT 184.12 24.065 184.33 24.135 ;
    RECT 184.12 26.225 184.33 26.295 ;
    RECT 184.12 26.945 184.33 27.015 ;
    RECT 184.505 13.98 184.775 14.05 ;
    RECT 184.505 16.87 184.775 16.94 ;
    RECT 184.505 19.035 184.775 19.105 ;
    RECT 184.505 19.75 184.775 19.82 ;
    RECT 184.505 20.47 184.775 20.54 ;
    RECT 184.505 21.915 184.775 21.985 ;
    RECT 184.505 22.63 184.775 22.7 ;
    RECT 184.505 23.35 184.775 23.42 ;
    RECT 184.505 24.79 184.775 24.86 ;
    RECT 184.505 25.51 184.775 25.58 ;
    RECT 184.915 14.7 184.985 14.77 ;
    RECT 184.915 14.7 184.985 14.77 ;
    RECT 184.915 34.155 184.985 34.225 ;
    RECT 185.115 33.435 185.185 33.505 ;
    RECT 185.315 30.555 185.385 30.625 ;
    RECT 185.515 27.675 185.585 27.745 ;
    RECT 185.515 31.99 185.585 32.06 ;
    RECT 185.715 25.51 185.785 25.58 ;
    RECT 185.715 31.27 185.785 31.34 ;
    RECT 185.91 22.63 185.98 22.7 ;
    RECT 185.91 32.71 185.98 32.78 ;
    RECT 186.11 19.03 186.18 19.1 ;
    RECT 186.11 19.75 186.18 19.82 ;
    RECT 186.11 29.835 186.18 29.905 ;
    RECT 186.31 16.87 186.38 16.94 ;
    RECT 186.31 29.115 186.38 29.185 ;
    RECT 186.51 13.98 186.58 14.05 ;
    RECT 186.51 28.39 186.58 28.46 ;
    RECT 186.73 20.47 186.8 20.54 ;
    RECT 186.73 21.195 186.8 21.265 ;
    RECT 186.73 21.915 186.8 21.985 ;
    RECT 186.73 23.35 186.8 23.42 ;
    RECT 186.73 24.79 186.8 24.86 ;
    RECT 187.045 13.98 187.255 14.05 ;
    RECT 187.045 16.87 187.255 16.94 ;
    RECT 187.045 18.31 187.255 18.38 ;
    RECT 187.045 19.03 187.255 19.1 ;
    RECT 187.045 19.75 187.255 19.82 ;
    RECT 187.045 22.63 187.255 22.7 ;
    RECT 187.045 25.515 187.255 25.585 ;
    RECT 187.045 27.675 187.255 27.745 ;
    RECT 187.045 28.395 187.255 28.465 ;
    RECT 187.045 29.115 187.255 29.185 ;
    RECT 187.045 29.835 187.255 29.905 ;
    RECT 187.045 30.555 187.255 30.625 ;
    RECT 187.045 31.28 187.255 31.35 ;
    RECT 187.045 32.0 187.255 32.07 ;
    RECT 187.045 32.72 187.255 32.79 ;
    RECT 187.045 33.435 187.255 33.505 ;
    RECT 187.46 14.7 187.67 14.77 ;
    RECT 187.46 16.87 187.67 16.94 ;
    RECT 187.46 18.315 187.67 18.385 ;
    RECT 187.46 19.035 187.685 19.105 ;
    RECT 187.46 19.755 187.67 19.825 ;
    RECT 187.46 21.195 187.7 21.265 ;
    RECT 187.46 22.63 187.695 22.7 ;
    RECT 187.46 25.51 187.69 25.58 ;
    RECT 187.46 34.155 187.67 34.225 ;
    RECT 187.465 13.98 187.705 14.05 ;
    RECT 187.47 30.555 187.705 30.625 ;
    RECT 187.47 31.28 187.705 31.35 ;
    RECT 187.47 32.0 187.705 32.07 ;
    RECT 187.47 32.72 187.705 32.79 ;
    RECT 187.47 33.435 187.705 33.505 ;
    RECT 187.475 29.115 187.705 29.185 ;
    RECT 187.475 29.835 187.705 29.905 ;
    RECT 187.495 27.675 187.705 27.745 ;
    RECT 187.495 28.395 187.705 28.465 ;
    RECT 187.835 20.47 187.905 20.54 ;
    RECT 187.835 20.47 187.905 20.54 ;
    RECT 187.835 21.915 187.905 21.985 ;
    RECT 187.835 21.915 187.905 21.985 ;
    RECT 187.835 23.35 187.905 23.42 ;
    RECT 187.835 23.35 187.905 23.42 ;
    RECT 187.835 24.79 187.905 24.86 ;
    RECT 187.835 24.79 187.905 24.86 ;
    RECT 188.025 28.395 188.095 28.465 ;
    RECT 188.215 29.11 188.285 29.18 ;
    RECT 188.42 29.835 188.49 29.905 ;
    RECT 188.62 32.71 188.69 32.78 ;
    RECT 188.82 31.275 188.89 31.345 ;
    RECT 189.02 31.99 189.09 32.06 ;
    RECT 189.22 30.555 189.29 30.625 ;
    RECT 189.415 33.43 189.485 33.5 ;
    RECT 189.62 20.47 189.855 20.54 ;
    RECT 189.62 21.915 189.855 21.985 ;
    RECT 189.62 22.63 189.855 22.7 ;
    RECT 189.62 23.35 189.855 23.42 ;
    RECT 189.62 25.51 189.87 25.58 ;
    RECT 189.625 24.79 189.875 24.86 ;
    RECT 189.635 14.695 189.87 14.765 ;
    RECT 189.635 19.035 189.87 19.105 ;
    RECT 190.04 13.98 190.25 14.05 ;
    RECT 190.04 16.87 190.25 16.94 ;
    RECT 190.04 18.315 190.25 18.385 ;
    RECT 190.04 19.755 190.25 19.825 ;
    RECT 190.04 22.63 190.25 22.7 ;
    RECT 190.04 34.155 190.25 34.225 ;
    RECT 190.76 20.47 190.83 20.54 ;
    RECT 190.76 21.915 190.83 21.985 ;
    RECT 190.76 23.35 190.83 23.42 ;
    RECT 190.99 21.19 191.26 21.26 ;
    RECT 190.99 22.63 191.23 22.7 ;
    RECT 191.01 13.98 191.22 14.05 ;
    RECT 191.01 24.795 191.22 24.865 ;
    RECT 191.02 24.065 191.23 24.135 ;
    RECT 191.02 25.515 191.23 25.585 ;
    RECT 191.02 26.225 191.23 26.295 ;
    RECT 191.02 26.945 191.23 27.015 ;
    RECT 191.485 22.63 191.555 22.7 ;
    RECT 191.485 24.79 191.555 24.86 ;
    RECT 191.485 25.51 191.555 25.58 ;
    RECT 191.49 13.265 191.56 13.335 ;
    RECT 191.49 27.67 191.56 27.74 ;
    RECT 191.51 13.99 191.58 14.06 ;
    RECT 191.52 21.19 191.59 21.26 ;
    RECT 191.81 20.47 192.08 20.54 ;
    RECT 191.81 21.915 192.08 21.985 ;
    RECT 191.81 23.35 192.075 23.42 ;
    RECT 191.82 22.63 192.08 22.7 ;
    RECT 191.82 27.67 192.08 27.74 ;
    RECT 191.835 24.79 192.08 24.86 ;
    RECT 191.855 13.265 192.08 13.335 ;
    RECT 191.855 13.98 192.08 14.05 ;
    RECT 191.855 21.19 192.08 21.26 ;
    RECT 191.855 25.51 192.08 25.58 ;
    RECT 192.82 13.985 193.09 14.055 ;
    RECT 192.825 11.51 193.085 11.58 ;
    RECT 192.85 11.84 193.06 11.91 ;
    RECT 192.85 13.27 193.06 13.34 ;
    RECT 192.85 15.435 193.06 15.505 ;
    RECT 192.85 16.155 193.06 16.225 ;
    RECT 192.85 16.87 193.06 16.94 ;
    RECT 192.85 18.315 193.06 18.385 ;
    RECT 192.85 19.03 193.06 19.1 ;
    RECT 192.85 19.755 193.06 19.825 ;
    RECT 192.85 20.47 193.06 20.54 ;
    RECT 192.85 21.915 193.06 21.985 ;
    RECT 192.85 23.355 193.06 23.425 ;
    RECT 192.85 25.515 193.06 25.585 ;
    RECT 192.85 27.675 193.06 27.745 ;
    RECT 192.88 17.59 193.09 17.66 ;
    RECT 193.565 12.555 193.835 12.625 ;
    RECT 193.565 13.985 193.835 14.055 ;
    RECT 193.57 11.835 193.83 11.905 ;
    RECT 193.57 14.7 193.83 14.77 ;
    RECT 193.57 29.11 193.78 29.18 ;
    RECT 193.57 29.83 193.78 29.9 ;
    RECT 193.57 30.55 193.83 30.62 ;
    RECT 193.57 31.275 193.83 31.345 ;
    RECT 193.57 31.995 193.83 32.065 ;
    RECT 193.57 32.715 193.83 32.785 ;
    RECT 193.57 33.43 193.83 33.5 ;
    RECT 193.595 24.065 193.805 24.135 ;
    RECT 193.595 26.225 193.805 26.295 ;
    RECT 193.595 26.945 193.805 27.015 ;
    RECT 193.62 15.435 193.83 15.505 ;
    RECT 193.62 17.595 193.83 17.665 ;
    RECT 193.62 20.475 193.83 20.545 ;
    RECT 193.62 21.915 193.83 21.985 ;
    RECT 193.62 23.355 193.83 23.425 ;
    RECT 193.62 25.515 193.83 25.585 ;
    RECT 193.62 27.675 193.83 27.745 ;
    RECT 193.625 16.155 193.835 16.225 ;
    RECT 194.015 26.225 194.085 26.295 ;
    RECT 194.015 26.945 194.085 27.015 ;
    RECT 194.015 27.675 194.085 27.745 ;
    RECT 194.015 29.11 194.085 29.18 ;
    RECT 194.015 29.83 194.085 29.9 ;
    RECT 194.015 30.55 194.085 30.62 ;
    RECT 194.015 31.275 194.085 31.345 ;
    RECT 194.015 31.995 194.085 32.065 ;
    RECT 194.015 32.715 194.085 32.785 ;
    RECT 194.015 33.43 194.085 33.5 ;
    RECT 194.015 34.155 194.085 34.225 ;
    RECT 194.505 11.835 194.765 11.905 ;
    RECT 194.505 12.55 194.765 12.62 ;
    RECT 194.505 13.985 194.765 14.055 ;
    RECT 194.505 14.7 194.765 14.77 ;
    RECT 194.505 15.435 194.765 15.505 ;
    RECT 194.505 16.15 194.765 16.22 ;
    RECT 194.505 17.59 194.765 17.66 ;
    RECT 194.505 23.35 194.765 23.42 ;
    RECT 194.505 26.225 194.765 26.295 ;
    RECT 194.505 26.945 194.765 27.015 ;
    RECT 194.505 27.675 194.765 27.745 ;
    RECT 194.505 29.11 194.765 29.18 ;
    RECT 194.505 29.83 194.765 29.9 ;
    RECT 194.505 30.55 194.765 30.62 ;
    RECT 194.505 31.275 194.765 31.345 ;
    RECT 194.505 31.995 194.765 32.065 ;
    RECT 194.505 32.715 194.765 32.785 ;
    RECT 194.505 33.43 194.765 33.5 ;
    RECT 194.505 34.15 194.765 34.22 ;
    RECT 194.535 13.27 194.745 13.34 ;
    RECT 194.535 16.87 194.745 16.94 ;
    RECT 194.535 18.315 194.745 18.385 ;
    RECT 194.535 19.03 194.745 19.1 ;
    RECT 194.535 19.755 194.745 19.825 ;
    RECT 195.63 11.835 195.84 11.905 ;
    RECT 195.63 12.55 195.84 12.62 ;
    RECT 195.63 13.265 195.84 13.335 ;
    RECT 195.63 13.985 195.84 14.055 ;
    RECT 195.63 14.715 195.84 14.785 ;
    RECT 195.63 15.435 195.84 15.505 ;
    RECT 195.63 16.15 195.84 16.22 ;
    RECT 195.63 16.87 195.84 16.94 ;
    RECT 195.63 17.59 195.84 17.66 ;
    RECT 195.63 18.31 195.84 18.38 ;
    RECT 195.63 19.035 195.84 19.105 ;
    RECT 195.63 19.755 195.84 19.825 ;
    RECT 195.63 22.63 195.84 22.7 ;
    RECT 195.63 23.35 195.84 23.42 ;
    RECT 195.63 24.795 195.84 24.865 ;
    RECT 195.63 26.225 195.84 26.295 ;
    RECT 195.63 26.945 195.84 27.015 ;
    RECT 195.63 27.675 195.84 27.745 ;
    RECT 195.63 28.39 195.84 28.46 ;
    RECT 195.63 29.11 195.84 29.18 ;
    RECT 195.63 29.83 195.84 29.9 ;
    RECT 195.63 30.55 195.84 30.62 ;
    RECT 195.63 31.275 195.84 31.345 ;
    RECT 195.63 31.995 195.84 32.065 ;
    RECT 195.63 32.715 195.84 32.785 ;
    RECT 195.63 33.43 195.84 33.5 ;
    RECT 195.63 34.15 195.84 34.22 ;
    RECT 197.465 12.01 198.255 12.08 ;
    RECT 197.465 12.73 198.255 12.8 ;
    RECT 197.465 13.445 198.255 13.515 ;
    RECT 197.465 14.17 198.255 14.24 ;
    RECT 197.465 14.89 198.255 14.96 ;
    RECT 197.465 15.61 198.255 15.68 ;
    RECT 197.465 16.325 198.255 16.395 ;
    RECT 197.465 17.05 198.255 17.12 ;
    RECT 197.465 17.77 198.255 17.84 ;
    RECT 197.465 18.485 198.255 18.555 ;
    RECT 197.465 19.21 198.255 19.28 ;
    RECT 197.465 19.93 198.255 20.0 ;
    RECT 197.465 20.65 198.255 20.72 ;
    RECT 197.465 21.37 198.255 21.44 ;
    RECT 197.465 22.09 198.255 22.16 ;
    RECT 197.465 22.81 198.255 22.88 ;
    RECT 197.465 23.53 198.255 23.6 ;
    RECT 197.465 24.25 198.255 24.32 ;
    RECT 197.465 24.97 198.255 25.04 ;
    RECT 197.465 25.69 198.255 25.76 ;
    RECT 197.465 26.41 198.255 26.48 ;
    RECT 197.465 27.13 198.255 27.2 ;
    RECT 197.465 27.845 198.255 27.915 ;
    RECT 197.465 28.565 198.255 28.635 ;
    RECT 197.465 29.29 198.255 29.36 ;
    RECT 197.465 30.01 198.255 30.08 ;
    RECT 197.465 30.73 198.255 30.8 ;
    RECT 197.465 31.45 198.255 31.52 ;
    RECT 197.465 32.17 198.255 32.24 ;
    RECT 197.465 32.885 198.255 32.955 ;
    RECT 197.465 33.605 198.255 33.675 ;
    RECT 197.465 34.33 198.255 34.4 ;
    RECT 199.245 11.565 199.515 34.675 ;
    RECT 199.245 32.445 199.515 32.515 ;
    RECT 192.85 39.915 193.06 39.985 ;
    RECT 180.81 39.912 181.02 39.982 ;
    RECT 193.595 19.752 193.805 19.822 ;
    RECT 188.225 49.272 188.295 49.342 ;
    RECT 193.595 19.032 193.805 19.102 ;
    RECT 193.595 18.312 193.805 18.382 ;
    RECT 193.595 16.872 193.805 16.942 ;
    RECT 185.715 48.552 185.785 48.622 ;
    RECT 188.225 42.792 188.295 42.862 ;
    RECT 186.31 39.192 186.38 39.262 ;
    RECT 175.75 40.005 175.96 40.075 ;
    RECT 185.715 47.832 185.785 47.902 ;
    RECT 188.225 42.072 188.295 42.142 ;
    RECT 192.85 47.835 193.06 47.905 ;
    RECT 180.81 47.832 181.02 47.902 ;
    RECT 198.605 39.285 198.815 39.355 ;
    RECT 175.75 47.925 175.96 47.995 ;
    RECT 192.85 39.195 193.06 39.265 ;
    RECT 186.31 38.472 186.38 38.542 ;
    RECT 175.75 19.845 175.96 19.915 ;
    RECT 180.81 39.192 181.02 39.262 ;
    RECT 175.75 19.125 175.96 19.195 ;
    RECT 175.75 18.405 175.96 18.475 ;
    RECT 175.75 39.285 175.96 39.355 ;
    RECT 185.715 47.112 185.785 47.182 ;
    RECT 175.75 17.685 175.96 17.755 ;
    RECT 198.605 47.205 198.815 47.275 ;
    RECT 175.75 16.965 175.96 17.035 ;
    RECT 192.85 47.115 193.06 47.185 ;
    RECT 175.75 16.245 175.96 16.315 ;
    RECT 175.75 15.525 175.96 15.595 ;
    RECT 180.81 47.112 181.02 47.182 ;
    RECT 186.31 37.752 186.38 37.822 ;
    RECT 174.56 59.105 174.63 59.175 ;
    RECT 175.16 59.105 175.37 59.175 ;
    RECT 175.515 60.125 175.585 60.195 ;
    RECT 176.355 59.56 177.095 59.63 ;
    RECT 177.375 59.27 177.585 59.34 ;
    RECT 177.835 60.125 178.045 60.195 ;
    RECT 178.23 59.27 178.44 59.34 ;
    RECT 179.88 59.27 180.09 59.34 ;
    RECT 180.44 60.125 180.65 60.195 ;
    RECT 180.81 59.7 181.02 59.77 ;
    RECT 181.225 60.125 181.295 60.195 ;
    RECT 181.835 60.125 182.045 60.195 ;
    RECT 182.565 60.125 182.775 60.195 ;
    RECT 183.085 59.7 183.295 59.77 ;
    RECT 184.12 59.7 184.33 59.77 ;
    RECT 184.535 60.125 184.745 60.195 ;
    RECT 184.915 59.27 184.985 59.34 ;
    RECT 186.695 60.125 186.905 60.195 ;
    RECT 187.46 59.27 187.67 59.34 ;
    RECT 187.835 60.125 187.905 60.195 ;
    RECT 189.655 60.125 189.865 60.195 ;
    RECT 190.04 59.27 190.25 59.34 ;
    RECT 190.745 60.125 190.815 60.195 ;
    RECT 191.02 59.7 191.23 59.77 ;
    RECT 191.49 59.415 191.56 59.485 ;
    RECT 191.84 60.125 192.05 60.195 ;
    RECT 192.85 59.27 193.06 59.34 ;
    RECT 193.595 59.7 193.805 59.77 ;
    RECT 194.535 59.27 194.745 59.34 ;
    RECT 195.055 60.125 195.265 60.195 ;
    RECT 196.185 59.27 196.255 59.34 ;
    RECT 196.43 60.125 196.64 60.195 ;
    RECT 196.81 59.27 197.02 59.34 ;
    RECT 197.465 59.56 198.255 59.63 ;
    RECT 198.99 60.125 199.06 60.195 ;
    RECT 199.245 59.105 199.515 59.175 ;
    RECT 199.885 60.125 200.095 60.195 ;
    RECT 198.605 38.565 198.815 38.635 ;
    RECT 192.85 38.475 193.06 38.545 ;
    RECT 180.81 38.472 181.02 38.542 ;
    RECT 188.225 55.752 188.295 55.822 ;
    RECT 175.75 14.805 175.96 14.875 ;
    RECT 175.75 14.085 175.96 14.155 ;
    RECT 175.75 13.365 175.96 13.435 ;
    RECT 175.75 12.645 175.96 12.715 ;
    RECT 175.75 47.205 175.96 47.275 ;
    RECT 175.75 11.925 175.96 11.995 ;
    RECT 198.605 59.267 198.815 59.337 ;
    RECT 193.595 59.267 193.805 59.337 ;
    RECT 175.75 38.565 175.96 38.635 ;
    RECT 198.605 46.485 198.815 46.555 ;
    RECT 186.51 37.032 186.58 37.102 ;
    RECT 192.85 46.395 193.06 46.465 ;
    RECT 180.81 46.392 181.02 46.462 ;
    RECT 198.605 37.845 198.815 37.915 ;
    RECT 192.85 37.755 193.06 37.825 ;
    RECT 180.81 37.752 181.02 37.822 ;
    RECT 188.225 55.032 188.295 55.102 ;
    RECT 192.85 59.7 193.06 59.77 ;
    RECT 191.02 59.267 191.23 59.337 ;
    RECT 186.51 36.312 186.58 36.382 ;
    RECT 175.75 46.485 175.96 46.555 ;
    RECT 175.75 37.845 175.96 37.915 ;
    RECT 190.04 59.7 190.25 59.77 ;
    RECT 184.915 59.7 184.985 59.77 ;
    RECT 184.12 59.267 184.33 59.337 ;
    RECT 198.605 45.765 198.815 45.835 ;
    RECT 183.085 59.267 183.295 59.337 ;
    RECT 192.85 45.675 193.06 45.745 ;
    RECT 180.81 59.267 181.02 59.337 ;
    RECT 180.81 45.672 181.02 45.742 ;
    RECT 198.605 37.125 198.815 37.195 ;
    RECT 188.225 54.312 188.295 54.382 ;
    RECT 192.85 37.035 193.06 37.105 ;
    RECT 179.88 59.7 180.09 59.77 ;
    RECT 175.75 59.267 175.96 59.337 ;
    RECT 175.75 45.765 175.96 45.835 ;
    RECT 180.81 37.032 181.02 37.102 ;
    RECT 175.75 37.125 175.96 37.195 ;
    RECT 198.605 45.045 198.815 45.115 ;
    RECT 192.85 44.955 193.06 45.025 ;
    RECT 188.225 53.592 188.295 53.662 ;
    RECT 180.81 44.952 181.02 45.022 ;
    RECT 198.605 36.405 198.815 36.475 ;
    RECT 192.85 36.315 193.06 36.385 ;
    RECT 188.225 52.872 188.295 52.942 ;
    RECT 175.75 45.045 175.96 45.115 ;
    RECT 180.81 36.312 181.02 36.382 ;
    RECT 175.75 36.405 175.96 36.475 ;
    RECT 198.605 44.325 198.815 44.395 ;
    RECT 192.85 44.235 193.06 44.305 ;
    RECT 198.605 35.685 198.815 35.755 ;
    RECT 192.85 35.595 193.06 35.665 ;
    RECT 195.63 59.557 195.84 59.627 ;
    RECT 188.225 52.152 188.295 52.222 ;
    RECT 178.79 59.557 179.0 59.627 ;
    RECT 180.81 44.232 181.02 44.302 ;
    RECT 175.75 44.325 175.96 44.395 ;
    RECT 180.81 35.592 181.02 35.662 ;
    RECT 175.75 35.685 175.96 35.755 ;
    RECT 198.605 43.605 198.815 43.675 ;
    RECT 192.85 43.515 193.06 43.585 ;
    RECT 198.605 34.965 198.815 35.035 ;
    RECT 192.85 34.875 193.06 34.945 ;
    RECT 188.425 58.652 188.495 58.722 ;
    RECT 188.225 51.432 188.295 51.502 ;
    RECT 188.225 48.552 188.295 48.622 ;
    RECT 180.81 43.512 181.02 43.582 ;
    RECT 198.605 54.405 198.815 54.475 ;
    RECT 192.85 54.315 193.06 54.385 ;
    RECT 175.75 43.605 175.96 43.675 ;
    RECT 188.225 57.192 188.295 57.262 ;
    RECT 180.81 54.312 181.02 54.382 ;
    RECT 198.605 42.885 198.815 42.955 ;
    RECT 180.81 34.152 181.02 34.222 ;
    RECT 192.85 42.795 193.06 42.865 ;
    RECT 180.81 29.117 181.02 29.187 ;
    RECT 175.75 54.405 175.96 54.475 ;
    RECT 188.225 47.832 188.295 47.902 ;
    RECT 180.81 42.792 181.02 42.862 ;
    RECT 198.605 53.685 198.815 53.755 ;
    RECT 192.85 53.595 193.06 53.665 ;
    RECT 175.75 42.885 175.96 42.955 ;
    RECT 180.81 53.592 181.02 53.662 ;
    RECT 198.605 58.745 198.815 58.815 ;
    RECT 192.85 58.655 193.06 58.725 ;
    RECT 198.605 42.165 198.815 42.235 ;
    RECT 192.85 42.075 193.06 42.145 ;
    RECT 175.75 53.685 175.96 53.755 ;
    RECT 188.225 47.112 188.295 47.182 ;
    RECT 180.81 19.032 181.02 19.102 ;
    RECT 180.81 58.652 181.02 58.722 ;
    RECT 180.81 18.312 181.02 18.382 ;
    RECT 180.81 14.697 181.02 14.767 ;
    RECT 175.75 58.745 175.96 58.815 ;
    RECT 180.81 13.982 181.02 14.052 ;
    RECT 180.81 42.072 181.02 42.142 ;
    RECT 198.605 52.965 198.815 53.035 ;
    RECT 192.85 52.875 193.06 52.945 ;
    RECT 175.75 42.165 175.96 42.235 ;
    RECT 180.81 52.872 181.02 52.942 ;
    RECT 188.225 46.392 188.295 46.462 ;
    RECT 198.605 57.285 198.815 57.355 ;
    RECT 192.85 57.195 193.06 57.265 ;
    RECT 175.75 34.245 175.96 34.315 ;
    RECT 175.75 33.525 175.96 33.595 ;
    RECT 175.75 32.805 175.96 32.875 ;
    RECT 175.75 52.965 175.96 53.035 ;
    RECT 180.81 57.192 181.02 57.262 ;
    RECT 175.75 57.285 175.96 57.355 ;
    RECT 198.605 52.245 198.815 52.315 ;
    RECT 192.85 52.155 193.06 52.225 ;
    RECT 175.75 32.085 175.96 32.155 ;
    RECT 175.75 31.365 175.96 31.435 ;
    RECT 180.81 52.152 181.02 52.222 ;
    RECT 175.75 30.645 175.96 30.715 ;
    RECT 198.605 56.565 198.815 56.635 ;
    RECT 192.85 56.475 193.06 56.545 ;
    RECT 198.605 41.445 198.815 41.515 ;
    RECT 175.75 52.245 175.96 52.315 ;
    RECT 195.63 58.087 195.84 58.157 ;
    RECT 178.79 58.087 179.0 58.157 ;
    RECT 175.75 29.925 175.96 29.995 ;
    RECT 180.81 56.472 181.02 56.542 ;
    RECT 175.75 29.205 175.96 29.275 ;
    RECT 175.75 56.565 175.96 56.635 ;
    RECT 175.75 28.485 175.96 28.555 ;
    RECT 198.605 51.525 198.815 51.595 ;
    RECT 192.85 51.435 193.06 51.505 ;
    RECT 175.75 27.765 175.96 27.835 ;
    RECT 175.75 27.045 175.96 27.115 ;
    RECT 180.81 51.432 181.02 51.502 ;
    RECT 374.13 4.055 374.2 4.125 ;
    RECT 373.93 4.455 374.0 4.525 ;
    RECT 373.94 5.33 374.01 5.54 ;
    RECT 373.94 3.235 374.01 3.445 ;
    RECT 374.36 11.065 374.43 11.135 ;
    RECT 374.15 11.325 374.22 11.395 ;
    RECT 373.94 9.12 374.01 9.33 ;
    RECT 227.3 4.455 227.51 4.525 ;
    RECT 216.42 7.28 216.63 7.35 ;
    RECT 216.42 6.385 216.63 6.455 ;
    RECT 250.54 4.455 250.75 4.525 ;
    RECT 366.74 3.235 366.95 3.445 ;
    RECT 366.74 5.33 366.95 5.54 ;
    RECT 366.74 9.12 366.95 9.33 ;
    RECT 366.31 4.845 366.38 4.915 ;
    RECT 366.31 9.43 366.38 9.5 ;
    RECT 365.33 9.765 365.54 9.835 ;
    RECT 364.87 2.585 365.08 2.795 ;
    RECT 364.87 5.86 365.08 6.07 ;
    RECT 364.87 6.385 365.08 6.455 ;
    RECT 364.87 7.28 365.08 7.35 ;
    RECT 306.06 4.055 306.27 4.125 ;
    RECT 363.42 3.235 363.63 3.445 ;
    RECT 363.42 5.33 363.63 5.54 ;
    RECT 363.42 9.12 363.63 9.33 ;
    RECT 362.99 4.845 363.06 4.915 ;
    RECT 362.99 9.43 363.06 9.5 ;
    RECT 362.01 9.765 362.22 9.835 ;
    RECT 361.55 2.585 361.76 2.795 ;
    RECT 361.55 5.86 361.76 6.07 ;
    RECT 361.55 6.385 361.76 6.455 ;
    RECT 361.55 7.28 361.76 7.35 ;
    RECT 246.3 4.055 246.51 4.125 ;
    RECT 360.1 3.235 360.31 3.445 ;
    RECT 360.1 5.33 360.31 5.54 ;
    RECT 360.1 9.12 360.31 9.33 ;
    RECT 359.67 4.845 359.74 4.915 ;
    RECT 359.67 9.43 359.74 9.5 ;
    RECT 358.69 9.765 358.9 9.835 ;
    RECT 358.23 2.585 358.44 2.795 ;
    RECT 358.23 5.86 358.44 6.07 ;
    RECT 358.23 6.385 358.44 6.455 ;
    RECT 358.23 7.28 358.44 7.35 ;
    RECT 356.78 3.235 356.99 3.445 ;
    RECT 356.78 5.33 356.99 5.54 ;
    RECT 356.78 9.12 356.99 9.33 ;
    RECT 356.35 4.845 356.42 4.915 ;
    RECT 356.35 9.43 356.42 9.5 ;
    RECT 355.37 9.765 355.58 9.835 ;
    RECT 354.91 2.585 355.12 2.795 ;
    RECT 354.91 5.86 355.12 6.07 ;
    RECT 354.91 6.385 355.12 6.455 ;
    RECT 354.91 7.28 355.12 7.35 ;
    RECT 353.46 3.235 353.67 3.445 ;
    RECT 353.46 5.33 353.67 5.54 ;
    RECT 353.46 9.12 353.67 9.33 ;
    RECT 353.03 4.845 353.1 4.915 ;
    RECT 353.03 9.43 353.1 9.5 ;
    RECT 352.05 9.765 352.26 9.835 ;
    RECT 351.59 2.585 351.8 2.795 ;
    RECT 351.59 5.86 351.8 6.07 ;
    RECT 351.59 6.385 351.8 6.455 ;
    RECT 351.59 7.28 351.8 7.35 ;
    RECT 350.14 3.235 350.35 3.445 ;
    RECT 350.14 5.33 350.35 5.54 ;
    RECT 350.14 9.12 350.35 9.33 ;
    RECT 349.71 4.845 349.78 4.915 ;
    RECT 349.71 9.43 349.78 9.5 ;
    RECT 348.73 9.765 348.94 9.835 ;
    RECT 348.27 2.585 348.48 2.795 ;
    RECT 348.27 5.86 348.48 6.07 ;
    RECT 348.27 6.385 348.48 6.455 ;
    RECT 348.27 7.28 348.48 7.35 ;
    RECT 346.82 3.235 347.03 3.445 ;
    RECT 346.82 5.33 347.03 5.54 ;
    RECT 346.82 9.12 347.03 9.33 ;
    RECT 346.39 4.845 346.46 4.915 ;
    RECT 346.39 9.43 346.46 9.5 ;
    RECT 345.41 9.765 345.62 9.835 ;
    RECT 344.95 2.585 345.16 2.795 ;
    RECT 344.95 5.86 345.16 6.07 ;
    RECT 344.95 6.385 345.16 6.455 ;
    RECT 344.95 7.28 345.16 7.35 ;
    RECT 343.5 3.235 343.71 3.445 ;
    RECT 343.5 5.33 343.71 5.54 ;
    RECT 343.5 9.12 343.71 9.33 ;
    RECT 343.07 4.845 343.14 4.915 ;
    RECT 343.07 9.43 343.14 9.5 ;
    RECT 342.09 9.765 342.3 9.835 ;
    RECT 341.63 2.585 341.84 2.795 ;
    RECT 341.63 5.86 341.84 6.07 ;
    RECT 341.63 6.385 341.84 6.455 ;
    RECT 341.63 7.28 341.84 7.35 ;
    RECT 340.18 3.235 340.39 3.445 ;
    RECT 340.18 5.33 340.39 5.54 ;
    RECT 340.18 9.12 340.39 9.33 ;
    RECT 339.75 4.845 339.82 4.915 ;
    RECT 339.75 9.43 339.82 9.5 ;
    RECT 338.77 9.765 338.98 9.835 ;
    RECT 338.31 2.585 338.52 2.795 ;
    RECT 338.31 5.86 338.52 6.07 ;
    RECT 338.31 6.385 338.52 6.455 ;
    RECT 338.31 7.28 338.52 7.35 ;
    RECT 336.86 3.235 337.07 3.445 ;
    RECT 336.86 5.33 337.07 5.54 ;
    RECT 336.86 9.12 337.07 9.33 ;
    RECT 336.43 4.845 336.5 4.915 ;
    RECT 336.43 9.43 336.5 9.5 ;
    RECT 335.45 9.765 335.66 9.835 ;
    RECT 334.99 2.585 335.2 2.795 ;
    RECT 334.99 5.86 335.2 6.07 ;
    RECT 334.99 6.385 335.2 6.455 ;
    RECT 334.99 7.28 335.2 7.35 ;
    RECT 252.94 7.28 253.15 7.35 ;
    RECT 352.54 7.28 352.75 7.35 ;
    RECT 252.94 6.385 253.15 6.455 ;
    RECT 352.54 6.385 352.75 6.455 ;
    RECT 252.94 5.86 253.15 6.07 ;
    RECT 352.54 5.86 352.75 6.07 ;
    RECT 252.94 2.585 253.15 2.795 ;
    RECT 216.42 5.86 216.63 6.07 ;
    RECT 352.54 2.585 352.75 2.795 ;
    RECT 343.5 4.455 343.71 4.525 ;
    RECT 216.42 2.585 216.63 2.795 ;
    RECT 223.98 4.455 224.19 4.525 ;
    RECT 333.54 3.235 333.75 3.445 ;
    RECT 333.54 5.33 333.75 5.54 ;
    RECT 333.54 9.12 333.75 9.33 ;
    RECT 333.11 4.845 333.18 4.915 ;
    RECT 333.11 9.43 333.18 9.5 ;
    RECT 332.13 9.765 332.34 9.835 ;
    RECT 331.67 2.585 331.88 2.795 ;
    RECT 331.67 5.86 331.88 6.07 ;
    RECT 331.67 6.385 331.88 6.455 ;
    RECT 331.67 7.28 331.88 7.35 ;
    RECT 330.22 3.235 330.43 3.445 ;
    RECT 330.22 5.33 330.43 5.54 ;
    RECT 330.22 9.12 330.43 9.33 ;
    RECT 329.79 4.845 329.86 4.915 ;
    RECT 329.79 9.43 329.86 9.5 ;
    RECT 328.81 9.765 329.02 9.835 ;
    RECT 328.35 2.585 328.56 2.795 ;
    RECT 328.35 5.86 328.56 6.07 ;
    RECT 328.35 6.385 328.56 6.455 ;
    RECT 328.35 7.28 328.56 7.35 ;
    RECT 326.9 3.235 327.11 3.445 ;
    RECT 326.9 5.33 327.11 5.54 ;
    RECT 326.9 9.12 327.11 9.33 ;
    RECT 326.47 4.845 326.54 4.915 ;
    RECT 326.47 9.43 326.54 9.5 ;
    RECT 325.49 9.765 325.7 9.835 ;
    RECT 325.03 2.585 325.24 2.795 ;
    RECT 325.03 5.86 325.24 6.07 ;
    RECT 325.03 6.385 325.24 6.455 ;
    RECT 325.03 7.28 325.24 7.35 ;
    RECT 323.58 3.235 323.79 3.445 ;
    RECT 323.58 5.33 323.79 5.54 ;
    RECT 323.58 9.12 323.79 9.33 ;
    RECT 323.15 4.845 323.22 4.915 ;
    RECT 323.15 9.43 323.22 9.5 ;
    RECT 322.17 9.765 322.38 9.835 ;
    RECT 321.71 2.585 321.92 2.795 ;
    RECT 321.71 5.86 321.92 6.07 ;
    RECT 321.71 6.385 321.92 6.455 ;
    RECT 321.71 7.28 321.92 7.35 ;
    RECT 320.26 3.235 320.47 3.445 ;
    RECT 320.26 5.33 320.47 5.54 ;
    RECT 320.26 9.12 320.47 9.33 ;
    RECT 319.83 4.845 319.9 4.915 ;
    RECT 319.83 9.43 319.9 9.5 ;
    RECT 318.85 9.765 319.06 9.835 ;
    RECT 318.39 2.585 318.6 2.795 ;
    RECT 318.39 5.86 318.6 6.07 ;
    RECT 318.39 6.385 318.6 6.455 ;
    RECT 318.39 7.28 318.6 7.35 ;
    RECT 302.74 4.055 302.95 4.125 ;
    RECT 247.22 4.455 247.43 4.525 ;
    RECT 316.94 3.235 317.15 3.445 ;
    RECT 316.94 5.33 317.15 5.54 ;
    RECT 316.94 9.12 317.15 9.33 ;
    RECT 316.51 4.845 316.58 4.915 ;
    RECT 316.51 9.43 316.58 9.5 ;
    RECT 315.53 9.765 315.74 9.835 ;
    RECT 315.07 2.585 315.28 2.795 ;
    RECT 315.07 5.86 315.28 6.07 ;
    RECT 315.07 6.385 315.28 6.455 ;
    RECT 315.07 7.28 315.28 7.35 ;
    RECT 242.98 4.055 243.19 4.125 ;
    RECT 313.62 3.235 313.83 3.445 ;
    RECT 313.62 5.33 313.83 5.54 ;
    RECT 313.62 9.12 313.83 9.33 ;
    RECT 313.19 4.845 313.26 4.915 ;
    RECT 313.19 9.43 313.26 9.5 ;
    RECT 312.21 9.765 312.42 9.835 ;
    RECT 311.75 2.585 311.96 2.795 ;
    RECT 311.75 5.86 311.96 6.07 ;
    RECT 311.75 6.385 311.96 6.455 ;
    RECT 311.75 7.28 311.96 7.35 ;
    RECT 310.3 3.235 310.51 3.445 ;
    RECT 310.3 5.33 310.51 5.54 ;
    RECT 310.3 9.12 310.51 9.33 ;
    RECT 309.87 4.845 309.94 4.915 ;
    RECT 309.87 9.43 309.94 9.5 ;
    RECT 308.89 9.765 309.1 9.835 ;
    RECT 308.43 2.585 308.64 2.795 ;
    RECT 308.43 5.86 308.64 6.07 ;
    RECT 308.43 6.385 308.64 6.455 ;
    RECT 308.43 7.28 308.64 7.35 ;
    RECT 339.26 7.28 339.47 7.35 ;
    RECT 306.98 3.235 307.19 3.445 ;
    RECT 306.98 5.33 307.19 5.54 ;
    RECT 306.98 9.12 307.19 9.33 ;
    RECT 306.55 4.845 306.62 4.915 ;
    RECT 306.55 9.43 306.62 9.5 ;
    RECT 305.57 9.765 305.78 9.835 ;
    RECT 305.11 2.585 305.32 2.795 ;
    RECT 305.11 5.86 305.32 6.07 ;
    RECT 305.11 6.385 305.32 6.455 ;
    RECT 305.11 7.28 305.32 7.35 ;
    RECT 339.26 6.385 339.47 6.455 ;
    RECT 303.66 3.235 303.87 3.445 ;
    RECT 303.66 5.33 303.87 5.54 ;
    RECT 303.66 9.12 303.87 9.33 ;
    RECT 303.23 4.845 303.3 4.915 ;
    RECT 303.23 9.43 303.3 9.5 ;
    RECT 302.25 9.765 302.46 9.835 ;
    RECT 301.79 2.585 302.0 2.795 ;
    RECT 301.79 5.86 302.0 6.07 ;
    RECT 301.79 6.385 302.0 6.455 ;
    RECT 301.79 7.28 302.0 7.35 ;
    RECT 339.26 5.86 339.47 6.07 ;
    RECT 339.26 2.585 339.47 2.795 ;
    RECT 249.62 7.28 249.83 7.35 ;
    RECT 249.62 6.385 249.83 6.455 ;
    RECT 349.22 7.28 349.43 7.35 ;
    RECT 213.1 7.28 213.31 7.35 ;
    RECT 349.22 6.385 349.43 6.455 ;
    RECT 213.1 6.385 213.31 6.455 ;
    RECT 340.18 4.455 340.39 4.525 ;
    RECT 213.1 5.86 213.31 6.07 ;
    RECT 213.1 2.585 213.31 2.795 ;
    RECT 233.94 3.235 234.15 3.445 ;
    RECT 233.94 5.33 234.15 5.54 ;
    RECT 233.94 9.12 234.15 9.33 ;
    RECT 233.51 4.845 233.58 4.915 ;
    RECT 233.51 9.43 233.58 9.5 ;
    RECT 232.53 9.765 232.74 9.835 ;
    RECT 232.07 2.585 232.28 2.795 ;
    RECT 232.07 5.86 232.28 6.07 ;
    RECT 232.07 6.385 232.28 6.455 ;
    RECT 232.07 7.28 232.28 7.35 ;
    RECT 230.62 3.235 230.83 3.445 ;
    RECT 230.62 5.33 230.83 5.54 ;
    RECT 230.62 9.12 230.83 9.33 ;
    RECT 230.19 4.845 230.26 4.915 ;
    RECT 230.19 9.43 230.26 9.5 ;
    RECT 229.21 9.765 229.42 9.835 ;
    RECT 228.75 2.585 228.96 2.795 ;
    RECT 228.75 5.86 228.96 6.07 ;
    RECT 228.75 6.385 228.96 6.455 ;
    RECT 228.75 7.28 228.96 7.35 ;
    RECT 227.3 3.235 227.51 3.445 ;
    RECT 227.3 5.33 227.51 5.54 ;
    RECT 227.3 9.12 227.51 9.33 ;
    RECT 226.87 4.845 226.94 4.915 ;
    RECT 226.87 9.43 226.94 9.5 ;
    RECT 225.89 9.765 226.1 9.835 ;
    RECT 225.43 2.585 225.64 2.795 ;
    RECT 225.43 5.86 225.64 6.07 ;
    RECT 225.43 6.385 225.64 6.455 ;
    RECT 225.43 7.28 225.64 7.35 ;
    RECT 223.98 3.235 224.19 3.445 ;
    RECT 223.98 5.33 224.19 5.54 ;
    RECT 223.98 9.12 224.19 9.33 ;
    RECT 223.55 4.845 223.62 4.915 ;
    RECT 223.55 9.43 223.62 9.5 ;
    RECT 222.57 9.765 222.78 9.835 ;
    RECT 222.11 2.585 222.32 2.795 ;
    RECT 222.11 5.86 222.32 6.07 ;
    RECT 222.11 6.385 222.32 6.455 ;
    RECT 222.11 7.28 222.32 7.35 ;
    RECT 220.66 3.235 220.87 3.445 ;
    RECT 220.66 5.33 220.87 5.54 ;
    RECT 220.66 9.12 220.87 9.33 ;
    RECT 220.23 4.845 220.3 4.915 ;
    RECT 220.23 9.43 220.3 9.5 ;
    RECT 219.25 9.765 219.46 9.835 ;
    RECT 218.79 2.585 219.0 2.795 ;
    RECT 218.79 5.86 219.0 6.07 ;
    RECT 218.79 6.385 219.0 6.455 ;
    RECT 218.79 7.28 219.0 7.35 ;
    RECT 300.34 3.235 300.55 3.445 ;
    RECT 300.34 5.33 300.55 5.54 ;
    RECT 300.34 9.12 300.55 9.33 ;
    RECT 299.91 4.845 299.98 4.915 ;
    RECT 299.91 9.43 299.98 9.5 ;
    RECT 298.93 9.765 299.14 9.835 ;
    RECT 298.47 2.585 298.68 2.795 ;
    RECT 298.47 5.86 298.68 6.07 ;
    RECT 298.47 6.385 298.68 6.455 ;
    RECT 298.47 7.28 298.68 7.35 ;
    RECT 233.02 4.055 233.23 4.125 ;
    RECT 217.34 3.235 217.55 3.445 ;
    RECT 217.34 5.33 217.55 5.54 ;
    RECT 217.34 9.12 217.55 9.33 ;
    RECT 216.91 4.845 216.98 4.915 ;
    RECT 216.91 9.43 216.98 9.5 ;
    RECT 215.93 9.765 216.14 9.835 ;
    RECT 215.47 2.585 215.68 2.795 ;
    RECT 215.47 5.86 215.68 6.07 ;
    RECT 215.47 6.385 215.68 6.455 ;
    RECT 215.47 7.28 215.68 7.35 ;
    RECT 297.02 3.235 297.23 3.445 ;
    RECT 297.02 5.33 297.23 5.54 ;
    RECT 297.02 9.12 297.23 9.33 ;
    RECT 296.59 4.845 296.66 4.915 ;
    RECT 296.59 9.43 296.66 9.5 ;
    RECT 295.61 9.765 295.82 9.835 ;
    RECT 295.15 2.585 295.36 2.795 ;
    RECT 295.15 5.86 295.36 6.07 ;
    RECT 295.15 6.385 295.36 6.455 ;
    RECT 295.15 7.28 295.36 7.35 ;
    RECT 214.02 3.235 214.23 3.445 ;
    RECT 214.02 5.33 214.23 5.54 ;
    RECT 214.02 9.12 214.23 9.33 ;
    RECT 213.59 4.845 213.66 4.915 ;
    RECT 213.59 9.43 213.66 9.5 ;
    RECT 212.61 9.765 212.82 9.835 ;
    RECT 212.15 2.585 212.36 2.795 ;
    RECT 212.15 5.86 212.36 6.07 ;
    RECT 212.15 6.385 212.36 6.455 ;
    RECT 212.15 7.28 212.36 7.35 ;
    RECT 293.7 3.235 293.91 3.445 ;
    RECT 293.7 5.33 293.91 5.54 ;
    RECT 293.7 9.12 293.91 9.33 ;
    RECT 293.27 4.845 293.34 4.915 ;
    RECT 293.27 9.43 293.34 9.5 ;
    RECT 292.29 9.765 292.5 9.835 ;
    RECT 291.83 2.585 292.04 2.795 ;
    RECT 291.83 5.86 292.04 6.07 ;
    RECT 291.83 6.385 292.04 6.455 ;
    RECT 291.83 7.28 292.04 7.35 ;
    RECT 210.7 3.235 210.91 3.445 ;
    RECT 210.7 5.33 210.91 5.54 ;
    RECT 210.7 9.12 210.91 9.33 ;
    RECT 210.27 4.845 210.34 4.915 ;
    RECT 210.27 9.43 210.34 9.5 ;
    RECT 209.29 9.765 209.5 9.835 ;
    RECT 208.83 2.585 209.04 2.795 ;
    RECT 208.83 5.86 209.04 6.07 ;
    RECT 208.83 6.385 209.04 6.455 ;
    RECT 208.83 7.28 209.04 7.35 ;
    RECT 290.38 3.235 290.59 3.445 ;
    RECT 290.38 5.33 290.59 5.54 ;
    RECT 290.38 9.12 290.59 9.33 ;
    RECT 289.95 4.845 290.02 4.915 ;
    RECT 289.95 9.43 290.02 9.5 ;
    RECT 288.97 9.765 289.18 9.835 ;
    RECT 288.51 2.585 288.72 2.795 ;
    RECT 288.51 5.86 288.72 6.07 ;
    RECT 288.51 6.385 288.72 6.455 ;
    RECT 288.51 7.28 288.72 7.35 ;
    RECT 207.38 3.235 207.59 3.445 ;
    RECT 207.38 5.33 207.59 5.54 ;
    RECT 207.38 9.12 207.59 9.33 ;
    RECT 206.95 4.845 207.02 4.915 ;
    RECT 206.95 9.43 207.02 9.5 ;
    RECT 205.97 9.765 206.18 9.835 ;
    RECT 205.51 2.585 205.72 2.795 ;
    RECT 205.51 5.86 205.72 6.07 ;
    RECT 205.51 6.385 205.72 6.455 ;
    RECT 205.51 7.28 205.72 7.35 ;
    RECT 287.06 3.235 287.27 3.445 ;
    RECT 287.06 5.33 287.27 5.54 ;
    RECT 287.06 9.12 287.27 9.33 ;
    RECT 286.63 4.845 286.7 4.915 ;
    RECT 286.63 9.43 286.7 9.5 ;
    RECT 285.65 9.765 285.86 9.835 ;
    RECT 285.19 2.585 285.4 2.795 ;
    RECT 285.19 5.86 285.4 6.07 ;
    RECT 285.19 6.385 285.4 6.455 ;
    RECT 285.19 7.28 285.4 7.35 ;
    RECT 283.74 3.235 283.95 3.445 ;
    RECT 283.74 5.33 283.95 5.54 ;
    RECT 283.74 9.12 283.95 9.33 ;
    RECT 283.31 4.845 283.38 4.915 ;
    RECT 283.31 9.43 283.38 9.5 ;
    RECT 282.33 9.765 282.54 9.835 ;
    RECT 281.87 2.585 282.08 2.795 ;
    RECT 281.87 5.86 282.08 6.07 ;
    RECT 281.87 6.385 282.08 6.455 ;
    RECT 281.87 7.28 282.08 7.35 ;
    RECT 280.42 3.235 280.63 3.445 ;
    RECT 280.42 5.33 280.63 5.54 ;
    RECT 280.42 9.12 280.63 9.33 ;
    RECT 279.99 4.845 280.06 4.915 ;
    RECT 279.99 9.43 280.06 9.5 ;
    RECT 279.01 9.765 279.22 9.835 ;
    RECT 278.55 2.585 278.76 2.795 ;
    RECT 278.55 5.86 278.76 6.07 ;
    RECT 278.55 6.385 278.76 6.455 ;
    RECT 278.55 7.28 278.76 7.35 ;
    RECT 277.1 3.235 277.31 3.445 ;
    RECT 277.1 5.33 277.31 5.54 ;
    RECT 277.1 9.12 277.31 9.33 ;
    RECT 276.67 4.845 276.74 4.915 ;
    RECT 276.67 9.43 276.74 9.5 ;
    RECT 275.69 9.765 275.9 9.835 ;
    RECT 275.23 2.585 275.44 2.795 ;
    RECT 275.23 5.86 275.44 6.07 ;
    RECT 275.23 6.385 275.44 6.455 ;
    RECT 275.23 7.28 275.44 7.35 ;
    RECT 273.78 3.235 273.99 3.445 ;
    RECT 273.78 5.33 273.99 5.54 ;
    RECT 273.78 9.12 273.99 9.33 ;
    RECT 273.35 4.845 273.42 4.915 ;
    RECT 273.35 9.43 273.42 9.5 ;
    RECT 272.37 9.765 272.58 9.835 ;
    RECT 271.91 2.585 272.12 2.795 ;
    RECT 271.91 5.86 272.12 6.07 ;
    RECT 271.91 6.385 272.12 6.455 ;
    RECT 271.91 7.28 272.12 7.35 ;
    RECT 270.46 3.235 270.67 3.445 ;
    RECT 270.46 5.33 270.67 5.54 ;
    RECT 270.46 9.12 270.67 9.33 ;
    RECT 270.03 4.845 270.1 4.915 ;
    RECT 270.03 9.43 270.1 9.5 ;
    RECT 269.05 9.765 269.26 9.835 ;
    RECT 268.59 2.585 268.8 2.795 ;
    RECT 268.59 5.86 268.8 6.07 ;
    RECT 268.59 6.385 268.8 6.455 ;
    RECT 268.59 7.28 268.8 7.35 ;
    RECT 239.66 4.055 239.87 4.125 ;
    RECT 249.62 5.86 249.83 6.07 ;
    RECT 349.22 5.86 349.43 6.07 ;
    RECT 249.62 2.585 249.83 2.795 ;
    RECT 335.94 7.28 336.15 7.35 ;
    RECT 349.22 2.585 349.43 2.795 ;
    RECT 335.94 6.385 336.15 6.455 ;
    RECT 335.94 5.86 336.15 6.07 ;
    RECT 335.94 2.585 336.15 2.795 ;
    RECT 220.66 4.455 220.87 4.525 ;
    RECT 299.42 7.28 299.63 7.35 ;
    RECT 299.42 6.385 299.63 6.455 ;
    RECT 209.78 7.28 209.99 7.35 ;
    RECT 336.86 4.455 337.07 4.525 ;
    RECT 209.78 6.385 209.99 6.455 ;
    RECT 267.14 3.235 267.35 3.445 ;
    RECT 267.14 5.33 267.35 5.54 ;
    RECT 267.14 9.12 267.35 9.33 ;
    RECT 266.71 4.845 266.78 4.915 ;
    RECT 266.71 9.43 266.78 9.5 ;
    RECT 265.73 9.765 265.94 9.835 ;
    RECT 265.27 2.585 265.48 2.795 ;
    RECT 265.27 5.86 265.48 6.07 ;
    RECT 265.27 6.385 265.48 6.455 ;
    RECT 265.27 7.28 265.48 7.35 ;
    RECT 209.78 5.86 209.99 6.07 ;
    RECT 243.9 4.455 244.11 4.525 ;
    RECT 263.82 3.235 264.03 3.445 ;
    RECT 263.82 5.33 264.03 5.54 ;
    RECT 263.82 9.12 264.03 9.33 ;
    RECT 263.39 4.845 263.46 4.915 ;
    RECT 263.39 9.43 263.46 9.5 ;
    RECT 262.41 9.765 262.62 9.835 ;
    RECT 261.95 2.585 262.16 2.795 ;
    RECT 261.95 5.86 262.16 6.07 ;
    RECT 261.95 6.385 262.16 6.455 ;
    RECT 261.95 7.28 262.16 7.35 ;
    RECT 209.78 2.585 209.99 2.795 ;
    RECT 260.5 3.235 260.71 3.445 ;
    RECT 260.5 5.33 260.71 5.54 ;
    RECT 260.5 9.12 260.71 9.33 ;
    RECT 260.07 4.845 260.14 4.915 ;
    RECT 260.07 9.43 260.14 9.5 ;
    RECT 259.09 9.765 259.3 9.835 ;
    RECT 258.63 2.585 258.84 2.795 ;
    RECT 258.63 5.86 258.84 6.07 ;
    RECT 258.63 6.385 258.84 6.455 ;
    RECT 258.63 7.28 258.84 7.35 ;
    RECT 365.82 4.055 366.03 4.125 ;
    RECT 257.18 3.235 257.39 3.445 ;
    RECT 257.18 5.33 257.39 5.54 ;
    RECT 257.18 9.12 257.39 9.33 ;
    RECT 256.75 4.845 256.82 4.915 ;
    RECT 256.75 9.43 256.82 9.5 ;
    RECT 255.77 9.765 255.98 9.835 ;
    RECT 255.31 2.585 255.52 2.795 ;
    RECT 255.31 5.86 255.52 6.07 ;
    RECT 255.31 6.385 255.52 6.455 ;
    RECT 255.31 7.28 255.52 7.35 ;
    RECT 253.86 3.235 254.07 3.445 ;
    RECT 253.86 5.33 254.07 5.54 ;
    RECT 253.86 9.12 254.07 9.33 ;
    RECT 253.43 4.845 253.5 4.915 ;
    RECT 253.43 9.43 253.5 9.5 ;
    RECT 252.45 9.765 252.66 9.835 ;
    RECT 251.99 2.585 252.2 2.795 ;
    RECT 251.99 5.86 252.2 6.07 ;
    RECT 251.99 6.385 252.2 6.455 ;
    RECT 251.99 7.28 252.2 7.35 ;
    RECT 229.7 4.055 229.91 4.125 ;
    RECT 250.54 3.235 250.75 3.445 ;
    RECT 250.54 5.33 250.75 5.54 ;
    RECT 250.54 9.12 250.75 9.33 ;
    RECT 250.11 4.845 250.18 4.915 ;
    RECT 250.11 9.43 250.18 9.5 ;
    RECT 249.13 9.765 249.34 9.835 ;
    RECT 248.67 2.585 248.88 2.795 ;
    RECT 248.67 5.86 248.88 6.07 ;
    RECT 248.67 6.385 248.88 6.455 ;
    RECT 248.67 7.28 248.88 7.35 ;
    RECT 247.22 3.235 247.43 3.445 ;
    RECT 247.22 5.33 247.43 5.54 ;
    RECT 247.22 9.12 247.43 9.33 ;
    RECT 246.79 4.845 246.86 4.915 ;
    RECT 246.79 9.43 246.86 9.5 ;
    RECT 245.81 9.765 246.02 9.835 ;
    RECT 245.35 2.585 245.56 2.795 ;
    RECT 245.35 5.86 245.56 6.07 ;
    RECT 245.35 6.385 245.56 6.455 ;
    RECT 245.35 7.28 245.56 7.35 ;
    RECT 243.9 3.235 244.11 3.445 ;
    RECT 243.9 5.33 244.11 5.54 ;
    RECT 243.9 9.12 244.11 9.33 ;
    RECT 243.47 4.845 243.54 4.915 ;
    RECT 243.47 9.43 243.54 9.5 ;
    RECT 242.49 9.765 242.7 9.835 ;
    RECT 242.03 2.585 242.24 2.795 ;
    RECT 242.03 5.86 242.24 6.07 ;
    RECT 242.03 6.385 242.24 6.455 ;
    RECT 242.03 7.28 242.24 7.35 ;
    RECT 240.58 3.235 240.79 3.445 ;
    RECT 240.58 5.33 240.79 5.54 ;
    RECT 240.58 9.12 240.79 9.33 ;
    RECT 240.15 4.845 240.22 4.915 ;
    RECT 240.15 9.43 240.22 9.5 ;
    RECT 239.17 9.765 239.38 9.835 ;
    RECT 238.71 2.585 238.92 2.795 ;
    RECT 238.71 5.86 238.92 6.07 ;
    RECT 238.71 6.385 238.92 6.455 ;
    RECT 238.71 7.28 238.92 7.35 ;
    RECT 237.26 3.235 237.47 3.445 ;
    RECT 237.26 5.33 237.47 5.54 ;
    RECT 237.26 9.12 237.47 9.33 ;
    RECT 236.83 4.845 236.9 4.915 ;
    RECT 236.83 9.43 236.9 9.5 ;
    RECT 235.85 9.765 236.06 9.835 ;
    RECT 235.39 2.585 235.6 2.795 ;
    RECT 235.39 5.86 235.6 6.07 ;
    RECT 235.39 6.385 235.6 6.455 ;
    RECT 235.39 7.28 235.6 7.35 ;
    RECT 300.34 4.455 300.55 4.525 ;
    RECT 236.34 4.055 236.55 4.125 ;
    RECT 246.3 7.28 246.51 7.35 ;
    RECT 246.3 6.385 246.51 6.455 ;
    RECT 246.3 5.86 246.51 6.07 ;
    RECT 299.42 5.86 299.63 6.07 ;
    RECT 246.3 2.585 246.51 2.795 ;
    RECT 299.42 2.585 299.63 2.795 ;
    RECT 217.34 4.455 217.55 4.525 ;
    RECT 362.5 4.055 362.71 4.125 ;
    RECT 240.58 4.455 240.79 4.525 ;
    RECT 226.38 4.055 226.59 4.125 ;
    RECT 297.02 4.455 297.23 4.525 ;
    RECT 296.1 7.28 296.31 7.35 ;
    RECT 242.98 7.28 243.19 7.35 ;
    RECT 296.1 6.385 296.31 6.455 ;
    RECT 242.98 6.385 243.19 6.455 ;
    RECT 206.46 7.28 206.67 7.35 ;
    RECT 296.1 5.86 296.31 6.07 ;
    RECT 242.98 5.86 243.19 6.07 ;
    RECT 206.46 6.385 206.67 6.455 ;
    RECT 296.1 2.585 296.31 2.795 ;
    RECT 242.98 2.585 243.19 2.795 ;
    RECT 206.46 5.86 206.67 6.07 ;
    RECT 206.46 2.585 206.67 2.795 ;
    RECT 214.02 4.455 214.23 4.525 ;
    RECT 359.18 4.055 359.39 4.125 ;
    RECT 299.42 4.055 299.63 4.125 ;
    RECT 223.06 4.055 223.27 4.125 ;
    RECT 237.26 4.455 237.47 4.525 ;
    RECT 293.7 4.455 293.91 4.525 ;
    RECT 292.78 7.28 292.99 7.35 ;
    RECT 292.78 6.385 292.99 6.455 ;
    RECT 203.14 7.28 203.35 7.35 ;
    RECT 292.78 5.86 292.99 6.07 ;
    RECT 203.14 6.385 203.35 6.455 ;
    RECT 292.78 2.585 292.99 2.795 ;
    RECT 332.62 7.28 332.83 7.35 ;
    RECT 203.14 5.86 203.35 6.07 ;
    RECT 332.62 6.385 332.83 6.455 ;
    RECT 203.14 2.585 203.35 2.795 ;
    RECT 355.86 4.055 356.07 4.125 ;
    RECT 296.1 4.055 296.31 4.125 ;
    RECT 219.74 4.055 219.95 4.125 ;
    RECT 373.38 3.235 373.59 3.445 ;
    RECT 373.38 5.33 373.59 5.54 ;
    RECT 373.38 9.12 373.59 9.33 ;
    RECT 372.95 4.845 373.02 4.915 ;
    RECT 372.95 9.43 373.02 9.5 ;
    RECT 371.97 9.765 372.18 9.835 ;
    RECT 371.51 2.585 371.72 2.795 ;
    RECT 371.51 5.86 371.72 6.07 ;
    RECT 371.51 6.385 371.72 6.455 ;
    RECT 371.51 7.28 371.72 7.35 ;
    RECT 239.66 7.28 239.87 7.35 ;
    RECT 239.66 6.385 239.87 6.455 ;
    RECT 239.66 5.86 239.87 6.07 ;
    RECT 239.66 2.585 239.87 2.795 ;
    RECT 204.06 3.235 204.27 3.445 ;
    RECT 204.06 5.33 204.27 5.54 ;
    RECT 204.06 9.12 204.27 9.33 ;
    RECT 203.63 4.845 203.7 4.915 ;
    RECT 203.63 9.43 203.7 9.5 ;
    RECT 202.65 9.765 202.86 9.835 ;
    RECT 202.19 2.585 202.4 2.795 ;
    RECT 202.19 5.86 202.4 6.07 ;
    RECT 202.19 6.385 202.4 6.455 ;
    RECT 202.19 7.28 202.4 7.35 ;
    RECT 332.62 5.86 332.83 6.07 ;
    RECT 332.62 2.585 332.83 2.795 ;
    RECT 290.38 4.455 290.59 4.525 ;
    RECT 277.1 4.455 277.31 4.525 ;
    RECT 333.54 4.455 333.75 4.525 ;
    RECT 210.7 4.455 210.91 4.525 ;
    RECT 352.54 4.055 352.75 4.125 ;
    RECT 292.78 4.055 292.99 4.125 ;
    RECT 216.42 4.055 216.63 4.125 ;
    RECT 289.46 7.28 289.67 7.35 ;
    RECT 236.34 7.28 236.55 7.35 ;
    RECT 289.46 6.385 289.67 6.455 ;
    RECT 236.34 6.385 236.55 6.455 ;
    RECT 289.46 5.86 289.67 6.07 ;
    RECT 236.34 5.86 236.55 6.07 ;
    RECT 289.46 2.585 289.67 2.795 ;
    RECT 329.3 7.28 329.51 7.35 ;
    RECT 236.34 2.585 236.55 2.795 ;
    RECT 329.3 6.385 329.51 6.455 ;
    RECT 329.3 5.86 329.51 6.07 ;
    RECT 329.3 2.585 329.51 2.795 ;
    RECT 273.78 4.455 273.99 4.525 ;
    RECT 330.22 4.455 330.43 4.525 ;
    RECT 207.38 4.455 207.59 4.525 ;
    RECT 349.22 4.055 349.43 4.125 ;
    RECT 289.46 4.055 289.67 4.125 ;
    RECT 213.1 4.055 213.31 4.125 ;
    RECT 287.06 4.455 287.27 4.525 ;
    RECT 286.14 7.28 286.35 7.35 ;
    RECT 286.14 6.385 286.35 6.455 ;
    RECT 286.14 5.86 286.35 6.07 ;
    RECT 325.98 7.28 326.19 7.35 ;
    RECT 286.14 2.585 286.35 2.795 ;
    RECT 325.98 6.385 326.19 6.455 ;
    RECT 325.98 5.86 326.19 6.07 ;
    RECT 325.98 2.585 326.19 2.795 ;
    RECT 270.46 4.455 270.67 4.525 ;
    RECT 326.9 4.455 327.11 4.525 ;
    RECT 204.06 4.455 204.27 4.525 ;
    RECT 345.9 4.055 346.11 4.125 ;
    RECT 286.14 4.055 286.35 4.125 ;
    RECT 209.78 4.055 209.99 4.125 ;
    RECT 372.46 7.28 372.67 7.35 ;
    RECT 372.46 6.385 372.67 6.455 ;
    RECT 372.46 5.86 372.67 6.07 ;
    RECT 372.46 2.585 372.67 2.795 ;
    RECT 283.74 4.455 283.95 4.525 ;
    RECT 282.82 7.28 283.03 7.35 ;
    RECT 282.82 6.385 283.03 6.455 ;
    RECT 323.58 4.455 323.79 4.525 ;
    RECT 342.58 4.055 342.79 4.125 ;
    RECT 282.82 4.055 283.03 4.125 ;
    RECT 206.46 4.055 206.67 4.125 ;
    RECT 282.82 5.86 283.03 6.07 ;
    RECT 282.82 2.585 283.03 2.795 ;
    RECT 322.66 7.28 322.87 7.35 ;
    RECT 322.66 6.385 322.87 6.455 ;
    RECT 369.14 7.28 369.35 7.35 ;
    RECT 322.66 5.86 322.87 6.07 ;
    RECT 369.14 6.385 369.35 6.455 ;
    RECT 322.66 2.585 322.87 2.795 ;
    RECT 369.14 5.86 369.35 6.07 ;
    RECT 280.42 4.455 280.63 4.525 ;
    RECT 369.14 2.585 369.35 2.795 ;
    RECT 366.74 4.455 366.95 4.525 ;
    RECT 332.62 4.055 332.83 4.125 ;
    RECT 373.38 4.455 373.59 4.525 ;
    RECT 339.26 4.055 339.47 4.125 ;
    RECT 279.5 4.055 279.71 4.125 ;
    RECT 203.14 4.055 203.35 4.125 ;
    RECT 279.5 7.28 279.71 7.35 ;
    RECT 279.5 6.385 279.71 6.455 ;
    RECT 279.5 5.86 279.71 6.07 ;
    RECT 279.5 2.585 279.71 2.795 ;
    RECT 319.34 7.28 319.55 7.35 ;
    RECT 319.34 6.385 319.55 6.455 ;
    RECT 319.34 5.86 319.55 6.07 ;
    RECT 319.34 2.585 319.55 2.795 ;
    RECT 363.42 4.455 363.63 4.525 ;
    RECT 329.3 4.055 329.51 4.125 ;
    RECT 233.02 7.28 233.23 7.35 ;
    RECT 233.02 6.385 233.23 6.455 ;
    RECT 370.06 4.455 370.27 4.525 ;
    RECT 320.26 4.455 320.47 4.525 ;
    RECT 335.94 4.055 336.15 4.125 ;
    RECT 276.18 4.055 276.39 4.125 ;
    RECT 276.18 7.28 276.39 7.35 ;
    RECT 276.18 6.385 276.39 6.455 ;
    RECT 276.18 5.86 276.39 6.07 ;
    RECT 276.18 2.585 276.39 2.795 ;
    RECT 316.02 7.28 316.23 7.35 ;
    RECT 316.02 6.385 316.23 6.455 ;
    RECT 233.02 5.86 233.23 6.07 ;
    RECT 233.02 2.585 233.23 2.795 ;
    RECT 325.98 4.055 326.19 4.125 ;
    RECT 360.1 4.455 360.31 4.525 ;
    RECT 266.22 4.055 266.43 4.125 ;
    RECT 267.14 4.455 267.35 4.525 ;
    RECT 316.94 4.455 317.15 4.525 ;
    RECT 316.02 5.86 316.23 6.07 ;
    RECT 316.02 2.585 316.23 2.795 ;
    RECT 272.86 4.055 273.07 4.125 ;
    RECT 266.22 7.28 266.43 7.35 ;
    RECT 266.22 6.385 266.43 6.455 ;
    RECT 365.82 7.28 366.03 7.35 ;
    RECT 229.7 7.28 229.91 7.35 ;
    RECT 365.82 6.385 366.03 6.455 ;
    RECT 229.7 6.385 229.91 6.455 ;
    RECT 229.7 5.86 229.91 6.07 ;
    RECT 229.7 2.585 229.91 2.795 ;
    RECT 322.66 4.055 322.87 4.125 ;
    RECT 262.9 4.055 263.11 4.125 ;
    RECT 356.78 4.455 356.99 4.525 ;
    RECT 263.82 4.455 264.03 4.525 ;
    RECT 266.22 5.86 266.43 6.07 ;
    RECT 266.22 2.585 266.43 2.795 ;
    RECT 272.86 7.28 273.07 7.35 ;
    RECT 272.86 6.385 273.07 6.455 ;
    RECT 313.62 4.455 313.83 4.525 ;
    RECT 272.86 5.86 273.07 6.07 ;
    RECT 272.86 2.585 273.07 2.795 ;
    RECT 312.7 7.28 312.91 7.35 ;
    RECT 269.54 4.055 269.75 4.125 ;
    RECT 312.7 6.385 312.91 6.455 ;
    RECT 312.7 5.86 312.91 6.07 ;
    RECT 365.82 5.86 366.03 6.07 ;
    RECT 312.7 2.585 312.91 2.795 ;
    RECT 365.82 2.585 366.03 2.795 ;
    RECT 226.38 7.28 226.59 7.35 ;
    RECT 226.38 6.385 226.59 6.455 ;
    RECT 319.34 4.055 319.55 4.125 ;
    RECT 226.38 5.86 226.59 6.07 ;
    RECT 259.58 4.055 259.79 4.125 ;
    RECT 226.38 2.585 226.59 2.795 ;
    RECT 260.5 4.455 260.71 4.525 ;
    RECT 262.9 7.28 263.11 7.35 ;
    RECT 262.9 6.385 263.11 6.455 ;
    RECT 262.9 5.86 263.11 6.07 ;
    RECT 262.9 2.585 263.11 2.795 ;
    RECT 269.54 7.28 269.75 7.35 ;
    RECT 269.54 6.385 269.75 6.455 ;
    RECT 269.54 5.86 269.75 6.07 ;
    RECT 309.38 7.28 309.59 7.35 ;
    RECT 269.54 2.585 269.75 2.795 ;
    RECT 362.5 7.28 362.71 7.35 ;
    RECT 309.38 6.385 309.59 6.455 ;
    RECT 362.5 6.385 362.71 6.455 ;
    RECT 309.38 5.86 309.59 6.07 ;
    RECT 362.5 5.86 362.71 6.07 ;
    RECT 309.38 2.585 309.59 2.795 ;
    RECT 362.5 2.585 362.71 2.795 ;
    RECT 353.46 4.455 353.67 4.525 ;
    RECT 316.02 4.055 316.23 4.125 ;
    RECT 256.26 4.055 256.47 4.125 ;
    RECT 310.3 4.455 310.51 4.525 ;
    RECT 257.18 4.455 257.39 4.525 ;
    RECT 259.58 7.28 259.79 7.35 ;
    RECT 259.58 6.385 259.79 6.455 ;
    RECT 259.58 5.86 259.79 6.07 ;
    RECT 259.58 2.585 259.79 2.795 ;
    RECT 233.94 4.455 234.15 4.525 ;
    RECT 359.18 7.28 359.39 7.35 ;
    RECT 223.06 7.28 223.27 7.35 ;
    RECT 359.18 6.385 359.39 6.455 ;
    RECT 223.06 6.385 223.27 6.455 ;
    RECT 359.18 5.86 359.39 6.07 ;
    RECT 223.06 5.86 223.27 6.07 ;
    RECT 359.18 2.585 359.39 2.795 ;
    RECT 223.06 2.585 223.27 2.795 ;
    RECT 350.14 4.455 350.35 4.525 ;
    RECT 345.9 7.28 346.11 7.35 ;
    RECT 372.46 4.055 372.67 4.125 ;
    RECT 345.9 6.385 346.11 6.455 ;
    RECT 312.7 4.055 312.91 4.125 ;
    RECT 345.9 5.86 346.11 6.07 ;
    RECT 252.94 4.055 253.15 4.125 ;
    RECT 345.9 2.585 346.11 2.795 ;
    RECT 306.98 4.455 307.19 4.525 ;
    RECT 306.06 7.28 306.27 7.35 ;
    RECT 306.06 6.385 306.27 6.455 ;
    RECT 306.06 5.86 306.27 6.07 ;
    RECT 306.06 2.585 306.27 2.795 ;
    RECT 230.62 4.455 230.83 4.525 ;
    RECT 219.74 7.28 219.95 7.35 ;
    RECT 219.74 6.385 219.95 6.455 ;
    RECT 219.74 5.86 219.95 6.07 ;
    RECT 219.74 2.585 219.95 2.795 ;
    RECT 346.82 4.455 347.03 4.525 ;
    RECT 253.86 4.455 254.07 4.525 ;
    RECT 369.14 4.055 369.35 4.125 ;
    RECT 309.38 4.055 309.59 4.125 ;
    RECT 249.62 4.055 249.83 4.125 ;
    RECT 342.58 7.28 342.79 7.35 ;
    RECT 342.58 6.385 342.79 6.455 ;
    RECT 342.58 5.86 342.79 6.07 ;
    RECT 342.58 2.585 342.79 2.795 ;
    RECT 303.66 4.455 303.87 4.525 ;
    RECT 256.26 7.28 256.47 7.35 ;
    RECT 302.74 7.28 302.95 7.35 ;
    RECT 256.26 6.385 256.47 6.455 ;
    RECT 355.86 7.28 356.07 7.35 ;
    RECT 302.74 6.385 302.95 6.455 ;
    RECT 256.26 5.86 256.47 6.07 ;
    RECT 355.86 6.385 356.07 6.455 ;
    RECT 370.06 3.235 370.27 3.445 ;
    RECT 370.06 5.33 370.27 5.54 ;
    RECT 370.06 9.12 370.27 9.33 ;
    RECT 369.63 4.845 369.7 4.915 ;
    RECT 369.63 9.43 369.7 9.5 ;
    RECT 368.65 9.765 368.86 9.835 ;
    RECT 368.19 2.585 368.4 2.795 ;
    RECT 368.19 5.86 368.4 6.07 ;
    RECT 368.19 6.385 368.4 6.455 ;
    RECT 368.19 7.28 368.4 7.35 ;
    RECT 302.74 5.86 302.95 6.07 ;
    RECT 256.26 2.585 256.47 2.795 ;
    RECT 355.86 5.86 356.07 6.07 ;
    RECT 302.74 2.585 302.95 2.795 ;
    RECT 355.86 2.585 356.07 2.795 ;
    RECT 316.02 0.915 316.23 1.125 ;
    RECT 362.5 2.055 362.71 2.125 ;
    RECT 362.5 1.742 362.71 1.812 ;
    RECT 311.75 1.24 311.96 1.31 ;
    RECT 362.5 0.915 362.71 1.125 ;
    RECT 358.23 1.24 358.44 1.31 ;
    RECT 312.7 2.055 312.91 2.125 ;
    RECT 312.7 1.742 312.91 1.812 ;
    RECT 312.7 0.915 312.91 1.125 ;
    RECT 359.18 2.055 359.39 2.125 ;
    RECT 359.18 1.742 359.39 1.812 ;
    RECT 308.43 1.24 308.64 1.31 ;
    RECT 359.18 0.915 359.39 1.125 ;
    RECT 354.91 1.24 355.12 1.31 ;
    RECT 355.86 2.055 356.07 2.125 ;
    RECT 355.86 1.742 356.07 1.812 ;
    RECT 355.86 0.915 356.07 1.125 ;
    RECT 226.38 2.055 226.59 2.125 ;
    RECT 226.38 1.742 226.59 1.812 ;
    RECT 226.38 0.915 226.59 1.125 ;
    RECT 351.59 1.24 351.8 1.31 ;
    RECT 352.54 2.055 352.75 2.125 ;
    RECT 352.54 1.742 352.75 1.812 ;
    RECT 371.51 1.24 371.72 1.31 ;
    RECT 372.46 2.055 372.67 2.125 ;
    RECT 372.46 1.742 372.67 1.812 ;
    RECT 222.11 1.24 222.32 1.31 ;
    RECT 372.46 0.915 372.67 1.125 ;
    RECT 223.06 2.055 223.27 2.125 ;
    RECT 223.06 1.742 223.27 1.812 ;
    RECT 223.06 0.915 223.27 1.125 ;
    RECT 352.54 0.915 352.75 1.125 ;
    RECT 348.27 1.24 348.48 1.31 ;
    RECT 349.22 2.055 349.43 2.125 ;
    RECT 349.22 1.742 349.43 1.812 ;
    RECT 368.19 1.24 368.4 1.31 ;
    RECT 369.14 2.055 369.35 2.125 ;
    RECT 369.14 1.742 369.35 1.812 ;
    RECT 218.79 1.24 219.0 1.31 ;
    RECT 219.74 2.055 219.95 2.125 ;
    RECT 219.74 1.742 219.95 1.812 ;
    RECT 349.22 0.915 349.43 1.125 ;
    RECT 369.14 0.915 369.35 1.125 ;
    RECT 219.74 0.915 219.95 1.125 ;
    RECT 215.47 1.24 215.68 1.31 ;
    RECT 216.42 2.055 216.63 2.125 ;
    RECT 216.42 1.742 216.63 1.812 ;
    RECT 251.99 1.24 252.2 1.31 ;
    RECT 252.94 2.055 253.15 2.125 ;
    RECT 252.94 1.742 253.15 1.812 ;
    RECT 216.42 0.915 216.63 1.125 ;
    RECT 252.94 0.915 253.15 1.125 ;
    RECT 212.15 1.24 212.36 1.31 ;
    RECT 248.67 1.24 248.88 1.31 ;
    RECT 249.62 2.055 249.83 2.125 ;
    RECT 249.62 1.742 249.83 1.812 ;
    RECT 213.1 2.055 213.31 2.125 ;
    RECT 213.1 1.742 213.31 1.812 ;
    RECT 213.1 0.915 213.31 1.125 ;
    RECT 249.62 0.915 249.83 1.125 ;
    RECT 208.83 1.24 209.04 1.31 ;
    RECT 245.35 1.24 245.56 1.31 ;
    RECT 209.78 2.055 209.99 2.125 ;
    RECT 209.78 1.742 209.99 1.812 ;
    RECT 209.78 0.915 209.99 1.125 ;
    RECT 246.3 2.055 246.51 2.125 ;
    RECT 246.3 1.742 246.51 1.812 ;
    RECT 246.3 0.915 246.51 1.125 ;
    RECT 242.03 1.24 242.24 1.31 ;
    RECT 205.51 1.24 205.72 1.31 ;
    RECT 206.46 2.055 206.67 2.125 ;
    RECT 206.46 1.742 206.67 1.812 ;
    RECT 206.46 0.915 206.67 1.125 ;
    RECT 242.98 2.055 243.19 2.125 ;
    RECT 242.98 1.742 243.19 1.812 ;
    RECT 242.98 0.915 243.19 1.125 ;
    RECT 309.38 2.055 309.59 2.125 ;
    RECT 309.38 1.742 309.59 1.812 ;
    RECT 309.38 0.915 309.59 1.125 ;
    RECT 202.19 1.24 202.4 1.31 ;
    RECT 203.14 2.055 203.35 2.125 ;
    RECT 203.14 1.742 203.35 1.812 ;
    RECT 238.71 1.24 238.92 1.31 ;
    RECT 239.66 2.055 239.87 2.125 ;
    RECT 239.66 1.742 239.87 1.812 ;
    RECT 239.66 0.915 239.87 1.125 ;
    RECT 203.14 0.915 203.35 1.125 ;
    RECT 305.11 1.24 305.32 1.31 ;
    RECT 306.06 2.055 306.27 2.125 ;
    RECT 306.06 1.742 306.27 1.812 ;
    RECT 306.06 0.915 306.27 1.125 ;
    RECT 235.39 1.24 235.6 1.31 ;
    RECT 236.34 2.055 236.55 2.125 ;
    RECT 236.34 1.742 236.55 1.812 ;
    RECT 301.79 1.24 302.0 1.31 ;
    RECT 302.74 2.055 302.95 2.125 ;
    RECT 302.74 1.742 302.95 1.812 ;
    RECT 236.34 0.915 236.55 1.125 ;
    RECT 364.87 1.24 365.08 1.31 ;
    RECT 365.82 2.055 366.03 2.125 ;
    RECT 365.82 1.742 366.03 1.812 ;
    RECT 282.82 0.915 283.03 1.125 ;
    RECT 302.74 0.915 302.95 1.125 ;
    RECT 278.55 1.24 278.76 1.31 ;
    RECT 279.5 2.055 279.71 2.125 ;
    RECT 279.5 1.742 279.71 1.812 ;
    RECT 279.5 0.915 279.71 1.125 ;
    RECT 334.99 1.24 335.2 1.31 ;
    RECT 232.07 1.24 232.28 1.31 ;
    RECT 335.94 2.055 336.15 2.125 ;
    RECT 335.94 1.742 336.15 1.812 ;
    RECT 233.02 2.055 233.23 2.125 ;
    RECT 233.02 1.742 233.23 1.812 ;
    RECT 275.23 1.24 275.44 1.31 ;
    RECT 335.94 0.915 336.15 1.125 ;
    RECT 233.02 0.915 233.23 1.125 ;
    RECT 370.06 1.41 370.27 1.62 ;
    RECT 369.63 1.005 369.9 2.125 ;
    RECT 369.14 1.24 369.35 1.31 ;
    RECT 368.19 0.915 368.4 2.125 ;
    RECT 276.18 2.055 276.39 2.125 ;
    RECT 276.18 1.742 276.39 1.812 ;
    RECT 276.18 0.915 276.39 1.125 ;
    RECT 228.75 1.24 228.96 1.31 ;
    RECT 366.74 1.41 366.95 1.62 ;
    RECT 366.31 1.005 366.58 2.125 ;
    RECT 365.82 1.24 366.03 1.31 ;
    RECT 364.87 0.915 365.08 2.125 ;
    RECT 363.42 1.41 363.63 1.62 ;
    RECT 362.99 1.005 363.26 2.125 ;
    RECT 362.5 1.24 362.71 1.31 ;
    RECT 361.55 0.915 361.76 2.125 ;
    RECT 265.27 1.24 265.48 1.31 ;
    RECT 360.1 1.41 360.31 1.62 ;
    RECT 359.67 1.005 359.94 2.125 ;
    RECT 359.18 1.24 359.39 1.31 ;
    RECT 358.23 0.915 358.44 2.125 ;
    RECT 356.78 1.41 356.99 1.62 ;
    RECT 356.35 1.005 356.62 2.125 ;
    RECT 355.86 1.24 356.07 1.31 ;
    RECT 354.91 0.915 355.12 2.125 ;
    RECT 353.46 1.41 353.67 1.62 ;
    RECT 353.03 1.005 353.3 2.125 ;
    RECT 352.54 1.24 352.75 1.31 ;
    RECT 351.59 0.915 351.8 2.125 ;
    RECT 266.22 2.055 266.43 2.125 ;
    RECT 350.14 1.41 350.35 1.62 ;
    RECT 349.71 1.005 349.98 2.125 ;
    RECT 349.22 1.24 349.43 1.31 ;
    RECT 348.27 0.915 348.48 2.125 ;
    RECT 266.22 1.742 266.43 1.812 ;
    RECT 346.82 1.41 347.03 1.62 ;
    RECT 346.39 1.005 346.66 2.125 ;
    RECT 345.9 1.24 346.11 1.31 ;
    RECT 344.95 0.915 345.16 2.125 ;
    RECT 343.5 1.41 343.71 1.62 ;
    RECT 343.07 1.005 343.34 2.125 ;
    RECT 342.58 1.24 342.79 1.31 ;
    RECT 341.63 0.915 341.84 2.125 ;
    RECT 340.18 1.41 340.39 1.62 ;
    RECT 339.75 1.005 340.02 2.125 ;
    RECT 339.26 1.24 339.47 1.31 ;
    RECT 338.31 0.915 338.52 2.125 ;
    RECT 336.86 1.41 337.07 1.62 ;
    RECT 336.43 1.005 336.7 2.125 ;
    RECT 335.94 1.24 336.15 1.31 ;
    RECT 334.99 0.915 335.2 2.125 ;
    RECT 229.7 2.055 229.91 2.125 ;
    RECT 229.7 1.742 229.91 1.812 ;
    RECT 229.7 0.915 229.91 1.125 ;
    RECT 266.22 0.915 266.43 1.125 ;
    RECT 333.54 1.41 333.75 1.62 ;
    RECT 333.11 1.005 333.38 2.125 ;
    RECT 332.62 1.24 332.83 1.31 ;
    RECT 331.67 0.915 331.88 2.125 ;
    RECT 271.91 1.24 272.12 1.31 ;
    RECT 330.22 1.41 330.43 1.62 ;
    RECT 329.79 1.005 330.06 2.125 ;
    RECT 329.3 1.24 329.51 1.31 ;
    RECT 328.35 0.915 328.56 2.125 ;
    RECT 326.9 1.41 327.11 1.62 ;
    RECT 326.47 1.005 326.74 2.125 ;
    RECT 325.98 1.24 326.19 1.31 ;
    RECT 325.03 0.915 325.24 2.125 ;
    RECT 323.58 1.41 323.79 1.62 ;
    RECT 323.15 1.005 323.42 2.125 ;
    RECT 322.66 1.24 322.87 1.31 ;
    RECT 321.71 0.915 321.92 2.125 ;
    RECT 272.86 2.055 273.07 2.125 ;
    RECT 320.26 1.41 320.47 1.62 ;
    RECT 319.83 1.005 320.1 2.125 ;
    RECT 319.34 1.24 319.55 1.31 ;
    RECT 318.39 0.915 318.6 2.125 ;
    RECT 272.86 1.742 273.07 1.812 ;
    RECT 316.94 1.41 317.15 1.62 ;
    RECT 316.51 1.005 316.78 2.125 ;
    RECT 316.02 1.24 316.23 1.31 ;
    RECT 315.07 0.915 315.28 2.125 ;
    RECT 313.62 1.41 313.83 1.62 ;
    RECT 313.19 1.005 313.46 2.125 ;
    RECT 312.7 1.24 312.91 1.31 ;
    RECT 311.75 0.915 311.96 2.125 ;
    RECT 310.3 1.41 310.51 1.62 ;
    RECT 309.87 1.005 310.14 2.125 ;
    RECT 309.38 1.24 309.59 1.31 ;
    RECT 308.43 0.915 308.64 2.125 ;
    RECT 306.98 1.41 307.19 1.62 ;
    RECT 306.55 1.005 306.82 2.125 ;
    RECT 306.06 1.24 306.27 1.31 ;
    RECT 305.11 0.915 305.32 2.125 ;
    RECT 272.86 0.915 273.07 1.125 ;
    RECT 303.66 1.41 303.87 1.62 ;
    RECT 303.23 1.005 303.5 2.125 ;
    RECT 302.74 1.24 302.95 1.31 ;
    RECT 301.79 0.915 302.0 2.125 ;
    RECT 225.43 1.24 225.64 1.31 ;
    RECT 261.95 1.24 262.16 1.31 ;
    RECT 300.34 1.41 300.55 1.62 ;
    RECT 299.91 1.005 300.18 2.125 ;
    RECT 299.42 1.24 299.63 1.31 ;
    RECT 298.47 0.915 298.68 2.125 ;
    RECT 297.02 1.41 297.23 1.62 ;
    RECT 296.59 1.005 296.86 2.125 ;
    RECT 296.1 1.24 296.31 1.31 ;
    RECT 295.15 0.915 295.36 2.125 ;
    RECT 293.7 1.41 293.91 1.62 ;
    RECT 293.27 1.005 293.54 2.125 ;
    RECT 292.78 1.24 292.99 1.31 ;
    RECT 291.83 0.915 292.04 2.125 ;
    RECT 290.38 1.41 290.59 1.62 ;
    RECT 289.95 1.005 290.22 2.125 ;
    RECT 289.46 1.24 289.67 1.31 ;
    RECT 288.51 0.915 288.72 2.125 ;
    RECT 287.06 1.41 287.27 1.62 ;
    RECT 286.63 1.005 286.9 2.125 ;
    RECT 286.14 1.24 286.35 1.31 ;
    RECT 285.19 0.915 285.4 2.125 ;
    RECT 283.74 1.41 283.95 1.62 ;
    RECT 283.31 1.005 283.58 2.125 ;
    RECT 282.82 1.24 283.03 1.31 ;
    RECT 281.87 0.915 282.08 2.125 ;
    RECT 280.42 1.41 280.63 1.62 ;
    RECT 279.99 1.005 280.26 2.125 ;
    RECT 279.5 1.24 279.71 1.31 ;
    RECT 278.55 0.915 278.76 2.125 ;
    RECT 277.1 1.41 277.31 1.62 ;
    RECT 276.67 1.005 276.94 2.125 ;
    RECT 276.18 1.24 276.39 1.31 ;
    RECT 275.23 0.915 275.44 2.125 ;
    RECT 273.78 1.41 273.99 1.62 ;
    RECT 273.35 1.005 273.62 2.125 ;
    RECT 272.86 1.24 273.07 1.31 ;
    RECT 271.91 0.915 272.12 2.125 ;
    RECT 270.46 1.41 270.67 1.62 ;
    RECT 270.03 1.005 270.3 2.125 ;
    RECT 269.54 1.24 269.75 1.31 ;
    RECT 268.59 0.915 268.8 2.125 ;
    RECT 262.9 2.055 263.11 2.125 ;
    RECT 262.9 1.742 263.11 1.812 ;
    RECT 262.9 0.915 263.11 1.125 ;
    RECT 268.59 1.24 268.8 1.31 ;
    RECT 269.54 2.055 269.75 2.125 ;
    RECT 269.54 1.742 269.75 1.812 ;
    RECT 267.14 1.41 267.35 1.62 ;
    RECT 266.71 1.005 266.98 2.125 ;
    RECT 266.22 1.24 266.43 1.31 ;
    RECT 265.27 0.915 265.48 2.125 ;
    RECT 263.82 1.41 264.03 1.62 ;
    RECT 263.39 1.005 263.66 2.125 ;
    RECT 262.9 1.24 263.11 1.31 ;
    RECT 261.95 0.915 262.16 2.125 ;
    RECT 260.5 1.41 260.71 1.62 ;
    RECT 260.07 1.005 260.34 2.125 ;
    RECT 259.58 1.24 259.79 1.31 ;
    RECT 258.63 0.915 258.84 2.125 ;
    RECT 257.18 1.41 257.39 1.62 ;
    RECT 256.75 1.005 257.02 2.125 ;
    RECT 256.26 1.24 256.47 1.31 ;
    RECT 255.31 0.915 255.52 2.125 ;
    RECT 253.86 1.41 254.07 1.62 ;
    RECT 253.43 1.005 253.7 2.125 ;
    RECT 252.94 1.24 253.15 1.31 ;
    RECT 251.99 0.915 252.2 2.125 ;
    RECT 258.63 1.24 258.84 1.31 ;
    RECT 250.54 1.41 250.75 1.62 ;
    RECT 250.11 1.005 250.38 2.125 ;
    RECT 249.62 1.24 249.83 1.31 ;
    RECT 248.67 0.915 248.88 2.125 ;
    RECT 247.22 1.41 247.43 1.62 ;
    RECT 246.79 1.005 247.06 2.125 ;
    RECT 246.3 1.24 246.51 1.31 ;
    RECT 245.35 0.915 245.56 2.125 ;
    RECT 243.9 1.41 244.11 1.62 ;
    RECT 243.47 1.005 243.74 2.125 ;
    RECT 242.98 1.24 243.19 1.31 ;
    RECT 242.03 0.915 242.24 2.125 ;
    RECT 240.58 1.41 240.79 1.62 ;
    RECT 240.15 1.005 240.42 2.125 ;
    RECT 239.66 1.24 239.87 1.31 ;
    RECT 238.71 0.915 238.92 2.125 ;
    RECT 237.26 1.41 237.47 1.62 ;
    RECT 236.83 1.005 237.1 2.125 ;
    RECT 236.34 1.24 236.55 1.31 ;
    RECT 235.39 0.915 235.6 2.125 ;
    RECT 269.54 0.915 269.75 1.125 ;
    RECT 259.58 2.055 259.79 2.125 ;
    RECT 259.58 1.742 259.79 1.812 ;
    RECT 259.58 0.915 259.79 1.125 ;
    RECT 255.31 1.24 255.52 1.31 ;
    RECT 256.26 2.055 256.47 2.125 ;
    RECT 256.26 1.742 256.47 1.812 ;
    RECT 256.26 0.915 256.47 1.125 ;
    RECT 373.38 1.41 373.59 1.62 ;
    RECT 372.95 1.005 373.22 2.125 ;
    RECT 372.46 1.24 372.67 1.31 ;
    RECT 371.51 0.915 371.72 2.125 ;
    RECT 298.47 1.24 298.68 1.31 ;
    RECT 204.06 1.41 204.27 1.62 ;
    RECT 203.63 1.005 203.9 2.125 ;
    RECT 203.14 1.24 203.35 1.31 ;
    RECT 202.19 0.915 202.4 2.125 ;
    RECT 299.42 2.055 299.63 2.125 ;
    RECT 299.42 1.742 299.63 1.812 ;
    RECT 233.94 1.41 234.15 1.62 ;
    RECT 233.51 1.005 233.78 2.125 ;
    RECT 233.02 1.24 233.23 1.31 ;
    RECT 232.07 0.915 232.28 2.125 ;
    RECT 230.62 1.41 230.83 1.62 ;
    RECT 230.19 1.005 230.46 2.125 ;
    RECT 229.7 1.24 229.91 1.31 ;
    RECT 228.75 0.915 228.96 2.125 ;
    RECT 227.3 1.41 227.51 1.62 ;
    RECT 226.87 1.005 227.14 2.125 ;
    RECT 226.38 1.24 226.59 1.31 ;
    RECT 225.43 0.915 225.64 2.125 ;
    RECT 223.98 1.41 224.19 1.62 ;
    RECT 223.55 1.005 223.82 2.125 ;
    RECT 223.06 1.24 223.27 1.31 ;
    RECT 222.11 0.915 222.32 2.125 ;
    RECT 220.66 1.41 220.87 1.62 ;
    RECT 220.23 1.005 220.5 2.125 ;
    RECT 219.74 1.24 219.95 1.31 ;
    RECT 218.79 0.915 219.0 2.125 ;
    RECT 217.34 1.41 217.55 1.62 ;
    RECT 216.91 1.005 217.18 2.125 ;
    RECT 216.42 1.24 216.63 1.31 ;
    RECT 215.47 0.915 215.68 2.125 ;
    RECT 214.02 1.41 214.23 1.62 ;
    RECT 213.59 1.005 213.86 2.125 ;
    RECT 213.1 1.24 213.31 1.31 ;
    RECT 212.15 0.915 212.36 2.125 ;
    RECT 210.7 1.41 210.91 1.62 ;
    RECT 210.27 1.005 210.54 2.125 ;
    RECT 209.78 1.24 209.99 1.31 ;
    RECT 208.83 0.915 209.04 2.125 ;
    RECT 207.38 1.41 207.59 1.62 ;
    RECT 206.95 1.005 207.22 2.125 ;
    RECT 206.46 1.24 206.67 1.31 ;
    RECT 205.51 0.915 205.72 2.125 ;
    RECT 299.42 0.915 299.63 1.125 ;
    RECT 295.15 1.24 295.36 1.31 ;
    RECT 296.1 2.055 296.31 2.125 ;
    RECT 296.1 1.742 296.31 1.812 ;
    RECT 331.67 1.24 331.88 1.31 ;
    RECT 296.1 0.915 296.31 1.125 ;
    RECT 332.62 2.055 332.83 2.125 ;
    RECT 332.62 1.742 332.83 1.812 ;
    RECT 291.83 1.24 292.04 1.31 ;
    RECT 332.62 0.915 332.83 1.125 ;
    RECT 292.78 2.055 292.99 2.125 ;
    RECT 292.78 1.742 292.99 1.812 ;
    RECT 328.35 1.24 328.56 1.31 ;
    RECT 292.78 0.915 292.99 1.125 ;
    RECT 329.3 2.055 329.51 2.125 ;
    RECT 329.3 1.742 329.51 1.812 ;
    RECT 329.3 0.915 329.51 1.125 ;
    RECT 288.51 1.24 288.72 1.31 ;
    RECT 289.46 2.055 289.67 2.125 ;
    RECT 289.46 1.742 289.67 1.812 ;
    RECT 325.03 1.24 325.24 1.31 ;
    RECT 289.46 0.915 289.67 1.125 ;
    RECT 344.95 1.24 345.16 1.31 ;
    RECT 325.98 2.055 326.19 2.125 ;
    RECT 325.98 1.742 326.19 1.812 ;
    RECT 345.9 2.055 346.11 2.125 ;
    RECT 345.9 1.742 346.11 1.812 ;
    RECT 325.98 0.915 326.19 1.125 ;
    RECT 345.9 0.915 346.11 1.125 ;
    RECT 285.19 1.24 285.4 1.31 ;
    RECT 286.14 2.055 286.35 2.125 ;
    RECT 286.14 1.742 286.35 1.812 ;
    RECT 341.63 1.24 341.84 1.31 ;
    RECT 321.71 1.24 321.92 1.31 ;
    RECT 286.14 0.915 286.35 1.125 ;
    RECT 322.66 2.055 322.87 2.125 ;
    RECT 322.66 1.742 322.87 1.812 ;
    RECT 342.58 2.055 342.79 2.125 ;
    RECT 342.58 1.742 342.79 1.812 ;
    RECT 322.66 0.915 322.87 1.125 ;
    RECT 342.58 0.915 342.79 1.125 ;
    RECT 281.87 1.24 282.08 1.31 ;
    RECT 282.82 2.055 283.03 2.125 ;
    RECT 282.82 1.742 283.03 1.812 ;
    RECT 318.39 1.24 318.6 1.31 ;
    RECT 319.34 2.055 319.55 2.125 ;
    RECT 338.31 1.24 338.52 1.31 ;
    RECT 319.34 1.742 319.55 1.812 ;
    RECT 339.26 2.055 339.47 2.125 ;
    RECT 339.26 1.742 339.47 1.812 ;
    RECT 339.26 0.915 339.47 1.125 ;
    RECT 319.34 0.915 319.55 1.125 ;
    RECT 315.07 1.24 315.28 1.31 ;
    RECT 365.82 0.915 366.03 1.125 ;
    RECT 316.02 2.055 316.23 2.125 ;
    RECT 316.02 1.742 316.23 1.812 ;
    RECT 361.55 1.24 361.76 1.31 ;
    RECT 245.81 10.805 246.02 10.875 ;
    RECT 222.57 11.065 222.78 11.135 ;
    RECT 355.37 10.805 355.58 10.875 ;
    RECT 342.58 11.325 342.79 11.395 ;
    RECT 322.17 11.065 322.38 11.135 ;
    RECT 295.61 10.805 295.82 10.875 ;
    RECT 343.04 11.325 343.25 11.395 ;
    RECT 262.41 11.065 262.62 11.135 ;
    RECT 305.57 10.805 305.78 10.875 ;
    RECT 286.14 11.325 286.35 11.395 ;
    RECT 286.6 11.325 286.81 11.395 ;
    RECT 242.49 10.805 242.7 10.875 ;
    RECT 216.42 11.325 216.63 11.395 ;
    RECT 216.88 11.325 217.09 11.395 ;
    RECT 332.62 11.325 332.83 11.395 ;
    RECT 333.08 11.325 333.29 11.395 ;
    RECT 352.05 10.805 352.26 10.875 ;
    RECT 292.29 10.805 292.5 10.875 ;
    RECT 339.26 11.325 339.47 11.395 ;
    RECT 259.09 11.065 259.3 11.135 ;
    RECT 339.72 11.325 339.93 11.395 ;
    RECT 302.25 10.805 302.46 10.875 ;
    RECT 219.25 11.065 219.46 11.135 ;
    RECT 213.1 11.325 213.31 11.395 ;
    RECT 213.56 11.325 213.77 11.395 ;
    RECT 318.85 11.065 319.06 11.135 ;
    RECT 329.3 11.325 329.51 11.395 ;
    RECT 329.76 11.325 329.97 11.395 ;
    RECT 282.82 11.325 283.03 11.395 ;
    RECT 283.28 11.325 283.49 11.395 ;
    RECT 348.73 10.805 348.94 10.875 ;
    RECT 288.97 10.805 289.18 10.875 ;
    RECT 255.77 11.065 255.98 11.135 ;
    RECT 335.94 11.325 336.15 11.395 ;
    RECT 336.4 11.325 336.61 11.395 ;
    RECT 239.17 10.805 239.38 10.875 ;
    RECT 215.93 11.065 216.14 11.135 ;
    RECT 365.33 11.065 365.54 11.135 ;
    RECT 209.78 11.325 209.99 11.395 ;
    RECT 315.53 11.065 315.74 11.135 ;
    RECT 210.24 11.325 210.45 11.395 ;
    RECT 325.98 11.325 326.19 11.395 ;
    RECT 326.44 11.325 326.65 11.395 ;
    RECT 279.5 11.325 279.71 11.395 ;
    RECT 279.96 11.325 280.17 11.395 ;
    RECT 345.41 10.805 345.62 10.875 ;
    RECT 285.65 10.805 285.86 10.875 ;
    RECT 235.85 10.805 236.06 10.875 ;
    RECT 373.375 10.545 373.595 10.615 ;
    RECT 370.055 10.545 370.275 10.615 ;
    RECT 212.61 11.065 212.82 11.135 ;
    RECT 362.01 11.065 362.22 11.135 ;
    RECT 371.97 11.065 372.18 11.135 ;
    RECT 312.21 11.065 312.42 11.135 ;
    RECT 206.46 11.325 206.67 11.395 ;
    RECT 252.45 11.065 252.66 11.135 ;
    RECT 206.92 11.325 207.13 11.395 ;
    RECT 322.66 11.325 322.87 11.395 ;
    RECT 323.12 11.325 323.33 11.395 ;
    RECT 366.735 10.545 366.955 10.615 ;
    RECT 363.415 10.545 363.635 10.615 ;
    RECT 276.18 11.325 276.39 11.395 ;
    RECT 360.095 10.545 360.315 10.615 ;
    RECT 276.64 11.325 276.85 11.395 ;
    RECT 356.775 10.545 356.995 10.615 ;
    RECT 353.455 10.545 353.675 10.615 ;
    RECT 350.135 10.545 350.355 10.615 ;
    RECT 346.815 10.545 347.035 10.615 ;
    RECT 343.495 10.545 343.715 10.615 ;
    RECT 342.09 10.805 342.3 10.875 ;
    RECT 340.175 10.545 340.395 10.615 ;
    RECT 282.33 10.805 282.54 10.875 ;
    RECT 336.855 10.545 337.075 10.615 ;
    RECT 209.29 11.065 209.5 11.135 ;
    RECT 266.22 11.325 266.43 11.395 ;
    RECT 266.68 11.325 266.89 11.395 ;
    RECT 358.69 11.065 358.9 11.135 ;
    RECT 368.65 11.065 368.86 11.135 ;
    RECT 308.89 11.065 309.1 11.135 ;
    RECT 249.13 11.065 249.34 11.135 ;
    RECT 333.535 10.545 333.755 10.615 ;
    RECT 203.14 11.325 203.35 11.395 ;
    RECT 330.215 10.545 330.435 10.615 ;
    RECT 203.6 11.325 203.81 11.395 ;
    RECT 326.895 10.545 327.115 10.615 ;
    RECT 323.575 10.545 323.795 10.615 ;
    RECT 319.34 11.325 319.55 11.395 ;
    RECT 320.255 10.545 320.475 10.615 ;
    RECT 319.8 11.325 320.01 11.395 ;
    RECT 316.935 10.545 317.155 10.615 ;
    RECT 313.615 10.545 313.835 10.615 ;
    RECT 272.86 11.325 273.07 11.395 ;
    RECT 310.295 10.545 310.515 10.615 ;
    RECT 273.32 11.325 273.53 11.395 ;
    RECT 306.975 10.545 307.195 10.615 ;
    RECT 303.655 10.545 303.875 10.615 ;
    RECT 232.53 10.805 232.74 10.875 ;
    RECT 279.01 10.805 279.22 10.875 ;
    RECT 372.46 11.325 372.67 11.395 ;
    RECT 372.92 11.325 373.13 11.395 ;
    RECT 205.97 11.065 206.18 11.135 ;
    RECT 262.9 11.325 263.11 11.395 ;
    RECT 263.36 11.325 263.57 11.395 ;
    RECT 355.37 11.065 355.58 11.135 ;
    RECT 300.335 10.545 300.555 10.615 ;
    RECT 297.015 10.545 297.235 10.615 ;
    RECT 293.695 10.545 293.915 10.615 ;
    RECT 305.57 11.065 305.78 11.135 ;
    RECT 338.77 10.805 338.98 10.875 ;
    RECT 290.375 10.545 290.595 10.615 ;
    RECT 245.81 11.065 246.02 11.135 ;
    RECT 287.055 10.545 287.275 10.615 ;
    RECT 283.735 10.545 283.955 10.615 ;
    RECT 280.415 10.545 280.635 10.615 ;
    RECT 277.095 10.545 277.315 10.615 ;
    RECT 273.775 10.545 273.995 10.615 ;
    RECT 270.455 10.545 270.675 10.615 ;
    RECT 269.54 11.325 269.75 11.395 ;
    RECT 270.0 11.325 270.21 11.395 ;
    RECT 229.21 10.805 229.42 10.875 ;
    RECT 275.69 10.805 275.9 10.875 ;
    RECT 369.14 11.325 369.35 11.395 ;
    RECT 316.02 11.325 316.23 11.395 ;
    RECT 369.6 11.325 369.81 11.395 ;
    RECT 316.48 11.325 316.69 11.395 ;
    RECT 202.65 11.065 202.86 11.135 ;
    RECT 267.135 10.545 267.355 10.615 ;
    RECT 263.815 10.545 264.035 10.615 ;
    RECT 260.495 10.545 260.715 10.615 ;
    RECT 259.58 11.325 259.79 11.395 ;
    RECT 257.175 10.545 257.395 10.615 ;
    RECT 260.04 11.325 260.25 11.395 ;
    RECT 253.855 10.545 254.075 10.615 ;
    RECT 250.535 10.545 250.755 10.615 ;
    RECT 247.215 10.545 247.435 10.615 ;
    RECT 302.25 11.065 302.46 11.135 ;
    RECT 335.45 10.805 335.66 10.875 ;
    RECT 243.895 10.545 244.115 10.615 ;
    RECT 242.49 11.065 242.7 11.135 ;
    RECT 240.575 10.545 240.795 10.615 ;
    RECT 237.255 10.545 237.475 10.615 ;
    RECT 225.89 10.805 226.1 10.875 ;
    RECT 352.05 11.065 352.26 11.135 ;
    RECT 312.7 11.325 312.91 11.395 ;
    RECT 313.16 11.325 313.37 11.395 ;
    RECT 256.26 11.325 256.47 11.395 ;
    RECT 256.72 11.325 256.93 11.395 ;
    RECT 239.17 11.065 239.38 11.135 ;
    RECT 272.37 10.805 272.58 10.875 ;
    RECT 222.57 10.805 222.78 10.875 ;
    RECT 348.73 11.065 348.94 11.135 ;
    RECT 309.38 11.325 309.59 11.395 ;
    RECT 309.84 11.325 310.05 11.395 ;
    RECT 252.94 11.325 253.15 11.395 ;
    RECT 253.4 11.325 253.61 11.395 ;
    RECT 235.85 11.065 236.06 11.135 ;
    RECT 269.05 10.805 269.26 10.875 ;
    RECT 219.25 10.805 219.46 10.875 ;
    RECT 345.41 11.065 345.62 11.135 ;
    RECT 306.06 11.325 306.27 11.395 ;
    RECT 306.52 11.325 306.73 11.395 ;
    RECT 332.13 10.805 332.34 10.875 ;
    RECT 298.93 11.065 299.14 11.135 ;
    RECT 215.93 10.805 216.14 10.875 ;
    RECT 342.09 11.065 342.3 11.135 ;
    RECT 249.62 11.325 249.83 11.395 ;
    RECT 250.08 11.325 250.29 11.395 ;
    RECT 365.82 11.325 366.03 11.395 ;
    RECT 302.74 11.325 302.95 11.395 ;
    RECT 366.28 11.325 366.49 11.395 ;
    RECT 303.2 11.325 303.41 11.395 ;
    RECT 295.61 11.065 295.82 11.135 ;
    RECT 328.81 10.805 329.02 10.875 ;
    RECT 212.61 10.805 212.82 10.875 ;
    RECT 338.77 11.065 338.98 11.135 ;
    RECT 246.3 11.325 246.51 11.395 ;
    RECT 246.76 11.325 246.97 11.395 ;
    RECT 233.935 10.545 234.155 10.615 ;
    RECT 230.615 10.545 230.835 10.615 ;
    RECT 227.295 10.545 227.515 10.615 ;
    RECT 362.5 11.325 362.71 11.395 ;
    RECT 223.975 10.545 224.195 10.615 ;
    RECT 362.96 11.325 363.17 11.395 ;
    RECT 220.655 10.545 220.875 10.615 ;
    RECT 217.335 10.545 217.555 10.615 ;
    RECT 214.015 10.545 214.235 10.615 ;
    RECT 210.695 10.545 210.915 10.615 ;
    RECT 207.375 10.545 207.595 10.615 ;
    RECT 204.055 10.545 204.275 10.615 ;
    RECT 292.29 11.065 292.5 11.135 ;
    RECT 325.49 10.805 325.7 10.875 ;
    RECT 265.73 10.805 265.94 10.875 ;
    RECT 209.29 10.805 209.5 10.875 ;
    RECT 335.45 11.065 335.66 11.135 ;
    RECT 275.69 11.065 275.9 11.135 ;
    RECT 242.98 11.325 243.19 11.395 ;
    RECT 243.44 11.325 243.65 11.395 ;
    RECT 359.18 11.325 359.39 11.395 ;
    RECT 359.64 11.325 359.85 11.395 ;
    RECT 288.97 11.065 289.18 11.135 ;
    RECT 322.17 10.805 322.38 10.875 ;
    RECT 262.41 10.805 262.62 10.875 ;
    RECT 233.02 11.325 233.23 11.395 ;
    RECT 233.48 11.325 233.69 11.395 ;
    RECT 272.37 11.065 272.58 11.135 ;
    RECT 239.66 11.325 239.87 11.395 ;
    RECT 240.12 11.325 240.33 11.395 ;
    RECT 355.86 11.325 356.07 11.395 ;
    RECT 356.32 11.325 356.53 11.395 ;
    RECT 205.97 10.805 206.18 10.875 ;
    RECT 318.85 10.805 319.06 10.875 ;
    RECT 259.09 10.805 259.3 10.875 ;
    RECT 229.7 11.325 229.91 11.395 ;
    RECT 230.16 11.325 230.37 11.395 ;
    RECT 269.05 11.065 269.26 11.135 ;
    RECT 299.42 11.325 299.63 11.395 ;
    RECT 236.34 11.325 236.55 11.395 ;
    RECT 299.88 11.325 300.09 11.395 ;
    RECT 236.8 11.325 237.01 11.395 ;
    RECT 285.65 11.065 285.86 11.135 ;
    RECT 352.54 11.325 352.75 11.395 ;
    RECT 202.65 10.805 202.86 10.875 ;
    RECT 353.0 11.325 353.21 11.395 ;
    RECT 315.53 10.805 315.74 10.875 ;
    RECT 255.77 10.805 255.98 10.875 ;
    RECT 232.53 11.065 232.74 11.135 ;
    RECT 226.38 11.325 226.59 11.395 ;
    RECT 226.84 11.325 227.05 11.395 ;
    RECT 332.13 11.065 332.34 11.135 ;
    RECT 365.33 10.805 365.54 10.875 ;
    RECT 296.1 11.325 296.31 11.395 ;
    RECT 296.56 11.325 296.77 11.395 ;
    RECT 282.33 11.065 282.54 11.135 ;
    RECT 312.21 10.805 312.42 10.875 ;
    RECT 252.45 10.805 252.66 10.875 ;
    RECT 229.21 11.065 229.42 11.135 ;
    RECT 223.06 11.325 223.27 11.395 ;
    RECT 223.52 11.325 223.73 11.395 ;
    RECT 349.22 11.325 349.43 11.395 ;
    RECT 349.68 11.325 349.89 11.395 ;
    RECT 362.01 10.805 362.22 10.875 ;
    RECT 328.81 11.065 329.02 11.135 ;
    RECT 371.97 10.805 372.18 10.875 ;
    RECT 292.78 11.325 292.99 11.395 ;
    RECT 279.01 11.065 279.22 11.135 ;
    RECT 293.24 11.325 293.45 11.395 ;
    RECT 308.89 10.805 309.1 10.875 ;
    RECT 249.13 10.805 249.34 10.875 ;
    RECT 225.89 11.065 226.1 11.135 ;
    RECT 219.74 11.325 219.95 11.395 ;
    RECT 220.2 11.325 220.41 11.395 ;
    RECT 345.9 11.325 346.11 11.395 ;
    RECT 358.69 10.805 358.9 10.875 ;
    RECT 346.36 11.325 346.57 11.395 ;
    RECT 325.49 11.065 325.7 11.135 ;
    RECT 298.93 10.805 299.14 10.875 ;
    RECT 265.73 11.065 265.94 11.135 ;
    RECT 368.65 10.805 368.86 10.875 ;
    RECT 289.46 11.325 289.67 11.395 ;
    RECT 289.92 11.325 290.13 11.395 ;
    RECT 177.375 3.342 177.585 3.412 ;
    RECT 175.16 5.125 175.37 5.195 ;
    RECT 175.16 3.342 175.37 3.412 ;
    RECT 174.56 11.325 174.63 11.395 ;
    RECT 185.25 10.232 185.32 10.302 ;
    RECT 199.28 10.077 199.49 10.147 ;
    RECT 199.28 6.385 199.49 6.455 ;
    RECT 199.28 5.295 199.49 5.365 ;
    RECT 182.27 9.29 182.34 9.5 ;
    RECT 174.56 10.062 174.63 10.272 ;
    RECT 174.56 5.125 174.63 5.195 ;
    RECT 174.56 3.342 174.63 3.412 ;
    RECT 174.56 1.727 174.63 1.797 ;
    RECT 182.27 4.87 182.34 4.94 ;
    RECT 182.27 4.62 182.34 4.69 ;
    RECT 199.28 2.585 199.49 2.795 ;
    RECT 182.27 3.182 182.34 3.252 ;
    RECT 198.605 10.342 198.815 10.412 ;
    RECT 182.27 1.495 182.34 1.565 ;
    RECT 181.835 5.945 182.045 6.155 ;
    RECT 198.605 5.72 198.815 5.79 ;
    RECT 198.605 4.607 198.815 4.677 ;
    RECT 198.605 4.11 198.815 4.32 ;
    RECT 196.81 8.135 197.02 8.205 ;
    RECT 196.81 6.385 197.02 6.455 ;
    RECT 196.81 5.295 197.02 5.365 ;
    RECT 196.81 2.585 197.02 2.795 ;
    RECT 196.81 1.48 197.02 1.55 ;
    RECT 196.185 8.135 196.255 8.205 ;
    RECT 196.185 6.385 196.255 6.455 ;
    RECT 196.185 5.295 196.255 5.365 ;
    RECT 196.185 2.585 196.255 2.795 ;
    RECT 194.535 8.135 194.745 8.205 ;
    RECT 194.535 5.295 194.745 5.365 ;
    RECT 194.535 2.585 194.745 2.795 ;
    RECT 193.595 5.72 193.805 5.79 ;
    RECT 193.595 4.11 193.805 4.32 ;
    RECT 192.85 8.135 193.06 8.205 ;
    RECT 192.85 6.105 193.06 6.175 ;
    RECT 192.85 5.295 193.06 5.365 ;
    RECT 192.85 2.585 193.06 2.795 ;
    RECT 191.02 4.11 191.23 4.32 ;
    RECT 190.04 6.105 190.25 6.175 ;
    RECT 190.04 5.295 190.25 5.365 ;
    RECT 190.04 2.585 190.25 2.795 ;
    RECT 200.815 10.545 200.885 10.615 ;
    RECT 200.815 9.205 200.885 9.415 ;
    RECT 200.815 5.33 200.885 5.54 ;
    RECT 200.815 3.235 200.885 3.445 ;
    RECT 187.46 5.295 187.67 5.365 ;
    RECT 187.46 2.585 187.67 2.795 ;
    RECT 200.815 1.41 200.885 1.62 ;
    RECT 199.885 0.752 200.095 0.822 ;
    RECT 199.702 1.852 199.772 1.922 ;
    RECT 198.99 2.255 199.06 2.325 ;
    RECT 196.43 2.255 196.64 2.325 ;
    RECT 184.915 5.295 184.985 5.365 ;
    RECT 184.915 2.585 184.985 2.795 ;
    RECT 184.12 4.11 184.33 4.32 ;
    RECT 183.085 4.11 183.295 4.32 ;
    RECT 195.055 2.255 195.265 2.325 ;
    RECT 191.84 2.255 192.05 2.325 ;
    RECT 181.455 5.295 181.665 5.365 ;
    RECT 181.455 2.585 181.665 2.795 ;
    RECT 180.81 7.922 181.02 7.992 ;
    RECT 191.49 9.29 191.56 9.5 ;
    RECT 191.49 7.562 191.56 7.632 ;
    RECT 191.49 4.87 191.56 4.94 ;
    RECT 191.49 3.182 191.56 3.252 ;
    RECT 191.49 1.03 191.56 1.1 ;
    RECT 180.81 4.11 181.02 4.32 ;
    RECT 180.81 1.19 181.02 1.26 ;
    RECT 179.88 2.585 180.09 2.795 ;
    RECT 178.23 2.585 178.44 2.795 ;
    RECT 177.375 2.585 177.585 2.795 ;
    RECT 190.745 2.255 190.815 2.325 ;
    RECT 189.655 2.255 189.865 2.325 ;
    RECT 186.695 2.255 186.905 2.325 ;
    RECT 173.735 2.385 173.805 2.455 ;
    RECT 173.735 4.455 173.805 4.525 ;
    RECT 173.735 4.455 173.805 4.525 ;
    RECT 173.735 10.315 173.805 10.385 ;
    RECT 173.945 1.73 174.015 1.8 ;
    RECT 173.945 3.575 174.015 3.645 ;
    RECT 173.945 4.055 174.015 4.125 ;
    RECT 173.945 11.325 174.015 11.395 ;
    RECT 174.155 9.09 174.225 9.16 ;
    RECT 174.155 9.09 174.225 9.16 ;
    RECT 174.155 11.065 174.225 11.135 ;
    RECT 174.56 11.565 174.63 11.635 ;
    RECT 174.775 6.61 174.845 6.68 ;
    RECT 174.925 1.4 174.995 1.47 ;
    RECT 174.925 5.475 174.995 5.545 ;
    RECT 175.16 4.11 175.37 4.32 ;
    RECT 175.16 10.125 175.37 10.195 ;
    RECT 175.515 1.75 175.585 1.82 ;
    RECT 175.515 3.185 175.585 3.255 ;
    RECT 175.515 4.715 175.585 4.785 ;
    RECT 175.515 4.87 175.585 4.94 ;
    RECT 175.515 9.29 175.585 9.36 ;
    RECT 175.515 9.43 175.585 9.5 ;
    RECT 175.515 10.545 175.585 10.615 ;
    RECT 175.725 1.58 175.795 1.65 ;
    RECT 175.725 1.58 175.985 1.65 ;
    RECT 175.735 2.585 175.965 2.795 ;
    RECT 175.735 6.385 175.98 6.455 ;
    RECT 175.75 1.055 175.96 1.125 ;
    RECT 175.915 1.58 175.985 1.65 ;
    RECT 176.345 10.81 176.575 10.88 ;
    RECT 176.875 10.81 177.105 10.88 ;
    RECT 177.345 1.235 177.615 1.305 ;
    RECT 177.36 7.915 177.6 7.985 ;
    RECT 177.365 4.11 177.575 4.32 ;
    RECT 177.81 4.885 178.075 4.955 ;
    RECT 177.815 1.605 178.075 1.675 ;
    RECT 177.825 9.29 178.055 9.5 ;
    RECT 177.835 1.925 178.045 1.995 ;
    RECT 177.835 3.185 178.045 3.255 ;
    RECT 177.835 5.295 178.045 5.365 ;
    RECT 177.835 8.14 178.045 8.21 ;
    RECT 178.23 1.235 178.44 1.305 ;
    RECT 178.23 4.11 178.44 4.32 ;
    RECT 178.23 7.885 178.44 7.955 ;
    RECT 178.765 9.765 179.025 10.165 ;
    RECT 179.175 4.575 179.385 4.645 ;
    RECT 179.315 5.29 179.385 5.36 ;
    RECT 179.5 6.035 179.71 6.105 ;
    RECT 179.87 7.915 180.1 7.985 ;
    RECT 179.87 10.15 180.1 10.36 ;
    RECT 179.88 1.19 180.09 1.26 ;
    RECT 179.88 4.11 180.09 4.32 ;
    RECT 180.44 1.925 180.65 1.995 ;
    RECT 180.44 3.185 180.65 3.255 ;
    RECT 180.44 4.62 180.65 4.94 ;
    RECT 180.44 7.56 180.65 7.63 ;
    RECT 180.44 9.29 180.65 9.5 ;
    RECT 180.505 5.985 180.575 6.195 ;
    RECT 180.79 1.64 180.86 1.71 ;
    RECT 180.79 1.64 181.04 1.71 ;
    RECT 180.79 5.935 180.86 6.005 ;
    RECT 180.79 5.935 181.04 6.005 ;
    RECT 180.8 9.955 181.03 10.165 ;
    RECT 180.81 2.585 181.02 2.795 ;
    RECT 180.97 1.64 181.04 1.71 ;
    RECT 180.97 5.935 181.04 6.005 ;
    RECT 181.225 1.925 181.295 1.995 ;
    RECT 181.225 3.185 181.295 3.255 ;
    RECT 181.225 4.62 181.295 4.69 ;
    RECT 181.225 4.87 181.295 4.94 ;
    RECT 181.225 6.125 181.295 6.195 ;
    RECT 181.225 7.56 181.295 7.63 ;
    RECT 181.225 9.29 181.295 9.5 ;
    RECT 181.455 1.19 181.665 1.26 ;
    RECT 181.455 4.11 181.665 4.32 ;
    RECT 181.455 7.915 181.665 7.985 ;
    RECT 181.825 9.29 182.055 9.5 ;
    RECT 181.835 1.495 182.045 1.565 ;
    RECT 181.835 1.925 182.045 1.995 ;
    RECT 181.835 3.185 182.045 3.255 ;
    RECT 181.835 4.62 182.045 4.945 ;
    RECT 181.835 7.56 182.045 7.63 ;
    RECT 182.27 5.945 182.34 6.155 ;
    RECT 182.545 9.29 182.795 9.5 ;
    RECT 182.555 4.62 182.785 4.945 ;
    RECT 182.565 1.495 182.775 1.565 ;
    RECT 182.565 3.185 182.775 3.255 ;
    RECT 183.055 5.295 183.125 5.365 ;
    RECT 183.055 5.295 183.325 5.365 ;
    RECT 183.06 8.135 183.325 8.205 ;
    RECT 183.065 2.585 183.315 2.795 ;
    RECT 183.255 5.295 183.325 5.365 ;
    RECT 183.255 8.135 183.325 8.205 ;
    RECT 183.49 1.34 183.56 1.41 ;
    RECT 183.49 10.225 183.56 10.295 ;
    RECT 183.715 3.345 183.785 3.415 ;
    RECT 183.715 5.125 183.785 5.195 ;
    RECT 183.715 5.125 183.785 5.195 ;
    RECT 183.715 10.715 183.785 10.785 ;
    RECT 183.715 10.715 183.785 10.785 ;
    RECT 184.1 5.295 184.17 5.365 ;
    RECT 184.1 5.295 184.35 5.365 ;
    RECT 184.115 2.585 184.335 2.795 ;
    RECT 184.12 8.135 184.33 8.205 ;
    RECT 184.28 5.295 184.35 5.365 ;
    RECT 184.515 4.62 184.765 4.945 ;
    RECT 184.525 9.29 184.755 9.5 ;
    RECT 184.535 3.185 184.745 3.255 ;
    RECT 184.915 4.11 184.985 4.32 ;
    RECT 184.92 7.705 184.99 7.775 ;
    RECT 185.25 7.56 185.32 7.63 ;
    RECT 185.42 1.78 185.82 1.85 ;
    RECT 185.42 8.135 185.49 8.205 ;
    RECT 185.75 7.705 185.82 7.775 ;
    RECT 186.14 1.495 186.21 1.565 ;
    RECT 186.14 10.235 186.21 10.305 ;
    RECT 186.695 1.03 186.905 1.1 ;
    RECT 186.695 3.185 186.905 3.255 ;
    RECT 186.695 4.875 186.905 4.945 ;
    RECT 186.695 7.565 186.905 7.635 ;
    RECT 186.765 9.29 186.835 9.5 ;
    RECT 187.435 4.11 187.695 4.32 ;
    RECT 188.625 1.64 188.95 1.71 ;
    RECT 188.645 6.43 188.915 6.5 ;
    RECT 189.64 4.885 189.88 4.955 ;
    RECT 189.64 9.29 189.88 9.5 ;
    RECT 189.655 1.03 189.865 1.1 ;
    RECT 189.655 3.185 189.865 3.255 ;
    RECT 189.655 4.43 189.865 4.5 ;
    RECT 189.655 7.565 189.865 7.635 ;
    RECT 190.04 4.11 190.25 4.32 ;
    RECT 190.745 1.03 190.815 1.1 ;
    RECT 190.745 3.185 190.815 3.255 ;
    RECT 190.745 4.87 190.815 4.94 ;
    RECT 190.745 7.565 190.815 7.635 ;
    RECT 190.745 9.29 190.815 9.5 ;
    RECT 190.99 5.295 191.06 5.365 ;
    RECT 190.99 5.295 191.26 5.365 ;
    RECT 190.99 6.105 191.06 6.175 ;
    RECT 190.99 6.105 191.26 6.175 ;
    RECT 191.01 2.585 191.24 2.795 ;
    RECT 191.02 8.135 191.23 8.205 ;
    RECT 191.19 5.295 191.26 5.365 ;
    RECT 191.19 6.105 191.26 6.175 ;
    RECT 191.485 2.255 191.555 2.325 ;
    RECT 191.83 4.875 192.06 4.945 ;
    RECT 191.83 9.29 192.06 9.5 ;
    RECT 191.84 1.03 192.05 1.1 ;
    RECT 191.84 3.185 192.05 3.255 ;
    RECT 191.84 7.565 192.05 7.635 ;
    RECT 192.85 5.72 193.06 5.79 ;
    RECT 192.855 4.11 193.065 4.32 ;
    RECT 193.21 1.185 193.28 1.255 ;
    RECT 193.21 9.91 193.42 9.98 ;
    RECT 193.565 5.295 193.635 5.365 ;
    RECT 193.565 5.295 193.835 5.365 ;
    RECT 193.565 6.595 193.635 6.665 ;
    RECT 193.565 6.595 193.835 6.665 ;
    RECT 193.565 9.08 193.635 9.15 ;
    RECT 193.565 9.08 193.835 9.15 ;
    RECT 193.585 2.585 193.815 2.795 ;
    RECT 193.595 6.105 193.805 6.175 ;
    RECT 193.595 8.135 193.805 8.205 ;
    RECT 193.595 10.085 193.805 10.295 ;
    RECT 193.765 5.295 193.835 5.365 ;
    RECT 193.765 6.595 193.835 6.665 ;
    RECT 193.765 9.08 193.835 9.15 ;
    RECT 194.015 3.345 194.085 3.415 ;
    RECT 194.015 5.125 194.085 5.195 ;
    RECT 194.015 5.125 194.085 5.195 ;
    RECT 194.515 10.085 194.77 10.295 ;
    RECT 194.535 4.11 194.745 4.32 ;
    RECT 194.535 5.72 194.745 5.79 ;
    RECT 195.025 5.98 195.3 6.05 ;
    RECT 195.025 6.595 195.3 6.665 ;
    RECT 195.04 4.875 195.28 4.945 ;
    RECT 195.04 9.29 195.28 9.5 ;
    RECT 195.055 1.03 195.265 1.1 ;
    RECT 195.055 3.185 195.265 3.255 ;
    RECT 195.055 7.565 195.265 7.85 ;
    RECT 195.63 9.765 195.84 9.835 ;
    RECT 195.63 11.07 195.84 11.28 ;
    RECT 196.185 4.61 196.255 4.68 ;
    RECT 196.185 5.72 196.255 5.79 ;
    RECT 196.19 4.11 196.26 4.18 ;
    RECT 196.19 4.11 196.26 4.18 ;
    RECT 196.19 4.25 196.26 4.32 ;
    RECT 196.19 4.25 196.26 4.32 ;
    RECT 196.2 10.085 196.27 10.155 ;
    RECT 196.2 10.085 196.27 10.155 ;
    RECT 196.2 10.225 196.27 10.295 ;
    RECT 196.2 10.225 196.27 10.295 ;
    RECT 196.43 1.03 196.64 1.1 ;
    RECT 196.43 3.185 196.64 3.255 ;
    RECT 196.43 4.87 196.64 4.94 ;
    RECT 196.43 5.98 196.64 6.05 ;
    RECT 196.43 7.565 196.64 7.85 ;
    RECT 196.43 9.29 196.64 9.5 ;
    RECT 196.78 7.965 197.05 8.035 ;
    RECT 196.78 10.085 197.05 10.295 ;
    RECT 196.81 4.11 197.02 4.32 ;
    RECT 196.81 4.61 197.02 4.68 ;
    RECT 196.81 5.72 197.02 5.79 ;
    RECT 197.225 3.345 197.295 3.415 ;
    RECT 197.225 5.13 197.295 5.2 ;
    RECT 197.465 11.1 197.675 11.17 ;
    RECT 198.045 11.1 198.115 11.17 ;
    RECT 198.045 11.1 198.255 11.17 ;
    RECT 198.185 11.1 198.255 11.17 ;
    RECT 198.185 11.1 198.255 11.17 ;
    RECT 198.4 6.62 198.47 6.69 ;
    RECT 198.605 1.48 198.675 1.55 ;
    RECT 198.605 1.48 198.815 1.55 ;
    RECT 198.605 2.585 198.675 2.655 ;
    RECT 198.605 2.585 198.675 2.655 ;
    RECT 198.605 2.585 198.815 2.795 ;
    RECT 198.605 2.725 198.675 2.795 ;
    RECT 198.605 2.725 198.675 2.795 ;
    RECT 198.605 5.295 198.675 5.365 ;
    RECT 198.605 5.295 198.675 5.365 ;
    RECT 198.605 5.295 198.815 5.365 ;
    RECT 198.605 6.385 198.675 6.455 ;
    RECT 198.605 6.385 198.675 6.455 ;
    RECT 198.605 6.385 198.815 6.455 ;
    RECT 198.605 8.135 198.675 8.205 ;
    RECT 198.605 8.135 198.815 8.205 ;
    RECT 198.605 10.08 198.675 10.15 ;
    RECT 198.605 10.08 198.815 10.15 ;
    RECT 198.745 1.48 198.815 1.55 ;
    RECT 198.745 2.585 198.815 2.655 ;
    RECT 198.745 2.585 198.815 2.655 ;
    RECT 198.745 2.725 198.815 2.795 ;
    RECT 198.745 2.725 198.815 2.795 ;
    RECT 198.745 5.295 198.815 5.365 ;
    RECT 198.745 5.295 198.815 5.365 ;
    RECT 198.745 6.385 198.815 6.455 ;
    RECT 198.745 6.385 198.815 6.455 ;
    RECT 198.745 8.135 198.815 8.205 ;
    RECT 198.745 10.08 198.815 10.15 ;
    RECT 198.99 1.03 199.06 1.1 ;
    RECT 198.99 3.18 199.06 3.25 ;
    RECT 198.99 3.18 199.06 3.25 ;
    RECT 198.99 9.29 199.06 9.36 ;
    RECT 198.99 9.29 199.06 9.36 ;
    RECT 198.99 9.43 199.06 9.5 ;
    RECT 198.99 9.43 199.06 9.5 ;
    RECT 198.99 10.545 199.06 10.615 ;
    RECT 198.995 4.875 199.065 4.945 ;
    RECT 198.995 4.875 199.065 4.945 ;
    RECT 199.26 4.11 199.47 4.32 ;
    RECT 199.265 4.61 199.475 4.68 ;
    RECT 199.275 10.34 199.485 10.41 ;
    RECT 199.295 5.855 199.365 6.115 ;
    RECT 199.705 9.915 199.775 9.985 ;
    RECT 199.885 3.18 200.095 3.25 ;
    RECT 199.885 4.875 200.095 4.945 ;
    RECT 199.885 9.29 200.095 9.5 ;
    RECT 199.885 10.545 200.095 10.615 ;
    RECT 200.395 11.065 200.465 11.135 ;
    RECT 200.4 9.095 200.47 9.165 ;
    RECT 200.4 9.095 200.47 9.165 ;
    RECT 200.595 5.665 200.665 5.735 ;
    RECT 200.595 5.665 200.665 5.735 ;
    RECT 200.605 3.59 200.675 3.66 ;
    RECT 200.605 4.055 200.675 4.125 ;
    RECT 200.605 11.325 200.675 11.395 ;
    RECT 200.81 0.75 200.88 0.82 ;
    RECT 200.815 4.455 200.885 4.525 ;
    RECT 200.815 4.455 200.885 4.525 ;
    RECT 200.815 10.315 200.885 10.385 ;
    RECT 175.75 10.062 175.96 10.272 ;
    RECT 175.75 4.11 175.96 4.32 ;
    RECT 175.16 6.385 175.37 6.455 ;
    RECT 184.535 2.255 184.745 2.325 ;
    RECT 182.565 2.255 182.775 2.325 ;
    RECT 181.835 2.255 182.045 2.325 ;
    RECT 181.225 8.14 181.295 8.21 ;
    RECT 181.225 2.255 181.295 2.325 ;
    RECT 175.16 2.585 175.37 2.795 ;
    RECT 175.16 0.915 175.37 1.125 ;
    RECT 174.56 6.385 174.63 6.455 ;
    RECT 180.44 8.14 180.65 8.21 ;
    RECT 180.44 2.255 180.65 2.325 ;
    RECT 174.56 2.585 174.63 2.795 ;
    RECT 199.28 5.125 199.49 5.195 ;
    RECT 174.56 0.915 174.63 1.125 ;
    RECT 199.28 3.342 199.49 3.412 ;
    RECT 197.222 4.607 197.292 4.677 ;
    RECT 177.835 2.255 178.045 2.325 ;
    RECT 197.222 4.11 197.292 4.32 ;
    RECT 196.81 5.125 197.02 5.195 ;
    RECT 196.81 3.342 197.02 3.412 ;
    RECT 196.185 5.125 196.255 5.195 ;
    RECT 196.185 3.342 196.255 3.412 ;
    RECT 194.535 5.125 194.745 5.195 ;
    RECT 194.535 3.342 194.745 3.412 ;
    RECT 194.015 5.72 194.085 5.79 ;
    RECT 175.515 2.255 175.585 2.325 ;
    RECT 173.735 10.545 173.805 10.615 ;
    RECT 173.735 9.205 173.805 9.415 ;
    RECT 173.735 5.33 173.805 5.54 ;
    RECT 173.735 3.235 173.805 3.445 ;
    RECT 194.015 4.11 194.085 4.32 ;
    RECT 192.85 5.125 193.06 5.195 ;
    RECT 192.85 3.342 193.06 3.412 ;
    RECT 190.04 5.125 190.25 5.195 ;
    RECT 190.04 3.342 190.25 3.412 ;
    RECT 200.395 9.765 200.465 9.835 ;
    RECT 173.735 1.41 173.805 1.62 ;
    RECT 187.46 5.125 187.67 5.195 ;
    RECT 174.155 9.765 174.225 9.835 ;
    RECT 187.46 3.342 187.67 3.412 ;
    RECT 184.915 5.125 184.985 5.195 ;
    RECT 184.915 3.342 184.985 3.412 ;
    RECT 183.715 4.11 183.785 4.32 ;
    RECT 181.455 10.717 181.665 10.787 ;
    RECT 181.455 5.125 181.665 5.195 ;
    RECT 181.455 3.342 181.665 3.412 ;
    RECT 179.88 5.125 180.09 5.195 ;
    RECT 179.88 3.342 180.09 3.412 ;
    RECT 176.885 9.765 177.095 9.835 ;
    RECT 176.355 9.765 176.565 9.835 ;
    RECT 198.045 9.765 198.255 9.835 ;
    RECT 197.465 9.765 197.675 9.835 ;
    RECT 178.23 10.647 178.44 10.717 ;
    RECT 178.23 5.125 178.44 5.195 ;
    RECT 178.23 3.342 178.44 3.412 ;
    RECT 177.375 10.647 177.585 10.717 ;
    RECT 177.375 5.125 177.585 5.195 ;
    RECT 102.5 1.24 102.71 1.31 ;
    RECT 97.31 1.41 97.52 1.62 ;
    RECT 97.68 1.005 97.95 2.125 ;
    RECT 98.23 1.24 98.44 1.31 ;
    RECT 99.18 0.915 99.39 2.125 ;
    RECT 93.99 1.41 94.2 1.62 ;
    RECT 94.36 1.005 94.63 2.125 ;
    RECT 94.91 1.24 95.12 1.31 ;
    RECT 95.86 0.915 96.07 2.125 ;
    RECT 101.55 2.055 101.76 2.125 ;
    RECT 90.67 1.41 90.88 1.62 ;
    RECT 91.04 1.005 91.31 2.125 ;
    RECT 91.59 1.24 91.8 1.31 ;
    RECT 92.54 0.915 92.75 2.125 ;
    RECT 87.35 1.41 87.56 1.62 ;
    RECT 87.72 1.005 87.99 2.125 ;
    RECT 88.27 1.24 88.48 1.31 ;
    RECT 89.22 0.915 89.43 2.125 ;
    RECT 5.27 0.915 5.48 1.125 ;
    RECT 84.03 1.41 84.24 1.62 ;
    RECT 84.4 1.005 84.67 2.125 ;
    RECT 84.95 1.24 85.16 1.31 ;
    RECT 85.9 0.915 86.11 2.125 ;
    RECT 80.71 1.41 80.92 1.62 ;
    RECT 81.08 1.005 81.35 2.125 ;
    RECT 81.63 1.24 81.84 1.31 ;
    RECT 82.58 0.915 82.79 2.125 ;
    RECT 77.39 1.41 77.6 1.62 ;
    RECT 77.76 1.005 78.03 2.125 ;
    RECT 78.31 1.24 78.52 1.31 ;
    RECT 79.26 0.915 79.47 2.125 ;
    RECT 74.07 1.41 74.28 1.62 ;
    RECT 74.44 1.005 74.71 2.125 ;
    RECT 74.99 1.24 75.2 1.31 ;
    RECT 75.94 0.915 76.15 2.125 ;
    RECT 70.75 1.41 70.96 1.62 ;
    RECT 71.12 1.005 71.39 2.125 ;
    RECT 71.67 1.24 71.88 1.31 ;
    RECT 72.62 0.915 72.83 2.125 ;
    RECT 67.43 1.41 67.64 1.62 ;
    RECT 67.8 1.005 68.07 2.125 ;
    RECT 68.35 1.24 68.56 1.31 ;
    RECT 69.3 0.915 69.51 2.125 ;
    RECT 16.18 1.24 16.39 1.31 ;
    RECT 101.55 1.742 101.76 1.812 ;
    RECT 119.1 1.24 119.31 1.31 ;
    RECT 101.55 0.915 101.76 1.125 ;
    RECT 118.15 2.055 118.36 2.125 ;
    RECT 64.11 1.41 64.32 1.62 ;
    RECT 64.48 1.005 64.75 2.125 ;
    RECT 65.03 1.24 65.24 1.31 ;
    RECT 65.98 0.915 66.19 2.125 ;
    RECT 60.79 1.41 61.0 1.62 ;
    RECT 61.16 1.005 61.43 2.125 ;
    RECT 61.71 1.24 61.92 1.31 ;
    RECT 62.66 0.915 62.87 2.125 ;
    RECT 57.47 1.41 57.68 1.62 ;
    RECT 57.84 1.005 58.11 2.125 ;
    RECT 58.39 1.24 58.6 1.31 ;
    RECT 59.34 0.915 59.55 2.125 ;
    RECT 54.15 1.41 54.36 1.62 ;
    RECT 54.52 1.005 54.79 2.125 ;
    RECT 55.07 1.24 55.28 1.31 ;
    RECT 56.02 0.915 56.23 2.125 ;
    RECT 158.94 1.24 159.15 1.31 ;
    RECT 50.83 1.41 51.04 1.62 ;
    RECT 51.2 1.005 51.47 2.125 ;
    RECT 51.75 1.24 51.96 1.31 ;
    RECT 52.7 0.915 52.91 2.125 ;
    RECT 15.23 2.055 15.44 2.125 ;
    RECT 47.51 1.41 47.72 1.62 ;
    RECT 47.88 1.005 48.15 2.125 ;
    RECT 48.43 1.24 48.64 1.31 ;
    RECT 49.38 0.915 49.59 2.125 ;
    RECT 15.23 1.742 15.44 1.812 ;
    RECT 44.19 1.41 44.4 1.62 ;
    RECT 44.56 1.005 44.83 2.125 ;
    RECT 45.11 1.24 45.32 1.31 ;
    RECT 46.06 0.915 46.27 2.125 ;
    RECT 157.99 2.055 158.2 2.125 ;
    RECT 79.26 1.24 79.47 1.31 ;
    RECT 40.87 1.41 41.08 1.62 ;
    RECT 41.24 1.005 41.51 2.125 ;
    RECT 41.79 1.24 42.0 1.31 ;
    RECT 42.74 0.915 42.95 2.125 ;
    RECT 157.99 1.742 158.2 1.812 ;
    RECT 37.55 1.41 37.76 1.62 ;
    RECT 37.92 1.005 38.19 2.125 ;
    RECT 38.47 1.24 38.68 1.31 ;
    RECT 39.42 0.915 39.63 2.125 ;
    RECT 34.23 1.41 34.44 1.62 ;
    RECT 34.6 1.005 34.87 2.125 ;
    RECT 35.15 1.24 35.36 1.31 ;
    RECT 36.1 0.915 36.31 2.125 ;
    RECT 78.31 2.055 78.52 2.125 ;
    RECT 15.23 0.915 15.44 1.125 ;
    RECT 78.31 1.742 78.52 1.812 ;
    RECT 78.31 0.915 78.52 1.125 ;
    RECT 118.15 1.742 118.36 1.812 ;
    RECT 118.15 0.915 118.36 1.125 ;
    RECT 157.99 0.915 158.2 1.125 ;
    RECT 115.78 1.24 115.99 1.31 ;
    RECT 155.62 1.24 155.83 1.31 ;
    RECT 154.67 2.055 154.88 2.125 ;
    RECT 154.67 1.742 154.88 1.812 ;
    RECT 114.83 2.055 115.04 2.125 ;
    RECT 114.83 1.742 115.04 1.812 ;
    RECT 132.38 1.24 132.59 1.31 ;
    RECT 114.83 0.915 115.04 1.125 ;
    RECT 154.67 0.915 154.88 1.125 ;
    RECT 152.3 1.24 152.51 1.31 ;
    RECT 151.35 2.055 151.56 2.125 ;
    RECT 112.46 1.24 112.67 1.31 ;
    RECT 111.51 2.055 111.72 2.125 ;
    RECT 111.51 1.742 111.72 1.812 ;
    RECT 111.51 0.915 111.72 1.125 ;
    RECT 151.35 1.742 151.56 1.812 ;
    RECT 151.35 0.915 151.56 1.125 ;
    RECT 48.43 2.055 48.64 2.125 ;
    RECT 48.43 1.742 48.64 1.812 ;
    RECT 65.98 1.24 66.19 1.31 ;
    RECT 48.43 0.915 48.64 1.125 ;
    RECT 65.03 2.055 65.24 2.125 ;
    RECT 65.03 1.742 65.24 1.812 ;
    RECT 65.03 0.915 65.24 1.125 ;
    RECT 2.9 1.24 3.11 1.31 ;
    RECT 32.78 1.24 32.99 1.31 ;
    RECT 148.98 1.24 149.19 1.31 ;
    RECT 1.95 2.055 2.16 2.125 ;
    RECT 109.14 1.24 109.35 1.31 ;
    RECT 108.19 2.055 108.4 2.125 ;
    RECT 108.19 1.742 108.4 1.812 ;
    RECT 148.03 2.055 148.24 2.125 ;
    RECT 1.95 1.742 2.16 1.812 ;
    RECT 31.83 2.055 32.04 2.125 ;
    RECT 148.03 1.742 148.24 1.812 ;
    RECT 31.83 1.742 32.04 1.812 ;
    RECT 165.58 1.24 165.79 1.31 ;
    RECT 1.95 0.915 2.16 1.125 ;
    RECT 148.03 0.915 148.24 1.125 ;
    RECT 31.83 0.915 32.04 1.125 ;
    RECT 108.19 0.915 108.4 1.125 ;
    RECT 164.63 2.055 164.84 2.125 ;
    RECT 164.63 1.742 164.84 1.812 ;
    RECT 164.63 0.915 164.84 1.125 ;
    RECT 12.86 1.24 13.07 1.31 ;
    RECT 11.91 2.055 12.12 2.125 ;
    RECT 11.91 1.742 12.12 1.812 ;
    RECT 46.06 1.24 46.27 1.31 ;
    RECT 11.91 0.915 12.12 1.125 ;
    RECT 45.11 2.055 45.32 2.125 ;
    RECT 45.11 1.742 45.32 1.812 ;
    RECT 45.11 0.915 45.32 1.125 ;
    RECT 62.66 1.24 62.87 1.31 ;
    RECT 61.71 2.055 61.92 2.125 ;
    RECT 61.71 1.742 61.92 1.812 ;
    RECT 61.71 0.915 61.92 1.125 ;
    RECT 21.87 0.915 22.08 1.125 ;
    RECT 105.82 1.24 106.03 1.31 ;
    RECT 104.87 2.055 105.08 2.125 ;
    RECT 104.87 1.742 105.08 1.812 ;
    RECT 145.66 1.24 145.87 1.31 ;
    RECT 29.46 1.24 29.67 1.31 ;
    RECT 144.71 2.055 144.92 2.125 ;
    RECT 28.51 2.055 28.72 2.125 ;
    RECT 144.71 1.742 144.92 1.812 ;
    RECT 28.51 1.742 28.72 1.812 ;
    RECT 144.71 0.915 144.92 1.125 ;
    RECT 28.51 0.915 28.72 1.125 ;
    RECT 162.26 1.24 162.47 1.31 ;
    RECT 161.31 2.055 161.52 2.125 ;
    RECT 161.31 1.742 161.52 1.812 ;
    RECT 161.31 0.915 161.52 1.125 ;
    RECT 42.74 1.24 42.95 1.31 ;
    RECT 41.79 2.055 42.0 2.125 ;
    RECT 41.79 1.742 42.0 1.812 ;
    RECT 99.18 1.24 99.39 1.31 ;
    RECT 59.34 1.24 59.55 1.31 ;
    RECT 41.79 0.915 42.0 1.125 ;
    RECT 58.39 2.055 58.6 2.125 ;
    RECT 58.39 1.742 58.6 1.812 ;
    RECT 98.23 2.055 98.44 2.125 ;
    RECT 98.23 1.742 98.44 1.812 ;
    RECT 98.23 0.915 98.44 1.125 ;
    RECT 58.39 0.915 58.6 1.125 ;
    RECT 142.34 1.24 142.55 1.31 ;
    RECT 26.14 1.24 26.35 1.31 ;
    RECT 141.39 2.055 141.6 2.125 ;
    RECT 25.19 2.055 25.4 2.125 ;
    RECT 141.39 1.742 141.6 1.812 ;
    RECT 25.19 1.742 25.4 1.812 ;
    RECT 25.19 0.915 25.4 1.125 ;
    RECT 141.39 0.915 141.6 1.125 ;
    RECT 39.42 1.24 39.63 1.31 ;
    RECT 38.47 2.055 38.68 2.125 ;
    RECT 38.47 1.742 38.68 1.812 ;
    RECT 56.02 1.24 56.23 1.31 ;
    RECT 38.47 0.915 38.68 1.125 ;
    RECT 55.07 2.055 55.28 2.125 ;
    RECT 55.07 1.742 55.28 1.812 ;
    RECT 95.86 1.24 96.07 1.31 ;
    RECT 94.91 2.055 95.12 2.125 ;
    RECT 94.91 1.742 95.12 1.812 ;
    RECT 94.91 0.915 95.12 1.125 ;
    RECT 55.07 0.915 55.28 1.125 ;
    RECT 22.82 1.24 23.03 1.31 ;
    RECT 139.02 1.24 139.23 1.31 ;
    RECT 21.87 2.055 22.08 2.125 ;
    RECT 138.07 2.055 138.28 2.125 ;
    RECT 21.87 1.742 22.08 1.812 ;
    RECT 138.07 1.742 138.28 1.812 ;
    RECT 138.07 0.915 138.28 1.125 ;
    RECT 36.1 1.24 36.31 1.31 ;
    RECT 35.15 2.055 35.36 2.125 ;
    RECT 75.94 1.24 76.15 1.31 ;
    RECT 74.99 2.055 75.2 2.125 ;
    RECT 74.99 1.742 75.2 1.812 ;
    RECT 35.15 1.742 35.36 1.812 ;
    RECT 52.7 1.24 52.91 1.31 ;
    RECT 35.15 0.915 35.36 1.125 ;
    RECT 51.75 2.055 51.96 2.125 ;
    RECT 92.54 1.24 92.75 1.31 ;
    RECT 74.99 0.915 75.2 1.125 ;
    RECT 91.59 2.055 91.8 2.125 ;
    RECT 91.59 1.742 91.8 1.812 ;
    RECT 131.43 2.055 131.64 2.125 ;
    RECT 131.43 1.742 131.64 1.812 ;
    RECT 9.54 1.24 9.75 1.31 ;
    RECT 51.75 1.742 51.96 1.812 ;
    RECT 131.43 0.915 131.64 1.125 ;
    RECT 8.59 2.055 8.8 2.125 ;
    RECT 8.59 1.742 8.8 1.812 ;
    RECT 51.75 0.915 51.96 1.125 ;
    RECT 91.59 0.915 91.8 1.125 ;
    RECT 135.7 1.24 135.91 1.31 ;
    RECT 134.75 2.055 134.96 2.125 ;
    RECT 8.59 0.915 8.8 1.125 ;
    RECT 19.5 1.24 19.71 1.31 ;
    RECT 18.55 2.055 18.76 2.125 ;
    RECT 134.75 1.742 134.96 1.812 ;
    RECT 134.75 0.915 134.96 1.125 ;
    RECT 18.55 1.742 18.76 1.812 ;
    RECT 18.55 0.915 18.76 1.125 ;
    RECT 72.62 1.24 72.83 1.31 ;
    RECT 71.67 2.055 71.88 2.125 ;
    RECT 71.67 1.742 71.88 1.812 ;
    RECT 49.38 1.24 49.59 1.31 ;
    RECT 89.22 1.24 89.43 1.31 ;
    RECT 71.67 0.915 71.88 1.125 ;
    RECT 88.27 2.055 88.48 2.125 ;
    RECT 88.27 1.742 88.48 1.812 ;
    RECT 129.06 1.24 129.27 1.31 ;
    RECT 128.11 2.055 128.32 2.125 ;
    RECT 128.11 1.742 128.32 1.812 ;
    RECT 128.11 0.915 128.32 1.125 ;
    RECT 88.27 0.915 88.48 1.125 ;
    RECT 172.22 1.24 172.43 1.31 ;
    RECT 171.27 2.055 171.48 2.125 ;
    RECT 171.27 1.742 171.48 1.812 ;
    RECT 171.27 0.915 171.48 1.125 ;
    RECT 69.3 1.24 69.51 1.31 ;
    RECT 68.35 2.055 68.56 2.125 ;
    RECT 68.35 1.742 68.56 1.812 ;
    RECT 85.9 1.24 86.11 1.31 ;
    RECT 68.35 0.915 68.56 1.125 ;
    RECT 84.95 2.055 85.16 2.125 ;
    RECT 125.74 1.24 125.95 1.31 ;
    RECT 124.79 2.055 125.0 2.125 ;
    RECT 124.79 1.742 125.0 1.812 ;
    RECT 84.95 1.742 85.16 1.812 ;
    RECT 84.95 0.915 85.16 1.125 ;
    RECT 170.35 1.41 170.56 1.62 ;
    RECT 170.72 1.005 170.99 2.125 ;
    RECT 171.27 1.24 171.48 1.31 ;
    RECT 172.22 0.915 172.43 2.125 ;
    RECT 124.79 0.915 125.0 1.125 ;
    RECT 1.03 1.41 1.24 1.62 ;
    RECT 1.4 1.005 1.67 2.125 ;
    RECT 1.95 1.24 2.16 1.31 ;
    RECT 2.9 0.915 3.11 2.125 ;
    RECT 168.9 1.24 169.11 1.31 ;
    RECT 167.95 2.055 168.16 2.125 ;
    RECT 30.91 1.41 31.12 1.62 ;
    RECT 31.28 1.005 31.55 2.125 ;
    RECT 31.83 1.24 32.04 1.31 ;
    RECT 32.78 0.915 32.99 2.125 ;
    RECT 27.59 1.41 27.8 1.62 ;
    RECT 27.96 1.005 28.23 2.125 ;
    RECT 28.51 1.24 28.72 1.31 ;
    RECT 29.46 0.915 29.67 2.125 ;
    RECT 24.27 1.41 24.48 1.62 ;
    RECT 24.64 1.005 24.91 2.125 ;
    RECT 25.19 1.24 25.4 1.31 ;
    RECT 26.14 0.915 26.35 2.125 ;
    RECT 20.95 1.41 21.16 1.62 ;
    RECT 21.32 1.005 21.59 2.125 ;
    RECT 21.87 1.24 22.08 1.31 ;
    RECT 22.82 0.915 23.03 2.125 ;
    RECT 17.63 1.41 17.84 1.62 ;
    RECT 18.0 1.005 18.27 2.125 ;
    RECT 18.55 1.24 18.76 1.31 ;
    RECT 19.5 0.915 19.71 2.125 ;
    RECT 14.31 1.41 14.52 1.62 ;
    RECT 14.68 1.005 14.95 2.125 ;
    RECT 15.23 1.24 15.44 1.31 ;
    RECT 16.18 0.915 16.39 2.125 ;
    RECT 10.99 1.41 11.2 1.62 ;
    RECT 11.36 1.005 11.63 2.125 ;
    RECT 11.91 1.24 12.12 1.31 ;
    RECT 12.86 0.915 13.07 2.125 ;
    RECT 7.67 1.41 7.88 1.62 ;
    RECT 8.04 1.005 8.31 2.125 ;
    RECT 8.59 1.24 8.8 1.31 ;
    RECT 9.54 0.915 9.75 2.125 ;
    RECT 4.35 1.41 4.56 1.62 ;
    RECT 4.72 1.005 4.99 2.125 ;
    RECT 5.27 1.24 5.48 1.31 ;
    RECT 6.22 0.915 6.43 2.125 ;
    RECT 167.95 1.742 168.16 1.812 ;
    RECT 167.95 0.915 168.16 1.125 ;
    RECT 82.58 1.24 82.79 1.31 ;
    RECT 122.42 1.24 122.63 1.31 ;
    RECT 104.87 0.915 105.08 1.125 ;
    RECT 121.47 2.055 121.68 2.125 ;
    RECT 121.47 1.742 121.68 1.812 ;
    RECT 167.03 1.41 167.24 1.62 ;
    RECT 167.4 1.005 167.67 2.125 ;
    RECT 167.95 1.24 168.16 1.31 ;
    RECT 168.9 0.915 169.11 2.125 ;
    RECT 81.63 2.055 81.84 2.125 ;
    RECT 81.63 1.742 81.84 1.812 ;
    RECT 81.63 0.915 81.84 1.125 ;
    RECT 163.71 1.41 163.92 1.62 ;
    RECT 164.08 1.005 164.35 2.125 ;
    RECT 164.63 1.24 164.84 1.31 ;
    RECT 165.58 0.915 165.79 2.125 ;
    RECT 121.47 0.915 121.68 1.125 ;
    RECT 160.39 1.41 160.6 1.62 ;
    RECT 160.76 1.005 161.03 2.125 ;
    RECT 161.31 1.24 161.52 1.31 ;
    RECT 162.26 0.915 162.47 2.125 ;
    RECT 157.07 1.41 157.28 1.62 ;
    RECT 157.44 1.005 157.71 2.125 ;
    RECT 157.99 1.24 158.2 1.31 ;
    RECT 158.94 0.915 159.15 2.125 ;
    RECT 153.75 1.41 153.96 1.62 ;
    RECT 154.12 1.005 154.39 2.125 ;
    RECT 154.67 1.24 154.88 1.31 ;
    RECT 155.62 0.915 155.83 2.125 ;
    RECT 150.43 1.41 150.64 1.62 ;
    RECT 150.8 1.005 151.07 2.125 ;
    RECT 151.35 1.24 151.56 1.31 ;
    RECT 152.3 0.915 152.51 2.125 ;
    RECT 147.11 1.41 147.32 1.62 ;
    RECT 147.48 1.005 147.75 2.125 ;
    RECT 148.03 1.24 148.24 1.31 ;
    RECT 148.98 0.915 149.19 2.125 ;
    RECT 143.79 1.41 144.0 1.62 ;
    RECT 144.16 1.005 144.43 2.125 ;
    RECT 144.71 1.24 144.92 1.31 ;
    RECT 145.66 0.915 145.87 2.125 ;
    RECT 140.47 1.41 140.68 1.62 ;
    RECT 140.84 1.005 141.11 2.125 ;
    RECT 141.39 1.24 141.6 1.31 ;
    RECT 142.34 0.915 142.55 2.125 ;
    RECT 137.15 1.41 137.36 1.62 ;
    RECT 137.52 1.005 137.79 2.125 ;
    RECT 138.07 1.24 138.28 1.31 ;
    RECT 139.02 0.915 139.23 2.125 ;
    RECT 133.83 1.41 134.04 1.62 ;
    RECT 134.2 1.005 134.47 2.125 ;
    RECT 134.75 1.24 134.96 1.31 ;
    RECT 135.7 0.915 135.91 2.125 ;
    RECT 130.51 1.41 130.72 1.62 ;
    RECT 130.88 1.005 131.15 2.125 ;
    RECT 131.43 1.24 131.64 1.31 ;
    RECT 132.38 0.915 132.59 2.125 ;
    RECT 127.19 1.41 127.4 1.62 ;
    RECT 127.56 1.005 127.83 2.125 ;
    RECT 128.11 1.24 128.32 1.31 ;
    RECT 129.06 0.915 129.27 2.125 ;
    RECT 123.87 1.41 124.08 1.62 ;
    RECT 124.24 1.005 124.51 2.125 ;
    RECT 124.79 1.24 125.0 1.31 ;
    RECT 125.74 0.915 125.95 2.125 ;
    RECT 120.55 1.41 120.76 1.62 ;
    RECT 120.92 1.005 121.19 2.125 ;
    RECT 121.47 1.24 121.68 1.31 ;
    RECT 122.42 0.915 122.63 2.125 ;
    RECT 117.23 1.41 117.44 1.62 ;
    RECT 117.6 1.005 117.87 2.125 ;
    RECT 118.15 1.24 118.36 1.31 ;
    RECT 119.1 0.915 119.31 2.125 ;
    RECT 6.22 1.24 6.43 1.31 ;
    RECT 113.91 1.41 114.12 1.62 ;
    RECT 114.28 1.005 114.55 2.125 ;
    RECT 114.83 1.24 115.04 1.31 ;
    RECT 115.78 0.915 115.99 2.125 ;
    RECT 110.59 1.41 110.8 1.62 ;
    RECT 110.96 1.005 111.23 2.125 ;
    RECT 111.51 1.24 111.72 1.31 ;
    RECT 112.46 0.915 112.67 2.125 ;
    RECT 107.27 1.41 107.48 1.62 ;
    RECT 107.64 1.005 107.91 2.125 ;
    RECT 108.19 1.24 108.4 1.31 ;
    RECT 109.14 0.915 109.35 2.125 ;
    RECT 5.27 2.055 5.48 2.125 ;
    RECT 103.95 1.41 104.16 1.62 ;
    RECT 104.32 1.005 104.59 2.125 ;
    RECT 104.87 1.24 105.08 1.31 ;
    RECT 105.82 0.915 106.03 2.125 ;
    RECT 5.27 1.742 5.48 1.812 ;
    RECT 100.63 1.41 100.84 1.62 ;
    RECT 101.0 1.005 101.27 2.125 ;
    RECT 101.55 1.24 101.76 1.31 ;
    RECT 102.5 0.915 102.71 2.125 ;
    RECT 55.07 11.325 55.28 11.395 ;
    RECT 72.16 10.805 72.37 10.875 ;
    RECT 38.96 11.065 39.17 11.135 ;
    RECT 22.36 10.805 22.57 10.875 ;
    RECT 148.52 11.065 148.73 11.135 ;
    RECT 54.61 11.325 54.82 11.395 ;
    RECT 108.19 11.325 108.4 11.395 ;
    RECT 107.73 11.325 107.94 11.395 ;
    RECT 68.84 10.805 69.05 10.875 ;
    RECT 35.64 11.065 35.85 11.135 ;
    RECT 19.04 10.805 19.25 10.875 ;
    RECT 145.2 11.065 145.41 11.135 ;
    RECT 51.75 11.325 51.96 11.395 ;
    RECT 51.29 11.325 51.5 11.395 ;
    RECT 131.92 10.805 132.13 10.875 ;
    RECT 104.87 11.325 105.08 11.395 ;
    RECT 98.72 11.065 98.93 11.135 ;
    RECT 104.41 11.325 104.62 11.395 ;
    RECT 164.63 11.325 164.84 11.395 ;
    RECT 141.88 11.065 142.09 11.135 ;
    RECT 164.17 11.325 164.38 11.395 ;
    RECT 48.43 11.325 48.64 11.395 ;
    RECT 47.97 11.325 48.18 11.395 ;
    RECT 128.6 10.805 128.81 10.875 ;
    RECT 15.72 10.805 15.93 10.875 ;
    RECT 101.55 11.325 101.76 11.395 ;
    RECT 101.09 11.325 101.3 11.395 ;
    RECT 138.56 11.065 138.77 11.135 ;
    RECT 161.31 11.325 161.52 11.395 ;
    RECT 160.85 11.325 161.06 11.395 ;
    RECT 45.11 11.325 45.32 11.395 ;
    RECT 44.65 11.325 44.86 11.395 ;
    RECT 170.345 10.545 170.565 10.615 ;
    RECT 167.025 10.545 167.245 10.615 ;
    RECT 95.4 11.065 95.61 11.135 ;
    RECT 125.28 10.805 125.49 10.875 ;
    RECT 12.4 10.805 12.61 10.875 ;
    RECT 65.52 10.805 65.73 10.875 ;
    RECT 163.705 10.545 163.925 10.615 ;
    RECT 160.385 10.545 160.605 10.615 ;
    RECT 157.065 10.545 157.285 10.615 ;
    RECT 153.745 10.545 153.965 10.615 ;
    RECT 150.425 10.545 150.645 10.615 ;
    RECT 147.105 10.545 147.325 10.615 ;
    RECT 143.785 10.545 144.005 10.615 ;
    RECT 135.24 11.065 135.45 11.135 ;
    RECT 140.465 10.545 140.685 10.615 ;
    RECT 75.48 11.065 75.69 11.135 ;
    RECT 137.145 10.545 137.365 10.615 ;
    RECT 157.99 11.325 158.2 11.395 ;
    RECT 133.825 10.545 134.045 10.615 ;
    RECT 157.53 11.325 157.74 11.395 ;
    RECT 41.79 11.325 42.0 11.395 ;
    RECT 41.33 11.325 41.54 11.395 ;
    RECT 92.08 11.065 92.29 11.135 ;
    RECT 121.96 10.805 122.17 10.875 ;
    RECT 9.08 10.805 9.29 10.875 ;
    RECT 62.2 10.805 62.41 10.875 ;
    RECT 130.505 10.545 130.725 10.615 ;
    RECT 127.185 10.545 127.405 10.615 ;
    RECT 123.865 10.545 124.085 10.615 ;
    RECT 120.545 10.545 120.765 10.615 ;
    RECT 117.225 10.545 117.445 10.615 ;
    RECT 113.905 10.545 114.125 10.615 ;
    RECT 110.585 10.545 110.805 10.615 ;
    RECT 107.265 10.545 107.485 10.615 ;
    RECT 103.945 10.545 104.165 10.615 ;
    RECT 31.83 11.325 32.04 11.395 ;
    RECT 100.625 10.545 100.845 10.615 ;
    RECT 31.37 11.325 31.58 11.395 ;
    RECT 72.16 11.065 72.37 11.135 ;
    RECT 154.67 11.325 154.88 11.395 ;
    RECT 38.47 11.325 38.68 11.395 ;
    RECT 88.76 11.065 88.97 11.135 ;
    RECT 118.64 10.805 118.85 10.875 ;
    RECT 5.76 10.805 5.97 10.875 ;
    RECT 97.305 10.545 97.525 10.615 ;
    RECT 93.985 10.545 94.205 10.615 ;
    RECT 90.665 10.545 90.885 10.615 ;
    RECT 58.88 10.805 59.09 10.875 ;
    RECT 87.345 10.545 87.565 10.615 ;
    RECT 84.025 10.545 84.245 10.615 ;
    RECT 154.21 11.325 154.42 11.395 ;
    RECT 80.705 10.545 80.925 10.615 ;
    RECT 77.385 10.545 77.605 10.615 ;
    RECT 38.01 11.325 38.22 11.395 ;
    RECT 74.065 10.545 74.285 10.615 ;
    RECT 70.745 10.545 70.965 10.615 ;
    RECT 67.425 10.545 67.645 10.615 ;
    RECT 28.51 11.325 28.72 11.395 ;
    RECT 28.05 11.325 28.26 11.395 ;
    RECT 68.84 11.065 69.05 11.135 ;
    RECT 98.23 11.325 98.44 11.395 ;
    RECT 97.77 11.325 97.98 11.395 ;
    RECT 85.44 11.065 85.65 11.135 ;
    RECT 64.105 10.545 64.325 10.615 ;
    RECT 2.44 10.805 2.65 10.875 ;
    RECT 60.785 10.545 61.005 10.615 ;
    RECT 57.465 10.545 57.685 10.615 ;
    RECT 54.145 10.545 54.365 10.615 ;
    RECT 50.825 10.545 51.045 10.615 ;
    RECT 47.505 10.545 47.725 10.615 ;
    RECT 44.185 10.545 44.405 10.615 ;
    RECT 55.56 10.805 55.77 10.875 ;
    RECT 40.865 10.545 41.085 10.615 ;
    RECT 37.545 10.545 37.765 10.615 ;
    RECT 151.35 11.325 151.56 11.395 ;
    RECT 34.225 10.545 34.445 10.615 ;
    RECT 150.89 11.325 151.1 11.395 ;
    RECT 35.15 11.325 35.36 11.395 ;
    RECT 34.69 11.325 34.9 11.395 ;
    RECT 165.12 10.805 165.33 10.875 ;
    RECT 32.32 11.065 32.53 11.135 ;
    RECT 25.19 11.325 25.4 11.395 ;
    RECT 24.73 11.325 24.94 11.395 ;
    RECT 131.92 11.065 132.13 11.135 ;
    RECT 94.91 11.325 95.12 11.395 ;
    RECT 94.45 11.325 94.66 11.395 ;
    RECT 115.32 10.805 115.53 10.875 ;
    RECT 82.12 11.065 82.33 11.135 ;
    RECT 52.24 10.805 52.45 10.875 ;
    RECT 148.03 11.325 148.24 11.395 ;
    RECT 147.57 11.325 147.78 11.395 ;
    RECT 161.8 10.805 162.01 10.875 ;
    RECT 171.76 10.805 171.97 10.875 ;
    RECT 21.87 11.325 22.08 11.395 ;
    RECT 91.59 11.325 91.8 11.395 ;
    RECT 112.0 10.805 112.21 10.875 ;
    RECT 91.13 11.325 91.34 11.395 ;
    RECT 78.8 11.065 79.01 11.135 ;
    RECT 29.0 11.065 29.21 11.135 ;
    RECT 21.41 11.325 21.62 11.395 ;
    RECT 128.6 11.065 128.81 11.135 ;
    RECT 144.71 11.325 144.92 11.395 ;
    RECT 144.25 11.325 144.46 11.395 ;
    RECT 158.48 10.805 158.69 10.875 ;
    RECT 168.44 10.805 168.65 10.875 ;
    RECT 65.52 11.065 65.73 11.135 ;
    RECT 98.72 10.805 98.93 10.875 ;
    RECT 108.68 10.805 108.89 10.875 ;
    RECT 88.27 11.325 88.48 11.395 ;
    RECT 48.92 10.805 49.13 10.875 ;
    RECT 25.68 11.065 25.89 11.135 ;
    RECT 18.55 11.325 18.76 11.395 ;
    RECT 18.09 11.325 18.3 11.395 ;
    RECT 125.28 11.065 125.49 11.135 ;
    RECT 141.39 11.325 141.6 11.395 ;
    RECT 155.16 10.805 155.37 10.875 ;
    RECT 140.93 11.325 141.14 11.395 ;
    RECT 87.81 11.325 88.02 11.395 ;
    RECT 95.4 10.805 95.61 10.875 ;
    RECT 105.36 10.805 105.57 10.875 ;
    RECT 45.6 10.805 45.81 10.875 ;
    RECT 22.36 11.065 22.57 11.135 ;
    RECT 15.23 11.325 15.44 11.395 ;
    RECT 14.77 11.325 14.98 11.395 ;
    RECT 121.96 11.065 122.17 11.135 ;
    RECT 131.43 11.325 131.64 11.395 ;
    RECT 62.2 11.065 62.41 11.135 ;
    RECT 130.97 11.325 131.18 11.395 ;
    RECT 151.84 10.805 152.05 10.875 ;
    RECT 138.07 11.325 138.28 11.395 ;
    RECT 84.95 11.325 85.16 11.395 ;
    RECT 84.49 11.325 84.7 11.395 ;
    RECT 92.08 10.805 92.29 10.875 ;
    RECT 102.04 10.805 102.25 10.875 ;
    RECT 42.28 10.805 42.49 10.875 ;
    RECT 30.905 10.545 31.125 10.615 ;
    RECT 27.585 10.545 27.805 10.615 ;
    RECT 24.265 10.545 24.485 10.615 ;
    RECT 20.945 10.545 21.165 10.615 ;
    RECT 19.04 11.065 19.25 11.135 ;
    RECT 17.625 10.545 17.845 10.615 ;
    RECT 14.305 10.545 14.525 10.615 ;
    RECT 10.985 10.545 11.205 10.615 ;
    RECT 7.665 10.545 7.885 10.615 ;
    RECT 4.345 10.545 4.565 10.615 ;
    RECT 11.91 11.325 12.12 11.395 ;
    RECT 1.025 10.545 1.245 10.615 ;
    RECT 11.45 11.325 11.66 11.395 ;
    RECT 118.64 11.065 118.85 11.135 ;
    RECT 58.88 11.065 59.09 11.135 ;
    RECT 128.11 11.325 128.32 11.395 ;
    RECT 137.61 11.325 137.82 11.395 ;
    RECT 127.65 11.325 127.86 11.395 ;
    RECT 81.63 11.325 81.84 11.395 ;
    RECT 81.17 11.325 81.38 11.395 ;
    RECT 88.76 10.805 88.97 10.875 ;
    RECT 38.96 10.805 39.17 10.875 ;
    RECT 148.52 10.805 148.73 10.875 ;
    RECT 15.72 11.065 15.93 11.135 ;
    RECT 165.12 11.065 165.33 11.135 ;
    RECT 115.32 11.065 115.53 11.135 ;
    RECT 8.59 11.325 8.8 11.395 ;
    RECT 55.56 11.065 55.77 11.135 ;
    RECT 8.13 11.325 8.34 11.395 ;
    RECT 134.75 11.325 134.96 11.395 ;
    RECT 134.29 11.325 134.5 11.395 ;
    RECT 124.79 11.325 125.0 11.395 ;
    RECT 124.33 11.325 124.54 11.395 ;
    RECT 78.31 11.325 78.52 11.395 ;
    RECT 77.85 11.325 78.06 11.395 ;
    RECT 85.44 10.805 85.65 10.875 ;
    RECT 35.64 10.805 35.85 10.875 ;
    RECT 145.2 10.805 145.41 10.875 ;
    RECT 12.4 11.065 12.61 11.135 ;
    RECT 171.76 11.065 171.97 11.135 ;
    RECT 112.0 11.065 112.21 11.135 ;
    RECT 52.24 11.065 52.45 11.135 ;
    RECT 5.27 11.325 5.48 11.395 ;
    RECT 121.47 11.325 121.68 11.395 ;
    RECT 74.99 11.325 75.2 11.395 ;
    RECT 74.53 11.325 74.74 11.395 ;
    RECT 161.8 11.065 162.01 11.135 ;
    RECT 141.88 10.805 142.09 10.875 ;
    RECT 4.81 11.325 5.02 11.395 ;
    RECT 121.01 11.325 121.22 11.395 ;
    RECT 9.08 11.065 9.29 11.135 ;
    RECT 65.03 11.325 65.24 11.395 ;
    RECT 64.57 11.325 64.78 11.395 ;
    RECT 168.44 11.065 168.65 11.135 ;
    RECT 108.68 11.065 108.89 11.135 ;
    RECT 48.92 11.065 49.13 11.135 ;
    RECT 82.12 10.805 82.33 10.875 ;
    RECT 71.67 11.325 71.88 11.395 ;
    RECT 32.32 10.805 32.53 10.875 ;
    RECT 158.48 11.065 158.69 11.135 ;
    RECT 138.56 10.805 138.77 10.875 ;
    RECT 1.95 11.325 2.16 11.395 ;
    RECT 1.49 11.325 1.7 11.395 ;
    RECT 171.27 11.325 171.48 11.395 ;
    RECT 118.15 11.325 118.36 11.395 ;
    RECT 117.69 11.325 117.9 11.395 ;
    RECT 5.76 11.065 5.97 11.135 ;
    RECT 61.71 11.325 61.92 11.395 ;
    RECT 71.21 11.325 71.42 11.395 ;
    RECT 61.25 11.325 61.46 11.395 ;
    RECT 105.36 11.065 105.57 11.135 ;
    RECT 45.6 11.065 45.81 11.135 ;
    RECT 78.8 10.805 79.01 10.875 ;
    RECT 170.81 11.325 171.02 11.395 ;
    RECT 29.0 10.805 29.21 10.875 ;
    RECT 155.16 11.065 155.37 11.135 ;
    RECT 135.24 10.805 135.45 10.875 ;
    RECT 114.83 11.325 115.04 11.395 ;
    RECT 2.44 11.065 2.65 11.135 ;
    RECT 114.37 11.325 114.58 11.395 ;
    RECT 68.35 11.325 68.56 11.395 ;
    RECT 58.39 11.325 58.6 11.395 ;
    RECT 67.89 11.325 68.1 11.395 ;
    RECT 57.93 11.325 58.14 11.395 ;
    RECT 102.04 11.065 102.25 11.135 ;
    RECT 75.48 10.805 75.69 10.875 ;
    RECT 42.28 11.065 42.49 11.135 ;
    RECT 167.95 11.325 168.16 11.395 ;
    RECT 167.49 11.325 167.7 11.395 ;
    RECT 25.68 10.805 25.89 10.875 ;
    RECT 151.84 11.065 152.05 11.135 ;
    RECT 111.51 11.325 111.72 11.395 ;
    RECT 111.05 11.325 111.26 11.395 ;
    RECT 0.42 4.055 0.49 4.125 ;
    RECT 0.62 4.455 0.69 4.525 ;
    RECT 0.61 5.33 0.68 5.54 ;
    RECT 0.61 3.235 0.68 3.445 ;
    RECT 0.19 11.065 0.26 11.135 ;
    RECT 0.4 11.325 0.47 11.395 ;
    RECT 0.61 9.12 0.68 9.33 ;
    RECT 15.23 4.055 15.44 4.125 ;
    RECT 91.59 6.385 91.8 6.455 ;
    RECT 91.59 5.86 91.8 6.07 ;
    RECT 91.59 2.585 91.8 2.795 ;
    RECT 151.35 4.055 151.56 4.125 ;
    RECT 64.11 3.235 64.32 3.445 ;
    RECT 64.11 5.33 64.32 5.54 ;
    RECT 64.11 9.12 64.32 9.33 ;
    RECT 64.68 4.845 64.75 4.915 ;
    RECT 64.68 9.43 64.75 9.5 ;
    RECT 65.52 9.765 65.73 9.835 ;
    RECT 65.98 2.585 66.19 2.795 ;
    RECT 65.98 5.86 66.19 6.07 ;
    RECT 65.98 6.385 66.19 6.455 ;
    RECT 65.98 7.28 66.19 7.35 ;
    RECT 60.79 3.235 61.0 3.445 ;
    RECT 60.79 5.33 61.0 5.54 ;
    RECT 60.79 9.12 61.0 9.33 ;
    RECT 61.36 4.845 61.43 4.915 ;
    RECT 61.36 9.43 61.43 9.5 ;
    RECT 62.2 9.765 62.41 9.835 ;
    RECT 62.66 2.585 62.87 2.795 ;
    RECT 62.66 5.86 62.87 6.07 ;
    RECT 62.66 6.385 62.87 6.455 ;
    RECT 62.66 7.28 62.87 7.35 ;
    RECT 57.47 3.235 57.68 3.445 ;
    RECT 57.47 5.33 57.68 5.54 ;
    RECT 57.47 9.12 57.68 9.33 ;
    RECT 58.04 4.845 58.11 4.915 ;
    RECT 58.04 9.43 58.11 9.5 ;
    RECT 58.88 9.765 59.09 9.835 ;
    RECT 59.34 2.585 59.55 2.795 ;
    RECT 59.34 5.86 59.55 6.07 ;
    RECT 59.34 6.385 59.55 6.455 ;
    RECT 59.34 7.28 59.55 7.35 ;
    RECT 121.47 7.28 121.68 7.35 ;
    RECT 151.35 7.28 151.56 7.35 ;
    RECT 54.15 3.235 54.36 3.445 ;
    RECT 54.15 5.33 54.36 5.54 ;
    RECT 54.15 9.12 54.36 9.33 ;
    RECT 54.72 4.845 54.79 4.915 ;
    RECT 54.72 9.43 54.79 9.5 ;
    RECT 55.56 9.765 55.77 9.835 ;
    RECT 56.02 2.585 56.23 2.795 ;
    RECT 56.02 5.86 56.23 6.07 ;
    RECT 56.02 6.385 56.23 6.455 ;
    RECT 56.02 7.28 56.23 7.35 ;
    RECT 121.47 6.385 121.68 6.455 ;
    RECT 151.35 6.385 151.56 6.455 ;
    RECT 50.83 3.235 51.04 3.445 ;
    RECT 50.83 5.33 51.04 5.54 ;
    RECT 50.83 9.12 51.04 9.33 ;
    RECT 51.4 4.845 51.47 4.915 ;
    RECT 51.4 9.43 51.47 9.5 ;
    RECT 52.24 9.765 52.45 9.835 ;
    RECT 52.7 2.585 52.91 2.795 ;
    RECT 52.7 5.86 52.91 6.07 ;
    RECT 52.7 6.385 52.91 6.455 ;
    RECT 52.7 7.28 52.91 7.35 ;
    RECT 121.47 5.86 121.68 6.07 ;
    RECT 151.35 5.86 151.56 6.07 ;
    RECT 123.87 4.455 124.08 4.525 ;
    RECT 47.51 3.235 47.72 3.445 ;
    RECT 47.51 5.33 47.72 5.54 ;
    RECT 47.51 9.12 47.72 9.33 ;
    RECT 48.08 4.845 48.15 4.915 ;
    RECT 48.08 9.43 48.15 9.5 ;
    RECT 48.92 9.765 49.13 9.835 ;
    RECT 49.38 2.585 49.59 2.795 ;
    RECT 49.38 5.86 49.59 6.07 ;
    RECT 49.38 6.385 49.59 6.455 ;
    RECT 49.38 7.28 49.59 7.35 ;
    RECT 93.99 4.455 94.2 4.525 ;
    RECT 121.47 2.585 121.68 2.795 ;
    RECT 44.19 3.235 44.4 3.445 ;
    RECT 44.19 5.33 44.4 5.54 ;
    RECT 44.19 9.12 44.4 9.33 ;
    RECT 44.76 4.845 44.83 4.915 ;
    RECT 44.76 9.43 44.83 9.5 ;
    RECT 45.6 9.765 45.81 9.835 ;
    RECT 46.06 2.585 46.27 2.795 ;
    RECT 46.06 5.86 46.27 6.07 ;
    RECT 46.06 6.385 46.27 6.455 ;
    RECT 46.06 7.28 46.27 7.35 ;
    RECT 40.87 3.235 41.08 3.445 ;
    RECT 40.87 5.33 41.08 5.54 ;
    RECT 40.87 9.12 41.08 9.33 ;
    RECT 41.44 4.845 41.51 4.915 ;
    RECT 41.44 9.43 41.51 9.5 ;
    RECT 42.28 9.765 42.49 9.835 ;
    RECT 42.74 2.585 42.95 2.795 ;
    RECT 42.74 5.86 42.95 6.07 ;
    RECT 42.74 6.385 42.95 6.455 ;
    RECT 42.74 7.28 42.95 7.35 ;
    RECT 37.55 3.235 37.76 3.445 ;
    RECT 37.55 5.33 37.76 5.54 ;
    RECT 37.55 9.12 37.76 9.33 ;
    RECT 38.12 4.845 38.19 4.915 ;
    RECT 38.12 9.43 38.19 9.5 ;
    RECT 38.96 9.765 39.17 9.835 ;
    RECT 39.42 2.585 39.63 2.795 ;
    RECT 39.42 5.86 39.63 6.07 ;
    RECT 39.42 6.385 39.63 6.455 ;
    RECT 39.42 7.28 39.63 7.35 ;
    RECT 34.23 3.235 34.44 3.445 ;
    RECT 34.23 5.33 34.44 5.54 ;
    RECT 34.23 9.12 34.44 9.33 ;
    RECT 34.8 4.845 34.87 4.915 ;
    RECT 34.8 9.43 34.87 9.5 ;
    RECT 35.64 9.765 35.85 9.835 ;
    RECT 36.1 2.585 36.31 2.795 ;
    RECT 36.1 5.86 36.31 6.07 ;
    RECT 36.1 6.385 36.31 6.455 ;
    RECT 36.1 7.28 36.31 7.35 ;
    RECT 100.63 4.455 100.84 4.525 ;
    RECT 74.99 4.055 75.2 4.125 ;
    RECT 27.59 4.455 27.8 4.525 ;
    RECT 50.83 4.455 51.04 4.525 ;
    RECT 151.35 2.585 151.56 2.795 ;
    RECT 18.55 7.28 18.76 7.35 ;
    RECT 1.95 4.055 2.16 4.125 ;
    RECT 18.55 6.385 18.76 6.455 ;
    RECT 18.55 5.86 18.76 6.07 ;
    RECT 55.07 4.055 55.28 4.125 ;
    RECT 48.43 7.28 48.64 7.35 ;
    RECT 48.43 6.385 48.64 6.455 ;
    RECT 131.43 4.055 131.64 4.125 ;
    RECT 48.43 5.86 48.64 6.07 ;
    RECT 48.43 2.585 48.64 2.795 ;
    RECT 78.31 7.28 78.52 7.35 ;
    RECT 78.31 6.385 78.52 6.455 ;
    RECT 18.55 2.585 18.76 2.795 ;
    RECT 78.31 5.86 78.52 6.07 ;
    RECT 78.31 2.585 78.52 2.795 ;
    RECT 138.07 4.055 138.28 4.125 ;
    RECT 163.71 4.455 163.92 4.525 ;
    RECT 120.55 4.455 120.76 4.525 ;
    RECT 80.71 4.455 80.92 4.525 ;
    RECT 108.19 7.28 108.4 7.35 ;
    RECT 118.15 4.055 118.36 4.125 ;
    RECT 170.35 4.455 170.56 4.525 ;
    RECT 30.91 3.235 31.12 3.445 ;
    RECT 30.91 5.33 31.12 5.54 ;
    RECT 30.91 9.12 31.12 9.33 ;
    RECT 31.48 4.845 31.55 4.915 ;
    RECT 31.48 9.43 31.55 9.5 ;
    RECT 32.32 9.765 32.53 9.835 ;
    RECT 32.78 2.585 32.99 2.795 ;
    RECT 32.78 5.86 32.99 6.07 ;
    RECT 32.78 6.385 32.99 6.455 ;
    RECT 32.78 7.28 32.99 7.35 ;
    RECT 27.59 3.235 27.8 3.445 ;
    RECT 27.59 5.33 27.8 5.54 ;
    RECT 27.59 9.12 27.8 9.33 ;
    RECT 28.16 4.845 28.23 4.915 ;
    RECT 28.16 9.43 28.23 9.5 ;
    RECT 29.0 9.765 29.21 9.835 ;
    RECT 29.46 2.585 29.67 2.795 ;
    RECT 29.46 5.86 29.67 6.07 ;
    RECT 29.46 6.385 29.67 6.455 ;
    RECT 29.46 7.28 29.67 7.35 ;
    RECT 24.27 3.235 24.48 3.445 ;
    RECT 24.27 5.33 24.48 5.54 ;
    RECT 24.27 9.12 24.48 9.33 ;
    RECT 24.84 4.845 24.91 4.915 ;
    RECT 24.84 9.43 24.91 9.5 ;
    RECT 25.68 9.765 25.89 9.835 ;
    RECT 26.14 2.585 26.35 2.795 ;
    RECT 26.14 5.86 26.35 6.07 ;
    RECT 26.14 6.385 26.35 6.455 ;
    RECT 26.14 7.28 26.35 7.35 ;
    RECT 14.31 4.455 14.52 4.525 ;
    RECT 37.55 4.455 37.76 4.525 ;
    RECT 20.95 3.235 21.16 3.445 ;
    RECT 20.95 5.33 21.16 5.54 ;
    RECT 20.95 9.12 21.16 9.33 ;
    RECT 21.52 4.845 21.59 4.915 ;
    RECT 21.52 9.43 21.59 9.5 ;
    RECT 22.36 9.765 22.57 9.835 ;
    RECT 22.82 2.585 23.03 2.795 ;
    RECT 22.82 5.86 23.03 6.07 ;
    RECT 22.82 6.385 23.03 6.455 ;
    RECT 22.82 7.28 23.03 7.35 ;
    RECT 17.63 3.235 17.84 3.445 ;
    RECT 17.63 5.33 17.84 5.54 ;
    RECT 17.63 9.12 17.84 9.33 ;
    RECT 18.2 4.845 18.27 4.915 ;
    RECT 18.2 9.43 18.27 9.5 ;
    RECT 19.04 9.765 19.25 9.835 ;
    RECT 19.5 2.585 19.71 2.795 ;
    RECT 19.5 5.86 19.71 6.07 ;
    RECT 19.5 6.385 19.71 6.455 ;
    RECT 19.5 7.28 19.71 7.35 ;
    RECT 14.31 3.235 14.52 3.445 ;
    RECT 14.31 5.33 14.52 5.54 ;
    RECT 14.31 9.12 14.52 9.33 ;
    RECT 14.88 4.845 14.95 4.915 ;
    RECT 14.88 9.43 14.95 9.5 ;
    RECT 15.72 9.765 15.93 9.835 ;
    RECT 16.18 2.585 16.39 2.795 ;
    RECT 16.18 5.86 16.39 6.07 ;
    RECT 16.18 6.385 16.39 6.455 ;
    RECT 16.18 7.28 16.39 7.35 ;
    RECT 10.99 3.235 11.2 3.445 ;
    RECT 10.99 5.33 11.2 5.54 ;
    RECT 10.99 9.12 11.2 9.33 ;
    RECT 11.56 4.845 11.63 4.915 ;
    RECT 11.56 9.43 11.63 9.5 ;
    RECT 12.4 9.765 12.61 9.835 ;
    RECT 12.86 2.585 13.07 2.795 ;
    RECT 12.86 5.86 13.07 6.07 ;
    RECT 12.86 6.385 13.07 6.455 ;
    RECT 12.86 7.28 13.07 7.35 ;
    RECT 41.79 4.055 42.0 4.125 ;
    RECT 7.67 3.235 7.88 3.445 ;
    RECT 7.67 5.33 7.88 5.54 ;
    RECT 7.67 9.12 7.88 9.33 ;
    RECT 8.24 4.845 8.31 4.915 ;
    RECT 8.24 9.43 8.31 9.5 ;
    RECT 9.08 9.765 9.29 9.835 ;
    RECT 9.54 2.585 9.75 2.795 ;
    RECT 9.54 5.86 9.75 6.07 ;
    RECT 9.54 6.385 9.75 6.455 ;
    RECT 9.54 7.28 9.75 7.35 ;
    RECT 4.35 3.235 4.56 3.445 ;
    RECT 4.35 5.33 4.56 5.54 ;
    RECT 4.35 9.12 4.56 9.33 ;
    RECT 4.92 4.845 4.99 4.915 ;
    RECT 4.92 9.43 4.99 9.5 ;
    RECT 5.76 9.765 5.97 9.835 ;
    RECT 6.22 2.585 6.43 2.795 ;
    RECT 6.22 5.86 6.43 6.07 ;
    RECT 6.22 6.385 6.43 6.455 ;
    RECT 6.22 7.28 6.43 7.35 ;
    RECT 138.07 7.28 138.28 7.35 ;
    RECT 108.19 6.385 108.4 6.455 ;
    RECT 138.07 6.385 138.28 6.455 ;
    RECT 108.19 5.86 108.4 6.07 ;
    RECT 138.07 5.86 138.28 6.07 ;
    RECT 108.19 2.585 108.4 2.795 ;
    RECT 138.07 2.585 138.28 2.795 ;
    RECT 167.95 7.28 168.16 7.35 ;
    RECT 131.43 7.28 131.64 7.35 ;
    RECT 167.95 6.385 168.16 6.455 ;
    RECT 160.39 4.455 160.6 4.525 ;
    RECT 131.43 6.385 131.64 6.455 ;
    RECT 167.95 5.86 168.16 6.07 ;
    RECT 117.23 4.455 117.44 4.525 ;
    RECT 131.43 5.86 131.64 6.07 ;
    RECT 131.43 2.585 131.64 2.795 ;
    RECT 98.23 4.055 98.44 4.125 ;
    RECT 161.31 7.28 161.52 7.35 ;
    RECT 161.31 6.385 161.52 6.455 ;
    RECT 161.31 5.86 161.52 6.07 ;
    RECT 5.27 7.28 5.48 7.35 ;
    RECT 161.31 2.585 161.52 2.795 ;
    RECT 5.27 6.385 5.48 6.455 ;
    RECT 35.15 7.28 35.36 7.35 ;
    RECT 5.27 5.86 5.48 6.07 ;
    RECT 35.15 6.385 35.36 6.455 ;
    RECT 5.27 2.585 5.48 2.795 ;
    RECT 35.15 5.86 35.36 6.07 ;
    RECT 25.19 4.055 25.4 4.125 ;
    RECT 104.87 4.055 105.08 4.125 ;
    RECT 167.95 2.585 168.16 2.795 ;
    RECT 58.39 7.28 58.6 7.35 ;
    RECT 161.31 4.055 161.52 4.125 ;
    RECT 167.03 4.455 167.24 4.525 ;
    RECT 60.79 4.455 61.0 4.525 ;
    RECT 84.95 4.055 85.16 4.125 ;
    RECT 157.07 4.455 157.28 4.525 ;
    RECT 113.91 4.455 114.12 4.525 ;
    RECT 28.51 7.28 28.72 7.35 ;
    RECT 35.15 2.585 35.36 2.795 ;
    RECT 28.51 6.385 28.72 6.455 ;
    RECT 28.51 5.86 28.72 6.07 ;
    RECT 28.51 2.585 28.72 2.795 ;
    RECT 67.43 4.455 67.64 4.525 ;
    RECT 167.95 4.055 168.16 4.125 ;
    RECT 11.91 4.055 12.12 4.125 ;
    RECT 58.39 6.385 58.6 6.455 ;
    RECT 58.39 5.86 58.6 6.07 ;
    RECT 58.39 2.585 58.6 2.795 ;
    RECT 1.03 4.455 1.24 4.525 ;
    RECT 88.27 7.28 88.48 7.35 ;
    RECT 148.03 4.055 148.24 4.125 ;
    RECT 88.27 6.385 88.48 6.455 ;
    RECT 88.27 5.86 88.48 6.07 ;
    RECT 88.27 2.585 88.48 2.795 ;
    RECT 65.03 4.055 65.24 4.125 ;
    RECT 118.15 7.28 118.36 7.35 ;
    RECT 118.15 6.385 118.36 6.455 ;
    RECT 90.67 4.455 90.88 4.525 ;
    RECT 118.15 5.86 118.36 6.07 ;
    RECT 71.67 4.055 71.88 4.125 ;
    RECT 24.27 4.455 24.48 4.525 ;
    RECT 47.51 4.455 47.72 4.525 ;
    RECT 148.03 7.28 148.24 7.35 ;
    RECT 153.75 4.455 153.96 4.525 ;
    RECT 148.03 6.385 148.24 6.455 ;
    RECT 110.59 4.455 110.8 4.525 ;
    RECT 148.03 5.86 148.24 6.07 ;
    RECT 118.15 2.585 118.36 2.795 ;
    RECT 148.03 2.585 148.24 2.795 ;
    RECT 51.75 4.055 51.96 4.125 ;
    RECT 128.11 4.055 128.32 4.125 ;
    RECT 45.11 7.28 45.32 7.35 ;
    RECT 45.11 6.385 45.32 6.455 ;
    RECT 45.11 5.86 45.32 6.07 ;
    RECT 45.11 2.585 45.32 2.795 ;
    RECT 15.23 7.28 15.44 7.35 ;
    RECT 15.23 6.385 15.44 6.455 ;
    RECT 74.99 7.28 75.2 7.35 ;
    RECT 134.75 4.055 134.96 4.125 ;
    RECT 15.23 5.86 15.44 6.07 ;
    RECT 15.23 2.585 15.44 2.795 ;
    RECT 150.43 4.455 150.64 4.525 ;
    RECT 107.27 4.455 107.48 4.525 ;
    RECT 114.83 4.055 115.04 4.125 ;
    RECT 74.99 6.385 75.2 6.455 ;
    RECT 74.99 5.86 75.2 6.07 ;
    RECT 74.99 2.585 75.2 2.795 ;
    RECT 38.47 4.055 38.68 4.125 ;
    RECT 77.39 4.455 77.6 4.525 ;
    RECT 104.87 7.28 105.08 7.35 ;
    RECT 134.75 7.28 134.96 7.35 ;
    RECT 104.87 6.385 105.08 6.455 ;
    RECT 134.75 6.385 134.96 6.455 ;
    RECT 104.87 5.86 105.08 6.07 ;
    RECT 134.75 5.86 134.96 6.07 ;
    RECT 104.87 2.585 105.08 2.795 ;
    RECT 147.11 4.455 147.32 4.525 ;
    RECT 98.23 7.28 98.44 7.35 ;
    RECT 128.11 7.28 128.32 7.35 ;
    RECT 103.95 4.455 104.16 4.525 ;
    RECT 10.99 4.455 11.2 4.525 ;
    RECT 98.23 6.385 98.44 6.455 ;
    RECT 128.11 6.385 128.32 6.455 ;
    RECT 34.23 4.455 34.44 4.525 ;
    RECT 98.23 5.86 98.44 6.07 ;
    RECT 128.11 5.86 128.32 6.07 ;
    RECT 98.23 2.585 98.44 2.795 ;
    RECT 128.11 2.585 128.32 2.795 ;
    RECT 94.91 4.055 95.12 4.125 ;
    RECT 134.75 2.585 134.96 2.795 ;
    RECT 157.99 7.28 158.2 7.35 ;
    RECT 1.95 7.28 2.16 7.35 ;
    RECT 1.95 6.385 2.16 6.455 ;
    RECT 1.95 5.86 2.16 6.07 ;
    RECT 21.87 4.055 22.08 4.125 ;
    RECT 101.55 4.055 101.76 4.125 ;
    RECT 157.99 4.055 158.2 4.125 ;
    RECT 57.47 4.455 57.68 4.525 ;
    RECT 157.99 6.385 158.2 6.455 ;
    RECT 81.63 4.055 81.84 4.125 ;
    RECT 157.99 5.86 158.2 6.07 ;
    RECT 157.99 2.585 158.2 2.795 ;
    RECT 1.95 2.585 2.16 2.795 ;
    RECT 25.19 7.28 25.4 7.35 ;
    RECT 55.07 7.28 55.28 7.35 ;
    RECT 55.07 6.385 55.28 6.455 ;
    RECT 55.07 5.86 55.28 6.07 ;
    RECT 55.07 2.585 55.28 2.795 ;
    RECT 143.79 4.455 144.0 4.525 ;
    RECT 144.71 4.055 144.92 4.125 ;
    RECT 25.19 6.385 25.4 6.455 ;
    RECT 25.19 5.86 25.4 6.07 ;
    RECT 84.95 7.28 85.16 7.35 ;
    RECT 25.19 2.585 25.4 2.795 ;
    RECT 84.95 6.385 85.16 6.455 ;
    RECT 84.95 5.86 85.16 6.07 ;
    RECT 8.59 4.055 8.8 4.125 ;
    RECT 61.71 4.055 61.92 4.125 ;
    RECT 68.35 4.055 68.56 4.125 ;
    RECT 84.95 2.585 85.16 2.795 ;
    RECT 140.47 4.455 140.68 4.525 ;
    RECT 114.83 7.28 115.04 7.35 ;
    RECT 144.71 7.28 144.92 7.35 ;
    RECT 87.35 4.455 87.56 4.525 ;
    RECT 114.83 6.385 115.04 6.455 ;
    RECT 144.71 6.385 144.92 6.455 ;
    RECT 114.83 5.86 115.04 6.07 ;
    RECT 144.71 5.86 144.92 6.07 ;
    RECT 114.83 2.585 115.04 2.795 ;
    RECT 144.71 2.585 144.92 2.795 ;
    RECT 48.43 4.055 48.64 4.125 ;
    RECT 124.79 4.055 125.0 4.125 ;
    RECT 20.95 4.455 21.16 4.525 ;
    RECT 44.19 4.455 44.4 4.525 ;
    RECT 41.79 7.28 42.0 7.35 ;
    RECT 11.91 7.28 12.12 7.35 ;
    RECT 11.91 6.385 12.12 6.455 ;
    RECT 11.91 5.86 12.12 6.07 ;
    RECT 11.91 2.585 12.12 2.795 ;
    RECT 137.15 4.455 137.36 4.525 ;
    RECT 170.35 3.235 170.56 3.445 ;
    RECT 170.35 5.33 170.56 5.54 ;
    RECT 170.35 9.12 170.56 9.33 ;
    RECT 170.92 4.845 170.99 4.915 ;
    RECT 170.92 9.43 170.99 9.5 ;
    RECT 171.76 9.765 171.97 9.835 ;
    RECT 172.22 2.585 172.43 2.795 ;
    RECT 172.22 5.86 172.43 6.07 ;
    RECT 172.22 6.385 172.43 6.455 ;
    RECT 172.22 7.28 172.43 7.35 ;
    RECT 111.51 4.055 111.72 4.125 ;
    RECT 1.03 3.235 1.24 3.445 ;
    RECT 1.03 5.33 1.24 5.54 ;
    RECT 1.03 9.12 1.24 9.33 ;
    RECT 1.6 4.845 1.67 4.915 ;
    RECT 1.6 9.43 1.67 9.5 ;
    RECT 2.44 9.765 2.65 9.835 ;
    RECT 2.9 2.585 3.11 2.795 ;
    RECT 2.9 5.86 3.11 6.07 ;
    RECT 2.9 6.385 3.11 6.455 ;
    RECT 2.9 7.28 3.11 7.35 ;
    RECT 71.67 7.28 71.88 7.35 ;
    RECT 41.79 6.385 42.0 6.455 ;
    RECT 71.67 6.385 71.88 6.455 ;
    RECT 41.79 5.86 42.0 6.07 ;
    RECT 71.67 5.86 71.88 6.07 ;
    RECT 41.79 2.585 42.0 2.795 ;
    RECT 71.67 2.585 71.88 2.795 ;
    RECT 35.15 4.055 35.36 4.125 ;
    RECT 31.83 4.055 32.04 4.125 ;
    RECT 74.07 4.455 74.28 4.525 ;
    RECT 101.55 7.28 101.76 7.35 ;
    RECT 101.55 6.385 101.76 6.455 ;
    RECT 65.03 7.28 65.24 7.35 ;
    RECT 101.55 5.86 101.76 6.07 ;
    RECT 65.03 6.385 65.24 6.455 ;
    RECT 65.03 5.86 65.24 6.07 ;
    RECT 65.03 2.585 65.24 2.795 ;
    RECT 7.67 4.455 7.88 4.525 ;
    RECT 94.91 7.28 95.12 7.35 ;
    RECT 124.79 7.28 125.0 7.35 ;
    RECT 94.91 6.385 95.12 6.455 ;
    RECT 94.91 5.86 95.12 6.07 ;
    RECT 91.59 4.055 91.8 4.125 ;
    RECT 94.91 2.585 95.12 2.795 ;
    RECT 101.55 2.585 101.76 2.795 ;
    RECT 18.55 4.055 18.76 4.125 ;
    RECT 133.83 4.455 134.04 4.525 ;
    RECT 154.67 4.055 154.88 4.125 ;
    RECT 78.31 4.055 78.52 4.125 ;
    RECT 154.67 7.28 154.88 7.35 ;
    RECT 124.79 6.385 125.0 6.455 ;
    RECT 154.67 6.385 154.88 6.455 ;
    RECT 124.79 5.86 125.0 6.07 ;
    RECT 154.67 5.86 154.88 6.07 ;
    RECT 124.79 2.585 125.0 2.795 ;
    RECT 154.67 2.585 154.88 2.795 ;
    RECT 97.31 4.455 97.52 4.525 ;
    RECT 51.75 7.28 51.96 7.35 ;
    RECT 51.75 6.385 51.96 6.455 ;
    RECT 30.91 4.455 31.12 4.525 ;
    RECT 51.75 5.86 51.96 6.07 ;
    RECT 54.15 4.455 54.36 4.525 ;
    RECT 21.87 7.28 22.08 7.35 ;
    RECT 21.87 6.385 22.08 6.455 ;
    RECT 21.87 5.86 22.08 6.07 ;
    RECT 21.87 2.585 22.08 2.795 ;
    RECT 5.27 4.055 5.48 4.125 ;
    RECT 58.39 4.055 58.6 4.125 ;
    RECT 51.75 2.585 51.96 2.795 ;
    RECT 81.63 7.28 81.84 7.35 ;
    RECT 81.63 6.385 81.84 6.455 ;
    RECT 81.63 5.86 81.84 6.07 ;
    RECT 167.03 3.235 167.24 3.445 ;
    RECT 167.03 5.33 167.24 5.54 ;
    RECT 167.03 9.12 167.24 9.33 ;
    RECT 167.6 4.845 167.67 4.915 ;
    RECT 167.6 9.43 167.67 9.5 ;
    RECT 168.44 9.765 168.65 9.835 ;
    RECT 168.9 2.585 169.11 2.795 ;
    RECT 168.9 5.86 169.11 6.07 ;
    RECT 168.9 6.385 169.11 6.455 ;
    RECT 168.9 7.28 169.11 7.35 ;
    RECT 81.63 2.585 81.84 2.795 ;
    RECT 141.39 4.055 141.6 4.125 ;
    RECT 84.03 4.455 84.24 4.525 ;
    RECT 111.51 7.28 111.72 7.35 ;
    RECT 141.39 7.28 141.6 7.35 ;
    RECT 111.51 6.385 111.72 6.455 ;
    RECT 45.11 4.055 45.32 4.125 ;
    RECT 111.51 5.86 111.72 6.07 ;
    RECT 111.51 2.585 111.72 2.795 ;
    RECT 121.47 4.055 121.68 4.125 ;
    RECT 163.71 3.235 163.92 3.445 ;
    RECT 163.71 5.33 163.92 5.54 ;
    RECT 163.71 9.12 163.92 9.33 ;
    RECT 164.28 4.845 164.35 4.915 ;
    RECT 164.28 9.43 164.35 9.5 ;
    RECT 165.12 9.765 165.33 9.835 ;
    RECT 165.58 2.585 165.79 2.795 ;
    RECT 165.58 5.86 165.79 6.07 ;
    RECT 165.58 6.385 165.79 6.455 ;
    RECT 165.58 7.28 165.79 7.35 ;
    RECT 160.39 3.235 160.6 3.445 ;
    RECT 160.39 5.33 160.6 5.54 ;
    RECT 160.39 9.12 160.6 9.33 ;
    RECT 160.96 4.845 161.03 4.915 ;
    RECT 160.96 9.43 161.03 9.5 ;
    RECT 161.8 9.765 162.01 9.835 ;
    RECT 162.26 2.585 162.47 2.795 ;
    RECT 162.26 5.86 162.47 6.07 ;
    RECT 162.26 6.385 162.47 6.455 ;
    RECT 162.26 7.28 162.47 7.35 ;
    RECT 17.63 4.455 17.84 4.525 ;
    RECT 157.07 3.235 157.28 3.445 ;
    RECT 157.07 5.33 157.28 5.54 ;
    RECT 157.07 9.12 157.28 9.33 ;
    RECT 157.64 4.845 157.71 4.915 ;
    RECT 157.64 9.43 157.71 9.5 ;
    RECT 158.48 9.765 158.69 9.835 ;
    RECT 158.94 2.585 159.15 2.795 ;
    RECT 158.94 5.86 159.15 6.07 ;
    RECT 158.94 6.385 159.15 6.455 ;
    RECT 158.94 7.28 159.15 7.35 ;
    RECT 153.75 3.235 153.96 3.445 ;
    RECT 153.75 5.33 153.96 5.54 ;
    RECT 153.75 9.12 153.96 9.33 ;
    RECT 154.32 4.845 154.39 4.915 ;
    RECT 154.32 9.43 154.39 9.5 ;
    RECT 155.16 9.765 155.37 9.835 ;
    RECT 155.62 2.585 155.83 2.795 ;
    RECT 155.62 5.86 155.83 6.07 ;
    RECT 155.62 6.385 155.83 6.455 ;
    RECT 155.62 7.28 155.83 7.35 ;
    RECT 40.87 4.455 41.08 4.525 ;
    RECT 150.43 3.235 150.64 3.445 ;
    RECT 150.43 5.33 150.64 5.54 ;
    RECT 150.43 9.12 150.64 9.33 ;
    RECT 151.0 4.845 151.07 4.915 ;
    RECT 151.0 9.43 151.07 9.5 ;
    RECT 151.84 9.765 152.05 9.835 ;
    RECT 152.3 2.585 152.51 2.795 ;
    RECT 152.3 5.86 152.51 6.07 ;
    RECT 152.3 6.385 152.51 6.455 ;
    RECT 152.3 7.28 152.51 7.35 ;
    RECT 147.11 3.235 147.32 3.445 ;
    RECT 147.11 5.33 147.32 5.54 ;
    RECT 147.11 9.12 147.32 9.33 ;
    RECT 147.68 4.845 147.75 4.915 ;
    RECT 147.68 9.43 147.75 9.5 ;
    RECT 148.52 9.765 148.73 9.835 ;
    RECT 148.98 2.585 149.19 2.795 ;
    RECT 148.98 5.86 149.19 6.07 ;
    RECT 148.98 6.385 149.19 6.455 ;
    RECT 148.98 7.28 149.19 7.35 ;
    RECT 143.79 3.235 144.0 3.445 ;
    RECT 143.79 5.33 144.0 5.54 ;
    RECT 143.79 9.12 144.0 9.33 ;
    RECT 144.36 4.845 144.43 4.915 ;
    RECT 144.36 9.43 144.43 9.5 ;
    RECT 145.2 9.765 145.41 9.835 ;
    RECT 145.66 2.585 145.87 2.795 ;
    RECT 145.66 5.86 145.87 6.07 ;
    RECT 145.66 6.385 145.87 6.455 ;
    RECT 145.66 7.28 145.87 7.35 ;
    RECT 140.47 3.235 140.68 3.445 ;
    RECT 140.47 5.33 140.68 5.54 ;
    RECT 140.47 9.12 140.68 9.33 ;
    RECT 141.04 4.845 141.11 4.915 ;
    RECT 141.04 9.43 141.11 9.5 ;
    RECT 141.88 9.765 142.09 9.835 ;
    RECT 142.34 2.585 142.55 2.795 ;
    RECT 142.34 5.86 142.55 6.07 ;
    RECT 142.34 6.385 142.55 6.455 ;
    RECT 142.34 7.28 142.55 7.35 ;
    RECT 137.15 3.235 137.36 3.445 ;
    RECT 137.15 5.33 137.36 5.54 ;
    RECT 137.15 9.12 137.36 9.33 ;
    RECT 137.72 4.845 137.79 4.915 ;
    RECT 137.72 9.43 137.79 9.5 ;
    RECT 138.56 9.765 138.77 9.835 ;
    RECT 139.02 2.585 139.23 2.795 ;
    RECT 139.02 5.86 139.23 6.07 ;
    RECT 139.02 6.385 139.23 6.455 ;
    RECT 139.02 7.28 139.23 7.35 ;
    RECT 133.83 3.235 134.04 3.445 ;
    RECT 133.83 5.33 134.04 5.54 ;
    RECT 133.83 9.12 134.04 9.33 ;
    RECT 134.4 4.845 134.47 4.915 ;
    RECT 134.4 9.43 134.47 9.5 ;
    RECT 135.24 9.765 135.45 9.835 ;
    RECT 135.7 2.585 135.91 2.795 ;
    RECT 135.7 5.86 135.91 6.07 ;
    RECT 135.7 6.385 135.91 6.455 ;
    RECT 135.7 7.28 135.91 7.35 ;
    RECT 141.39 6.385 141.6 6.455 ;
    RECT 141.39 5.86 141.6 6.07 ;
    RECT 141.39 2.585 141.6 2.795 ;
    RECT 8.59 7.28 8.8 7.35 ;
    RECT 171.27 7.28 171.48 7.35 ;
    RECT 171.27 6.385 171.48 6.455 ;
    RECT 171.27 5.86 171.48 6.07 ;
    RECT 171.27 2.585 171.48 2.795 ;
    RECT 130.51 4.455 130.72 4.525 ;
    RECT 130.51 3.235 130.72 3.445 ;
    RECT 130.51 5.33 130.72 5.54 ;
    RECT 130.51 9.12 130.72 9.33 ;
    RECT 131.08 4.845 131.15 4.915 ;
    RECT 131.08 9.43 131.15 9.5 ;
    RECT 131.92 9.765 132.13 9.835 ;
    RECT 132.38 2.585 132.59 2.795 ;
    RECT 132.38 5.86 132.59 6.07 ;
    RECT 132.38 6.385 132.59 6.455 ;
    RECT 132.38 7.28 132.59 7.35 ;
    RECT 127.19 3.235 127.4 3.445 ;
    RECT 127.19 5.33 127.4 5.54 ;
    RECT 127.19 9.12 127.4 9.33 ;
    RECT 127.76 4.845 127.83 4.915 ;
    RECT 127.76 9.43 127.83 9.5 ;
    RECT 128.6 9.765 128.81 9.835 ;
    RECT 129.06 2.585 129.27 2.795 ;
    RECT 129.06 5.86 129.27 6.07 ;
    RECT 129.06 6.385 129.27 6.455 ;
    RECT 129.06 7.28 129.27 7.35 ;
    RECT 123.87 3.235 124.08 3.445 ;
    RECT 123.87 5.33 124.08 5.54 ;
    RECT 123.87 9.12 124.08 9.33 ;
    RECT 124.44 4.845 124.51 4.915 ;
    RECT 124.44 9.43 124.51 9.5 ;
    RECT 125.28 9.765 125.49 9.835 ;
    RECT 125.74 2.585 125.95 2.795 ;
    RECT 125.74 5.86 125.95 6.07 ;
    RECT 125.74 6.385 125.95 6.455 ;
    RECT 125.74 7.28 125.95 7.35 ;
    RECT 164.63 7.28 164.84 7.35 ;
    RECT 120.55 3.235 120.76 3.445 ;
    RECT 120.55 5.33 120.76 5.54 ;
    RECT 120.55 9.12 120.76 9.33 ;
    RECT 121.12 4.845 121.19 4.915 ;
    RECT 121.12 9.43 121.19 9.5 ;
    RECT 121.96 9.765 122.17 9.835 ;
    RECT 122.42 2.585 122.63 2.795 ;
    RECT 122.42 5.86 122.63 6.07 ;
    RECT 122.42 6.385 122.63 6.455 ;
    RECT 122.42 7.28 122.63 7.35 ;
    RECT 164.63 6.385 164.84 6.455 ;
    RECT 117.23 3.235 117.44 3.445 ;
    RECT 117.23 5.33 117.44 5.54 ;
    RECT 117.23 9.12 117.44 9.33 ;
    RECT 117.8 4.845 117.87 4.915 ;
    RECT 117.8 9.43 117.87 9.5 ;
    RECT 118.64 9.765 118.85 9.835 ;
    RECT 119.1 2.585 119.31 2.795 ;
    RECT 119.1 5.86 119.31 6.07 ;
    RECT 119.1 6.385 119.31 6.455 ;
    RECT 119.1 7.28 119.31 7.35 ;
    RECT 164.63 5.86 164.84 6.07 ;
    RECT 113.91 3.235 114.12 3.445 ;
    RECT 113.91 5.33 114.12 5.54 ;
    RECT 113.91 9.12 114.12 9.33 ;
    RECT 114.48 4.845 114.55 4.915 ;
    RECT 114.48 9.43 114.55 9.5 ;
    RECT 115.32 9.765 115.53 9.835 ;
    RECT 115.78 2.585 115.99 2.795 ;
    RECT 115.78 5.86 115.99 6.07 ;
    RECT 115.78 6.385 115.99 6.455 ;
    RECT 115.78 7.28 115.99 7.35 ;
    RECT 164.63 2.585 164.84 2.795 ;
    RECT 8.59 6.385 8.8 6.455 ;
    RECT 110.59 3.235 110.8 3.445 ;
    RECT 110.59 5.33 110.8 5.54 ;
    RECT 110.59 9.12 110.8 9.33 ;
    RECT 111.16 4.845 111.23 4.915 ;
    RECT 111.16 9.43 111.23 9.5 ;
    RECT 112.0 9.765 112.21 9.835 ;
    RECT 112.46 2.585 112.67 2.795 ;
    RECT 112.46 5.86 112.67 6.07 ;
    RECT 112.46 6.385 112.67 6.455 ;
    RECT 112.46 7.28 112.67 7.35 ;
    RECT 38.47 7.28 38.68 7.35 ;
    RECT 68.35 7.28 68.56 7.35 ;
    RECT 8.59 5.86 8.8 6.07 ;
    RECT 107.27 3.235 107.48 3.445 ;
    RECT 107.27 5.33 107.48 5.54 ;
    RECT 107.27 9.12 107.48 9.33 ;
    RECT 107.84 4.845 107.91 4.915 ;
    RECT 107.84 9.43 107.91 9.5 ;
    RECT 108.68 9.765 108.89 9.835 ;
    RECT 109.14 2.585 109.35 2.795 ;
    RECT 109.14 5.86 109.35 6.07 ;
    RECT 109.14 6.385 109.35 6.455 ;
    RECT 109.14 7.28 109.35 7.35 ;
    RECT 38.47 6.385 38.68 6.455 ;
    RECT 68.35 6.385 68.56 6.455 ;
    RECT 8.59 2.585 8.8 2.795 ;
    RECT 103.95 3.235 104.16 3.445 ;
    RECT 103.95 5.33 104.16 5.54 ;
    RECT 103.95 9.12 104.16 9.33 ;
    RECT 104.52 4.845 104.59 4.915 ;
    RECT 104.52 9.43 104.59 9.5 ;
    RECT 105.36 9.765 105.57 9.835 ;
    RECT 105.82 2.585 106.03 2.795 ;
    RECT 105.82 5.86 106.03 6.07 ;
    RECT 105.82 6.385 106.03 6.455 ;
    RECT 105.82 7.28 106.03 7.35 ;
    RECT 38.47 5.86 38.68 6.07 ;
    RECT 68.35 5.86 68.56 6.07 ;
    RECT 100.63 3.235 100.84 3.445 ;
    RECT 100.63 5.33 100.84 5.54 ;
    RECT 100.63 9.12 100.84 9.33 ;
    RECT 101.2 4.845 101.27 4.915 ;
    RECT 101.2 9.43 101.27 9.5 ;
    RECT 102.04 9.765 102.25 9.835 ;
    RECT 102.5 2.585 102.71 2.795 ;
    RECT 102.5 5.86 102.71 6.07 ;
    RECT 102.5 6.385 102.71 6.455 ;
    RECT 102.5 7.28 102.71 7.35 ;
    RECT 38.47 2.585 38.68 2.795 ;
    RECT 28.51 4.055 28.72 4.125 ;
    RECT 70.75 4.455 70.96 4.525 ;
    RECT 108.19 4.055 108.4 4.125 ;
    RECT 61.71 7.28 61.92 7.35 ;
    RECT 61.71 6.385 61.92 6.455 ;
    RECT 61.71 5.86 61.92 6.07 ;
    RECT 61.71 2.585 61.92 2.795 ;
    RECT 64.11 4.455 64.32 4.525 ;
    RECT 164.63 4.055 164.84 4.125 ;
    RECT 4.35 4.455 4.56 4.525 ;
    RECT 31.83 7.28 32.04 7.35 ;
    RECT 127.19 4.455 127.4 4.525 ;
    RECT 68.35 2.585 68.56 2.795 ;
    RECT 88.27 4.055 88.48 4.125 ;
    RECT 31.83 6.385 32.04 6.455 ;
    RECT 97.31 3.235 97.52 3.445 ;
    RECT 97.31 5.33 97.52 5.54 ;
    RECT 97.31 9.12 97.52 9.33 ;
    RECT 97.88 4.845 97.95 4.915 ;
    RECT 97.88 9.43 97.95 9.5 ;
    RECT 98.72 9.765 98.93 9.835 ;
    RECT 99.18 2.585 99.39 2.795 ;
    RECT 99.18 5.86 99.39 6.07 ;
    RECT 99.18 6.385 99.39 6.455 ;
    RECT 99.18 7.28 99.39 7.35 ;
    RECT 91.59 7.28 91.8 7.35 ;
    RECT 31.83 5.86 32.04 6.07 ;
    RECT 93.99 3.235 94.2 3.445 ;
    RECT 93.99 5.33 94.2 5.54 ;
    RECT 93.99 9.12 94.2 9.33 ;
    RECT 94.56 4.845 94.63 4.915 ;
    RECT 94.56 9.43 94.63 9.5 ;
    RECT 95.4 9.765 95.61 9.835 ;
    RECT 95.86 2.585 96.07 2.795 ;
    RECT 95.86 5.86 96.07 6.07 ;
    RECT 95.86 6.385 96.07 6.455 ;
    RECT 95.86 7.28 96.07 7.35 ;
    RECT 31.83 2.585 32.04 2.795 ;
    RECT 90.67 3.235 90.88 3.445 ;
    RECT 90.67 5.33 90.88 5.54 ;
    RECT 90.67 9.12 90.88 9.33 ;
    RECT 91.24 4.845 91.31 4.915 ;
    RECT 91.24 9.43 91.31 9.5 ;
    RECT 92.08 9.765 92.29 9.835 ;
    RECT 92.54 2.585 92.75 2.795 ;
    RECT 92.54 5.86 92.75 6.07 ;
    RECT 92.54 6.385 92.75 6.455 ;
    RECT 92.54 7.28 92.75 7.35 ;
    RECT 87.35 3.235 87.56 3.445 ;
    RECT 87.35 5.33 87.56 5.54 ;
    RECT 87.35 9.12 87.56 9.33 ;
    RECT 87.92 4.845 87.99 4.915 ;
    RECT 87.92 9.43 87.99 9.5 ;
    RECT 88.76 9.765 88.97 9.835 ;
    RECT 89.22 2.585 89.43 2.795 ;
    RECT 89.22 5.86 89.43 6.07 ;
    RECT 89.22 6.385 89.43 6.455 ;
    RECT 89.22 7.28 89.43 7.35 ;
    RECT 84.03 3.235 84.24 3.445 ;
    RECT 84.03 5.33 84.24 5.54 ;
    RECT 84.03 9.12 84.24 9.33 ;
    RECT 84.6 4.845 84.67 4.915 ;
    RECT 84.6 9.43 84.67 9.5 ;
    RECT 85.44 9.765 85.65 9.835 ;
    RECT 85.9 2.585 86.11 2.795 ;
    RECT 85.9 5.86 86.11 6.07 ;
    RECT 85.9 6.385 86.11 6.455 ;
    RECT 85.9 7.28 86.11 7.35 ;
    RECT 80.71 3.235 80.92 3.445 ;
    RECT 80.71 5.33 80.92 5.54 ;
    RECT 80.71 9.12 80.92 9.33 ;
    RECT 81.28 4.845 81.35 4.915 ;
    RECT 81.28 9.43 81.35 9.5 ;
    RECT 82.12 9.765 82.33 9.835 ;
    RECT 82.58 2.585 82.79 2.795 ;
    RECT 82.58 5.86 82.79 6.07 ;
    RECT 82.58 6.385 82.79 6.455 ;
    RECT 82.58 7.28 82.79 7.35 ;
    RECT 77.39 3.235 77.6 3.445 ;
    RECT 77.39 5.33 77.6 5.54 ;
    RECT 77.39 9.12 77.6 9.33 ;
    RECT 77.96 4.845 78.03 4.915 ;
    RECT 77.96 9.43 78.03 9.5 ;
    RECT 78.8 9.765 79.01 9.835 ;
    RECT 79.26 2.585 79.47 2.795 ;
    RECT 79.26 5.86 79.47 6.07 ;
    RECT 79.26 6.385 79.47 6.455 ;
    RECT 79.26 7.28 79.47 7.35 ;
    RECT 74.07 3.235 74.28 3.445 ;
    RECT 74.07 5.33 74.28 5.54 ;
    RECT 74.07 9.12 74.28 9.33 ;
    RECT 74.64 4.845 74.71 4.915 ;
    RECT 74.64 9.43 74.71 9.5 ;
    RECT 75.48 9.765 75.69 9.835 ;
    RECT 75.94 2.585 76.15 2.795 ;
    RECT 75.94 5.86 76.15 6.07 ;
    RECT 75.94 6.385 76.15 6.455 ;
    RECT 75.94 7.28 76.15 7.35 ;
    RECT 70.75 3.235 70.96 3.445 ;
    RECT 70.75 5.33 70.96 5.54 ;
    RECT 70.75 9.12 70.96 9.33 ;
    RECT 71.32 4.845 71.39 4.915 ;
    RECT 71.32 9.43 71.39 9.5 ;
    RECT 72.16 9.765 72.37 9.835 ;
    RECT 72.62 2.585 72.83 2.795 ;
    RECT 72.62 5.86 72.83 6.07 ;
    RECT 72.62 6.385 72.83 6.455 ;
    RECT 72.62 7.28 72.83 7.35 ;
    RECT 67.43 3.235 67.64 3.445 ;
    RECT 67.43 5.33 67.64 5.54 ;
    RECT 67.43 9.12 67.64 9.33 ;
    RECT 68.0 4.845 68.07 4.915 ;
    RECT 68.0 9.43 68.07 9.5 ;
    RECT 68.84 9.765 69.05 9.835 ;
    RECT 69.3 2.585 69.51 2.795 ;
    RECT 69.3 5.86 69.51 6.07 ;
    RECT 69.3 6.385 69.51 6.455 ;
    RECT 69.3 7.28 69.51 7.35 ;
    RECT 171.27 4.055 171.48 4.125 ;
    RECT 266.685 61.05 266.895 61.12 ;
    RECT 266.21 61.05 266.42 61.12 ;
    RECT 265.725 60.77 265.935 60.84 ;
    RECT 263.365 61.05 263.575 61.12 ;
    RECT 262.89 61.05 263.1 61.12 ;
    RECT 262.405 60.77 262.615 60.84 ;
    RECT 260.045 61.05 260.255 61.12 ;
    RECT 259.57 61.05 259.78 61.12 ;
    RECT 259.085 60.77 259.295 60.84 ;
    RECT 256.725 61.05 256.935 61.12 ;
    RECT 256.25 61.05 256.46 61.12 ;
    RECT 255.765 60.77 255.975 60.84 ;
    RECT 253.405 61.05 253.615 61.12 ;
    RECT 252.93 61.05 253.14 61.12 ;
    RECT 252.445 60.77 252.655 60.84 ;
    RECT 250.085 61.05 250.295 61.12 ;
    RECT 249.61 61.05 249.82 61.12 ;
    RECT 249.125 60.77 249.335 60.84 ;
    RECT 246.765 61.05 246.975 61.12 ;
    RECT 246.29 61.05 246.5 61.12 ;
    RECT 245.805 60.77 246.015 60.84 ;
    RECT 243.445 61.05 243.655 61.12 ;
    RECT 242.97 61.05 243.18 61.12 ;
    RECT 242.485 60.77 242.695 60.84 ;
    RECT 240.125 61.05 240.335 61.12 ;
    RECT 239.65 61.05 239.86 61.12 ;
    RECT 239.165 60.77 239.375 60.84 ;
    RECT 236.805 61.05 237.015 61.12 ;
    RECT 236.33 61.05 236.54 61.12 ;
    RECT 235.845 60.77 236.055 60.84 ;
    RECT 170.805 61.05 171.015 61.12 ;
    RECT 171.28 61.05 171.49 61.12 ;
    RECT 171.765 60.77 171.975 60.84 ;
    RECT 167.485 61.05 167.695 61.12 ;
    RECT 167.96 61.05 168.17 61.12 ;
    RECT 168.445 60.77 168.655 60.84 ;
    RECT 164.165 61.05 164.375 61.12 ;
    RECT 164.64 61.05 164.85 61.12 ;
    RECT 165.125 60.77 165.335 60.84 ;
    RECT 160.845 61.05 161.055 61.12 ;
    RECT 161.32 61.05 161.53 61.12 ;
    RECT 161.805 60.77 162.015 60.84 ;
    RECT 157.525 61.05 157.735 61.12 ;
    RECT 158.0 61.05 158.21 61.12 ;
    RECT 158.485 60.77 158.695 60.84 ;
    RECT 154.205 61.05 154.415 61.12 ;
    RECT 154.68 61.05 154.89 61.12 ;
    RECT 155.165 60.77 155.375 60.84 ;
    RECT 150.885 61.05 151.095 61.12 ;
    RECT 151.36 61.05 151.57 61.12 ;
    RECT 151.845 60.77 152.055 60.84 ;
    RECT 147.565 61.05 147.775 61.12 ;
    RECT 148.04 61.05 148.25 61.12 ;
    RECT 148.525 60.77 148.735 60.84 ;
    RECT 144.245 61.05 144.455 61.12 ;
    RECT 144.72 61.05 144.93 61.12 ;
    RECT 145.205 60.77 145.415 60.84 ;
    RECT 140.925 61.05 141.135 61.12 ;
    RECT 141.4 61.05 141.61 61.12 ;
    RECT 141.885 60.77 142.095 60.84 ;
    RECT 137.605 61.05 137.815 61.12 ;
    RECT 138.08 61.05 138.29 61.12 ;
    RECT 138.565 60.77 138.775 60.84 ;
    RECT 134.285 61.05 134.495 61.12 ;
    RECT 134.76 61.05 134.97 61.12 ;
    RECT 135.245 60.77 135.455 60.84 ;
    RECT 176.885 60.79 177.095 60.86 ;
    RECT 176.355 60.79 176.565 60.86 ;
    RECT 130.965 61.05 131.175 61.12 ;
    RECT 131.44 61.05 131.65 61.12 ;
    RECT 131.925 60.77 132.135 60.84 ;
    RECT 127.645 61.05 127.855 61.12 ;
    RECT 128.12 61.05 128.33 61.12 ;
    RECT 128.605 60.77 128.815 60.84 ;
    RECT 124.325 61.05 124.535 61.12 ;
    RECT 124.8 61.05 125.01 61.12 ;
    RECT 125.285 60.77 125.495 60.84 ;
    RECT 121.005 61.05 121.215 61.12 ;
    RECT 121.48 61.05 121.69 61.12 ;
    RECT 121.965 60.77 122.175 60.84 ;
    RECT 117.685 61.05 117.895 61.12 ;
    RECT 118.16 61.05 118.37 61.12 ;
    RECT 118.645 60.77 118.855 60.84 ;
    RECT 114.365 61.05 114.575 61.12 ;
    RECT 114.84 61.05 115.05 61.12 ;
    RECT 115.325 60.77 115.535 60.84 ;
    RECT 111.045 61.05 111.255 61.12 ;
    RECT 111.52 61.05 111.73 61.12 ;
    RECT 112.005 60.77 112.215 60.84 ;
    RECT 107.725 61.05 107.935 61.12 ;
    RECT 108.2 61.05 108.41 61.12 ;
    RECT 108.685 60.77 108.895 60.84 ;
    RECT 233.485 61.05 233.695 61.12 ;
    RECT 233.01 61.05 233.22 61.12 ;
    RECT 232.525 60.77 232.735 60.84 ;
    RECT 104.405 61.05 104.615 61.12 ;
    RECT 104.88 61.05 105.09 61.12 ;
    RECT 105.365 60.77 105.575 60.84 ;
    RECT 230.165 61.05 230.375 61.12 ;
    RECT 229.69 61.05 229.9 61.12 ;
    RECT 229.205 60.77 229.415 60.84 ;
    RECT 101.085 61.05 101.295 61.12 ;
    RECT 101.56 61.05 101.77 61.12 ;
    RECT 102.045 60.77 102.255 60.84 ;
    RECT 226.845 61.05 227.055 61.12 ;
    RECT 226.37 61.05 226.58 61.12 ;
    RECT 225.885 60.77 226.095 60.84 ;
    RECT 223.525 61.05 223.735 61.12 ;
    RECT 223.05 61.05 223.26 61.12 ;
    RECT 222.565 60.77 222.775 60.84 ;
    RECT 220.205 61.05 220.415 61.12 ;
    RECT 219.73 61.05 219.94 61.12 ;
    RECT 219.245 60.77 219.455 60.84 ;
    RECT 216.885 61.05 217.095 61.12 ;
    RECT 216.41 61.05 216.62 61.12 ;
    RECT 215.925 60.77 216.135 60.84 ;
    RECT 213.565 61.05 213.775 61.12 ;
    RECT 213.09 61.05 213.3 61.12 ;
    RECT 212.605 60.77 212.815 60.84 ;
    RECT 210.245 61.05 210.455 61.12 ;
    RECT 209.77 61.05 209.98 61.12 ;
    RECT 209.285 60.77 209.495 60.84 ;
    RECT 206.925 61.05 207.135 61.12 ;
    RECT 206.45 61.05 206.66 61.12 ;
    RECT 205.965 60.77 206.175 60.84 ;
    RECT 203.605 61.05 203.815 61.12 ;
    RECT 203.13 61.05 203.34 61.12 ;
    RECT 202.645 60.77 202.855 60.84 ;
    RECT 97.765 61.05 97.975 61.12 ;
    RECT 98.24 61.05 98.45 61.12 ;
    RECT 98.725 60.77 98.935 60.84 ;
    RECT 198.605 61.062 198.815 61.132 ;
    RECT 94.445 61.05 94.655 61.12 ;
    RECT 94.92 61.05 95.13 61.12 ;
    RECT 95.405 60.77 95.615 60.84 ;
    RECT 91.125 61.05 91.335 61.12 ;
    RECT 91.6 61.05 91.81 61.12 ;
    RECT 92.085 60.77 92.295 60.84 ;
    RECT 193.595 61.062 193.805 61.132 ;
    RECT 87.805 61.05 88.015 61.12 ;
    RECT 88.28 61.05 88.49 61.12 ;
    RECT 88.765 60.77 88.975 60.84 ;
    RECT 84.485 61.05 84.695 61.12 ;
    RECT 84.96 61.05 85.17 61.12 ;
    RECT 85.445 60.77 85.655 60.84 ;
    RECT 81.165 61.05 81.375 61.12 ;
    RECT 81.64 61.05 81.85 61.12 ;
    RECT 82.125 60.77 82.335 60.84 ;
    RECT 77.845 61.05 78.055 61.12 ;
    RECT 78.32 61.05 78.53 61.12 ;
    RECT 78.805 60.77 79.015 60.84 ;
    RECT 0.4 61.07 0.47 61.14 ;
    RECT 184.12 61.062 184.33 61.132 ;
    RECT 74.525 61.05 74.735 61.12 ;
    RECT 75.0 61.05 75.21 61.12 ;
    RECT 75.485 60.77 75.695 60.84 ;
    RECT 71.205 61.05 71.415 61.12 ;
    RECT 71.68 61.05 71.89 61.12 ;
    RECT 72.165 60.77 72.375 60.84 ;
    RECT 183.085 61.062 183.295 61.132 ;
    RECT 67.885 61.05 68.095 61.12 ;
    RECT 68.36 61.05 68.57 61.12 ;
    RECT 68.845 60.77 69.055 60.84 ;
    RECT 0.19 60.79 0.26 60.86 ;
    RECT 64.565 61.05 64.775 61.12 ;
    RECT 65.04 61.05 65.25 61.12 ;
    RECT 65.525 60.77 65.735 60.84 ;
    RECT 198.045 60.79 198.255 60.86 ;
    RECT 61.245 61.05 61.455 61.12 ;
    RECT 61.72 61.05 61.93 61.12 ;
    RECT 62.205 60.77 62.415 60.84 ;
    RECT 197.465 60.79 197.675 60.86 ;
    RECT 57.925 61.05 58.135 61.12 ;
    RECT 58.4 61.05 58.61 61.12 ;
    RECT 58.885 60.77 59.095 60.84 ;
    RECT 54.605 61.05 54.815 61.12 ;
    RECT 55.08 61.05 55.29 61.12 ;
    RECT 55.565 60.77 55.775 60.84 ;
    RECT 51.285 61.05 51.495 61.12 ;
    RECT 51.76 61.05 51.97 61.12 ;
    RECT 52.245 60.77 52.455 60.84 ;
    RECT 47.965 61.05 48.175 61.12 ;
    RECT 48.44 61.05 48.65 61.12 ;
    RECT 48.925 60.77 49.135 60.84 ;
    RECT 44.645 61.05 44.855 61.12 ;
    RECT 45.12 61.05 45.33 61.12 ;
    RECT 45.605 60.77 45.815 60.84 ;
    RECT 41.325 61.05 41.535 61.12 ;
    RECT 41.8 61.05 42.01 61.12 ;
    RECT 42.285 60.77 42.495 60.84 ;
    RECT 38.005 61.05 38.215 61.12 ;
    RECT 38.48 61.05 38.69 61.12 ;
    RECT 38.965 60.77 39.175 60.84 ;
    RECT 34.685 61.05 34.895 61.12 ;
    RECT 35.16 61.05 35.37 61.12 ;
    RECT 35.645 60.77 35.855 60.84 ;
    RECT 175.75 61.062 175.96 61.132 ;
    RECT 372.925 61.05 373.135 61.12 ;
    RECT 372.45 61.05 372.66 61.12 ;
    RECT 371.965 60.77 372.175 60.84 ;
    RECT 369.605 61.05 369.815 61.12 ;
    RECT 369.13 61.05 369.34 61.12 ;
    RECT 368.645 60.77 368.855 60.84 ;
    RECT 366.285 61.05 366.495 61.12 ;
    RECT 365.81 61.05 366.02 61.12 ;
    RECT 365.325 60.77 365.535 60.84 ;
    RECT 362.965 61.05 363.175 61.12 ;
    RECT 362.49 61.05 362.7 61.12 ;
    RECT 362.005 60.77 362.215 60.84 ;
    RECT 359.645 61.05 359.855 61.12 ;
    RECT 359.17 61.05 359.38 61.12 ;
    RECT 358.685 60.77 358.895 60.84 ;
    RECT 31.365 61.05 31.575 61.12 ;
    RECT 31.84 61.05 32.05 61.12 ;
    RECT 32.325 60.77 32.535 60.84 ;
    RECT 356.325 61.05 356.535 61.12 ;
    RECT 355.85 61.05 356.06 61.12 ;
    RECT 355.365 60.77 355.575 60.84 ;
    RECT 28.045 61.05 28.255 61.12 ;
    RECT 28.52 61.05 28.73 61.12 ;
    RECT 29.005 60.77 29.215 60.84 ;
    RECT 353.005 61.05 353.215 61.12 ;
    RECT 352.53 61.05 352.74 61.12 ;
    RECT 352.045 60.77 352.255 60.84 ;
    RECT 24.725 61.05 24.935 61.12 ;
    RECT 25.2 61.05 25.41 61.12 ;
    RECT 25.685 60.77 25.895 60.84 ;
    RECT 349.685 61.05 349.895 61.12 ;
    RECT 349.21 61.05 349.42 61.12 ;
    RECT 348.725 60.77 348.935 60.84 ;
    RECT 21.405 61.05 21.615 61.12 ;
    RECT 21.88 61.05 22.09 61.12 ;
    RECT 22.365 60.77 22.575 60.84 ;
    RECT 346.365 61.05 346.575 61.12 ;
    RECT 345.89 61.05 346.1 61.12 ;
    RECT 345.405 60.77 345.615 60.84 ;
    RECT 18.085 61.05 18.295 61.12 ;
    RECT 18.56 61.05 18.77 61.12 ;
    RECT 19.045 60.77 19.255 60.84 ;
    RECT 343.045 61.05 343.255 61.12 ;
    RECT 342.57 61.05 342.78 61.12 ;
    RECT 342.085 60.77 342.295 60.84 ;
    RECT 14.765 61.05 14.975 61.12 ;
    RECT 15.24 61.05 15.45 61.12 ;
    RECT 15.725 60.77 15.935 60.84 ;
    RECT 339.725 61.05 339.935 61.12 ;
    RECT 339.25 61.05 339.46 61.12 ;
    RECT 338.765 60.77 338.975 60.84 ;
    RECT 11.445 61.05 11.655 61.12 ;
    RECT 11.92 61.05 12.13 61.12 ;
    RECT 12.405 60.77 12.615 60.84 ;
    RECT 336.405 61.05 336.615 61.12 ;
    RECT 335.93 61.05 336.14 61.12 ;
    RECT 335.445 60.77 335.655 60.84 ;
    RECT 8.125 61.05 8.335 61.12 ;
    RECT 8.6 61.05 8.81 61.12 ;
    RECT 9.085 60.77 9.295 60.84 ;
    RECT 4.805 61.05 5.015 61.12 ;
    RECT 5.28 61.05 5.49 61.12 ;
    RECT 5.765 60.77 5.975 60.84 ;
    RECT 1.485 61.05 1.695 61.12 ;
    RECT 1.96 61.05 2.17 61.12 ;
    RECT 2.445 60.77 2.655 60.84 ;
    RECT 174.56 61.07 174.63 61.14 ;
    RECT 174.85 60.79 174.92 60.86 ;
    RECT 175.16 61.07 175.37 61.14 ;
    RECT 177.375 61.07 177.585 61.14 ;
    RECT 178.23 61.07 178.44 61.14 ;
    RECT 178.79 60.79 179.0 60.86 ;
    RECT 179.88 61.07 180.09 61.14 ;
    RECT 184.92 61.07 184.99 61.14 ;
    RECT 187.46 61.07 187.67 61.14 ;
    RECT 190.04 61.07 190.25 61.14 ;
    RECT 192.85 61.065 193.06 61.135 ;
    RECT 194.535 61.07 194.745 61.14 ;
    RECT 195.63 60.79 195.84 60.86 ;
    RECT 196.19 61.07 196.26 61.14 ;
    RECT 196.81 61.07 197.02 61.14 ;
    RECT 199.28 61.07 199.49 61.14 ;
    RECT 374.15 61.07 374.22 61.14 ;
    RECT 374.36 60.79 374.43 60.86 ;
    RECT 333.085 61.05 333.295 61.12 ;
    RECT 332.61 61.05 332.82 61.12 ;
    RECT 332.125 60.77 332.335 60.84 ;
    RECT 329.765 61.05 329.975 61.12 ;
    RECT 329.29 61.05 329.5 61.12 ;
    RECT 328.805 60.77 329.015 60.84 ;
    RECT 326.445 61.05 326.655 61.12 ;
    RECT 325.97 61.05 326.18 61.12 ;
    RECT 325.485 60.77 325.695 60.84 ;
    RECT 323.125 61.05 323.335 61.12 ;
    RECT 322.65 61.05 322.86 61.12 ;
    RECT 322.165 60.77 322.375 60.84 ;
    RECT 319.805 61.05 320.015 61.12 ;
    RECT 319.33 61.05 319.54 61.12 ;
    RECT 318.845 60.77 319.055 60.84 ;
    RECT 316.485 61.05 316.695 61.12 ;
    RECT 316.01 61.05 316.22 61.12 ;
    RECT 315.525 60.77 315.735 60.84 ;
    RECT 313.165 61.05 313.375 61.12 ;
    RECT 312.69 61.05 312.9 61.12 ;
    RECT 312.205 60.77 312.415 60.84 ;
    RECT 309.845 61.05 310.055 61.12 ;
    RECT 309.37 61.05 309.58 61.12 ;
    RECT 308.885 60.77 309.095 60.84 ;
    RECT 306.525 61.05 306.735 61.12 ;
    RECT 306.05 61.05 306.26 61.12 ;
    RECT 305.565 60.77 305.775 60.84 ;
    RECT 303.205 61.05 303.415 61.12 ;
    RECT 302.73 61.05 302.94 61.12 ;
    RECT 302.245 60.77 302.455 60.84 ;
    RECT 299.885 61.05 300.095 61.12 ;
    RECT 299.41 61.05 299.62 61.12 ;
    RECT 298.925 60.77 299.135 60.84 ;
    RECT 296.565 61.05 296.775 61.12 ;
    RECT 296.09 61.05 296.3 61.12 ;
    RECT 295.605 60.77 295.815 60.84 ;
    RECT 293.245 61.05 293.455 61.12 ;
    RECT 292.77 61.05 292.98 61.12 ;
    RECT 292.285 60.77 292.495 60.84 ;
    RECT 289.925 61.05 290.135 61.12 ;
    RECT 289.45 61.05 289.66 61.12 ;
    RECT 288.965 60.77 289.175 60.84 ;
    RECT 286.605 61.05 286.815 61.12 ;
    RECT 286.13 61.05 286.34 61.12 ;
    RECT 285.645 60.77 285.855 60.84 ;
    RECT 283.285 61.05 283.495 61.12 ;
    RECT 282.81 61.05 283.02 61.12 ;
    RECT 282.325 60.77 282.535 60.84 ;
    RECT 279.965 61.05 280.175 61.12 ;
    RECT 279.49 61.05 279.7 61.12 ;
    RECT 279.005 60.77 279.215 60.84 ;
    RECT 276.645 61.05 276.855 61.12 ;
    RECT 276.17 61.05 276.38 61.12 ;
    RECT 275.685 60.77 275.895 60.84 ;
    RECT 273.325 61.05 273.535 61.12 ;
    RECT 272.85 61.05 273.06 61.12 ;
    RECT 272.365 60.77 272.575 60.84 ;
    RECT 270.005 61.05 270.215 61.12 ;
    RECT 269.53 61.05 269.74 61.12 ;
    RECT 269.045 60.77 269.255 60.84 ;
    LAYER M4 DESIGNRULEWIDTH 0.165 ;
    RECT 59.305 0.37 59.585 0.695 ;
    RECT 55.985 0.37 56.265 0.695 ;
    RECT 52.665 0.37 52.945 0.695 ;
    RECT 49.345 0.37 49.625 0.695 ;
    RECT 331.635 0.37 331.915 0.695 ;
    RECT 46.025 0.37 46.305 0.695 ;
    RECT 328.315 0.37 328.595 0.695 ;
    RECT 42.705 0.37 42.985 0.695 ;
    RECT 324.995 0.37 325.275 0.695 ;
    RECT 39.385 0.37 39.665 0.695 ;
    RECT 321.675 0.37 321.955 0.695 ;
    RECT 36.065 0.37 36.345 0.695 ;
    RECT 318.355 0.37 318.635 0.695 ;
    RECT 315.035 0.37 315.315 0.695 ;
    RECT 311.715 0.37 311.995 0.695 ;
    RECT 308.395 0.37 308.675 0.695 ;
    RECT 305.075 0.37 305.355 0.695 ;
    RECT 173.565 0.0 173.645 0.695 ;
    RECT 174.315 0.0 174.45 0.695 ;
    RECT 174.74 0.0 175.09 0.695 ;
    RECT 175.675 0.0 177.24 0.695 ;
    RECT 178.51 0.0 178.665 0.695 ;
    RECT 179.125 0.32 179.75 0.695 ;
    RECT 179.125 0.0 179.36 0.32 ;
    RECT 180.22 0.0 180.37 0.695 ;
    RECT 180.72 0.0 181.115 0.695 ;
    RECT 181.405 0.0 181.725 0.695 ;
    RECT 182.155 0.0 182.435 0.695 ;
    RECT 182.905 0.0 183.605 0.695 ;
    RECT 183.895 0.0 184.405 0.695 ;
    RECT 185.075 0.0 186.625 0.695 ;
    RECT 186.975 0.0 187.325 0.695 ;
    RECT 187.805 0.0 189.52 0.695 ;
    RECT 190.32 0.0 190.64 0.695 ;
    RECT 190.92 0.0 191.38 0.695 ;
    RECT 192.18 0.0 193.905 0.695 ;
    RECT 194.195 0.0 194.4 0.695 ;
    RECT 195.4 0.0 195.56 0.695 ;
    RECT 195.91 0.0 196.08 0.695 ;
    RECT 197.15 0.0 198.885 0.695 ;
    RECT 199.625 0.0 199.815 0.695 ;
    RECT 200.165 0.0 200.305 0.695 ;
    RECT 200.975 0.0 201.055 0.695 ;
    RECT 301.755 0.37 302.035 0.695 ;
    RECT 232.035 0.37 232.315 0.695 ;
    RECT 228.715 0.37 228.995 0.695 ;
    RECT 298.435 0.37 298.715 0.695 ;
    RECT 225.395 0.37 225.675 0.695 ;
    RECT 295.115 0.37 295.395 0.695 ;
    RECT 222.075 0.37 222.355 0.695 ;
    RECT 291.795 0.37 292.075 0.695 ;
    RECT 218.755 0.37 219.035 0.695 ;
    RECT 288.475 0.37 288.755 0.695 ;
    RECT 215.435 0.37 215.715 0.695 ;
    RECT 285.155 0.37 285.435 0.695 ;
    RECT 212.115 0.37 212.395 0.695 ;
    RECT 281.835 0.37 282.115 0.695 ;
    RECT 208.795 0.37 209.075 0.695 ;
    RECT 278.515 0.37 278.795 0.695 ;
    RECT 172.185 0.37 172.465 0.695 ;
    RECT 205.475 0.37 205.755 0.695 ;
    RECT 275.195 0.37 275.475 0.695 ;
    RECT 168.865 0.37 169.145 0.695 ;
    RECT 202.155 0.37 202.435 0.695 ;
    RECT 271.875 0.37 272.155 0.695 ;
    RECT 268.555 0.37 268.835 0.695 ;
    RECT 165.545 0.37 165.825 0.695 ;
    RECT 162.225 0.37 162.505 0.695 ;
    RECT 265.235 0.37 265.515 0.695 ;
    RECT 158.905 0.37 159.185 0.695 ;
    RECT 261.915 0.37 262.195 0.695 ;
    RECT 155.585 0.37 155.865 0.695 ;
    RECT 258.595 0.37 258.875 0.695 ;
    RECT 152.265 0.37 152.545 0.695 ;
    RECT 255.275 0.37 255.555 0.695 ;
    RECT 148.945 0.37 149.225 0.695 ;
    RECT 251.955 0.37 252.235 0.695 ;
    RECT 145.625 0.37 145.905 0.695 ;
    RECT 248.635 0.37 248.915 0.695 ;
    RECT 142.305 0.37 142.585 0.695 ;
    RECT 245.315 0.37 245.595 0.695 ;
    RECT 138.985 0.37 139.265 0.695 ;
    RECT 241.995 0.37 242.275 0.695 ;
    RECT 135.665 0.37 135.945 0.695 ;
    RECT 238.675 0.37 238.955 0.695 ;
    RECT 32.745 0.37 33.025 0.695 ;
    RECT 235.355 0.37 235.635 0.695 ;
    RECT 29.425 0.37 29.705 0.695 ;
    RECT 26.105 0.37 26.385 0.695 ;
    RECT 22.785 0.37 23.065 0.695 ;
    RECT 19.465 0.37 19.745 0.695 ;
    RECT 16.145 0.37 16.425 0.695 ;
    RECT 12.825 0.37 13.105 0.695 ;
    RECT 9.505 0.37 9.785 0.695 ;
    RECT 6.185 0.37 6.465 0.695 ;
    RECT 2.865 0.37 3.145 0.695 ;
    RECT 132.345 0.37 132.625 0.695 ;
    RECT 129.025 0.37 129.305 0.695 ;
    RECT 125.705 0.37 125.985 0.695 ;
    RECT 122.385 0.37 122.665 0.695 ;
    RECT 119.065 0.37 119.345 0.695 ;
    RECT 115.745 0.37 116.025 0.695 ;
    RECT 112.425 0.37 112.705 0.695 ;
    RECT 109.105 0.37 109.385 0.695 ;
    RECT 105.785 0.37 106.065 0.695 ;
    RECT 102.465 0.37 102.745 0.695 ;
    RECT 371.475 0.37 371.755 0.695 ;
    RECT 368.155 0.37 368.435 0.695 ;
    RECT 99.145 0.37 99.425 0.695 ;
    RECT 95.825 0.37 96.105 0.695 ;
    RECT 92.505 0.37 92.785 0.695 ;
    RECT 89.185 0.37 89.465 0.695 ;
    RECT 85.865 0.37 86.145 0.695 ;
    RECT 364.835 0.37 365.115 0.695 ;
    RECT 82.545 0.37 82.825 0.695 ;
    RECT 361.515 0.37 361.795 0.695 ;
    RECT 79.225 0.37 79.505 0.695 ;
    RECT 358.195 0.37 358.475 0.695 ;
    RECT 75.905 0.37 76.185 0.695 ;
    RECT 354.875 0.37 355.155 0.695 ;
    RECT 72.585 0.37 72.865 0.695 ;
    RECT 351.555 0.37 351.835 0.695 ;
    RECT 69.265 0.37 69.545 0.695 ;
    RECT 348.235 0.37 348.515 0.695 ;
    RECT 344.915 0.37 345.195 0.695 ;
    RECT 341.595 0.37 341.875 0.695 ;
    RECT 338.275 0.37 338.555 0.695 ;
    RECT 334.955 0.37 335.235 0.695 ;
    RECT 65.945 0.37 66.225 0.695 ;
    RECT 62.625 0.37 62.905 0.695 ;
    RECT 174.33 56.96 174.45 57.68 ;
    RECT 174.74 56.96 175.09 57.68 ;
    RECT 175.675 56.96 177.24 57.68 ;
    RECT 178.51 56.96 178.665 57.68 ;
    RECT 179.125 56.96 179.75 57.68 ;
    RECT 180.22 56.96 180.37 57.68 ;
    RECT 180.72 56.96 181.115 57.68 ;
    RECT 181.405 56.96 181.725 57.68 ;
    RECT 182.155 56.96 182.435 57.68 ;
    RECT 182.905 56.96 183.605 57.68 ;
    RECT 183.895 56.96 184.405 57.68 ;
    RECT 185.075 56.96 186.625 57.68 ;
    RECT 186.975 56.96 187.325 57.68 ;
    RECT 187.98 56.96 189.52 57.68 ;
    RECT 190.32 56.96 190.64 57.68 ;
    RECT 190.92 56.96 191.38 57.68 ;
    RECT 192.18 56.96 192.72 57.68 ;
    RECT 193.19 56.96 193.905 57.68 ;
    RECT 194.195 56.96 194.4 57.68 ;
    RECT 195.4 56.96 195.56 57.68 ;
    RECT 195.91 56.96 196.08 57.68 ;
    RECT 197.15 56.96 198.885 57.68 ;
    RECT 199.625 56.96 199.815 57.68 ;
    RECT 200.165 56.96 200.29 57.68 ;
    RECT 174.33 56.24 174.45 56.96 ;
    RECT 174.74 56.24 175.09 56.96 ;
    RECT 175.675 56.24 177.24 56.96 ;
    RECT 178.51 56.24 178.665 56.96 ;
    RECT 179.125 56.24 179.75 56.96 ;
    RECT 180.22 56.24 180.37 56.96 ;
    RECT 180.72 56.24 181.115 56.96 ;
    RECT 181.405 56.24 181.725 56.96 ;
    RECT 182.155 56.24 182.435 56.96 ;
    RECT 182.905 56.24 183.605 56.96 ;
    RECT 183.895 56.24 184.405 56.96 ;
    RECT 185.075 56.24 186.625 56.96 ;
    RECT 186.975 56.24 187.325 56.96 ;
    RECT 187.98 56.24 189.52 56.96 ;
    RECT 190.32 56.24 190.64 56.96 ;
    RECT 190.92 56.24 191.38 56.96 ;
    RECT 192.18 56.24 192.72 56.96 ;
    RECT 193.19 56.24 193.905 56.96 ;
    RECT 194.195 56.24 194.4 56.96 ;
    RECT 195.4 56.24 195.56 56.96 ;
    RECT 195.91 56.24 196.08 56.96 ;
    RECT 197.15 56.24 198.885 56.96 ;
    RECT 199.625 56.24 199.815 56.96 ;
    RECT 200.165 56.24 200.29 56.96 ;
    RECT 174.33 55.52 174.45 56.24 ;
    RECT 174.74 55.52 175.09 56.24 ;
    RECT 175.675 55.52 177.24 56.24 ;
    RECT 178.51 55.52 178.665 56.24 ;
    RECT 179.125 55.52 179.75 56.24 ;
    RECT 180.22 55.52 180.37 56.24 ;
    RECT 180.72 55.52 181.115 56.24 ;
    RECT 181.405 55.52 181.725 56.24 ;
    RECT 182.155 55.52 182.435 56.24 ;
    RECT 182.905 55.52 183.605 56.24 ;
    RECT 183.895 55.52 184.405 56.24 ;
    RECT 185.075 55.52 186.625 56.24 ;
    RECT 186.975 55.52 187.325 56.24 ;
    RECT 187.98 55.52 189.52 56.24 ;
    RECT 190.32 55.52 190.64 56.24 ;
    RECT 190.92 55.52 191.38 56.24 ;
    RECT 192.18 55.52 192.72 56.24 ;
    RECT 193.19 55.52 193.905 56.24 ;
    RECT 194.195 55.52 194.4 56.24 ;
    RECT 195.4 55.52 195.56 56.24 ;
    RECT 195.91 55.52 196.08 56.24 ;
    RECT 197.15 55.52 198.885 56.24 ;
    RECT 199.625 55.52 199.815 56.24 ;
    RECT 200.165 55.52 200.29 56.24 ;
    RECT 174.33 54.8 174.45 55.52 ;
    RECT 174.74 54.8 175.09 55.52 ;
    RECT 175.675 54.8 177.24 55.52 ;
    RECT 178.51 54.8 178.665 55.52 ;
    RECT 179.125 54.8 179.75 55.52 ;
    RECT 180.22 54.8 180.37 55.52 ;
    RECT 180.72 54.8 181.115 55.52 ;
    RECT 181.405 54.8 181.725 55.52 ;
    RECT 182.155 54.8 182.435 55.52 ;
    RECT 182.905 54.8 183.605 55.52 ;
    RECT 183.895 54.8 184.405 55.52 ;
    RECT 185.075 54.8 186.625 55.52 ;
    RECT 186.975 54.8 187.325 55.52 ;
    RECT 187.98 54.8 189.52 55.52 ;
    RECT 190.32 54.8 190.64 55.52 ;
    RECT 190.92 54.8 191.38 55.52 ;
    RECT 192.18 54.8 192.72 55.52 ;
    RECT 193.19 54.8 193.905 55.52 ;
    RECT 194.195 54.8 194.4 55.52 ;
    RECT 195.4 54.8 195.56 55.52 ;
    RECT 195.91 54.8 196.08 55.52 ;
    RECT 197.15 54.8 198.885 55.52 ;
    RECT 199.625 54.8 199.815 55.52 ;
    RECT 200.165 54.8 200.29 55.52 ;
    RECT 174.33 54.08 174.45 54.8 ;
    RECT 174.74 54.08 175.09 54.8 ;
    RECT 175.675 54.08 177.24 54.8 ;
    RECT 178.51 54.08 178.665 54.8 ;
    RECT 179.125 54.08 179.75 54.8 ;
    RECT 180.22 54.08 180.37 54.8 ;
    RECT 180.72 54.08 181.115 54.8 ;
    RECT 181.405 54.08 181.725 54.8 ;
    RECT 182.155 54.08 182.435 54.8 ;
    RECT 182.905 54.08 183.605 54.8 ;
    RECT 183.895 54.08 184.405 54.8 ;
    RECT 185.075 54.08 186.625 54.8 ;
    RECT 186.975 54.08 187.325 54.8 ;
    RECT 187.98 54.08 189.52 54.8 ;
    RECT 190.32 54.08 190.64 54.8 ;
    RECT 190.92 54.08 191.38 54.8 ;
    RECT 192.18 54.08 192.72 54.8 ;
    RECT 193.19 54.08 193.905 54.8 ;
    RECT 194.195 54.08 194.4 54.8 ;
    RECT 195.4 54.08 195.56 54.8 ;
    RECT 195.91 54.08 196.08 54.8 ;
    RECT 197.15 54.08 198.885 54.8 ;
    RECT 199.625 54.08 199.815 54.8 ;
    RECT 200.165 54.08 200.29 54.8 ;
    RECT 174.33 53.36 174.45 54.08 ;
    RECT 174.74 53.36 175.09 54.08 ;
    RECT 175.675 53.36 177.24 54.08 ;
    RECT 178.51 53.36 178.665 54.08 ;
    RECT 179.125 53.36 179.75 54.08 ;
    RECT 180.22 53.36 180.37 54.08 ;
    RECT 180.72 53.36 181.115 54.08 ;
    RECT 181.405 53.36 181.725 54.08 ;
    RECT 182.155 53.36 182.435 54.08 ;
    RECT 182.905 53.36 183.605 54.08 ;
    RECT 183.895 53.36 184.405 54.08 ;
    RECT 185.075 53.36 186.625 54.08 ;
    RECT 186.975 53.36 187.325 54.08 ;
    RECT 187.98 53.36 189.52 54.08 ;
    RECT 190.32 53.36 190.64 54.08 ;
    RECT 190.92 53.36 191.38 54.08 ;
    RECT 192.18 53.36 192.72 54.08 ;
    RECT 193.19 53.36 193.905 54.08 ;
    RECT 194.195 53.36 194.4 54.08 ;
    RECT 195.4 53.36 195.56 54.08 ;
    RECT 195.91 53.36 196.08 54.08 ;
    RECT 197.15 53.36 198.885 54.08 ;
    RECT 199.625 53.36 199.815 54.08 ;
    RECT 200.165 53.36 200.29 54.08 ;
    RECT 174.33 52.64 174.45 53.36 ;
    RECT 174.74 52.64 175.09 53.36 ;
    RECT 175.675 52.64 177.24 53.36 ;
    RECT 178.51 52.64 178.665 53.36 ;
    RECT 179.125 52.64 179.75 53.36 ;
    RECT 180.22 52.64 180.37 53.36 ;
    RECT 180.72 52.64 181.115 53.36 ;
    RECT 181.405 52.64 181.725 53.36 ;
    RECT 182.155 52.64 182.435 53.36 ;
    RECT 182.905 52.64 183.605 53.36 ;
    RECT 183.895 52.64 184.405 53.36 ;
    RECT 185.075 52.64 186.625 53.36 ;
    RECT 186.975 52.64 187.325 53.36 ;
    RECT 187.98 52.64 189.52 53.36 ;
    RECT 190.32 52.64 190.64 53.36 ;
    RECT 190.92 52.64 191.38 53.36 ;
    RECT 192.18 52.64 192.72 53.36 ;
    RECT 193.19 52.64 193.905 53.36 ;
    RECT 194.195 52.64 194.4 53.36 ;
    RECT 195.4 52.64 195.56 53.36 ;
    RECT 195.91 52.64 196.08 53.36 ;
    RECT 197.15 52.64 198.885 53.36 ;
    RECT 199.625 52.64 199.815 53.36 ;
    RECT 200.165 52.64 200.29 53.36 ;
    RECT 174.33 51.92 174.45 52.64 ;
    RECT 174.74 51.92 175.09 52.64 ;
    RECT 175.675 51.92 177.24 52.64 ;
    RECT 178.51 51.92 178.665 52.64 ;
    RECT 179.125 51.92 179.75 52.64 ;
    RECT 180.22 51.92 180.37 52.64 ;
    RECT 180.72 51.92 181.115 52.64 ;
    RECT 181.405 51.92 181.725 52.64 ;
    RECT 182.155 51.92 182.435 52.64 ;
    RECT 182.905 51.92 183.605 52.64 ;
    RECT 183.895 51.92 184.405 52.64 ;
    RECT 185.075 51.92 186.625 52.64 ;
    RECT 186.975 51.92 187.325 52.64 ;
    RECT 187.98 51.92 189.52 52.64 ;
    RECT 190.32 51.92 190.64 52.64 ;
    RECT 190.92 51.92 191.38 52.64 ;
    RECT 192.18 51.92 192.72 52.64 ;
    RECT 193.19 51.92 193.905 52.64 ;
    RECT 194.195 51.92 194.4 52.64 ;
    RECT 195.4 51.92 195.56 52.64 ;
    RECT 195.91 51.92 196.08 52.64 ;
    RECT 197.15 51.92 198.885 52.64 ;
    RECT 199.625 51.92 199.815 52.64 ;
    RECT 200.165 51.92 200.29 52.64 ;
    RECT 174.33 51.2 174.45 51.92 ;
    RECT 174.74 51.2 175.09 51.92 ;
    RECT 175.675 51.2 177.24 51.92 ;
    RECT 178.51 51.2 178.665 51.92 ;
    RECT 179.125 51.2 179.75 51.92 ;
    RECT 180.22 51.2 180.37 51.92 ;
    RECT 180.72 51.2 181.115 51.92 ;
    RECT 181.405 51.2 181.725 51.92 ;
    RECT 182.155 51.2 182.435 51.92 ;
    RECT 182.905 51.2 183.605 51.92 ;
    RECT 183.895 51.2 184.405 51.92 ;
    RECT 185.075 51.2 186.625 51.92 ;
    RECT 186.975 51.2 187.325 51.92 ;
    RECT 187.98 51.2 189.52 51.92 ;
    RECT 190.32 51.2 190.64 51.92 ;
    RECT 190.92 51.2 191.38 51.92 ;
    RECT 192.18 51.2 192.72 51.92 ;
    RECT 193.19 51.2 193.905 51.92 ;
    RECT 194.195 51.2 194.4 51.92 ;
    RECT 195.4 51.2 195.56 51.92 ;
    RECT 195.91 51.2 196.08 51.92 ;
    RECT 197.15 51.2 198.885 51.92 ;
    RECT 199.625 51.2 199.815 51.92 ;
    RECT 200.165 51.2 200.29 51.92 ;
    RECT 174.33 50.48 174.45 51.2 ;
    RECT 174.74 50.48 175.09 51.2 ;
    RECT 175.675 50.48 177.24 51.2 ;
    RECT 178.51 50.48 178.665 51.2 ;
    RECT 179.125 50.48 179.75 51.2 ;
    RECT 180.22 50.48 180.37 51.2 ;
    RECT 180.72 50.48 181.115 51.2 ;
    RECT 181.405 50.48 181.725 51.2 ;
    RECT 182.155 50.48 182.435 51.2 ;
    RECT 182.905 50.48 183.605 51.2 ;
    RECT 183.895 50.48 184.405 51.2 ;
    RECT 185.075 50.48 186.625 51.2 ;
    RECT 186.975 50.48 187.325 51.2 ;
    RECT 187.98 50.48 189.52 51.2 ;
    RECT 190.32 50.48 190.64 51.2 ;
    RECT 190.92 50.48 191.38 51.2 ;
    RECT 192.18 50.48 192.72 51.2 ;
    RECT 193.19 50.48 193.905 51.2 ;
    RECT 194.195 50.48 194.4 51.2 ;
    RECT 195.4 50.48 195.56 51.2 ;
    RECT 195.91 50.48 196.08 51.2 ;
    RECT 197.15 50.48 198.885 51.2 ;
    RECT 199.625 50.48 199.815 51.2 ;
    RECT 200.165 50.48 200.29 51.2 ;
    RECT 174.33 49.76 174.45 50.48 ;
    RECT 174.74 49.76 175.09 50.48 ;
    RECT 175.675 49.76 177.24 50.48 ;
    RECT 178.51 49.76 178.665 50.48 ;
    RECT 179.125 49.76 179.75 50.48 ;
    RECT 180.22 49.76 180.37 50.48 ;
    RECT 180.72 49.76 181.115 50.48 ;
    RECT 181.405 49.76 181.725 50.48 ;
    RECT 182.155 49.76 182.435 50.48 ;
    RECT 182.905 49.76 183.605 50.48 ;
    RECT 183.895 49.76 184.405 50.48 ;
    RECT 185.075 49.76 186.625 50.48 ;
    RECT 186.975 49.76 187.325 50.48 ;
    RECT 187.98 49.76 189.52 50.48 ;
    RECT 190.32 49.76 190.64 50.48 ;
    RECT 190.92 49.76 191.38 50.48 ;
    RECT 192.18 49.76 192.72 50.48 ;
    RECT 193.19 49.76 193.905 50.48 ;
    RECT 194.195 49.76 194.4 50.48 ;
    RECT 195.4 49.76 195.56 50.48 ;
    RECT 195.91 49.76 196.08 50.48 ;
    RECT 197.15 49.76 198.885 50.48 ;
    RECT 199.625 49.76 199.815 50.48 ;
    RECT 200.165 49.76 200.29 50.48 ;
    RECT 174.33 49.04 174.45 49.76 ;
    RECT 174.74 49.04 175.09 49.76 ;
    RECT 175.675 49.04 177.24 49.76 ;
    RECT 178.51 49.04 178.665 49.76 ;
    RECT 179.125 49.04 179.75 49.76 ;
    RECT 180.22 49.04 180.37 49.76 ;
    RECT 180.72 49.04 181.115 49.76 ;
    RECT 181.405 49.04 181.725 49.76 ;
    RECT 182.155 49.04 182.435 49.76 ;
    RECT 182.905 49.04 183.605 49.76 ;
    RECT 183.895 49.04 184.405 49.76 ;
    RECT 185.075 49.04 186.625 49.76 ;
    RECT 186.975 49.04 187.325 49.76 ;
    RECT 187.98 49.04 189.52 49.76 ;
    RECT 190.32 49.04 190.64 49.76 ;
    RECT 190.92 49.04 191.38 49.76 ;
    RECT 192.18 49.04 192.72 49.76 ;
    RECT 193.19 49.04 193.905 49.76 ;
    RECT 194.195 49.04 194.4 49.76 ;
    RECT 195.4 49.04 195.56 49.76 ;
    RECT 195.91 49.04 196.08 49.76 ;
    RECT 197.15 49.04 198.885 49.76 ;
    RECT 199.625 49.04 199.815 49.76 ;
    RECT 200.165 49.04 200.29 49.76 ;
    RECT 174.33 58.42 174.45 59.14 ;
    RECT 174.74 58.42 175.09 59.14 ;
    RECT 175.675 58.42 177.24 59.14 ;
    RECT 178.51 58.42 178.665 59.14 ;
    RECT 179.125 58.42 179.75 59.14 ;
    RECT 180.22 58.42 180.37 59.14 ;
    RECT 180.72 58.42 181.115 59.14 ;
    RECT 181.405 58.42 181.725 59.14 ;
    RECT 182.155 58.42 182.435 59.14 ;
    RECT 182.905 58.42 183.605 59.14 ;
    RECT 183.895 58.42 184.405 59.14 ;
    RECT 185.075 58.42 186.625 59.14 ;
    RECT 186.975 58.42 187.325 59.14 ;
    RECT 187.98 58.42 189.52 59.14 ;
    RECT 190.32 58.42 190.64 59.14 ;
    RECT 190.92 58.42 191.38 59.14 ;
    RECT 192.18 58.42 192.72 59.14 ;
    RECT 193.19 58.42 193.905 59.14 ;
    RECT 194.195 58.42 194.4 59.14 ;
    RECT 195.4 58.42 195.56 59.14 ;
    RECT 195.91 58.42 196.08 59.14 ;
    RECT 197.15 58.42 198.885 59.14 ;
    RECT 199.625 58.42 199.815 59.14 ;
    RECT 200.165 58.42 200.29 59.14 ;
    RECT 174.33 48.32 174.45 49.04 ;
    RECT 174.74 48.32 175.09 49.04 ;
    RECT 175.675 48.32 177.24 49.04 ;
    RECT 178.51 48.32 178.665 49.04 ;
    RECT 179.125 48.32 179.75 49.04 ;
    RECT 180.22 48.32 180.37 49.04 ;
    RECT 180.72 48.32 181.115 49.04 ;
    RECT 181.405 48.32 181.725 49.04 ;
    RECT 182.155 48.32 182.435 49.04 ;
    RECT 182.905 48.32 183.605 49.04 ;
    RECT 183.895 48.32 184.405 49.04 ;
    RECT 185.075 48.32 186.625 49.04 ;
    RECT 186.975 48.32 187.325 49.04 ;
    RECT 187.98 48.32 189.52 49.04 ;
    RECT 190.32 48.32 190.64 49.04 ;
    RECT 190.92 48.32 191.38 49.04 ;
    RECT 192.18 48.32 192.72 49.04 ;
    RECT 193.19 48.32 193.905 49.04 ;
    RECT 194.195 48.32 194.4 49.04 ;
    RECT 195.4 48.32 195.56 49.04 ;
    RECT 195.91 48.32 196.08 49.04 ;
    RECT 197.15 48.32 198.885 49.04 ;
    RECT 199.625 48.32 199.815 49.04 ;
    RECT 200.165 48.32 200.29 49.04 ;
    RECT 174.33 47.6 174.45 48.32 ;
    RECT 174.74 47.6 175.09 48.32 ;
    RECT 175.675 47.6 177.24 48.32 ;
    RECT 178.51 47.6 178.665 48.32 ;
    RECT 179.125 47.6 179.75 48.32 ;
    RECT 180.22 47.6 180.37 48.32 ;
    RECT 180.72 47.6 181.115 48.32 ;
    RECT 181.405 47.6 181.725 48.32 ;
    RECT 182.155 47.6 182.435 48.32 ;
    RECT 182.905 47.6 183.605 48.32 ;
    RECT 183.895 47.6 184.405 48.32 ;
    RECT 185.075 47.6 186.625 48.32 ;
    RECT 186.975 47.6 187.325 48.32 ;
    RECT 187.98 47.6 189.52 48.32 ;
    RECT 190.32 47.6 190.64 48.32 ;
    RECT 190.92 47.6 191.38 48.32 ;
    RECT 192.18 47.6 192.72 48.32 ;
    RECT 193.19 47.6 193.905 48.32 ;
    RECT 194.195 47.6 194.4 48.32 ;
    RECT 195.4 47.6 195.56 48.32 ;
    RECT 195.91 47.6 196.08 48.32 ;
    RECT 197.15 47.6 198.885 48.32 ;
    RECT 199.625 47.6 199.815 48.32 ;
    RECT 200.165 47.6 200.29 48.32 ;
    RECT 174.33 46.88 174.45 47.6 ;
    RECT 174.74 46.88 175.09 47.6 ;
    RECT 175.675 46.88 177.24 47.6 ;
    RECT 178.51 46.88 178.665 47.6 ;
    RECT 179.125 46.88 179.75 47.6 ;
    RECT 180.22 46.88 180.37 47.6 ;
    RECT 180.72 46.88 181.115 47.6 ;
    RECT 181.405 46.88 181.725 47.6 ;
    RECT 182.155 46.88 182.435 47.6 ;
    RECT 182.905 46.88 183.605 47.6 ;
    RECT 183.895 46.88 184.405 47.6 ;
    RECT 185.075 46.88 186.625 47.6 ;
    RECT 186.975 46.88 187.325 47.6 ;
    RECT 187.98 46.88 189.52 47.6 ;
    RECT 190.32 46.88 190.64 47.6 ;
    RECT 190.92 46.88 191.38 47.6 ;
    RECT 192.18 46.88 192.72 47.6 ;
    RECT 193.19 46.88 193.905 47.6 ;
    RECT 194.195 46.88 194.4 47.6 ;
    RECT 195.4 46.88 195.56 47.6 ;
    RECT 195.91 46.88 196.08 47.6 ;
    RECT 197.15 46.88 198.885 47.6 ;
    RECT 199.625 46.88 199.815 47.6 ;
    RECT 200.165 46.88 200.29 47.6 ;
    RECT 174.33 46.16 174.45 46.88 ;
    RECT 174.74 46.16 175.09 46.88 ;
    RECT 175.675 46.16 177.24 46.88 ;
    RECT 178.51 46.16 178.665 46.88 ;
    RECT 179.125 46.16 179.75 46.88 ;
    RECT 180.22 46.16 180.37 46.88 ;
    RECT 180.72 46.16 181.115 46.88 ;
    RECT 181.405 46.16 181.725 46.88 ;
    RECT 182.155 46.16 182.435 46.88 ;
    RECT 182.905 46.16 183.605 46.88 ;
    RECT 183.895 46.16 184.405 46.88 ;
    RECT 185.075 46.16 186.625 46.88 ;
    RECT 186.975 46.16 187.325 46.88 ;
    RECT 187.98 46.16 189.52 46.88 ;
    RECT 190.32 46.16 190.64 46.88 ;
    RECT 190.92 46.16 191.38 46.88 ;
    RECT 192.18 46.16 192.72 46.88 ;
    RECT 193.19 46.16 193.905 46.88 ;
    RECT 194.195 46.16 194.4 46.88 ;
    RECT 195.4 46.16 195.56 46.88 ;
    RECT 195.91 46.16 196.08 46.88 ;
    RECT 197.15 46.16 198.885 46.88 ;
    RECT 199.625 46.16 199.815 46.88 ;
    RECT 200.165 46.16 200.29 46.88 ;
    RECT 174.33 45.44 174.45 46.16 ;
    RECT 174.74 45.44 175.09 46.16 ;
    RECT 175.675 45.44 177.24 46.16 ;
    RECT 178.51 45.44 178.665 46.16 ;
    RECT 179.125 45.44 179.75 46.16 ;
    RECT 180.22 45.44 180.37 46.16 ;
    RECT 180.72 45.44 181.115 46.16 ;
    RECT 181.405 45.44 181.725 46.16 ;
    RECT 182.155 45.44 182.435 46.16 ;
    RECT 182.905 45.44 183.605 46.16 ;
    RECT 183.895 45.44 184.405 46.16 ;
    RECT 185.075 45.44 186.625 46.16 ;
    RECT 186.975 45.44 187.325 46.16 ;
    RECT 187.98 45.44 189.52 46.16 ;
    RECT 190.32 45.44 190.64 46.16 ;
    RECT 190.92 45.44 191.38 46.16 ;
    RECT 192.18 45.44 192.72 46.16 ;
    RECT 193.19 45.44 193.905 46.16 ;
    RECT 194.195 45.44 194.4 46.16 ;
    RECT 195.4 45.44 195.56 46.16 ;
    RECT 195.91 45.44 196.08 46.16 ;
    RECT 197.15 45.44 198.885 46.16 ;
    RECT 199.625 45.44 199.815 46.16 ;
    RECT 200.165 45.44 200.29 46.16 ;
    RECT 174.33 44.72 174.45 45.44 ;
    RECT 174.74 44.72 175.09 45.44 ;
    RECT 175.675 44.72 177.24 45.44 ;
    RECT 178.51 44.72 178.665 45.44 ;
    RECT 179.125 44.72 179.75 45.44 ;
    RECT 180.22 44.72 180.37 45.44 ;
    RECT 180.72 44.72 181.115 45.44 ;
    RECT 181.405 44.72 181.725 45.44 ;
    RECT 182.155 44.72 182.435 45.44 ;
    RECT 182.905 44.72 183.605 45.44 ;
    RECT 183.895 44.72 184.405 45.44 ;
    RECT 185.075 44.72 186.625 45.44 ;
    RECT 186.975 44.72 187.325 45.44 ;
    RECT 187.98 44.72 189.52 45.44 ;
    RECT 190.32 44.72 190.64 45.44 ;
    RECT 190.92 44.72 191.38 45.44 ;
    RECT 192.18 44.72 192.72 45.44 ;
    RECT 193.19 44.72 193.905 45.44 ;
    RECT 194.195 44.72 194.4 45.44 ;
    RECT 195.4 44.72 195.56 45.44 ;
    RECT 195.91 44.72 196.08 45.44 ;
    RECT 197.15 44.72 198.885 45.44 ;
    RECT 199.625 44.72 199.815 45.44 ;
    RECT 200.165 44.72 200.29 45.44 ;
    RECT 174.33 44.0 174.45 44.72 ;
    RECT 174.74 44.0 175.09 44.72 ;
    RECT 175.675 44.0 177.24 44.72 ;
    RECT 178.51 44.0 178.665 44.72 ;
    RECT 179.125 44.0 179.75 44.72 ;
    RECT 180.22 44.0 180.37 44.72 ;
    RECT 180.72 44.0 181.115 44.72 ;
    RECT 181.405 44.0 181.725 44.72 ;
    RECT 182.155 44.0 182.435 44.72 ;
    RECT 182.905 44.0 183.605 44.72 ;
    RECT 183.895 44.0 184.405 44.72 ;
    RECT 185.075 44.0 186.625 44.72 ;
    RECT 186.975 44.0 187.325 44.72 ;
    RECT 187.98 44.0 189.52 44.72 ;
    RECT 190.32 44.0 190.64 44.72 ;
    RECT 190.92 44.0 191.38 44.72 ;
    RECT 192.18 44.0 192.72 44.72 ;
    RECT 193.19 44.0 193.905 44.72 ;
    RECT 194.195 44.0 194.4 44.72 ;
    RECT 195.4 44.0 195.56 44.72 ;
    RECT 195.91 44.0 196.08 44.72 ;
    RECT 197.15 44.0 198.885 44.72 ;
    RECT 199.625 44.0 199.815 44.72 ;
    RECT 200.165 44.0 200.29 44.72 ;
    RECT 174.33 43.28 174.45 44.0 ;
    RECT 174.74 43.28 175.09 44.0 ;
    RECT 175.675 43.28 177.24 44.0 ;
    RECT 178.51 43.28 178.665 44.0 ;
    RECT 179.125 43.28 179.75 44.0 ;
    RECT 180.22 43.28 180.37 44.0 ;
    RECT 180.72 43.28 181.115 44.0 ;
    RECT 181.405 43.28 181.725 44.0 ;
    RECT 182.155 43.28 182.435 44.0 ;
    RECT 182.905 43.28 183.605 44.0 ;
    RECT 183.895 43.28 184.405 44.0 ;
    RECT 185.075 43.28 186.625 44.0 ;
    RECT 186.975 43.28 187.325 44.0 ;
    RECT 187.98 43.28 189.52 44.0 ;
    RECT 190.32 43.28 190.64 44.0 ;
    RECT 190.92 43.28 191.38 44.0 ;
    RECT 192.18 43.28 192.72 44.0 ;
    RECT 193.19 43.28 193.905 44.0 ;
    RECT 194.195 43.28 194.4 44.0 ;
    RECT 195.4 43.28 195.56 44.0 ;
    RECT 195.91 43.28 196.08 44.0 ;
    RECT 197.15 43.28 198.885 44.0 ;
    RECT 199.625 43.28 199.815 44.0 ;
    RECT 200.165 43.28 200.29 44.0 ;
    RECT 174.33 42.56 174.45 43.28 ;
    RECT 174.74 42.56 175.09 43.28 ;
    RECT 175.675 42.56 177.24 43.28 ;
    RECT 178.51 42.56 178.665 43.28 ;
    RECT 179.125 42.56 179.75 43.28 ;
    RECT 180.22 42.56 180.37 43.28 ;
    RECT 180.72 42.56 181.115 43.28 ;
    RECT 181.405 42.56 181.725 43.28 ;
    RECT 182.155 42.56 182.435 43.28 ;
    RECT 182.905 42.56 183.605 43.28 ;
    RECT 183.895 42.56 184.405 43.28 ;
    RECT 185.075 42.56 186.625 43.28 ;
    RECT 186.975 42.56 187.325 43.28 ;
    RECT 187.98 42.56 189.52 43.28 ;
    RECT 190.32 42.56 190.64 43.28 ;
    RECT 190.92 42.56 191.38 43.28 ;
    RECT 192.18 42.56 192.72 43.28 ;
    RECT 193.19 42.56 193.905 43.28 ;
    RECT 194.195 42.56 194.4 43.28 ;
    RECT 195.4 42.56 195.56 43.28 ;
    RECT 195.91 42.56 196.08 43.28 ;
    RECT 197.15 42.56 198.885 43.28 ;
    RECT 199.625 42.56 199.815 43.28 ;
    RECT 200.165 42.56 200.29 43.28 ;
    RECT 174.33 41.84 174.45 42.56 ;
    RECT 174.74 41.84 175.09 42.56 ;
    RECT 175.675 41.84 177.24 42.56 ;
    RECT 178.51 41.84 178.665 42.56 ;
    RECT 179.125 41.84 179.75 42.56 ;
    RECT 180.22 41.84 180.37 42.56 ;
    RECT 180.72 41.84 181.115 42.56 ;
    RECT 181.405 41.84 181.725 42.56 ;
    RECT 182.155 41.84 182.435 42.56 ;
    RECT 182.905 41.84 183.605 42.56 ;
    RECT 183.895 41.84 184.405 42.56 ;
    RECT 185.075 41.84 186.625 42.56 ;
    RECT 186.975 41.84 187.325 42.56 ;
    RECT 187.98 41.84 189.52 42.56 ;
    RECT 190.32 41.84 190.64 42.56 ;
    RECT 190.92 41.84 191.38 42.56 ;
    RECT 192.18 41.84 192.72 42.56 ;
    RECT 193.19 41.84 193.905 42.56 ;
    RECT 194.195 41.84 194.4 42.56 ;
    RECT 195.4 41.84 195.56 42.56 ;
    RECT 195.91 41.84 196.08 42.56 ;
    RECT 197.15 41.84 198.885 42.56 ;
    RECT 199.625 41.84 199.815 42.56 ;
    RECT 200.165 41.84 200.29 42.56 ;
    RECT 174.33 57.68 174.45 58.42 ;
    RECT 174.74 57.68 175.09 58.42 ;
    RECT 175.675 57.68 177.24 58.42 ;
    RECT 178.51 57.68 178.665 58.42 ;
    RECT 179.125 57.68 179.75 58.42 ;
    RECT 180.22 57.68 180.37 58.42 ;
    RECT 180.72 57.68 181.115 58.42 ;
    RECT 181.405 57.68 181.725 58.42 ;
    RECT 182.155 57.68 182.435 58.42 ;
    RECT 182.905 57.68 183.605 58.42 ;
    RECT 183.895 57.68 184.405 58.42 ;
    RECT 184.875 57.68 186.625 58.42 ;
    RECT 186.975 57.68 187.325 58.42 ;
    RECT 187.98 57.68 189.52 58.42 ;
    RECT 190.32 57.68 190.64 58.42 ;
    RECT 190.92 57.68 191.38 58.42 ;
    RECT 192.18 57.68 192.72 58.42 ;
    RECT 193.19 57.68 193.905 58.42 ;
    RECT 194.195 57.68 194.4 58.42 ;
    RECT 195.4 57.68 195.56 58.42 ;
    RECT 195.91 57.68 196.08 58.42 ;
    RECT 197.15 57.68 198.885 58.42 ;
    RECT 199.625 57.68 199.815 58.42 ;
    RECT 200.165 57.68 200.29 58.42 ;
    RECT 174.33 41.12 174.45 41.84 ;
    RECT 174.74 41.12 175.09 41.84 ;
    RECT 175.675 41.12 177.24 41.84 ;
    RECT 178.51 41.12 178.665 41.84 ;
    RECT 179.125 41.12 179.75 41.84 ;
    RECT 180.22 41.12 180.37 41.84 ;
    RECT 180.72 41.12 181.115 41.84 ;
    RECT 181.405 41.12 181.725 41.84 ;
    RECT 182.155 41.12 182.435 41.84 ;
    RECT 182.905 41.12 183.605 41.84 ;
    RECT 183.895 41.12 184.405 41.84 ;
    RECT 185.075 41.12 186.625 41.84 ;
    RECT 186.975 41.12 187.325 41.84 ;
    RECT 187.98 41.12 189.52 41.84 ;
    RECT 190.32 41.12 190.64 41.84 ;
    RECT 190.92 41.12 191.38 41.84 ;
    RECT 192.18 41.12 192.72 41.84 ;
    RECT 193.19 41.12 193.905 41.84 ;
    RECT 194.195 41.12 194.4 41.84 ;
    RECT 195.4 41.12 195.56 41.84 ;
    RECT 195.91 41.12 196.08 41.84 ;
    RECT 197.15 41.12 198.885 41.84 ;
    RECT 199.625 41.12 199.815 41.84 ;
    RECT 200.165 41.12 200.29 41.84 ;
    RECT 174.33 40.4 174.45 41.12 ;
    RECT 174.74 40.4 175.09 41.12 ;
    RECT 175.675 40.4 177.24 41.12 ;
    RECT 178.51 40.4 178.665 41.12 ;
    RECT 179.125 40.4 179.75 41.12 ;
    RECT 180.22 40.4 180.37 41.12 ;
    RECT 180.72 40.4 181.115 41.12 ;
    RECT 181.405 40.4 181.725 41.12 ;
    RECT 182.155 40.4 182.435 41.12 ;
    RECT 182.905 40.4 183.605 41.12 ;
    RECT 183.895 40.4 184.405 41.12 ;
    RECT 185.075 40.4 186.625 41.12 ;
    RECT 186.975 40.4 187.325 41.12 ;
    RECT 187.98 40.4 189.52 41.12 ;
    RECT 190.32 40.4 190.64 41.12 ;
    RECT 190.92 40.4 191.38 41.12 ;
    RECT 192.18 40.4 192.72 41.12 ;
    RECT 193.19 40.4 193.905 41.12 ;
    RECT 194.195 40.4 194.4 41.12 ;
    RECT 195.4 40.4 195.56 41.12 ;
    RECT 195.91 40.4 196.08 41.12 ;
    RECT 197.15 40.4 198.885 41.12 ;
    RECT 199.625 40.4 199.815 41.12 ;
    RECT 200.165 40.4 200.29 41.12 ;
    RECT 174.33 39.68 174.45 40.4 ;
    RECT 174.74 39.68 175.09 40.4 ;
    RECT 175.675 39.68 177.24 40.4 ;
    RECT 178.51 39.68 178.665 40.4 ;
    RECT 179.125 39.68 179.75 40.4 ;
    RECT 180.22 39.68 180.37 40.4 ;
    RECT 180.72 39.68 181.115 40.4 ;
    RECT 181.405 39.68 181.725 40.4 ;
    RECT 182.155 39.68 182.435 40.4 ;
    RECT 182.905 39.68 183.605 40.4 ;
    RECT 183.895 39.68 184.405 40.4 ;
    RECT 185.075 39.68 186.625 40.4 ;
    RECT 186.975 39.68 187.325 40.4 ;
    RECT 187.98 39.68 189.52 40.4 ;
    RECT 190.32 39.68 190.64 40.4 ;
    RECT 190.92 39.68 191.38 40.4 ;
    RECT 192.18 39.68 192.72 40.4 ;
    RECT 193.19 39.68 193.905 40.4 ;
    RECT 194.195 39.68 194.4 40.4 ;
    RECT 195.4 39.68 195.56 40.4 ;
    RECT 195.91 39.68 196.08 40.4 ;
    RECT 197.15 39.68 198.885 40.4 ;
    RECT 199.625 39.68 199.815 40.4 ;
    RECT 200.165 39.68 200.29 40.4 ;
    RECT 174.33 38.96 174.45 39.68 ;
    RECT 174.74 38.96 175.09 39.68 ;
    RECT 175.675 38.96 177.24 39.68 ;
    RECT 178.51 38.96 178.665 39.68 ;
    RECT 179.125 38.96 179.75 39.68 ;
    RECT 180.22 38.96 180.37 39.68 ;
    RECT 180.72 38.96 181.115 39.68 ;
    RECT 181.405 38.96 181.725 39.68 ;
    RECT 182.155 38.96 182.435 39.68 ;
    RECT 182.905 38.96 183.605 39.68 ;
    RECT 183.895 38.96 184.405 39.68 ;
    RECT 185.075 38.96 186.625 39.68 ;
    RECT 186.975 38.96 187.325 39.68 ;
    RECT 187.98 38.96 189.52 39.68 ;
    RECT 190.32 38.96 190.64 39.68 ;
    RECT 190.92 38.96 191.38 39.68 ;
    RECT 192.18 38.96 192.72 39.68 ;
    RECT 193.19 38.96 193.905 39.68 ;
    RECT 194.195 38.96 194.4 39.68 ;
    RECT 195.4 38.96 195.56 39.68 ;
    RECT 195.91 38.96 196.08 39.68 ;
    RECT 197.15 38.96 198.885 39.68 ;
    RECT 199.625 38.96 199.815 39.68 ;
    RECT 200.165 38.96 200.29 39.68 ;
    RECT 174.33 38.24 174.45 38.96 ;
    RECT 174.74 38.24 175.09 38.96 ;
    RECT 175.675 38.24 177.24 38.96 ;
    RECT 178.51 38.24 178.665 38.96 ;
    RECT 179.125 38.24 179.75 38.96 ;
    RECT 180.22 38.24 180.37 38.96 ;
    RECT 180.72 38.24 181.115 38.96 ;
    RECT 181.405 38.24 181.725 38.96 ;
    RECT 182.155 38.24 182.435 38.96 ;
    RECT 182.905 38.24 183.605 38.96 ;
    RECT 183.895 38.24 184.405 38.96 ;
    RECT 185.075 38.24 186.625 38.96 ;
    RECT 186.975 38.24 187.325 38.96 ;
    RECT 187.98 38.24 189.52 38.96 ;
    RECT 190.32 38.24 190.64 38.96 ;
    RECT 190.92 38.24 191.38 38.96 ;
    RECT 192.18 38.24 192.72 38.96 ;
    RECT 193.19 38.24 193.905 38.96 ;
    RECT 194.195 38.24 194.4 38.96 ;
    RECT 195.4 38.24 195.56 38.96 ;
    RECT 195.91 38.24 196.08 38.96 ;
    RECT 197.15 38.24 198.885 38.96 ;
    RECT 199.625 38.24 199.815 38.96 ;
    RECT 200.165 38.24 200.29 38.96 ;
    RECT 174.33 37.52 174.45 38.24 ;
    RECT 174.74 37.52 175.09 38.24 ;
    RECT 175.675 37.52 177.24 38.24 ;
    RECT 178.51 37.52 178.665 38.24 ;
    RECT 179.125 37.52 179.75 38.24 ;
    RECT 180.22 37.52 180.37 38.24 ;
    RECT 180.72 37.52 181.115 38.24 ;
    RECT 181.405 37.52 181.725 38.24 ;
    RECT 182.155 37.52 182.435 38.24 ;
    RECT 182.905 37.52 183.605 38.24 ;
    RECT 183.895 37.52 184.405 38.24 ;
    RECT 185.075 37.52 186.625 38.24 ;
    RECT 186.975 37.52 187.325 38.24 ;
    RECT 187.98 37.52 189.52 38.24 ;
    RECT 190.32 37.52 190.64 38.24 ;
    RECT 190.92 37.52 191.38 38.24 ;
    RECT 192.18 37.52 192.72 38.24 ;
    RECT 193.19 37.52 193.905 38.24 ;
    RECT 194.195 37.52 194.4 38.24 ;
    RECT 195.4 37.52 195.56 38.24 ;
    RECT 195.91 37.52 196.08 38.24 ;
    RECT 197.15 37.52 198.885 38.24 ;
    RECT 199.625 37.52 199.815 38.24 ;
    RECT 200.165 37.52 200.29 38.24 ;
    RECT 174.33 36.8 174.45 37.52 ;
    RECT 174.74 36.8 175.09 37.52 ;
    RECT 175.675 36.8 177.24 37.52 ;
    RECT 178.51 36.8 178.665 37.52 ;
    RECT 179.125 36.8 179.75 37.52 ;
    RECT 180.22 36.8 180.37 37.52 ;
    RECT 180.72 36.8 181.115 37.52 ;
    RECT 181.405 36.8 181.725 37.52 ;
    RECT 182.155 36.8 182.435 37.52 ;
    RECT 182.905 36.8 183.605 37.52 ;
    RECT 183.895 36.8 184.405 37.52 ;
    RECT 185.075 36.8 186.625 37.52 ;
    RECT 186.975 36.8 187.325 37.52 ;
    RECT 187.98 36.8 189.52 37.52 ;
    RECT 190.32 36.8 190.64 37.52 ;
    RECT 190.92 36.8 191.38 37.52 ;
    RECT 192.18 36.8 192.72 37.52 ;
    RECT 193.19 36.8 193.905 37.52 ;
    RECT 194.195 36.8 194.4 37.52 ;
    RECT 195.4 36.8 195.56 37.52 ;
    RECT 195.91 36.8 196.08 37.52 ;
    RECT 197.15 36.8 198.885 37.52 ;
    RECT 199.625 36.8 199.815 37.52 ;
    RECT 200.165 36.8 200.29 37.52 ;
    RECT 174.33 36.08 174.45 36.8 ;
    RECT 174.74 36.08 175.09 36.8 ;
    RECT 175.675 36.08 177.24 36.8 ;
    RECT 178.51 36.08 178.665 36.8 ;
    RECT 179.125 36.08 179.75 36.8 ;
    RECT 180.22 36.08 180.37 36.8 ;
    RECT 180.72 36.08 181.115 36.8 ;
    RECT 181.405 36.08 181.725 36.8 ;
    RECT 182.155 36.08 182.435 36.8 ;
    RECT 182.905 36.08 183.605 36.8 ;
    RECT 183.895 36.08 184.405 36.8 ;
    RECT 185.075 36.08 186.625 36.8 ;
    RECT 186.975 36.08 187.325 36.8 ;
    RECT 187.98 36.08 189.52 36.8 ;
    RECT 190.32 36.08 190.64 36.8 ;
    RECT 190.92 36.08 191.38 36.8 ;
    RECT 192.18 36.08 192.72 36.8 ;
    RECT 193.19 36.08 193.905 36.8 ;
    RECT 194.195 36.08 194.4 36.8 ;
    RECT 195.4 36.08 195.56 36.8 ;
    RECT 195.91 36.08 196.08 36.8 ;
    RECT 197.15 36.08 198.885 36.8 ;
    RECT 199.625 36.08 199.815 36.8 ;
    RECT 200.165 36.08 200.29 36.8 ;
    RECT 174.33 35.36 174.45 36.08 ;
    RECT 174.74 35.36 175.09 36.08 ;
    RECT 175.675 35.36 177.24 36.08 ;
    RECT 178.51 35.36 178.665 36.08 ;
    RECT 179.125 35.36 179.75 36.08 ;
    RECT 180.22 35.36 180.37 36.08 ;
    RECT 180.72 35.36 181.115 36.08 ;
    RECT 181.405 35.36 181.725 36.08 ;
    RECT 182.155 35.36 182.435 36.08 ;
    RECT 182.905 35.36 183.605 36.08 ;
    RECT 183.895 35.36 184.405 36.08 ;
    RECT 185.075 35.36 186.625 36.08 ;
    RECT 186.975 35.36 187.325 36.08 ;
    RECT 187.98 35.36 189.52 36.08 ;
    RECT 190.32 35.36 190.64 36.08 ;
    RECT 190.92 35.36 191.38 36.08 ;
    RECT 192.18 35.36 192.72 36.08 ;
    RECT 193.19 35.36 193.905 36.08 ;
    RECT 194.195 35.36 194.4 36.08 ;
    RECT 195.4 35.36 195.56 36.08 ;
    RECT 195.91 35.36 196.08 36.08 ;
    RECT 197.15 35.36 198.885 36.08 ;
    RECT 199.625 35.36 199.815 36.08 ;
    RECT 200.165 35.36 200.29 36.08 ;
    RECT 174.33 34.64 174.45 35.36 ;
    RECT 174.74 34.64 175.09 35.36 ;
    RECT 175.675 34.64 177.24 35.36 ;
    RECT 178.51 34.64 178.665 35.36 ;
    RECT 179.125 34.64 179.75 35.36 ;
    RECT 180.22 34.64 180.37 35.36 ;
    RECT 180.72 34.64 181.115 35.36 ;
    RECT 181.405 34.64 181.725 35.36 ;
    RECT 182.155 34.64 182.435 35.36 ;
    RECT 182.905 34.64 183.605 35.36 ;
    RECT 183.895 34.64 184.405 35.36 ;
    RECT 185.075 34.64 186.625 35.36 ;
    RECT 186.975 34.64 187.325 35.36 ;
    RECT 187.98 34.64 189.52 35.36 ;
    RECT 190.32 34.64 190.64 35.36 ;
    RECT 190.92 34.64 191.38 35.36 ;
    RECT 192.18 34.64 192.72 35.36 ;
    RECT 193.19 34.64 193.905 35.36 ;
    RECT 194.195 34.64 194.4 35.36 ;
    RECT 195.4 34.64 195.56 35.36 ;
    RECT 195.91 34.64 196.08 35.36 ;
    RECT 197.15 34.64 198.885 35.36 ;
    RECT 199.625 34.64 199.815 35.36 ;
    RECT 200.165 34.64 200.29 35.36 ;
    RECT 174.33 11.6 174.45 34.64 ;
    RECT 174.74 11.6 175.09 34.64 ;
    RECT 175.675 11.6 177.24 34.64 ;
    RECT 178.51 11.6 178.665 34.64 ;
    RECT 179.125 11.6 179.75 34.64 ;
    RECT 180.22 11.6 180.37 34.64 ;
    RECT 180.72 11.6 181.115 34.64 ;
    RECT 181.405 29.31 181.725 34.64 ;
    RECT 182.155 11.6 182.435 34.64 ;
    RECT 182.905 11.6 183.605 34.64 ;
    RECT 183.895 11.6 184.405 34.64 ;
    RECT 184.875 12.39 185.075 23.5 ;
    RECT 184.875 24.775 185.075 25.66 ;
    RECT 184.875 27.655 185.075 33.58 ;
    RECT 185.075 11.6 185.1 34.64 ;
    RECT 185.1 11.6 185.2 34.785 ;
    RECT 185.2 11.6 185.3 34.64 ;
    RECT 185.3 11.6 185.4 34.785 ;
    RECT 185.4 11.6 185.5 34.64 ;
    RECT 185.5 11.6 185.6 34.785 ;
    RECT 185.6 11.6 185.7 34.64 ;
    RECT 185.7 11.6 185.8 34.785 ;
    RECT 185.8 11.6 185.895 34.64 ;
    RECT 185.895 11.6 185.995 34.785 ;
    RECT 185.995 11.6 186.095 34.64 ;
    RECT 186.095 11.6 186.195 34.785 ;
    RECT 186.195 11.6 186.295 34.64 ;
    RECT 186.295 11.6 186.395 34.785 ;
    RECT 186.395 11.6 186.495 34.64 ;
    RECT 186.495 11.6 186.595 34.785 ;
    RECT 186.595 11.6 186.625 34.64 ;
    RECT 186.975 11.6 187.325 34.64 ;
    RECT 187.805 11.6 187.98 33.58 ;
    RECT 187.98 11.6 188.01 34.64 ;
    RECT 188.01 11.6 188.11 34.785 ;
    RECT 188.11 11.6 188.21 34.64 ;
    RECT 188.21 11.6 188.31 34.785 ;
    RECT 188.31 11.6 188.41 34.64 ;
    RECT 188.41 11.6 188.51 34.785 ;
    RECT 188.51 11.6 188.605 34.64 ;
    RECT 188.605 11.6 188.705 34.785 ;
    RECT 188.705 11.6 188.805 34.64 ;
    RECT 188.805 11.6 188.905 34.785 ;
    RECT 188.905 11.6 189.005 34.64 ;
    RECT 189.005 11.6 189.105 34.785 ;
    RECT 189.105 11.6 189.205 34.64 ;
    RECT 189.205 11.6 189.305 34.785 ;
    RECT 189.305 11.6 189.4 34.64 ;
    RECT 189.4 11.6 189.5 34.785 ;
    RECT 189.5 11.6 189.52 34.64 ;
    RECT 190.32 11.6 190.64 34.64 ;
    RECT 190.92 11.6 191.38 34.64 ;
    RECT 192.18 11.6 192.72 34.64 ;
    RECT 193.19 11.6 193.905 34.64 ;
    RECT 194.195 11.6 194.4 34.64 ;
    RECT 195.4 11.6 195.56 34.64 ;
    RECT 195.91 11.6 196.08 34.64 ;
    RECT 197.15 11.6 198.885 34.64 ;
    RECT 199.625 11.6 199.815 34.64 ;
    RECT 200.165 11.6 200.29 34.64 ;
    RECT 174.33 59.14 174.45 60.67 ;
    RECT 174.74 59.14 175.09 60.105 ;
    RECT 175.675 59.14 177.24 60.67 ;
    RECT 178.51 59.14 178.665 60.67 ;
    RECT 179.125 59.14 179.75 60.67 ;
    RECT 180.22 59.14 180.37 60.67 ;
    RECT 180.72 59.14 181.115 60.67 ;
    RECT 181.405 59.14 181.725 60.67 ;
    RECT 182.155 59.14 182.435 60.67 ;
    RECT 182.905 59.14 183.605 60.67 ;
    RECT 183.895 59.14 184.405 60.67 ;
    RECT 185.075 59.14 185.1 60.67 ;
    RECT 185.1 59.115 185.2 60.67 ;
    RECT 185.2 59.14 186.625 60.67 ;
    RECT 186.975 59.14 187.325 60.67 ;
    RECT 187.98 59.14 189.52 60.67 ;
    RECT 190.32 59.14 190.64 60.67 ;
    RECT 190.92 59.14 191.38 60.67 ;
    RECT 192.18 59.14 192.72 60.67 ;
    RECT 193.19 59.14 193.905 60.67 ;
    RECT 194.195 59.14 194.4 60.67 ;
    RECT 195.4 59.14 195.56 60.67 ;
    RECT 195.91 59.14 196.08 60.67 ;
    RECT 197.15 59.14 198.885 60.67 ;
    RECT 199.625 59.14 199.815 60.67 ;
    RECT 200.165 59.14 200.29 60.67 ;
    RECT 366.31 4.77 366.38 9.56 ;
    RECT 364.835 2.31 365.115 8.3 ;
    RECT 362.99 4.77 363.06 9.56 ;
    RECT 361.515 2.31 361.795 8.3 ;
    RECT 359.67 4.77 359.74 9.56 ;
    RECT 358.195 2.31 358.475 8.3 ;
    RECT 356.35 4.77 356.42 9.56 ;
    RECT 354.875 2.31 355.155 8.3 ;
    RECT 353.03 4.77 353.1 9.56 ;
    RECT 351.555 2.31 351.835 8.3 ;
    RECT 349.71 4.77 349.78 9.56 ;
    RECT 348.235 2.31 348.515 8.3 ;
    RECT 346.39 4.77 346.46 9.56 ;
    RECT 344.915 2.31 345.195 8.3 ;
    RECT 343.07 4.77 343.14 9.56 ;
    RECT 341.595 2.31 341.875 8.3 ;
    RECT 339.75 4.77 339.82 9.56 ;
    RECT 338.275 2.31 338.555 8.3 ;
    RECT 336.43 4.77 336.5 9.56 ;
    RECT 334.955 2.31 335.235 8.3 ;
    RECT 333.11 4.77 333.18 9.56 ;
    RECT 331.635 2.31 331.915 8.3 ;
    RECT 329.79 4.77 329.86 9.56 ;
    RECT 328.315 2.31 328.595 8.3 ;
    RECT 326.47 4.77 326.54 9.56 ;
    RECT 324.995 2.31 325.275 8.3 ;
    RECT 323.15 4.77 323.22 9.56 ;
    RECT 321.675 2.31 321.955 8.3 ;
    RECT 319.83 4.77 319.9 9.56 ;
    RECT 318.355 2.31 318.635 8.3 ;
    RECT 316.51 4.77 316.58 9.56 ;
    RECT 315.035 2.31 315.315 8.3 ;
    RECT 313.19 4.77 313.26 9.56 ;
    RECT 311.715 2.31 311.995 8.3 ;
    RECT 309.87 4.77 309.94 9.56 ;
    RECT 308.395 2.31 308.675 8.3 ;
    RECT 306.55 4.77 306.62 9.56 ;
    RECT 305.075 2.31 305.355 8.3 ;
    RECT 303.23 4.77 303.3 9.56 ;
    RECT 301.755 2.31 302.035 8.3 ;
    RECT 233.51 4.77 233.58 9.56 ;
    RECT 232.035 2.31 232.315 8.3 ;
    RECT 230.19 4.77 230.26 9.56 ;
    RECT 228.715 2.31 228.995 8.3 ;
    RECT 226.87 4.77 226.94 9.56 ;
    RECT 225.395 2.31 225.675 8.3 ;
    RECT 223.55 4.77 223.62 9.56 ;
    RECT 222.075 2.31 222.355 8.3 ;
    RECT 220.23 4.77 220.3 9.56 ;
    RECT 218.755 2.31 219.035 8.3 ;
    RECT 299.91 4.77 299.98 9.56 ;
    RECT 298.435 2.31 298.715 8.3 ;
    RECT 216.91 4.77 216.98 9.56 ;
    RECT 215.435 2.31 215.715 8.3 ;
    RECT 296.59 4.77 296.66 9.56 ;
    RECT 295.115 2.31 295.395 8.3 ;
    RECT 213.59 4.77 213.66 9.56 ;
    RECT 212.115 2.31 212.395 8.3 ;
    RECT 293.27 4.77 293.34 9.56 ;
    RECT 291.795 2.31 292.075 8.3 ;
    RECT 210.27 4.77 210.34 9.56 ;
    RECT 208.795 2.31 209.075 8.3 ;
    RECT 289.95 4.77 290.02 9.56 ;
    RECT 288.475 2.31 288.755 8.3 ;
    RECT 206.95 4.77 207.02 9.56 ;
    RECT 205.475 2.31 205.755 8.3 ;
    RECT 286.63 4.77 286.7 9.56 ;
    RECT 285.155 2.31 285.435 8.3 ;
    RECT 283.31 4.77 283.38 9.56 ;
    RECT 281.835 2.31 282.115 8.3 ;
    RECT 279.99 4.77 280.06 9.56 ;
    RECT 278.515 2.31 278.795 8.3 ;
    RECT 276.67 4.77 276.74 9.56 ;
    RECT 275.195 2.31 275.475 8.3 ;
    RECT 273.35 4.77 273.42 9.56 ;
    RECT 271.875 2.31 272.155 8.3 ;
    RECT 270.03 4.77 270.1 9.56 ;
    RECT 268.555 2.31 268.835 8.3 ;
    RECT 266.71 4.77 266.78 9.56 ;
    RECT 265.235 2.31 265.515 8.3 ;
    RECT 263.39 4.77 263.46 9.56 ;
    RECT 261.915 2.31 262.195 8.3 ;
    RECT 260.07 4.77 260.14 9.56 ;
    RECT 258.595 2.31 258.875 8.3 ;
    RECT 256.75 4.77 256.82 9.56 ;
    RECT 255.275 2.31 255.555 8.3 ;
    RECT 253.43 4.77 253.5 9.56 ;
    RECT 251.955 2.31 252.235 8.3 ;
    RECT 250.11 4.77 250.18 9.56 ;
    RECT 248.635 2.31 248.915 8.3 ;
    RECT 246.79 4.77 246.86 9.56 ;
    RECT 245.315 2.31 245.595 8.3 ;
    RECT 243.47 4.77 243.54 9.56 ;
    RECT 241.995 2.31 242.275 8.3 ;
    RECT 240.15 4.77 240.22 9.56 ;
    RECT 238.675 2.31 238.955 8.3 ;
    RECT 236.83 4.77 236.9 9.56 ;
    RECT 235.355 2.31 235.635 8.3 ;
    RECT 372.95 4.77 373.02 9.56 ;
    RECT 371.475 2.31 371.755 8.3 ;
    RECT 203.63 4.77 203.7 9.56 ;
    RECT 202.155 2.31 202.435 8.3 ;
    RECT 369.63 4.77 369.7 9.56 ;
    RECT 368.155 2.31 368.435 8.3 ;
    RECT 369.63 0.895 369.9 2.195 ;
    RECT 368.155 0.695 368.435 2.31 ;
    RECT 366.31 0.895 366.58 2.195 ;
    RECT 364.835 0.695 365.115 2.31 ;
    RECT 362.99 0.895 363.26 2.195 ;
    RECT 361.515 0.695 361.795 2.31 ;
    RECT 359.67 0.895 359.94 2.195 ;
    RECT 358.195 0.695 358.475 2.31 ;
    RECT 356.35 0.895 356.62 2.195 ;
    RECT 354.875 0.695 355.155 2.31 ;
    RECT 353.03 0.895 353.3 2.195 ;
    RECT 351.555 0.695 351.835 2.31 ;
    RECT 349.71 0.895 349.98 2.195 ;
    RECT 348.235 0.695 348.515 2.31 ;
    RECT 346.39 0.895 346.66 2.195 ;
    RECT 344.915 0.695 345.195 2.31 ;
    RECT 343.07 0.895 343.34 2.195 ;
    RECT 341.595 0.695 341.875 2.31 ;
    RECT 339.75 0.895 340.02 2.195 ;
    RECT 338.275 0.695 338.555 2.31 ;
    RECT 336.43 0.895 336.7 2.195 ;
    RECT 334.955 0.695 335.235 2.31 ;
    RECT 333.11 0.895 333.38 2.195 ;
    RECT 331.635 0.695 331.915 2.31 ;
    RECT 329.79 0.895 330.06 2.195 ;
    RECT 328.315 0.695 328.595 2.31 ;
    RECT 326.47 0.895 326.74 2.195 ;
    RECT 324.995 0.695 325.275 2.31 ;
    RECT 323.15 0.895 323.42 2.195 ;
    RECT 321.675 0.695 321.955 2.31 ;
    RECT 319.83 0.895 320.1 2.195 ;
    RECT 318.355 0.695 318.635 2.31 ;
    RECT 316.51 0.895 316.78 2.195 ;
    RECT 315.035 0.695 315.315 2.31 ;
    RECT 313.19 0.895 313.46 2.195 ;
    RECT 311.715 0.695 311.995 2.31 ;
    RECT 309.87 0.895 310.14 2.195 ;
    RECT 308.395 0.695 308.675 2.31 ;
    RECT 306.55 0.895 306.82 2.195 ;
    RECT 305.075 0.695 305.355 2.31 ;
    RECT 303.23 0.895 303.5 2.195 ;
    RECT 301.755 0.695 302.035 2.31 ;
    RECT 299.91 0.895 300.18 2.195 ;
    RECT 298.435 0.695 298.715 2.31 ;
    RECT 296.59 0.895 296.86 2.195 ;
    RECT 295.115 0.695 295.395 2.31 ;
    RECT 293.27 0.895 293.54 2.195 ;
    RECT 291.795 0.695 292.075 2.31 ;
    RECT 289.95 0.895 290.22 2.195 ;
    RECT 288.475 0.695 288.755 2.31 ;
    RECT 286.63 0.895 286.9 2.195 ;
    RECT 285.155 0.695 285.435 2.31 ;
    RECT 283.31 0.895 283.58 2.195 ;
    RECT 281.835 0.695 282.115 2.31 ;
    RECT 279.99 0.895 280.26 2.195 ;
    RECT 278.515 0.695 278.795 2.31 ;
    RECT 276.67 0.895 276.94 2.195 ;
    RECT 275.195 0.695 275.475 2.31 ;
    RECT 273.35 0.895 273.62 2.195 ;
    RECT 271.875 0.695 272.155 2.31 ;
    RECT 270.03 0.895 270.3 2.195 ;
    RECT 268.555 0.695 268.835 2.31 ;
    RECT 266.71 0.895 266.98 2.195 ;
    RECT 265.235 0.695 265.515 2.31 ;
    RECT 263.39 0.895 263.66 2.195 ;
    RECT 261.915 0.695 262.195 2.31 ;
    RECT 260.07 0.895 260.34 2.195 ;
    RECT 258.595 0.695 258.875 2.31 ;
    RECT 256.75 0.895 257.02 2.195 ;
    RECT 255.275 0.695 255.555 2.31 ;
    RECT 253.43 0.895 253.7 2.195 ;
    RECT 251.955 0.695 252.235 2.31 ;
    RECT 250.11 0.895 250.38 2.195 ;
    RECT 248.635 0.695 248.915 2.31 ;
    RECT 246.79 0.895 247.06 2.195 ;
    RECT 245.315 0.695 245.595 2.31 ;
    RECT 243.47 0.895 243.74 2.195 ;
    RECT 241.995 0.695 242.275 2.31 ;
    RECT 240.15 0.895 240.42 2.195 ;
    RECT 238.675 0.695 238.955 2.31 ;
    RECT 236.83 0.895 237.1 2.195 ;
    RECT 235.355 0.695 235.635 2.31 ;
    RECT 372.95 0.895 373.22 2.195 ;
    RECT 371.475 0.695 371.755 2.31 ;
    RECT 203.63 0.895 203.9 2.195 ;
    RECT 202.155 0.695 202.435 2.31 ;
    RECT 233.51 0.895 233.78 2.195 ;
    RECT 232.035 0.695 232.315 2.31 ;
    RECT 230.19 0.895 230.46 2.195 ;
    RECT 228.715 0.695 228.995 2.31 ;
    RECT 226.87 0.895 227.14 2.195 ;
    RECT 225.395 0.695 225.675 2.31 ;
    RECT 223.55 0.895 223.82 2.195 ;
    RECT 222.075 0.695 222.355 2.31 ;
    RECT 220.23 0.895 220.5 2.195 ;
    RECT 218.755 0.695 219.035 2.31 ;
    RECT 216.91 0.895 217.18 2.195 ;
    RECT 215.435 0.695 215.715 2.31 ;
    RECT 213.59 0.895 213.86 2.195 ;
    RECT 212.115 0.695 212.395 2.31 ;
    RECT 210.27 0.895 210.54 2.195 ;
    RECT 208.795 0.695 209.075 2.31 ;
    RECT 206.95 0.895 207.22 2.195 ;
    RECT 205.475 0.695 205.755 2.31 ;
    RECT 173.565 0.695 173.645 11.6 ;
    RECT 174.315 0.695 174.45 11.6 ;
    RECT 174.74 0.695 175.09 11.6 ;
    RECT 175.675 0.695 175.725 11.6 ;
    RECT 175.725 0.695 175.985 11.635 ;
    RECT 175.985 0.695 176.325 11.6 ;
    RECT 176.595 0.695 176.855 11.6 ;
    RECT 177.125 0.695 177.24 11.6 ;
    RECT 178.51 0.695 178.665 11.6 ;
    RECT 179.125 0.695 179.75 11.6 ;
    RECT 180.22 0.695 180.37 11.6 ;
    RECT 180.72 0.695 180.79 11.6 ;
    RECT 180.79 0.695 181.04 11.635 ;
    RECT 181.04 0.695 181.115 11.6 ;
    RECT 182.155 0.695 182.435 11.6 ;
    RECT 182.905 0.695 183.055 11.6 ;
    RECT 183.055 0.695 183.325 11.635 ;
    RECT 183.325 0.695 183.605 11.6 ;
    RECT 183.895 0.695 184.1 11.6 ;
    RECT 184.1 0.695 184.35 11.635 ;
    RECT 184.35 0.695 184.405 11.6 ;
    RECT 185.075 0.695 186.625 11.6 ;
    RECT 186.975 0.695 187.325 11.6 ;
    RECT 187.805 0.695 189.52 11.6 ;
    RECT 190.32 0.695 190.64 11.6 ;
    RECT 190.92 0.695 190.99 11.6 ;
    RECT 190.99 0.695 191.26 11.635 ;
    RECT 191.26 0.695 191.38 11.6 ;
    RECT 192.18 0.695 192.72 11.6 ;
    RECT 192.72 0.695 193.19 1.62 ;
    RECT 193.19 0.695 193.565 11.6 ;
    RECT 193.565 0.695 193.835 11.635 ;
    RECT 193.835 0.695 193.905 11.6 ;
    RECT 194.195 0.695 194.4 11.6 ;
    RECT 195.4 0.695 195.56 11.6 ;
    RECT 195.91 0.695 196.08 11.6 ;
    RECT 197.15 0.695 197.37 3.185 ;
    RECT 197.15 5.375 197.37 11.6 ;
    RECT 197.37 0.695 197.435 11.6 ;
    RECT 197.705 0.695 198.045 11.6 ;
    RECT 198.255 0.695 198.605 11.6 ;
    RECT 198.605 0.695 198.815 11.635 ;
    RECT 198.815 0.695 198.885 11.6 ;
    RECT 199.625 0.695 199.815 11.6 ;
    RECT 200.165 0.695 200.305 11.6 ;
    RECT 200.975 0.695 201.055 11.6 ;
    RECT 97.68 0.895 97.95 2.195 ;
    RECT 99.145 0.695 99.425 2.31 ;
    RECT 94.36 0.895 94.63 2.195 ;
    RECT 95.825 0.695 96.105 2.31 ;
    RECT 91.04 0.895 91.31 2.195 ;
    RECT 92.505 0.695 92.785 2.31 ;
    RECT 87.72 0.895 87.99 2.195 ;
    RECT 89.185 0.695 89.465 2.31 ;
    RECT 84.4 0.895 84.67 2.195 ;
    RECT 85.865 0.695 86.145 2.31 ;
    RECT 81.08 0.895 81.35 2.195 ;
    RECT 82.545 0.695 82.825 2.31 ;
    RECT 77.76 0.895 78.03 2.195 ;
    RECT 79.225 0.695 79.505 2.31 ;
    RECT 74.44 0.895 74.71 2.195 ;
    RECT 75.905 0.695 76.185 2.31 ;
    RECT 71.12 0.895 71.39 2.195 ;
    RECT 72.585 0.695 72.865 2.31 ;
    RECT 67.8 0.895 68.07 2.195 ;
    RECT 69.265 0.695 69.545 2.31 ;
    RECT 64.48 0.895 64.75 2.195 ;
    RECT 65.945 0.695 66.225 2.31 ;
    RECT 61.16 0.895 61.43 2.195 ;
    RECT 62.625 0.695 62.905 2.31 ;
    RECT 57.84 0.895 58.11 2.195 ;
    RECT 59.305 0.695 59.585 2.31 ;
    RECT 54.52 0.895 54.79 2.195 ;
    RECT 55.985 0.695 56.265 2.31 ;
    RECT 51.2 0.895 51.47 2.195 ;
    RECT 52.665 0.695 52.945 2.31 ;
    RECT 47.88 0.895 48.15 2.195 ;
    RECT 49.345 0.695 49.625 2.31 ;
    RECT 44.56 0.895 44.83 2.195 ;
    RECT 46.025 0.695 46.305 2.31 ;
    RECT 41.24 0.895 41.51 2.195 ;
    RECT 42.705 0.695 42.985 2.31 ;
    RECT 37.92 0.895 38.19 2.195 ;
    RECT 39.385 0.695 39.665 2.31 ;
    RECT 34.6 0.895 34.87 2.195 ;
    RECT 36.065 0.695 36.345 2.31 ;
    RECT 170.72 0.895 170.99 2.195 ;
    RECT 172.185 0.695 172.465 2.31 ;
    RECT 1.4 0.895 1.67 2.195 ;
    RECT 2.865 0.695 3.145 2.31 ;
    RECT 31.28 0.895 31.55 2.195 ;
    RECT 32.745 0.695 33.025 2.31 ;
    RECT 27.96 0.895 28.23 2.195 ;
    RECT 29.425 0.695 29.705 2.31 ;
    RECT 24.64 0.895 24.91 2.195 ;
    RECT 26.105 0.695 26.385 2.31 ;
    RECT 21.32 0.895 21.59 2.195 ;
    RECT 22.785 0.695 23.065 2.31 ;
    RECT 18.0 0.895 18.27 2.195 ;
    RECT 19.465 0.695 19.745 2.31 ;
    RECT 14.68 0.895 14.95 2.195 ;
    RECT 16.145 0.695 16.425 2.31 ;
    RECT 11.36 0.895 11.63 2.195 ;
    RECT 12.825 0.695 13.105 2.31 ;
    RECT 8.04 0.895 8.31 2.195 ;
    RECT 9.505 0.695 9.785 2.31 ;
    RECT 4.72 0.895 4.99 2.195 ;
    RECT 6.185 0.695 6.465 2.31 ;
    RECT 167.4 0.895 167.67 2.195 ;
    RECT 168.865 0.695 169.145 2.31 ;
    RECT 164.08 0.895 164.35 2.195 ;
    RECT 165.545 0.695 165.825 2.31 ;
    RECT 160.76 0.895 161.03 2.195 ;
    RECT 162.225 0.695 162.505 2.31 ;
    RECT 157.44 0.895 157.71 2.195 ;
    RECT 158.905 0.695 159.185 2.31 ;
    RECT 154.12 0.895 154.39 2.195 ;
    RECT 155.585 0.695 155.865 2.31 ;
    RECT 150.8 0.895 151.07 2.195 ;
    RECT 152.265 0.695 152.545 2.31 ;
    RECT 147.48 0.895 147.75 2.195 ;
    RECT 148.945 0.695 149.225 2.31 ;
    RECT 144.16 0.895 144.43 2.195 ;
    RECT 145.625 0.695 145.905 2.31 ;
    RECT 140.84 0.895 141.11 2.195 ;
    RECT 142.305 0.695 142.585 2.31 ;
    RECT 137.52 0.895 137.79 2.195 ;
    RECT 138.985 0.695 139.265 2.31 ;
    RECT 134.2 0.895 134.47 2.195 ;
    RECT 135.665 0.695 135.945 2.31 ;
    RECT 130.88 0.895 131.15 2.195 ;
    RECT 132.345 0.695 132.625 2.31 ;
    RECT 127.56 0.895 127.83 2.195 ;
    RECT 129.025 0.695 129.305 2.31 ;
    RECT 124.24 0.895 124.51 2.195 ;
    RECT 125.705 0.695 125.985 2.31 ;
    RECT 120.92 0.895 121.19 2.195 ;
    RECT 122.385 0.695 122.665 2.31 ;
    RECT 117.6 0.895 117.87 2.195 ;
    RECT 119.065 0.695 119.345 2.31 ;
    RECT 114.28 0.895 114.55 2.195 ;
    RECT 115.745 0.695 116.025 2.31 ;
    RECT 110.96 0.895 111.23 2.195 ;
    RECT 112.425 0.695 112.705 2.31 ;
    RECT 107.64 0.895 107.91 2.195 ;
    RECT 109.105 0.695 109.385 2.31 ;
    RECT 104.32 0.895 104.59 2.195 ;
    RECT 105.785 0.695 106.065 2.31 ;
    RECT 101.0 0.895 101.27 2.195 ;
    RECT 102.465 0.695 102.745 2.31 ;
    RECT 64.68 4.77 64.75 9.56 ;
    RECT 65.945 2.31 66.225 8.3 ;
    RECT 61.36 4.77 61.43 9.56 ;
    RECT 62.625 2.31 62.905 8.3 ;
    RECT 58.04 4.77 58.11 9.56 ;
    RECT 59.305 2.31 59.585 8.3 ;
    RECT 54.72 4.77 54.79 9.56 ;
    RECT 55.985 2.31 56.265 8.3 ;
    RECT 51.4 4.77 51.47 9.56 ;
    RECT 52.665 2.31 52.945 8.3 ;
    RECT 48.08 4.77 48.15 9.56 ;
    RECT 49.345 2.31 49.625 8.3 ;
    RECT 44.76 4.77 44.83 9.56 ;
    RECT 46.025 2.31 46.305 8.3 ;
    RECT 41.44 4.77 41.51 9.56 ;
    RECT 42.705 2.31 42.985 8.3 ;
    RECT 38.12 4.77 38.19 9.56 ;
    RECT 39.385 2.31 39.665 8.3 ;
    RECT 34.8 4.77 34.87 9.56 ;
    RECT 36.065 2.31 36.345 8.3 ;
    RECT 31.48 4.77 31.55 9.56 ;
    RECT 32.745 2.31 33.025 8.3 ;
    RECT 28.16 4.77 28.23 9.56 ;
    RECT 29.425 2.31 29.705 8.3 ;
    RECT 24.84 4.77 24.91 9.56 ;
    RECT 26.105 2.31 26.385 8.3 ;
    RECT 21.52 4.77 21.59 9.56 ;
    RECT 22.785 2.31 23.065 8.3 ;
    RECT 18.2 4.77 18.27 9.56 ;
    RECT 19.465 2.31 19.745 8.3 ;
    RECT 14.88 4.77 14.95 9.56 ;
    RECT 16.145 2.31 16.425 8.3 ;
    RECT 11.56 4.77 11.63 9.56 ;
    RECT 12.825 2.31 13.105 8.3 ;
    RECT 8.24 4.77 8.31 9.56 ;
    RECT 9.505 2.31 9.785 8.3 ;
    RECT 4.92 4.77 4.99 9.56 ;
    RECT 6.185 2.31 6.465 8.3 ;
    RECT 170.92 4.77 170.99 9.56 ;
    RECT 172.185 2.31 172.465 8.3 ;
    RECT 1.6 4.77 1.67 9.56 ;
    RECT 2.865 2.31 3.145 8.3 ;
    RECT 167.6 4.77 167.67 9.56 ;
    RECT 168.865 2.31 169.145 8.3 ;
    RECT 164.28 4.77 164.35 9.56 ;
    RECT 165.545 2.31 165.825 8.3 ;
    RECT 160.96 4.77 161.03 9.56 ;
    RECT 162.225 2.31 162.505 8.3 ;
    RECT 157.64 4.77 157.71 9.56 ;
    RECT 158.905 2.31 159.185 8.3 ;
    RECT 154.32 4.77 154.39 9.56 ;
    RECT 155.585 2.31 155.865 8.3 ;
    RECT 151.0 4.77 151.07 9.56 ;
    RECT 152.265 2.31 152.545 8.3 ;
    RECT 147.68 4.77 147.75 9.56 ;
    RECT 148.945 2.31 149.225 8.3 ;
    RECT 144.36 4.77 144.43 9.56 ;
    RECT 145.625 2.31 145.905 8.3 ;
    RECT 141.04 4.77 141.11 9.56 ;
    RECT 142.305 2.31 142.585 8.3 ;
    RECT 137.72 4.77 137.79 9.56 ;
    RECT 138.985 2.31 139.265 8.3 ;
    RECT 134.4 4.77 134.47 9.56 ;
    RECT 135.665 2.31 135.945 8.3 ;
    RECT 131.08 4.77 131.15 9.56 ;
    RECT 132.345 2.31 132.625 8.3 ;
    RECT 127.76 4.77 127.83 9.56 ;
    RECT 129.025 2.31 129.305 8.3 ;
    RECT 124.44 4.77 124.51 9.56 ;
    RECT 125.705 2.31 125.985 8.3 ;
    RECT 121.12 4.77 121.19 9.56 ;
    RECT 122.385 2.31 122.665 8.3 ;
    RECT 117.8 4.77 117.87 9.56 ;
    RECT 119.065 2.31 119.345 8.3 ;
    RECT 114.48 4.77 114.55 9.56 ;
    RECT 115.745 2.31 116.025 8.3 ;
    RECT 111.16 4.77 111.23 9.56 ;
    RECT 112.425 2.31 112.705 8.3 ;
    RECT 107.84 4.77 107.91 9.56 ;
    RECT 109.105 2.31 109.385 8.3 ;
    RECT 104.52 4.77 104.59 9.56 ;
    RECT 105.785 2.31 106.065 8.3 ;
    RECT 101.2 4.77 101.27 9.56 ;
    RECT 102.465 2.31 102.745 8.3 ;
    RECT 97.88 4.77 97.95 9.56 ;
    RECT 99.145 2.31 99.425 8.3 ;
    RECT 94.56 4.77 94.63 9.56 ;
    RECT 95.825 2.31 96.105 8.3 ;
    RECT 91.24 4.77 91.31 9.56 ;
    RECT 92.505 2.31 92.785 8.3 ;
    RECT 87.92 4.77 87.99 9.56 ;
    RECT 89.185 2.31 89.465 8.3 ;
    RECT 84.6 4.77 84.67 9.56 ;
    RECT 85.865 2.31 86.145 8.3 ;
    RECT 81.28 4.77 81.35 9.56 ;
    RECT 82.545 2.31 82.825 8.3 ;
    RECT 77.96 4.77 78.03 9.56 ;
    RECT 79.225 2.31 79.505 8.3 ;
    RECT 74.64 4.77 74.71 9.56 ;
    RECT 75.905 2.31 76.185 8.3 ;
    RECT 71.32 4.77 71.39 9.56 ;
    RECT 72.585 2.31 72.865 8.3 ;
    RECT 68.0 4.77 68.07 9.56 ;
    RECT 69.265 2.31 69.545 8.3 ;
    RECT 173.565 60.67 173.645 61.255 ;
    RECT 174.315 60.67 174.45 61.255 ;
    RECT 174.74 61.06 175.09 61.255 ;
    RECT 175.675 60.67 177.24 61.255 ;
    RECT 178.51 60.67 178.665 61.255 ;
    RECT 179.125 60.67 179.75 61.255 ;
    RECT 180.22 60.67 180.37 61.255 ;
    RECT 180.72 60.67 181.115 61.255 ;
    RECT 181.405 60.67 181.725 61.255 ;
    RECT 182.155 60.67 182.435 61.255 ;
    RECT 182.905 60.67 183.605 61.255 ;
    RECT 183.895 60.67 184.405 61.255 ;
    RECT 185.075 60.67 186.625 61.255 ;
    RECT 186.975 60.67 187.325 61.255 ;
    RECT 187.805 60.67 189.52 61.255 ;
    RECT 190.32 60.67 190.64 61.255 ;
    RECT 190.92 60.67 191.38 61.255 ;
    RECT 192.18 60.67 192.72 61.255 ;
    RECT 193.19 60.67 193.905 61.255 ;
    RECT 194.195 60.67 194.4 61.255 ;
    RECT 195.4 60.67 195.56 61.255 ;
    RECT 195.91 60.67 196.08 61.255 ;
    RECT 197.15 60.67 198.885 61.255 ;
    RECT 199.625 60.67 199.815 61.255 ;
    RECT 200.165 60.67 200.305 61.255 ;
    RECT 200.975 60.67 201.055 61.255 ;
    #obstructions of filtered out pwrgnd shapes
    RECT 303.165 33.12 303.445 34.0 ;
    RECT 372.885 33.12 373.165 34.0 ;
    RECT 369.565 33.12 369.845 34.0 ;
    RECT 299.845 33.12 300.125 34.0 ;
    RECT 296.525 33.12 296.805 34.0 ;
    RECT 293.205 33.12 293.485 34.0 ;
    RECT 289.885 33.12 290.165 34.0 ;
    RECT 286.565 33.12 286.845 34.0 ;
    RECT 283.245 33.12 283.525 34.0 ;
    RECT 279.925 33.12 280.205 34.0 ;
    RECT 276.605 33.12 276.885 34.0 ;
    RECT 273.285 33.12 273.565 34.0 ;
    RECT 269.965 33.12 270.245 34.0 ;
    RECT 233.445 33.12 233.725 34.0 ;
    RECT 230.125 33.12 230.405 34.0 ;
    RECT 366.245 33.12 366.525 34.0 ;
    RECT 226.805 33.12 227.085 34.0 ;
    RECT 362.925 33.12 363.205 34.0 ;
    RECT 223.485 33.12 223.765 34.0 ;
    RECT 359.605 33.12 359.885 34.0 ;
    RECT 220.165 33.12 220.445 34.0 ;
    RECT 356.285 33.12 356.565 34.0 ;
    RECT 352.965 33.12 353.245 34.0 ;
    RECT 216.845 33.12 217.125 34.0 ;
    RECT 349.645 33.12 349.925 34.0 ;
    RECT 213.525 33.12 213.805 34.0 ;
    RECT 346.325 33.12 346.605 34.0 ;
    RECT 210.205 33.12 210.485 34.0 ;
    RECT 343.005 33.12 343.285 34.0 ;
    RECT 206.885 33.12 207.165 34.0 ;
    RECT 339.685 33.12 339.965 34.0 ;
    RECT 203.565 33.12 203.845 34.0 ;
    RECT 336.365 33.12 336.645 34.0 ;
    RECT 266.645 33.12 266.925 34.0 ;
    RECT 263.325 33.12 263.605 34.0 ;
    RECT 260.005 33.12 260.285 34.0 ;
    RECT 256.685 33.12 256.965 34.0 ;
    RECT 253.365 33.12 253.645 34.0 ;
    RECT 250.045 33.12 250.325 34.0 ;
    RECT 246.725 33.12 247.005 34.0 ;
    RECT 243.405 33.12 243.685 34.0 ;
    RECT 240.085 33.12 240.365 34.0 ;
    RECT 236.765 33.12 237.045 34.0 ;
    RECT 333.045 33.12 333.325 34.0 ;
    RECT 329.725 33.12 330.005 34.0 ;
    RECT 326.405 33.12 326.685 34.0 ;
    RECT 323.085 33.12 323.365 34.0 ;
    RECT 319.765 33.12 320.045 34.0 ;
    RECT 316.445 33.12 316.725 34.0 ;
    RECT 313.125 33.12 313.405 34.0 ;
    RECT 309.805 33.12 310.085 34.0 ;
    RECT 306.485 33.12 306.765 34.0 ;
    RECT 303.165 18.0 303.445 18.88 ;
    RECT 372.885 18.0 373.165 18.88 ;
    RECT 369.565 18.0 369.845 18.88 ;
    RECT 299.845 18.0 300.125 18.88 ;
    RECT 296.525 18.0 296.805 18.88 ;
    RECT 293.205 18.0 293.485 18.88 ;
    RECT 289.885 18.0 290.165 18.88 ;
    RECT 286.565 18.0 286.845 18.88 ;
    RECT 283.245 18.0 283.525 18.88 ;
    RECT 279.925 18.0 280.205 18.88 ;
    RECT 276.605 18.0 276.885 18.88 ;
    RECT 273.285 18.0 273.565 18.88 ;
    RECT 269.965 18.0 270.245 18.88 ;
    RECT 233.445 18.0 233.725 18.88 ;
    RECT 230.125 18.0 230.405 18.88 ;
    RECT 366.245 18.0 366.525 18.88 ;
    RECT 226.805 18.0 227.085 18.88 ;
    RECT 362.925 18.0 363.205 18.88 ;
    RECT 223.485 18.0 223.765 18.88 ;
    RECT 359.605 18.0 359.885 18.88 ;
    RECT 220.165 18.0 220.445 18.88 ;
    RECT 356.285 18.0 356.565 18.88 ;
    RECT 352.965 18.0 353.245 18.88 ;
    RECT 216.845 18.0 217.125 18.88 ;
    RECT 349.645 18.0 349.925 18.88 ;
    RECT 213.525 18.0 213.805 18.88 ;
    RECT 346.325 18.0 346.605 18.88 ;
    RECT 210.205 18.0 210.485 18.88 ;
    RECT 343.005 18.0 343.285 18.88 ;
    RECT 206.885 18.0 207.165 18.88 ;
    RECT 339.685 18.0 339.965 18.88 ;
    RECT 203.565 18.0 203.845 18.88 ;
    RECT 336.365 18.0 336.645 18.88 ;
    RECT 266.645 18.0 266.925 18.88 ;
    RECT 263.325 18.0 263.605 18.88 ;
    RECT 260.005 18.0 260.285 18.88 ;
    RECT 256.685 18.0 256.965 18.88 ;
    RECT 253.365 18.0 253.645 18.88 ;
    RECT 250.045 18.0 250.325 18.88 ;
    RECT 246.725 18.0 247.005 18.88 ;
    RECT 243.405 18.0 243.685 18.88 ;
    RECT 240.085 18.0 240.365 18.88 ;
    RECT 236.765 18.0 237.045 18.88 ;
    RECT 333.045 18.0 333.325 18.88 ;
    RECT 329.725 18.0 330.005 18.88 ;
    RECT 326.405 18.0 326.685 18.88 ;
    RECT 323.085 18.0 323.365 18.88 ;
    RECT 319.765 18.0 320.045 18.88 ;
    RECT 316.445 18.0 316.725 18.88 ;
    RECT 313.125 18.0 313.405 18.88 ;
    RECT 309.805 18.0 310.085 18.88 ;
    RECT 306.485 18.0 306.765 18.88 ;
    RECT 303.165 17.28 303.445 18.16 ;
    RECT 372.885 17.28 373.165 18.16 ;
    RECT 369.565 17.28 369.845 18.16 ;
    RECT 299.845 17.28 300.125 18.16 ;
    RECT 296.525 17.28 296.805 18.16 ;
    RECT 293.205 17.28 293.485 18.16 ;
    RECT 289.885 17.28 290.165 18.16 ;
    RECT 286.565 17.28 286.845 18.16 ;
    RECT 283.245 17.28 283.525 18.16 ;
    RECT 279.925 17.28 280.205 18.16 ;
    RECT 276.605 17.28 276.885 18.16 ;
    RECT 273.285 17.28 273.565 18.16 ;
    RECT 269.965 17.28 270.245 18.16 ;
    RECT 233.445 17.28 233.725 18.16 ;
    RECT 230.125 17.28 230.405 18.16 ;
    RECT 366.245 17.28 366.525 18.16 ;
    RECT 226.805 17.28 227.085 18.16 ;
    RECT 362.925 17.28 363.205 18.16 ;
    RECT 223.485 17.28 223.765 18.16 ;
    RECT 359.605 17.28 359.885 18.16 ;
    RECT 220.165 17.28 220.445 18.16 ;
    RECT 356.285 17.28 356.565 18.16 ;
    RECT 352.965 17.28 353.245 18.16 ;
    RECT 216.845 17.28 217.125 18.16 ;
    RECT 349.645 17.28 349.925 18.16 ;
    RECT 213.525 17.28 213.805 18.16 ;
    RECT 346.325 17.28 346.605 18.16 ;
    RECT 210.205 17.28 210.485 18.16 ;
    RECT 343.005 17.28 343.285 18.16 ;
    RECT 206.885 17.28 207.165 18.16 ;
    RECT 339.685 17.28 339.965 18.16 ;
    RECT 203.565 17.28 203.845 18.16 ;
    RECT 336.365 17.28 336.645 18.16 ;
    RECT 266.645 17.28 266.925 18.16 ;
    RECT 263.325 17.28 263.605 18.16 ;
    RECT 260.005 17.28 260.285 18.16 ;
    RECT 256.685 17.28 256.965 18.16 ;
    RECT 253.365 17.28 253.645 18.16 ;
    RECT 250.045 17.28 250.325 18.16 ;
    RECT 246.725 17.28 247.005 18.16 ;
    RECT 243.405 17.28 243.685 18.16 ;
    RECT 240.085 17.28 240.365 18.16 ;
    RECT 236.765 17.28 237.045 18.16 ;
    RECT 333.045 17.28 333.325 18.16 ;
    RECT 329.725 17.28 330.005 18.16 ;
    RECT 326.405 17.28 326.685 18.16 ;
    RECT 323.085 17.28 323.365 18.16 ;
    RECT 319.765 17.28 320.045 18.16 ;
    RECT 316.445 17.28 316.725 18.16 ;
    RECT 313.125 17.28 313.405 18.16 ;
    RECT 309.805 17.28 310.085 18.16 ;
    RECT 306.485 17.28 306.765 18.16 ;
    RECT 303.165 16.56 303.445 17.44 ;
    RECT 372.885 16.56 373.165 17.44 ;
    RECT 369.565 16.56 369.845 17.44 ;
    RECT 299.845 16.56 300.125 17.44 ;
    RECT 296.525 16.56 296.805 17.44 ;
    RECT 293.205 16.56 293.485 17.44 ;
    RECT 289.885 16.56 290.165 17.44 ;
    RECT 286.565 16.56 286.845 17.44 ;
    RECT 283.245 16.56 283.525 17.44 ;
    RECT 279.925 16.56 280.205 17.44 ;
    RECT 276.605 16.56 276.885 17.44 ;
    RECT 273.285 16.56 273.565 17.44 ;
    RECT 269.965 16.56 270.245 17.44 ;
    RECT 233.445 16.56 233.725 17.44 ;
    RECT 230.125 16.56 230.405 17.44 ;
    RECT 366.245 16.56 366.525 17.44 ;
    RECT 226.805 16.56 227.085 17.44 ;
    RECT 362.925 16.56 363.205 17.44 ;
    RECT 223.485 16.56 223.765 17.44 ;
    RECT 359.605 16.56 359.885 17.44 ;
    RECT 220.165 16.56 220.445 17.44 ;
    RECT 356.285 16.56 356.565 17.44 ;
    RECT 352.965 16.56 353.245 17.44 ;
    RECT 216.845 16.56 217.125 17.44 ;
    RECT 349.645 16.56 349.925 17.44 ;
    RECT 213.525 16.56 213.805 17.44 ;
    RECT 346.325 16.56 346.605 17.44 ;
    RECT 210.205 16.56 210.485 17.44 ;
    RECT 343.005 16.56 343.285 17.44 ;
    RECT 206.885 16.56 207.165 17.44 ;
    RECT 339.685 16.56 339.965 17.44 ;
    RECT 203.565 16.56 203.845 17.44 ;
    RECT 336.365 16.56 336.645 17.44 ;
    RECT 266.645 16.56 266.925 17.44 ;
    RECT 263.325 16.56 263.605 17.44 ;
    RECT 260.005 16.56 260.285 17.44 ;
    RECT 256.685 16.56 256.965 17.44 ;
    RECT 253.365 16.56 253.645 17.44 ;
    RECT 250.045 16.56 250.325 17.44 ;
    RECT 246.725 16.56 247.005 17.44 ;
    RECT 243.405 16.56 243.685 17.44 ;
    RECT 240.085 16.56 240.365 17.44 ;
    RECT 236.765 16.56 237.045 17.44 ;
    RECT 333.045 16.56 333.325 17.44 ;
    RECT 329.725 16.56 330.005 17.44 ;
    RECT 326.405 16.56 326.685 17.44 ;
    RECT 323.085 16.56 323.365 17.44 ;
    RECT 319.765 16.56 320.045 17.44 ;
    RECT 316.445 16.56 316.725 17.44 ;
    RECT 313.125 16.56 313.405 17.44 ;
    RECT 309.805 16.56 310.085 17.44 ;
    RECT 306.485 16.56 306.765 17.44 ;
    RECT 303.165 32.4 303.445 33.28 ;
    RECT 372.885 32.4 373.165 33.28 ;
    RECT 369.565 32.4 369.845 33.28 ;
    RECT 299.845 32.4 300.125 33.28 ;
    RECT 296.525 32.4 296.805 33.28 ;
    RECT 293.205 32.4 293.485 33.28 ;
    RECT 289.885 32.4 290.165 33.28 ;
    RECT 286.565 32.4 286.845 33.28 ;
    RECT 283.245 32.4 283.525 33.28 ;
    RECT 279.925 32.4 280.205 33.28 ;
    RECT 276.605 32.4 276.885 33.28 ;
    RECT 273.285 32.4 273.565 33.28 ;
    RECT 269.965 32.4 270.245 33.28 ;
    RECT 233.445 32.4 233.725 33.28 ;
    RECT 230.125 32.4 230.405 33.28 ;
    RECT 366.245 32.4 366.525 33.28 ;
    RECT 226.805 32.4 227.085 33.28 ;
    RECT 362.925 32.4 363.205 33.28 ;
    RECT 223.485 32.4 223.765 33.28 ;
    RECT 359.605 32.4 359.885 33.28 ;
    RECT 220.165 32.4 220.445 33.28 ;
    RECT 356.285 32.4 356.565 33.28 ;
    RECT 352.965 32.4 353.245 33.28 ;
    RECT 216.845 32.4 217.125 33.28 ;
    RECT 349.645 32.4 349.925 33.28 ;
    RECT 213.525 32.4 213.805 33.28 ;
    RECT 346.325 32.4 346.605 33.28 ;
    RECT 210.205 32.4 210.485 33.28 ;
    RECT 343.005 32.4 343.285 33.28 ;
    RECT 206.885 32.4 207.165 33.28 ;
    RECT 339.685 32.4 339.965 33.28 ;
    RECT 203.565 32.4 203.845 33.28 ;
    RECT 336.365 32.4 336.645 33.28 ;
    RECT 266.645 32.4 266.925 33.28 ;
    RECT 263.325 32.4 263.605 33.28 ;
    RECT 260.005 32.4 260.285 33.28 ;
    RECT 256.685 32.4 256.965 33.28 ;
    RECT 253.365 32.4 253.645 33.28 ;
    RECT 250.045 32.4 250.325 33.28 ;
    RECT 246.725 32.4 247.005 33.28 ;
    RECT 243.405 32.4 243.685 33.28 ;
    RECT 240.085 32.4 240.365 33.28 ;
    RECT 236.765 32.4 237.045 33.28 ;
    RECT 333.045 32.4 333.325 33.28 ;
    RECT 329.725 32.4 330.005 33.28 ;
    RECT 326.405 32.4 326.685 33.28 ;
    RECT 323.085 32.4 323.365 33.28 ;
    RECT 319.765 32.4 320.045 33.28 ;
    RECT 316.445 32.4 316.725 33.28 ;
    RECT 313.125 32.4 313.405 33.28 ;
    RECT 309.805 32.4 310.085 33.28 ;
    RECT 306.485 32.4 306.765 33.28 ;
    RECT 303.165 15.84 303.445 16.72 ;
    RECT 372.885 15.84 373.165 16.72 ;
    RECT 369.565 15.84 369.845 16.72 ;
    RECT 299.845 15.84 300.125 16.72 ;
    RECT 296.525 15.84 296.805 16.72 ;
    RECT 293.205 15.84 293.485 16.72 ;
    RECT 289.885 15.84 290.165 16.72 ;
    RECT 286.565 15.84 286.845 16.72 ;
    RECT 283.245 15.84 283.525 16.72 ;
    RECT 279.925 15.84 280.205 16.72 ;
    RECT 276.605 15.84 276.885 16.72 ;
    RECT 273.285 15.84 273.565 16.72 ;
    RECT 269.965 15.84 270.245 16.72 ;
    RECT 233.445 15.84 233.725 16.72 ;
    RECT 230.125 15.84 230.405 16.72 ;
    RECT 366.245 15.84 366.525 16.72 ;
    RECT 226.805 15.84 227.085 16.72 ;
    RECT 362.925 15.84 363.205 16.72 ;
    RECT 223.485 15.84 223.765 16.72 ;
    RECT 359.605 15.84 359.885 16.72 ;
    RECT 220.165 15.84 220.445 16.72 ;
    RECT 356.285 15.84 356.565 16.72 ;
    RECT 352.965 15.84 353.245 16.72 ;
    RECT 216.845 15.84 217.125 16.72 ;
    RECT 349.645 15.84 349.925 16.72 ;
    RECT 213.525 15.84 213.805 16.72 ;
    RECT 346.325 15.84 346.605 16.72 ;
    RECT 210.205 15.84 210.485 16.72 ;
    RECT 343.005 15.84 343.285 16.72 ;
    RECT 206.885 15.84 207.165 16.72 ;
    RECT 339.685 15.84 339.965 16.72 ;
    RECT 203.565 15.84 203.845 16.72 ;
    RECT 336.365 15.84 336.645 16.72 ;
    RECT 266.645 15.84 266.925 16.72 ;
    RECT 263.325 15.84 263.605 16.72 ;
    RECT 260.005 15.84 260.285 16.72 ;
    RECT 256.685 15.84 256.965 16.72 ;
    RECT 253.365 15.84 253.645 16.72 ;
    RECT 250.045 15.84 250.325 16.72 ;
    RECT 246.725 15.84 247.005 16.72 ;
    RECT 243.405 15.84 243.685 16.72 ;
    RECT 240.085 15.84 240.365 16.72 ;
    RECT 236.765 15.84 237.045 16.72 ;
    RECT 333.045 15.84 333.325 16.72 ;
    RECT 329.725 15.84 330.005 16.72 ;
    RECT 326.405 15.84 326.685 16.72 ;
    RECT 323.085 15.84 323.365 16.72 ;
    RECT 319.765 15.84 320.045 16.72 ;
    RECT 316.445 15.84 316.725 16.72 ;
    RECT 313.125 15.84 313.405 16.72 ;
    RECT 309.805 15.84 310.085 16.72 ;
    RECT 306.485 15.84 306.765 16.72 ;
    RECT 303.165 31.68 303.445 32.56 ;
    RECT 372.885 31.68 373.165 32.56 ;
    RECT 369.565 31.68 369.845 32.56 ;
    RECT 299.845 31.68 300.125 32.56 ;
    RECT 296.525 31.68 296.805 32.56 ;
    RECT 293.205 31.68 293.485 32.56 ;
    RECT 289.885 31.68 290.165 32.56 ;
    RECT 286.565 31.68 286.845 32.56 ;
    RECT 283.245 31.68 283.525 32.56 ;
    RECT 279.925 31.68 280.205 32.56 ;
    RECT 276.605 31.68 276.885 32.56 ;
    RECT 273.285 31.68 273.565 32.56 ;
    RECT 269.965 31.68 270.245 32.56 ;
    RECT 233.445 31.68 233.725 32.56 ;
    RECT 230.125 31.68 230.405 32.56 ;
    RECT 366.245 31.68 366.525 32.56 ;
    RECT 226.805 31.68 227.085 32.56 ;
    RECT 362.925 31.68 363.205 32.56 ;
    RECT 223.485 31.68 223.765 32.56 ;
    RECT 359.605 31.68 359.885 32.56 ;
    RECT 220.165 31.68 220.445 32.56 ;
    RECT 356.285 31.68 356.565 32.56 ;
    RECT 352.965 31.68 353.245 32.56 ;
    RECT 216.845 31.68 217.125 32.56 ;
    RECT 349.645 31.68 349.925 32.56 ;
    RECT 213.525 31.68 213.805 32.56 ;
    RECT 346.325 31.68 346.605 32.56 ;
    RECT 210.205 31.68 210.485 32.56 ;
    RECT 343.005 31.68 343.285 32.56 ;
    RECT 206.885 31.68 207.165 32.56 ;
    RECT 339.685 31.68 339.965 32.56 ;
    RECT 203.565 31.68 203.845 32.56 ;
    RECT 336.365 31.68 336.645 32.56 ;
    RECT 266.645 31.68 266.925 32.56 ;
    RECT 263.325 31.68 263.605 32.56 ;
    RECT 260.005 31.68 260.285 32.56 ;
    RECT 256.685 31.68 256.965 32.56 ;
    RECT 253.365 31.68 253.645 32.56 ;
    RECT 250.045 31.68 250.325 32.56 ;
    RECT 246.725 31.68 247.005 32.56 ;
    RECT 243.405 31.68 243.685 32.56 ;
    RECT 240.085 31.68 240.365 32.56 ;
    RECT 236.765 31.68 237.045 32.56 ;
    RECT 333.045 31.68 333.325 32.56 ;
    RECT 329.725 31.68 330.005 32.56 ;
    RECT 326.405 31.68 326.685 32.56 ;
    RECT 323.085 31.68 323.365 32.56 ;
    RECT 319.765 31.68 320.045 32.56 ;
    RECT 316.445 31.68 316.725 32.56 ;
    RECT 313.125 31.68 313.405 32.56 ;
    RECT 309.805 31.68 310.085 32.56 ;
    RECT 306.485 31.68 306.765 32.56 ;
    RECT 303.165 15.12 303.445 16.0 ;
    RECT 372.885 15.12 373.165 16.0 ;
    RECT 369.565 15.12 369.845 16.0 ;
    RECT 299.845 15.12 300.125 16.0 ;
    RECT 296.525 15.12 296.805 16.0 ;
    RECT 293.205 15.12 293.485 16.0 ;
    RECT 289.885 15.12 290.165 16.0 ;
    RECT 286.565 15.12 286.845 16.0 ;
    RECT 283.245 15.12 283.525 16.0 ;
    RECT 279.925 15.12 280.205 16.0 ;
    RECT 276.605 15.12 276.885 16.0 ;
    RECT 273.285 15.12 273.565 16.0 ;
    RECT 269.965 15.12 270.245 16.0 ;
    RECT 233.445 15.12 233.725 16.0 ;
    RECT 230.125 15.12 230.405 16.0 ;
    RECT 366.245 15.12 366.525 16.0 ;
    RECT 226.805 15.12 227.085 16.0 ;
    RECT 362.925 15.12 363.205 16.0 ;
    RECT 223.485 15.12 223.765 16.0 ;
    RECT 359.605 15.12 359.885 16.0 ;
    RECT 220.165 15.12 220.445 16.0 ;
    RECT 356.285 15.12 356.565 16.0 ;
    RECT 352.965 15.12 353.245 16.0 ;
    RECT 216.845 15.12 217.125 16.0 ;
    RECT 349.645 15.12 349.925 16.0 ;
    RECT 213.525 15.12 213.805 16.0 ;
    RECT 346.325 15.12 346.605 16.0 ;
    RECT 210.205 15.12 210.485 16.0 ;
    RECT 343.005 15.12 343.285 16.0 ;
    RECT 206.885 15.12 207.165 16.0 ;
    RECT 339.685 15.12 339.965 16.0 ;
    RECT 203.565 15.12 203.845 16.0 ;
    RECT 336.365 15.12 336.645 16.0 ;
    RECT 266.645 15.12 266.925 16.0 ;
    RECT 263.325 15.12 263.605 16.0 ;
    RECT 260.005 15.12 260.285 16.0 ;
    RECT 256.685 15.12 256.965 16.0 ;
    RECT 253.365 15.12 253.645 16.0 ;
    RECT 250.045 15.12 250.325 16.0 ;
    RECT 246.725 15.12 247.005 16.0 ;
    RECT 243.405 15.12 243.685 16.0 ;
    RECT 240.085 15.12 240.365 16.0 ;
    RECT 236.765 15.12 237.045 16.0 ;
    RECT 333.045 15.12 333.325 16.0 ;
    RECT 329.725 15.12 330.005 16.0 ;
    RECT 326.405 15.12 326.685 16.0 ;
    RECT 323.085 15.12 323.365 16.0 ;
    RECT 319.765 15.12 320.045 16.0 ;
    RECT 316.445 15.12 316.725 16.0 ;
    RECT 313.125 15.12 313.405 16.0 ;
    RECT 309.805 15.12 310.085 16.0 ;
    RECT 306.485 15.12 306.765 16.0 ;
    RECT 303.165 30.96 303.445 31.84 ;
    RECT 372.885 30.96 373.165 31.84 ;
    RECT 369.565 30.96 369.845 31.84 ;
    RECT 299.845 30.96 300.125 31.84 ;
    RECT 296.525 30.96 296.805 31.84 ;
    RECT 293.205 30.96 293.485 31.84 ;
    RECT 289.885 30.96 290.165 31.84 ;
    RECT 286.565 30.96 286.845 31.84 ;
    RECT 283.245 30.96 283.525 31.84 ;
    RECT 279.925 30.96 280.205 31.84 ;
    RECT 276.605 30.96 276.885 31.84 ;
    RECT 273.285 30.96 273.565 31.84 ;
    RECT 269.965 30.96 270.245 31.84 ;
    RECT 233.445 30.96 233.725 31.84 ;
    RECT 230.125 30.96 230.405 31.84 ;
    RECT 366.245 30.96 366.525 31.84 ;
    RECT 226.805 30.96 227.085 31.84 ;
    RECT 362.925 30.96 363.205 31.84 ;
    RECT 223.485 30.96 223.765 31.84 ;
    RECT 359.605 30.96 359.885 31.84 ;
    RECT 220.165 30.96 220.445 31.84 ;
    RECT 356.285 30.96 356.565 31.84 ;
    RECT 352.965 30.96 353.245 31.84 ;
    RECT 216.845 30.96 217.125 31.84 ;
    RECT 349.645 30.96 349.925 31.84 ;
    RECT 213.525 30.96 213.805 31.84 ;
    RECT 346.325 30.96 346.605 31.84 ;
    RECT 210.205 30.96 210.485 31.84 ;
    RECT 343.005 30.96 343.285 31.84 ;
    RECT 206.885 30.96 207.165 31.84 ;
    RECT 339.685 30.96 339.965 31.84 ;
    RECT 203.565 30.96 203.845 31.84 ;
    RECT 336.365 30.96 336.645 31.84 ;
    RECT 266.645 30.96 266.925 31.84 ;
    RECT 263.325 30.96 263.605 31.84 ;
    RECT 260.005 30.96 260.285 31.84 ;
    RECT 256.685 30.96 256.965 31.84 ;
    RECT 253.365 30.96 253.645 31.84 ;
    RECT 250.045 30.96 250.325 31.84 ;
    RECT 246.725 30.96 247.005 31.84 ;
    RECT 243.405 30.96 243.685 31.84 ;
    RECT 240.085 30.96 240.365 31.84 ;
    RECT 236.765 30.96 237.045 31.84 ;
    RECT 333.045 30.96 333.325 31.84 ;
    RECT 329.725 30.96 330.005 31.84 ;
    RECT 326.405 30.96 326.685 31.84 ;
    RECT 323.085 30.96 323.365 31.84 ;
    RECT 319.765 30.96 320.045 31.84 ;
    RECT 316.445 30.96 316.725 31.84 ;
    RECT 313.125 30.96 313.405 31.84 ;
    RECT 309.805 30.96 310.085 31.84 ;
    RECT 306.485 30.96 306.765 31.84 ;
    RECT 303.165 14.4 303.445 15.28 ;
    RECT 372.885 14.4 373.165 15.28 ;
    RECT 369.565 14.4 369.845 15.28 ;
    RECT 299.845 14.4 300.125 15.28 ;
    RECT 296.525 14.4 296.805 15.28 ;
    RECT 293.205 14.4 293.485 15.28 ;
    RECT 289.885 14.4 290.165 15.28 ;
    RECT 286.565 14.4 286.845 15.28 ;
    RECT 283.245 14.4 283.525 15.28 ;
    RECT 279.925 14.4 280.205 15.28 ;
    RECT 276.605 14.4 276.885 15.28 ;
    RECT 273.285 14.4 273.565 15.28 ;
    RECT 269.965 14.4 270.245 15.28 ;
    RECT 233.445 14.4 233.725 15.28 ;
    RECT 230.125 14.4 230.405 15.28 ;
    RECT 366.245 14.4 366.525 15.28 ;
    RECT 226.805 14.4 227.085 15.28 ;
    RECT 362.925 14.4 363.205 15.28 ;
    RECT 223.485 14.4 223.765 15.28 ;
    RECT 359.605 14.4 359.885 15.28 ;
    RECT 220.165 14.4 220.445 15.28 ;
    RECT 356.285 14.4 356.565 15.28 ;
    RECT 352.965 14.4 353.245 15.28 ;
    RECT 216.845 14.4 217.125 15.28 ;
    RECT 349.645 14.4 349.925 15.28 ;
    RECT 213.525 14.4 213.805 15.28 ;
    RECT 346.325 14.4 346.605 15.28 ;
    RECT 210.205 14.4 210.485 15.28 ;
    RECT 343.005 14.4 343.285 15.28 ;
    RECT 206.885 14.4 207.165 15.28 ;
    RECT 339.685 14.4 339.965 15.28 ;
    RECT 203.565 14.4 203.845 15.28 ;
    RECT 336.365 14.4 336.645 15.28 ;
    RECT 266.645 14.4 266.925 15.28 ;
    RECT 263.325 14.4 263.605 15.28 ;
    RECT 260.005 14.4 260.285 15.28 ;
    RECT 256.685 14.4 256.965 15.28 ;
    RECT 253.365 14.4 253.645 15.28 ;
    RECT 250.045 14.4 250.325 15.28 ;
    RECT 246.725 14.4 247.005 15.28 ;
    RECT 243.405 14.4 243.685 15.28 ;
    RECT 240.085 14.4 240.365 15.28 ;
    RECT 236.765 14.4 237.045 15.28 ;
    RECT 333.045 14.4 333.325 15.28 ;
    RECT 329.725 14.4 330.005 15.28 ;
    RECT 326.405 14.4 326.685 15.28 ;
    RECT 323.085 14.4 323.365 15.28 ;
    RECT 319.765 14.4 320.045 15.28 ;
    RECT 316.445 14.4 316.725 15.28 ;
    RECT 313.125 14.4 313.405 15.28 ;
    RECT 309.805 14.4 310.085 15.28 ;
    RECT 306.485 14.4 306.765 15.28 ;
    RECT 303.165 30.24 303.445 31.12 ;
    RECT 372.885 30.24 373.165 31.12 ;
    RECT 369.565 30.24 369.845 31.12 ;
    RECT 299.845 30.24 300.125 31.12 ;
    RECT 296.525 30.24 296.805 31.12 ;
    RECT 293.205 30.24 293.485 31.12 ;
    RECT 289.885 30.24 290.165 31.12 ;
    RECT 286.565 30.24 286.845 31.12 ;
    RECT 283.245 30.24 283.525 31.12 ;
    RECT 279.925 30.24 280.205 31.12 ;
    RECT 276.605 30.24 276.885 31.12 ;
    RECT 273.285 30.24 273.565 31.12 ;
    RECT 269.965 30.24 270.245 31.12 ;
    RECT 233.445 30.24 233.725 31.12 ;
    RECT 230.125 30.24 230.405 31.12 ;
    RECT 366.245 30.24 366.525 31.12 ;
    RECT 226.805 30.24 227.085 31.12 ;
    RECT 362.925 30.24 363.205 31.12 ;
    RECT 223.485 30.24 223.765 31.12 ;
    RECT 359.605 30.24 359.885 31.12 ;
    RECT 220.165 30.24 220.445 31.12 ;
    RECT 356.285 30.24 356.565 31.12 ;
    RECT 352.965 30.24 353.245 31.12 ;
    RECT 216.845 30.24 217.125 31.12 ;
    RECT 349.645 30.24 349.925 31.12 ;
    RECT 213.525 30.24 213.805 31.12 ;
    RECT 346.325 30.24 346.605 31.12 ;
    RECT 210.205 30.24 210.485 31.12 ;
    RECT 343.005 30.24 343.285 31.12 ;
    RECT 206.885 30.24 207.165 31.12 ;
    RECT 339.685 30.24 339.965 31.12 ;
    RECT 203.565 30.24 203.845 31.12 ;
    RECT 336.365 30.24 336.645 31.12 ;
    RECT 266.645 30.24 266.925 31.12 ;
    RECT 263.325 30.24 263.605 31.12 ;
    RECT 260.005 30.24 260.285 31.12 ;
    RECT 256.685 30.24 256.965 31.12 ;
    RECT 253.365 30.24 253.645 31.12 ;
    RECT 250.045 30.24 250.325 31.12 ;
    RECT 246.725 30.24 247.005 31.12 ;
    RECT 243.405 30.24 243.685 31.12 ;
    RECT 240.085 30.24 240.365 31.12 ;
    RECT 236.765 30.24 237.045 31.12 ;
    RECT 333.045 30.24 333.325 31.12 ;
    RECT 329.725 30.24 330.005 31.12 ;
    RECT 326.405 30.24 326.685 31.12 ;
    RECT 323.085 30.24 323.365 31.12 ;
    RECT 319.765 30.24 320.045 31.12 ;
    RECT 316.445 30.24 316.725 31.12 ;
    RECT 313.125 30.24 313.405 31.12 ;
    RECT 309.805 30.24 310.085 31.12 ;
    RECT 306.485 30.24 306.765 31.12 ;
    RECT 303.165 13.68 303.445 14.56 ;
    RECT 372.885 13.68 373.165 14.56 ;
    RECT 369.565 13.68 369.845 14.56 ;
    RECT 299.845 13.68 300.125 14.56 ;
    RECT 296.525 13.68 296.805 14.56 ;
    RECT 293.205 13.68 293.485 14.56 ;
    RECT 289.885 13.68 290.165 14.56 ;
    RECT 286.565 13.68 286.845 14.56 ;
    RECT 283.245 13.68 283.525 14.56 ;
    RECT 279.925 13.68 280.205 14.56 ;
    RECT 276.605 13.68 276.885 14.56 ;
    RECT 273.285 13.68 273.565 14.56 ;
    RECT 269.965 13.68 270.245 14.56 ;
    RECT 233.445 13.68 233.725 14.56 ;
    RECT 230.125 13.68 230.405 14.56 ;
    RECT 366.245 13.68 366.525 14.56 ;
    RECT 226.805 13.68 227.085 14.56 ;
    RECT 362.925 13.68 363.205 14.56 ;
    RECT 223.485 13.68 223.765 14.56 ;
    RECT 359.605 13.68 359.885 14.56 ;
    RECT 220.165 13.68 220.445 14.56 ;
    RECT 356.285 13.68 356.565 14.56 ;
    RECT 352.965 13.68 353.245 14.56 ;
    RECT 216.845 13.68 217.125 14.56 ;
    RECT 349.645 13.68 349.925 14.56 ;
    RECT 213.525 13.68 213.805 14.56 ;
    RECT 346.325 13.68 346.605 14.56 ;
    RECT 210.205 13.68 210.485 14.56 ;
    RECT 343.005 13.68 343.285 14.56 ;
    RECT 206.885 13.68 207.165 14.56 ;
    RECT 339.685 13.68 339.965 14.56 ;
    RECT 203.565 13.68 203.845 14.56 ;
    RECT 336.365 13.68 336.645 14.56 ;
    RECT 266.645 13.68 266.925 14.56 ;
    RECT 263.325 13.68 263.605 14.56 ;
    RECT 260.005 13.68 260.285 14.56 ;
    RECT 256.685 13.68 256.965 14.56 ;
    RECT 253.365 13.68 253.645 14.56 ;
    RECT 250.045 13.68 250.325 14.56 ;
    RECT 246.725 13.68 247.005 14.56 ;
    RECT 243.405 13.68 243.685 14.56 ;
    RECT 240.085 13.68 240.365 14.56 ;
    RECT 236.765 13.68 237.045 14.56 ;
    RECT 333.045 13.68 333.325 14.56 ;
    RECT 329.725 13.68 330.005 14.56 ;
    RECT 326.405 13.68 326.685 14.56 ;
    RECT 323.085 13.68 323.365 14.56 ;
    RECT 319.765 13.68 320.045 14.56 ;
    RECT 316.445 13.68 316.725 14.56 ;
    RECT 313.125 13.68 313.405 14.56 ;
    RECT 309.805 13.68 310.085 14.56 ;
    RECT 306.485 13.68 306.765 14.56 ;
    RECT 303.165 29.52 303.445 30.4 ;
    RECT 372.885 29.52 373.165 30.4 ;
    RECT 369.565 29.52 369.845 30.4 ;
    RECT 299.845 29.52 300.125 30.4 ;
    RECT 296.525 29.52 296.805 30.4 ;
    RECT 293.205 29.52 293.485 30.4 ;
    RECT 289.885 29.52 290.165 30.4 ;
    RECT 286.565 29.52 286.845 30.4 ;
    RECT 283.245 29.52 283.525 30.4 ;
    RECT 279.925 29.52 280.205 30.4 ;
    RECT 276.605 29.52 276.885 30.4 ;
    RECT 273.285 29.52 273.565 30.4 ;
    RECT 269.965 29.52 270.245 30.4 ;
    RECT 233.445 29.52 233.725 30.4 ;
    RECT 230.125 29.52 230.405 30.4 ;
    RECT 366.245 29.52 366.525 30.4 ;
    RECT 226.805 29.52 227.085 30.4 ;
    RECT 362.925 29.52 363.205 30.4 ;
    RECT 223.485 29.52 223.765 30.4 ;
    RECT 359.605 29.52 359.885 30.4 ;
    RECT 220.165 29.52 220.445 30.4 ;
    RECT 356.285 29.52 356.565 30.4 ;
    RECT 352.965 29.52 353.245 30.4 ;
    RECT 216.845 29.52 217.125 30.4 ;
    RECT 349.645 29.52 349.925 30.4 ;
    RECT 213.525 29.52 213.805 30.4 ;
    RECT 346.325 29.52 346.605 30.4 ;
    RECT 210.205 29.52 210.485 30.4 ;
    RECT 343.005 29.52 343.285 30.4 ;
    RECT 206.885 29.52 207.165 30.4 ;
    RECT 339.685 29.52 339.965 30.4 ;
    RECT 203.565 29.52 203.845 30.4 ;
    RECT 336.365 29.52 336.645 30.4 ;
    RECT 266.645 29.52 266.925 30.4 ;
    RECT 263.325 29.52 263.605 30.4 ;
    RECT 260.005 29.52 260.285 30.4 ;
    RECT 256.685 29.52 256.965 30.4 ;
    RECT 253.365 29.52 253.645 30.4 ;
    RECT 250.045 29.52 250.325 30.4 ;
    RECT 246.725 29.52 247.005 30.4 ;
    RECT 243.405 29.52 243.685 30.4 ;
    RECT 240.085 29.52 240.365 30.4 ;
    RECT 236.765 29.52 237.045 30.4 ;
    RECT 333.045 29.52 333.325 30.4 ;
    RECT 329.725 29.52 330.005 30.4 ;
    RECT 326.405 29.52 326.685 30.4 ;
    RECT 323.085 29.52 323.365 30.4 ;
    RECT 319.765 29.52 320.045 30.4 ;
    RECT 316.445 29.52 316.725 30.4 ;
    RECT 313.125 29.52 313.405 30.4 ;
    RECT 309.805 29.52 310.085 30.4 ;
    RECT 306.485 29.52 306.765 30.4 ;
    RECT 303.165 12.96 303.445 13.84 ;
    RECT 372.885 12.96 373.165 13.84 ;
    RECT 369.565 12.96 369.845 13.84 ;
    RECT 299.845 12.96 300.125 13.84 ;
    RECT 296.525 12.96 296.805 13.84 ;
    RECT 293.205 12.96 293.485 13.84 ;
    RECT 289.885 12.96 290.165 13.84 ;
    RECT 286.565 12.96 286.845 13.84 ;
    RECT 283.245 12.96 283.525 13.84 ;
    RECT 279.925 12.96 280.205 13.84 ;
    RECT 276.605 12.96 276.885 13.84 ;
    RECT 273.285 12.96 273.565 13.84 ;
    RECT 269.965 12.96 270.245 13.84 ;
    RECT 233.445 12.96 233.725 13.84 ;
    RECT 230.125 12.96 230.405 13.84 ;
    RECT 366.245 12.96 366.525 13.84 ;
    RECT 226.805 12.96 227.085 13.84 ;
    RECT 362.925 12.96 363.205 13.84 ;
    RECT 223.485 12.96 223.765 13.84 ;
    RECT 359.605 12.96 359.885 13.84 ;
    RECT 220.165 12.96 220.445 13.84 ;
    RECT 356.285 12.96 356.565 13.84 ;
    RECT 352.965 12.96 353.245 13.84 ;
    RECT 216.845 12.96 217.125 13.84 ;
    RECT 349.645 12.96 349.925 13.84 ;
    RECT 213.525 12.96 213.805 13.84 ;
    RECT 346.325 12.96 346.605 13.84 ;
    RECT 210.205 12.96 210.485 13.84 ;
    RECT 343.005 12.96 343.285 13.84 ;
    RECT 206.885 12.96 207.165 13.84 ;
    RECT 339.685 12.96 339.965 13.84 ;
    RECT 203.565 12.96 203.845 13.84 ;
    RECT 336.365 12.96 336.645 13.84 ;
    RECT 266.645 12.96 266.925 13.84 ;
    RECT 263.325 12.96 263.605 13.84 ;
    RECT 260.005 12.96 260.285 13.84 ;
    RECT 256.685 12.96 256.965 13.84 ;
    RECT 253.365 12.96 253.645 13.84 ;
    RECT 250.045 12.96 250.325 13.84 ;
    RECT 246.725 12.96 247.005 13.84 ;
    RECT 243.405 12.96 243.685 13.84 ;
    RECT 240.085 12.96 240.365 13.84 ;
    RECT 236.765 12.96 237.045 13.84 ;
    RECT 333.045 12.96 333.325 13.84 ;
    RECT 329.725 12.96 330.005 13.84 ;
    RECT 326.405 12.96 326.685 13.84 ;
    RECT 323.085 12.96 323.365 13.84 ;
    RECT 319.765 12.96 320.045 13.84 ;
    RECT 316.445 12.96 316.725 13.84 ;
    RECT 313.125 12.96 313.405 13.84 ;
    RECT 309.805 12.96 310.085 13.84 ;
    RECT 306.485 12.96 306.765 13.84 ;
    RECT 303.165 28.8 303.445 29.68 ;
    RECT 372.885 28.8 373.165 29.68 ;
    RECT 369.565 28.8 369.845 29.68 ;
    RECT 299.845 28.8 300.125 29.68 ;
    RECT 296.525 28.8 296.805 29.68 ;
    RECT 293.205 28.8 293.485 29.68 ;
    RECT 289.885 28.8 290.165 29.68 ;
    RECT 286.565 28.8 286.845 29.68 ;
    RECT 283.245 28.8 283.525 29.68 ;
    RECT 279.925 28.8 280.205 29.68 ;
    RECT 276.605 28.8 276.885 29.68 ;
    RECT 273.285 28.8 273.565 29.68 ;
    RECT 269.965 28.8 270.245 29.68 ;
    RECT 233.445 28.8 233.725 29.68 ;
    RECT 230.125 28.8 230.405 29.68 ;
    RECT 366.245 28.8 366.525 29.68 ;
    RECT 226.805 28.8 227.085 29.68 ;
    RECT 362.925 28.8 363.205 29.68 ;
    RECT 223.485 28.8 223.765 29.68 ;
    RECT 359.605 28.8 359.885 29.68 ;
    RECT 220.165 28.8 220.445 29.68 ;
    RECT 356.285 28.8 356.565 29.68 ;
    RECT 352.965 28.8 353.245 29.68 ;
    RECT 216.845 28.8 217.125 29.68 ;
    RECT 349.645 28.8 349.925 29.68 ;
    RECT 213.525 28.8 213.805 29.68 ;
    RECT 346.325 28.8 346.605 29.68 ;
    RECT 210.205 28.8 210.485 29.68 ;
    RECT 343.005 28.8 343.285 29.68 ;
    RECT 206.885 28.8 207.165 29.68 ;
    RECT 339.685 28.8 339.965 29.68 ;
    RECT 203.565 28.8 203.845 29.68 ;
    RECT 336.365 28.8 336.645 29.68 ;
    RECT 266.645 28.8 266.925 29.68 ;
    RECT 263.325 28.8 263.605 29.68 ;
    RECT 260.005 28.8 260.285 29.68 ;
    RECT 256.685 28.8 256.965 29.68 ;
    RECT 253.365 28.8 253.645 29.68 ;
    RECT 250.045 28.8 250.325 29.68 ;
    RECT 246.725 28.8 247.005 29.68 ;
    RECT 243.405 28.8 243.685 29.68 ;
    RECT 240.085 28.8 240.365 29.68 ;
    RECT 236.765 28.8 237.045 29.68 ;
    RECT 333.045 28.8 333.325 29.68 ;
    RECT 329.725 28.8 330.005 29.68 ;
    RECT 326.405 28.8 326.685 29.68 ;
    RECT 323.085 28.8 323.365 29.68 ;
    RECT 319.765 28.8 320.045 29.68 ;
    RECT 316.445 28.8 316.725 29.68 ;
    RECT 313.125 28.8 313.405 29.68 ;
    RECT 309.805 28.8 310.085 29.68 ;
    RECT 306.485 28.8 306.765 29.68 ;
    RECT 303.165 12.24 303.445 13.12 ;
    RECT 372.885 12.24 373.165 13.12 ;
    RECT 369.565 12.24 369.845 13.12 ;
    RECT 299.845 12.24 300.125 13.12 ;
    RECT 296.525 12.24 296.805 13.12 ;
    RECT 293.205 12.24 293.485 13.12 ;
    RECT 289.885 12.24 290.165 13.12 ;
    RECT 286.565 12.24 286.845 13.12 ;
    RECT 283.245 12.24 283.525 13.12 ;
    RECT 279.925 12.24 280.205 13.12 ;
    RECT 276.605 12.24 276.885 13.12 ;
    RECT 273.285 12.24 273.565 13.12 ;
    RECT 269.965 12.24 270.245 13.12 ;
    RECT 233.445 12.24 233.725 13.12 ;
    RECT 230.125 12.24 230.405 13.12 ;
    RECT 366.245 12.24 366.525 13.12 ;
    RECT 226.805 12.24 227.085 13.12 ;
    RECT 362.925 12.24 363.205 13.12 ;
    RECT 223.485 12.24 223.765 13.12 ;
    RECT 359.605 12.24 359.885 13.12 ;
    RECT 220.165 12.24 220.445 13.12 ;
    RECT 356.285 12.24 356.565 13.12 ;
    RECT 352.965 12.24 353.245 13.12 ;
    RECT 216.845 12.24 217.125 13.12 ;
    RECT 349.645 12.24 349.925 13.12 ;
    RECT 213.525 12.24 213.805 13.12 ;
    RECT 346.325 12.24 346.605 13.12 ;
    RECT 210.205 12.24 210.485 13.12 ;
    RECT 343.005 12.24 343.285 13.12 ;
    RECT 206.885 12.24 207.165 13.12 ;
    RECT 339.685 12.24 339.965 13.12 ;
    RECT 203.565 12.24 203.845 13.12 ;
    RECT 336.365 12.24 336.645 13.12 ;
    RECT 266.645 12.24 266.925 13.12 ;
    RECT 263.325 12.24 263.605 13.12 ;
    RECT 260.005 12.24 260.285 13.12 ;
    RECT 256.685 12.24 256.965 13.12 ;
    RECT 253.365 12.24 253.645 13.12 ;
    RECT 250.045 12.24 250.325 13.12 ;
    RECT 246.725 12.24 247.005 13.12 ;
    RECT 243.405 12.24 243.685 13.12 ;
    RECT 240.085 12.24 240.365 13.12 ;
    RECT 236.765 12.24 237.045 13.12 ;
    RECT 333.045 12.24 333.325 13.12 ;
    RECT 329.725 12.24 330.005 13.12 ;
    RECT 326.405 12.24 326.685 13.12 ;
    RECT 323.085 12.24 323.365 13.12 ;
    RECT 319.765 12.24 320.045 13.12 ;
    RECT 316.445 12.24 316.725 13.12 ;
    RECT 313.125 12.24 313.405 13.12 ;
    RECT 309.805 12.24 310.085 13.12 ;
    RECT 306.485 12.24 306.765 13.12 ;
    RECT 303.165 28.08 303.445 28.96 ;
    RECT 372.885 28.08 373.165 28.96 ;
    RECT 369.565 28.08 369.845 28.96 ;
    RECT 299.845 28.08 300.125 28.96 ;
    RECT 296.525 28.08 296.805 28.96 ;
    RECT 293.205 28.08 293.485 28.96 ;
    RECT 289.885 28.08 290.165 28.96 ;
    RECT 286.565 28.08 286.845 28.96 ;
    RECT 283.245 28.08 283.525 28.96 ;
    RECT 279.925 28.08 280.205 28.96 ;
    RECT 276.605 28.08 276.885 28.96 ;
    RECT 273.285 28.08 273.565 28.96 ;
    RECT 269.965 28.08 270.245 28.96 ;
    RECT 233.445 28.08 233.725 28.96 ;
    RECT 230.125 28.08 230.405 28.96 ;
    RECT 366.245 28.08 366.525 28.96 ;
    RECT 226.805 28.08 227.085 28.96 ;
    RECT 362.925 28.08 363.205 28.96 ;
    RECT 223.485 28.08 223.765 28.96 ;
    RECT 359.605 28.08 359.885 28.96 ;
    RECT 220.165 28.08 220.445 28.96 ;
    RECT 356.285 28.08 356.565 28.96 ;
    RECT 352.965 28.08 353.245 28.96 ;
    RECT 216.845 28.08 217.125 28.96 ;
    RECT 349.645 28.08 349.925 28.96 ;
    RECT 213.525 28.08 213.805 28.96 ;
    RECT 346.325 28.08 346.605 28.96 ;
    RECT 210.205 28.08 210.485 28.96 ;
    RECT 343.005 28.08 343.285 28.96 ;
    RECT 206.885 28.08 207.165 28.96 ;
    RECT 339.685 28.08 339.965 28.96 ;
    RECT 203.565 28.08 203.845 28.96 ;
    RECT 336.365 28.08 336.645 28.96 ;
    RECT 266.645 28.08 266.925 28.96 ;
    RECT 263.325 28.08 263.605 28.96 ;
    RECT 260.005 28.08 260.285 28.96 ;
    RECT 256.685 28.08 256.965 28.96 ;
    RECT 253.365 28.08 253.645 28.96 ;
    RECT 250.045 28.08 250.325 28.96 ;
    RECT 246.725 28.08 247.005 28.96 ;
    RECT 243.405 28.08 243.685 28.96 ;
    RECT 240.085 28.08 240.365 28.96 ;
    RECT 236.765 28.08 237.045 28.96 ;
    RECT 333.045 28.08 333.325 28.96 ;
    RECT 329.725 28.08 330.005 28.96 ;
    RECT 326.405 28.08 326.685 28.96 ;
    RECT 323.085 28.08 323.365 28.96 ;
    RECT 319.765 28.08 320.045 28.96 ;
    RECT 316.445 28.08 316.725 28.96 ;
    RECT 313.125 28.08 313.405 28.96 ;
    RECT 309.805 28.08 310.085 28.96 ;
    RECT 306.485 28.08 306.765 28.96 ;
    RECT 303.165 27.36 303.445 28.24 ;
    RECT 372.885 27.36 373.165 28.24 ;
    RECT 369.565 27.36 369.845 28.24 ;
    RECT 299.845 27.36 300.125 28.24 ;
    RECT 296.525 27.36 296.805 28.24 ;
    RECT 293.205 27.36 293.485 28.24 ;
    RECT 289.885 27.36 290.165 28.24 ;
    RECT 286.565 27.36 286.845 28.24 ;
    RECT 283.245 27.36 283.525 28.24 ;
    RECT 279.925 27.36 280.205 28.24 ;
    RECT 276.605 27.36 276.885 28.24 ;
    RECT 273.285 27.36 273.565 28.24 ;
    RECT 269.965 27.36 270.245 28.24 ;
    RECT 233.445 27.36 233.725 28.24 ;
    RECT 230.125 27.36 230.405 28.24 ;
    RECT 366.245 27.36 366.525 28.24 ;
    RECT 226.805 27.36 227.085 28.24 ;
    RECT 362.925 27.36 363.205 28.24 ;
    RECT 223.485 27.36 223.765 28.24 ;
    RECT 359.605 27.36 359.885 28.24 ;
    RECT 220.165 27.36 220.445 28.24 ;
    RECT 356.285 27.36 356.565 28.24 ;
    RECT 352.965 27.36 353.245 28.24 ;
    RECT 216.845 27.36 217.125 28.24 ;
    RECT 349.645 27.36 349.925 28.24 ;
    RECT 213.525 27.36 213.805 28.24 ;
    RECT 346.325 27.36 346.605 28.24 ;
    RECT 210.205 27.36 210.485 28.24 ;
    RECT 343.005 27.36 343.285 28.24 ;
    RECT 206.885 27.36 207.165 28.24 ;
    RECT 339.685 27.36 339.965 28.24 ;
    RECT 203.565 27.36 203.845 28.24 ;
    RECT 336.365 27.36 336.645 28.24 ;
    RECT 266.645 27.36 266.925 28.24 ;
    RECT 263.325 27.36 263.605 28.24 ;
    RECT 260.005 27.36 260.285 28.24 ;
    RECT 256.685 27.36 256.965 28.24 ;
    RECT 253.365 27.36 253.645 28.24 ;
    RECT 250.045 27.36 250.325 28.24 ;
    RECT 246.725 27.36 247.005 28.24 ;
    RECT 243.405 27.36 243.685 28.24 ;
    RECT 240.085 27.36 240.365 28.24 ;
    RECT 236.765 27.36 237.045 28.24 ;
    RECT 333.045 27.36 333.325 28.24 ;
    RECT 329.725 27.36 330.005 28.24 ;
    RECT 326.405 27.36 326.685 28.24 ;
    RECT 323.085 27.36 323.365 28.24 ;
    RECT 319.765 27.36 320.045 28.24 ;
    RECT 316.445 27.36 316.725 28.24 ;
    RECT 313.125 27.36 313.405 28.24 ;
    RECT 309.805 27.36 310.085 28.24 ;
    RECT 306.485 27.36 306.765 28.24 ;
    RECT 303.165 26.64 303.445 27.52 ;
    RECT 372.885 26.64 373.165 27.52 ;
    RECT 369.565 26.64 369.845 27.52 ;
    RECT 299.845 26.64 300.125 27.52 ;
    RECT 296.525 26.64 296.805 27.52 ;
    RECT 293.205 26.64 293.485 27.52 ;
    RECT 289.885 26.64 290.165 27.52 ;
    RECT 286.565 26.64 286.845 27.52 ;
    RECT 283.245 26.64 283.525 27.52 ;
    RECT 279.925 26.64 280.205 27.52 ;
    RECT 276.605 26.64 276.885 27.52 ;
    RECT 273.285 26.64 273.565 27.52 ;
    RECT 269.965 26.64 270.245 27.52 ;
    RECT 233.445 26.64 233.725 27.52 ;
    RECT 230.125 26.64 230.405 27.52 ;
    RECT 366.245 26.64 366.525 27.52 ;
    RECT 226.805 26.64 227.085 27.52 ;
    RECT 362.925 26.64 363.205 27.52 ;
    RECT 223.485 26.64 223.765 27.52 ;
    RECT 359.605 26.64 359.885 27.52 ;
    RECT 220.165 26.64 220.445 27.52 ;
    RECT 356.285 26.64 356.565 27.52 ;
    RECT 352.965 26.64 353.245 27.52 ;
    RECT 216.845 26.64 217.125 27.52 ;
    RECT 349.645 26.64 349.925 27.52 ;
    RECT 213.525 26.64 213.805 27.52 ;
    RECT 346.325 26.64 346.605 27.52 ;
    RECT 210.205 26.64 210.485 27.52 ;
    RECT 343.005 26.64 343.285 27.52 ;
    RECT 206.885 26.64 207.165 27.52 ;
    RECT 339.685 26.64 339.965 27.52 ;
    RECT 203.565 26.64 203.845 27.52 ;
    RECT 336.365 26.64 336.645 27.52 ;
    RECT 266.645 26.64 266.925 27.52 ;
    RECT 263.325 26.64 263.605 27.52 ;
    RECT 260.005 26.64 260.285 27.52 ;
    RECT 256.685 26.64 256.965 27.52 ;
    RECT 253.365 26.64 253.645 27.52 ;
    RECT 250.045 26.64 250.325 27.52 ;
    RECT 246.725 26.64 247.005 27.52 ;
    RECT 243.405 26.64 243.685 27.52 ;
    RECT 240.085 26.64 240.365 27.52 ;
    RECT 236.765 26.64 237.045 27.52 ;
    RECT 333.045 26.64 333.325 27.52 ;
    RECT 329.725 26.64 330.005 27.52 ;
    RECT 326.405 26.64 326.685 27.52 ;
    RECT 323.085 26.64 323.365 27.52 ;
    RECT 319.765 26.64 320.045 27.52 ;
    RECT 316.445 26.64 316.725 27.52 ;
    RECT 313.125 26.64 313.405 27.52 ;
    RECT 309.805 26.64 310.085 27.52 ;
    RECT 306.485 26.64 306.765 27.52 ;
    RECT 303.165 25.92 303.445 26.8 ;
    RECT 372.885 25.92 373.165 26.8 ;
    RECT 369.565 25.92 369.845 26.8 ;
    RECT 299.845 25.92 300.125 26.8 ;
    RECT 296.525 25.92 296.805 26.8 ;
    RECT 293.205 25.92 293.485 26.8 ;
    RECT 289.885 25.92 290.165 26.8 ;
    RECT 286.565 25.92 286.845 26.8 ;
    RECT 283.245 25.92 283.525 26.8 ;
    RECT 279.925 25.92 280.205 26.8 ;
    RECT 276.605 25.92 276.885 26.8 ;
    RECT 273.285 25.92 273.565 26.8 ;
    RECT 269.965 25.92 270.245 26.8 ;
    RECT 233.445 25.92 233.725 26.8 ;
    RECT 230.125 25.92 230.405 26.8 ;
    RECT 366.245 25.92 366.525 26.8 ;
    RECT 226.805 25.92 227.085 26.8 ;
    RECT 362.925 25.92 363.205 26.8 ;
    RECT 223.485 25.92 223.765 26.8 ;
    RECT 359.605 25.92 359.885 26.8 ;
    RECT 220.165 25.92 220.445 26.8 ;
    RECT 356.285 25.92 356.565 26.8 ;
    RECT 352.965 25.92 353.245 26.8 ;
    RECT 216.845 25.92 217.125 26.8 ;
    RECT 349.645 25.92 349.925 26.8 ;
    RECT 213.525 25.92 213.805 26.8 ;
    RECT 346.325 25.92 346.605 26.8 ;
    RECT 210.205 25.92 210.485 26.8 ;
    RECT 343.005 25.92 343.285 26.8 ;
    RECT 206.885 25.92 207.165 26.8 ;
    RECT 339.685 25.92 339.965 26.8 ;
    RECT 203.565 25.92 203.845 26.8 ;
    RECT 336.365 25.92 336.645 26.8 ;
    RECT 266.645 25.92 266.925 26.8 ;
    RECT 263.325 25.92 263.605 26.8 ;
    RECT 260.005 25.92 260.285 26.8 ;
    RECT 256.685 25.92 256.965 26.8 ;
    RECT 253.365 25.92 253.645 26.8 ;
    RECT 250.045 25.92 250.325 26.8 ;
    RECT 246.725 25.92 247.005 26.8 ;
    RECT 243.405 25.92 243.685 26.8 ;
    RECT 240.085 25.92 240.365 26.8 ;
    RECT 236.765 25.92 237.045 26.8 ;
    RECT 333.045 25.92 333.325 26.8 ;
    RECT 329.725 25.92 330.005 26.8 ;
    RECT 326.405 25.92 326.685 26.8 ;
    RECT 323.085 25.92 323.365 26.8 ;
    RECT 319.765 25.92 320.045 26.8 ;
    RECT 316.445 25.92 316.725 26.8 ;
    RECT 313.125 25.92 313.405 26.8 ;
    RECT 309.805 25.92 310.085 26.8 ;
    RECT 306.485 25.92 306.765 26.8 ;
    RECT 303.165 35.28 303.445 36.16 ;
    RECT 372.885 35.28 373.165 36.16 ;
    RECT 369.565 35.28 369.845 36.16 ;
    RECT 299.845 35.28 300.125 36.16 ;
    RECT 296.525 35.28 296.805 36.16 ;
    RECT 293.205 35.28 293.485 36.16 ;
    RECT 289.885 35.28 290.165 36.16 ;
    RECT 286.565 35.28 286.845 36.16 ;
    RECT 283.245 35.28 283.525 36.16 ;
    RECT 279.925 35.28 280.205 36.16 ;
    RECT 276.605 35.28 276.885 36.16 ;
    RECT 273.285 35.28 273.565 36.16 ;
    RECT 269.965 35.28 270.245 36.16 ;
    RECT 233.445 35.28 233.725 36.16 ;
    RECT 230.125 35.28 230.405 36.16 ;
    RECT 366.245 35.28 366.525 36.16 ;
    RECT 226.805 35.28 227.085 36.16 ;
    RECT 362.925 35.28 363.205 36.16 ;
    RECT 223.485 35.28 223.765 36.16 ;
    RECT 359.605 35.28 359.885 36.16 ;
    RECT 220.165 35.28 220.445 36.16 ;
    RECT 356.285 35.28 356.565 36.16 ;
    RECT 352.965 35.28 353.245 36.16 ;
    RECT 216.845 35.28 217.125 36.16 ;
    RECT 349.645 35.28 349.925 36.16 ;
    RECT 213.525 35.28 213.805 36.16 ;
    RECT 346.325 35.28 346.605 36.16 ;
    RECT 210.205 35.28 210.485 36.16 ;
    RECT 343.005 35.28 343.285 36.16 ;
    RECT 206.885 35.28 207.165 36.16 ;
    RECT 339.685 35.28 339.965 36.16 ;
    RECT 203.565 35.28 203.845 36.16 ;
    RECT 336.365 35.28 336.645 36.16 ;
    RECT 266.645 35.28 266.925 36.16 ;
    RECT 263.325 35.28 263.605 36.16 ;
    RECT 260.005 35.28 260.285 36.16 ;
    RECT 256.685 35.28 256.965 36.16 ;
    RECT 253.365 35.28 253.645 36.16 ;
    RECT 250.045 35.28 250.325 36.16 ;
    RECT 246.725 35.28 247.005 36.16 ;
    RECT 243.405 35.28 243.685 36.16 ;
    RECT 240.085 35.28 240.365 36.16 ;
    RECT 236.765 35.28 237.045 36.16 ;
    RECT 333.045 35.28 333.325 36.16 ;
    RECT 329.725 35.28 330.005 36.16 ;
    RECT 326.405 35.28 326.685 36.16 ;
    RECT 323.085 35.28 323.365 36.16 ;
    RECT 319.765 35.28 320.045 36.16 ;
    RECT 316.445 35.28 316.725 36.16 ;
    RECT 313.125 35.28 313.405 36.16 ;
    RECT 309.805 35.28 310.085 36.16 ;
    RECT 306.485 35.28 306.765 36.16 ;
    RECT 233.445 59.14 233.725 60.67 ;
    RECT 230.125 59.14 230.405 60.67 ;
    RECT 226.805 59.14 227.085 60.67 ;
    RECT 223.485 59.14 223.765 60.67 ;
    RECT 220.165 59.14 220.445 60.67 ;
    RECT 216.845 59.14 217.125 60.67 ;
    RECT 213.525 59.14 213.805 60.67 ;
    RECT 210.205 59.14 210.485 60.67 ;
    RECT 206.885 59.14 207.165 60.67 ;
    RECT 203.565 59.14 203.845 60.67 ;
    RECT 372.885 59.14 373.165 60.67 ;
    RECT 369.565 59.14 369.845 60.67 ;
    RECT 366.245 59.14 366.525 60.67 ;
    RECT 362.925 59.14 363.205 60.67 ;
    RECT 359.605 59.14 359.885 60.67 ;
    RECT 356.285 59.14 356.565 60.67 ;
    RECT 352.965 59.14 353.245 60.67 ;
    RECT 349.645 59.14 349.925 60.67 ;
    RECT 346.325 59.14 346.605 60.67 ;
    RECT 343.005 59.14 343.285 60.67 ;
    RECT 339.685 59.14 339.965 60.67 ;
    RECT 336.365 59.14 336.645 60.67 ;
    RECT 333.045 59.14 333.325 60.67 ;
    RECT 329.725 59.14 330.005 60.67 ;
    RECT 326.405 59.14 326.685 60.67 ;
    RECT 323.085 59.14 323.365 60.67 ;
    RECT 319.765 59.14 320.045 60.67 ;
    RECT 316.445 59.14 316.725 60.67 ;
    RECT 313.125 59.14 313.405 60.67 ;
    RECT 309.805 59.14 310.085 60.67 ;
    RECT 306.485 59.14 306.765 60.67 ;
    RECT 303.165 59.14 303.445 60.67 ;
    RECT 299.845 59.14 300.125 60.67 ;
    RECT 296.525 59.14 296.805 60.67 ;
    RECT 293.205 59.14 293.485 60.67 ;
    RECT 289.885 59.14 290.165 60.67 ;
    RECT 286.565 59.14 286.845 60.67 ;
    RECT 283.245 59.14 283.525 60.67 ;
    RECT 279.925 59.14 280.205 60.67 ;
    RECT 276.605 59.14 276.885 60.67 ;
    RECT 273.285 59.14 273.565 60.67 ;
    RECT 269.965 59.14 270.245 60.67 ;
    RECT 266.645 59.14 266.925 60.67 ;
    RECT 263.325 59.14 263.605 60.67 ;
    RECT 260.005 59.14 260.285 60.67 ;
    RECT 256.685 59.14 256.965 60.67 ;
    RECT 253.365 59.14 253.645 60.67 ;
    RECT 250.045 59.14 250.325 60.67 ;
    RECT 246.725 59.14 247.005 60.67 ;
    RECT 243.405 59.14 243.685 60.67 ;
    RECT 240.085 59.14 240.365 60.67 ;
    RECT 236.765 59.14 237.045 60.67 ;
    RECT 303.165 25.2 303.445 26.08 ;
    RECT 372.885 25.2 373.165 26.08 ;
    RECT 369.565 25.2 369.845 26.08 ;
    RECT 299.845 25.2 300.125 26.08 ;
    RECT 296.525 25.2 296.805 26.08 ;
    RECT 293.205 25.2 293.485 26.08 ;
    RECT 289.885 25.2 290.165 26.08 ;
    RECT 286.565 25.2 286.845 26.08 ;
    RECT 283.245 25.2 283.525 26.08 ;
    RECT 279.925 25.2 280.205 26.08 ;
    RECT 276.605 25.2 276.885 26.08 ;
    RECT 273.285 25.2 273.565 26.08 ;
    RECT 269.965 25.2 270.245 26.08 ;
    RECT 233.445 25.2 233.725 26.08 ;
    RECT 230.125 25.2 230.405 26.08 ;
    RECT 366.245 25.2 366.525 26.08 ;
    RECT 226.805 25.2 227.085 26.08 ;
    RECT 362.925 25.2 363.205 26.08 ;
    RECT 223.485 25.2 223.765 26.08 ;
    RECT 359.605 25.2 359.885 26.08 ;
    RECT 220.165 25.2 220.445 26.08 ;
    RECT 356.285 25.2 356.565 26.08 ;
    RECT 352.965 25.2 353.245 26.08 ;
    RECT 216.845 25.2 217.125 26.08 ;
    RECT 349.645 25.2 349.925 26.08 ;
    RECT 213.525 25.2 213.805 26.08 ;
    RECT 346.325 25.2 346.605 26.08 ;
    RECT 210.205 25.2 210.485 26.08 ;
    RECT 343.005 25.2 343.285 26.08 ;
    RECT 206.885 25.2 207.165 26.08 ;
    RECT 339.685 25.2 339.965 26.08 ;
    RECT 203.565 25.2 203.845 26.08 ;
    RECT 336.365 25.2 336.645 26.08 ;
    RECT 266.645 25.2 266.925 26.08 ;
    RECT 263.325 25.2 263.605 26.08 ;
    RECT 260.005 25.2 260.285 26.08 ;
    RECT 256.685 25.2 256.965 26.08 ;
    RECT 253.365 25.2 253.645 26.08 ;
    RECT 250.045 25.2 250.325 26.08 ;
    RECT 246.725 25.2 247.005 26.08 ;
    RECT 243.405 25.2 243.685 26.08 ;
    RECT 240.085 25.2 240.365 26.08 ;
    RECT 236.765 25.2 237.045 26.08 ;
    RECT 333.045 25.2 333.325 26.08 ;
    RECT 329.725 25.2 330.005 26.08 ;
    RECT 326.405 25.2 326.685 26.08 ;
    RECT 323.085 25.2 323.365 26.08 ;
    RECT 319.765 25.2 320.045 26.08 ;
    RECT 316.445 25.2 316.725 26.08 ;
    RECT 313.125 25.2 313.405 26.08 ;
    RECT 309.805 25.2 310.085 26.08 ;
    RECT 306.485 25.2 306.765 26.08 ;
    RECT 303.165 24.48 303.445 25.36 ;
    RECT 372.885 24.48 373.165 25.36 ;
    RECT 369.565 24.48 369.845 25.36 ;
    RECT 299.845 24.48 300.125 25.36 ;
    RECT 296.525 24.48 296.805 25.36 ;
    RECT 293.205 24.48 293.485 25.36 ;
    RECT 289.885 24.48 290.165 25.36 ;
    RECT 286.565 24.48 286.845 25.36 ;
    RECT 283.245 24.48 283.525 25.36 ;
    RECT 279.925 24.48 280.205 25.36 ;
    RECT 276.605 24.48 276.885 25.36 ;
    RECT 273.285 24.48 273.565 25.36 ;
    RECT 269.965 24.48 270.245 25.36 ;
    RECT 233.445 24.48 233.725 25.36 ;
    RECT 230.125 24.48 230.405 25.36 ;
    RECT 366.245 24.48 366.525 25.36 ;
    RECT 226.805 24.48 227.085 25.36 ;
    RECT 362.925 24.48 363.205 25.36 ;
    RECT 223.485 24.48 223.765 25.36 ;
    RECT 359.605 24.48 359.885 25.36 ;
    RECT 220.165 24.48 220.445 25.36 ;
    RECT 356.285 24.48 356.565 25.36 ;
    RECT 352.965 24.48 353.245 25.36 ;
    RECT 216.845 24.48 217.125 25.36 ;
    RECT 349.645 24.48 349.925 25.36 ;
    RECT 213.525 24.48 213.805 25.36 ;
    RECT 346.325 24.48 346.605 25.36 ;
    RECT 210.205 24.48 210.485 25.36 ;
    RECT 343.005 24.48 343.285 25.36 ;
    RECT 206.885 24.48 207.165 25.36 ;
    RECT 339.685 24.48 339.965 25.36 ;
    RECT 203.565 24.48 203.845 25.36 ;
    RECT 336.365 24.48 336.645 25.36 ;
    RECT 266.645 24.48 266.925 25.36 ;
    RECT 263.325 24.48 263.605 25.36 ;
    RECT 260.005 24.48 260.285 25.36 ;
    RECT 256.685 24.48 256.965 25.36 ;
    RECT 253.365 24.48 253.645 25.36 ;
    RECT 250.045 24.48 250.325 25.36 ;
    RECT 246.725 24.48 247.005 25.36 ;
    RECT 243.405 24.48 243.685 25.36 ;
    RECT 240.085 24.48 240.365 25.36 ;
    RECT 236.765 24.48 237.045 25.36 ;
    RECT 333.045 24.48 333.325 25.36 ;
    RECT 329.725 24.48 330.005 25.36 ;
    RECT 326.405 24.48 326.685 25.36 ;
    RECT 323.085 24.48 323.365 25.36 ;
    RECT 319.765 24.48 320.045 25.36 ;
    RECT 316.445 24.48 316.725 25.36 ;
    RECT 313.125 24.48 313.405 25.36 ;
    RECT 309.805 24.48 310.085 25.36 ;
    RECT 306.485 24.48 306.765 25.36 ;
    RECT 303.165 23.76 303.445 24.64 ;
    RECT 372.885 23.76 373.165 24.64 ;
    RECT 369.565 23.76 369.845 24.64 ;
    RECT 299.845 23.76 300.125 24.64 ;
    RECT 296.525 23.76 296.805 24.64 ;
    RECT 293.205 23.76 293.485 24.64 ;
    RECT 289.885 23.76 290.165 24.64 ;
    RECT 286.565 23.76 286.845 24.64 ;
    RECT 283.245 23.76 283.525 24.64 ;
    RECT 279.925 23.76 280.205 24.64 ;
    RECT 276.605 23.76 276.885 24.64 ;
    RECT 273.285 23.76 273.565 24.64 ;
    RECT 269.965 23.76 270.245 24.64 ;
    RECT 233.445 23.76 233.725 24.64 ;
    RECT 230.125 23.76 230.405 24.64 ;
    RECT 366.245 23.76 366.525 24.64 ;
    RECT 226.805 23.76 227.085 24.64 ;
    RECT 362.925 23.76 363.205 24.64 ;
    RECT 223.485 23.76 223.765 24.64 ;
    RECT 359.605 23.76 359.885 24.64 ;
    RECT 220.165 23.76 220.445 24.64 ;
    RECT 356.285 23.76 356.565 24.64 ;
    RECT 352.965 23.76 353.245 24.64 ;
    RECT 216.845 23.76 217.125 24.64 ;
    RECT 349.645 23.76 349.925 24.64 ;
    RECT 213.525 23.76 213.805 24.64 ;
    RECT 346.325 23.76 346.605 24.64 ;
    RECT 210.205 23.76 210.485 24.64 ;
    RECT 343.005 23.76 343.285 24.64 ;
    RECT 206.885 23.76 207.165 24.64 ;
    RECT 339.685 23.76 339.965 24.64 ;
    RECT 203.565 23.76 203.845 24.64 ;
    RECT 336.365 23.76 336.645 24.64 ;
    RECT 266.645 23.76 266.925 24.64 ;
    RECT 263.325 23.76 263.605 24.64 ;
    RECT 260.005 23.76 260.285 24.64 ;
    RECT 256.685 23.76 256.965 24.64 ;
    RECT 253.365 23.76 253.645 24.64 ;
    RECT 250.045 23.76 250.325 24.64 ;
    RECT 246.725 23.76 247.005 24.64 ;
    RECT 243.405 23.76 243.685 24.64 ;
    RECT 240.085 23.76 240.365 24.64 ;
    RECT 236.765 23.76 237.045 24.64 ;
    RECT 333.045 23.76 333.325 24.64 ;
    RECT 329.725 23.76 330.005 24.64 ;
    RECT 326.405 23.76 326.685 24.64 ;
    RECT 323.085 23.76 323.365 24.64 ;
    RECT 319.765 23.76 320.045 24.64 ;
    RECT 316.445 23.76 316.725 24.64 ;
    RECT 313.125 23.76 313.405 24.64 ;
    RECT 309.805 23.76 310.085 24.64 ;
    RECT 306.485 23.76 306.765 24.64 ;
    RECT 303.165 23.04 303.445 23.92 ;
    RECT 372.885 23.04 373.165 23.92 ;
    RECT 369.565 23.04 369.845 23.92 ;
    RECT 299.845 23.04 300.125 23.92 ;
    RECT 296.525 23.04 296.805 23.92 ;
    RECT 293.205 23.04 293.485 23.92 ;
    RECT 289.885 23.04 290.165 23.92 ;
    RECT 286.565 23.04 286.845 23.92 ;
    RECT 283.245 23.04 283.525 23.92 ;
    RECT 279.925 23.04 280.205 23.92 ;
    RECT 276.605 23.04 276.885 23.92 ;
    RECT 273.285 23.04 273.565 23.92 ;
    RECT 269.965 23.04 270.245 23.92 ;
    RECT 233.445 23.04 233.725 23.92 ;
    RECT 230.125 23.04 230.405 23.92 ;
    RECT 366.245 23.04 366.525 23.92 ;
    RECT 226.805 23.04 227.085 23.92 ;
    RECT 362.925 23.04 363.205 23.92 ;
    RECT 223.485 23.04 223.765 23.92 ;
    RECT 359.605 23.04 359.885 23.92 ;
    RECT 220.165 23.04 220.445 23.92 ;
    RECT 356.285 23.04 356.565 23.92 ;
    RECT 352.965 23.04 353.245 23.92 ;
    RECT 216.845 23.04 217.125 23.92 ;
    RECT 349.645 23.04 349.925 23.92 ;
    RECT 213.525 23.04 213.805 23.92 ;
    RECT 346.325 23.04 346.605 23.92 ;
    RECT 210.205 23.04 210.485 23.92 ;
    RECT 343.005 23.04 343.285 23.92 ;
    RECT 206.885 23.04 207.165 23.92 ;
    RECT 339.685 23.04 339.965 23.92 ;
    RECT 203.565 23.04 203.845 23.92 ;
    RECT 336.365 23.04 336.645 23.92 ;
    RECT 266.645 23.04 266.925 23.92 ;
    RECT 263.325 23.04 263.605 23.92 ;
    RECT 260.005 23.04 260.285 23.92 ;
    RECT 256.685 23.04 256.965 23.92 ;
    RECT 253.365 23.04 253.645 23.92 ;
    RECT 250.045 23.04 250.325 23.92 ;
    RECT 246.725 23.04 247.005 23.92 ;
    RECT 243.405 23.04 243.685 23.92 ;
    RECT 240.085 23.04 240.365 23.92 ;
    RECT 236.765 23.04 237.045 23.92 ;
    RECT 333.045 23.04 333.325 23.92 ;
    RECT 329.725 23.04 330.005 23.92 ;
    RECT 326.405 23.04 326.685 23.92 ;
    RECT 323.085 23.04 323.365 23.92 ;
    RECT 319.765 23.04 320.045 23.92 ;
    RECT 316.445 23.04 316.725 23.92 ;
    RECT 313.125 23.04 313.405 23.92 ;
    RECT 309.805 23.04 310.085 23.92 ;
    RECT 306.485 23.04 306.765 23.92 ;
    RECT 303.165 22.32 303.445 23.2 ;
    RECT 372.885 22.32 373.165 23.2 ;
    RECT 369.565 22.32 369.845 23.2 ;
    RECT 299.845 22.32 300.125 23.2 ;
    RECT 296.525 22.32 296.805 23.2 ;
    RECT 293.205 22.32 293.485 23.2 ;
    RECT 289.885 22.32 290.165 23.2 ;
    RECT 286.565 22.32 286.845 23.2 ;
    RECT 283.245 22.32 283.525 23.2 ;
    RECT 279.925 22.32 280.205 23.2 ;
    RECT 276.605 22.32 276.885 23.2 ;
    RECT 273.285 22.32 273.565 23.2 ;
    RECT 269.965 22.32 270.245 23.2 ;
    RECT 233.445 22.32 233.725 23.2 ;
    RECT 230.125 22.32 230.405 23.2 ;
    RECT 366.245 22.32 366.525 23.2 ;
    RECT 226.805 22.32 227.085 23.2 ;
    RECT 362.925 22.32 363.205 23.2 ;
    RECT 223.485 22.32 223.765 23.2 ;
    RECT 359.605 22.32 359.885 23.2 ;
    RECT 220.165 22.32 220.445 23.2 ;
    RECT 356.285 22.32 356.565 23.2 ;
    RECT 352.965 22.32 353.245 23.2 ;
    RECT 216.845 22.32 217.125 23.2 ;
    RECT 349.645 22.32 349.925 23.2 ;
    RECT 213.525 22.32 213.805 23.2 ;
    RECT 346.325 22.32 346.605 23.2 ;
    RECT 210.205 22.32 210.485 23.2 ;
    RECT 343.005 22.32 343.285 23.2 ;
    RECT 206.885 22.32 207.165 23.2 ;
    RECT 339.685 22.32 339.965 23.2 ;
    RECT 203.565 22.32 203.845 23.2 ;
    RECT 336.365 22.32 336.645 23.2 ;
    RECT 266.645 22.32 266.925 23.2 ;
    RECT 263.325 22.32 263.605 23.2 ;
    RECT 260.005 22.32 260.285 23.2 ;
    RECT 256.685 22.32 256.965 23.2 ;
    RECT 253.365 22.32 253.645 23.2 ;
    RECT 250.045 22.32 250.325 23.2 ;
    RECT 246.725 22.32 247.005 23.2 ;
    RECT 243.405 22.32 243.685 23.2 ;
    RECT 240.085 22.32 240.365 23.2 ;
    RECT 236.765 22.32 237.045 23.2 ;
    RECT 333.045 22.32 333.325 23.2 ;
    RECT 329.725 22.32 330.005 23.2 ;
    RECT 326.405 22.32 326.685 23.2 ;
    RECT 323.085 22.32 323.365 23.2 ;
    RECT 319.765 22.32 320.045 23.2 ;
    RECT 316.445 22.32 316.725 23.2 ;
    RECT 313.125 22.32 313.405 23.2 ;
    RECT 309.805 22.32 310.085 23.2 ;
    RECT 306.485 22.32 306.765 23.2 ;
    RECT 303.165 21.6 303.445 22.48 ;
    RECT 372.885 21.6 373.165 22.48 ;
    RECT 369.565 21.6 369.845 22.48 ;
    RECT 299.845 21.6 300.125 22.48 ;
    RECT 296.525 21.6 296.805 22.48 ;
    RECT 293.205 21.6 293.485 22.48 ;
    RECT 289.885 21.6 290.165 22.48 ;
    RECT 286.565 21.6 286.845 22.48 ;
    RECT 283.245 21.6 283.525 22.48 ;
    RECT 279.925 21.6 280.205 22.48 ;
    RECT 276.605 21.6 276.885 22.48 ;
    RECT 273.285 21.6 273.565 22.48 ;
    RECT 269.965 21.6 270.245 22.48 ;
    RECT 233.445 21.6 233.725 22.48 ;
    RECT 230.125 21.6 230.405 22.48 ;
    RECT 366.245 21.6 366.525 22.48 ;
    RECT 226.805 21.6 227.085 22.48 ;
    RECT 362.925 21.6 363.205 22.48 ;
    RECT 223.485 21.6 223.765 22.48 ;
    RECT 359.605 21.6 359.885 22.48 ;
    RECT 220.165 21.6 220.445 22.48 ;
    RECT 356.285 21.6 356.565 22.48 ;
    RECT 352.965 21.6 353.245 22.48 ;
    RECT 216.845 21.6 217.125 22.48 ;
    RECT 349.645 21.6 349.925 22.48 ;
    RECT 213.525 21.6 213.805 22.48 ;
    RECT 346.325 21.6 346.605 22.48 ;
    RECT 210.205 21.6 210.485 22.48 ;
    RECT 343.005 21.6 343.285 22.48 ;
    RECT 206.885 21.6 207.165 22.48 ;
    RECT 339.685 21.6 339.965 22.48 ;
    RECT 203.565 21.6 203.845 22.48 ;
    RECT 336.365 21.6 336.645 22.48 ;
    RECT 266.645 21.6 266.925 22.48 ;
    RECT 263.325 21.6 263.605 22.48 ;
    RECT 260.005 21.6 260.285 22.48 ;
    RECT 256.685 21.6 256.965 22.48 ;
    RECT 253.365 21.6 253.645 22.48 ;
    RECT 250.045 21.6 250.325 22.48 ;
    RECT 246.725 21.6 247.005 22.48 ;
    RECT 243.405 21.6 243.685 22.48 ;
    RECT 240.085 21.6 240.365 22.48 ;
    RECT 236.765 21.6 237.045 22.48 ;
    RECT 333.045 21.6 333.325 22.48 ;
    RECT 329.725 21.6 330.005 22.48 ;
    RECT 326.405 21.6 326.685 22.48 ;
    RECT 323.085 21.6 323.365 22.48 ;
    RECT 319.765 21.6 320.045 22.48 ;
    RECT 316.445 21.6 316.725 22.48 ;
    RECT 313.125 21.6 313.405 22.48 ;
    RECT 309.805 21.6 310.085 22.48 ;
    RECT 306.485 21.6 306.765 22.48 ;
    RECT 303.165 20.88 303.445 21.76 ;
    RECT 372.885 20.88 373.165 21.76 ;
    RECT 369.565 20.88 369.845 21.76 ;
    RECT 299.845 20.88 300.125 21.76 ;
    RECT 296.525 20.88 296.805 21.76 ;
    RECT 293.205 20.88 293.485 21.76 ;
    RECT 289.885 20.88 290.165 21.76 ;
    RECT 286.565 20.88 286.845 21.76 ;
    RECT 283.245 20.88 283.525 21.76 ;
    RECT 279.925 20.88 280.205 21.76 ;
    RECT 276.605 20.88 276.885 21.76 ;
    RECT 273.285 20.88 273.565 21.76 ;
    RECT 269.965 20.88 270.245 21.76 ;
    RECT 233.445 20.88 233.725 21.76 ;
    RECT 230.125 20.88 230.405 21.76 ;
    RECT 366.245 20.88 366.525 21.76 ;
    RECT 226.805 20.88 227.085 21.76 ;
    RECT 362.925 20.88 363.205 21.76 ;
    RECT 223.485 20.88 223.765 21.76 ;
    RECT 359.605 20.88 359.885 21.76 ;
    RECT 220.165 20.88 220.445 21.76 ;
    RECT 356.285 20.88 356.565 21.76 ;
    RECT 352.965 20.88 353.245 21.76 ;
    RECT 216.845 20.88 217.125 21.76 ;
    RECT 349.645 20.88 349.925 21.76 ;
    RECT 213.525 20.88 213.805 21.76 ;
    RECT 346.325 20.88 346.605 21.76 ;
    RECT 210.205 20.88 210.485 21.76 ;
    RECT 343.005 20.88 343.285 21.76 ;
    RECT 206.885 20.88 207.165 21.76 ;
    RECT 339.685 20.88 339.965 21.76 ;
    RECT 203.565 20.88 203.845 21.76 ;
    RECT 336.365 20.88 336.645 21.76 ;
    RECT 266.645 20.88 266.925 21.76 ;
    RECT 263.325 20.88 263.605 21.76 ;
    RECT 260.005 20.88 260.285 21.76 ;
    RECT 256.685 20.88 256.965 21.76 ;
    RECT 253.365 20.88 253.645 21.76 ;
    RECT 250.045 20.88 250.325 21.76 ;
    RECT 246.725 20.88 247.005 21.76 ;
    RECT 243.405 20.88 243.685 21.76 ;
    RECT 240.085 20.88 240.365 21.76 ;
    RECT 236.765 20.88 237.045 21.76 ;
    RECT 333.045 20.88 333.325 21.76 ;
    RECT 329.725 20.88 330.005 21.76 ;
    RECT 326.405 20.88 326.685 21.76 ;
    RECT 323.085 20.88 323.365 21.76 ;
    RECT 319.765 20.88 320.045 21.76 ;
    RECT 316.445 20.88 316.725 21.76 ;
    RECT 313.125 20.88 313.405 21.76 ;
    RECT 309.805 20.88 310.085 21.76 ;
    RECT 306.485 20.88 306.765 21.76 ;
    RECT 303.165 34.56 303.445 35.44 ;
    RECT 372.885 34.56 373.165 35.44 ;
    RECT 369.565 34.56 369.845 35.44 ;
    RECT 299.845 34.56 300.125 35.44 ;
    RECT 296.525 34.56 296.805 35.44 ;
    RECT 293.205 34.56 293.485 35.44 ;
    RECT 289.885 34.56 290.165 35.44 ;
    RECT 286.565 34.56 286.845 35.44 ;
    RECT 283.245 34.56 283.525 35.44 ;
    RECT 279.925 34.56 280.205 35.44 ;
    RECT 276.605 34.56 276.885 35.44 ;
    RECT 273.285 34.56 273.565 35.44 ;
    RECT 269.965 34.56 270.245 35.44 ;
    RECT 233.445 34.56 233.725 35.44 ;
    RECT 230.125 34.56 230.405 35.44 ;
    RECT 366.245 34.56 366.525 35.44 ;
    RECT 226.805 34.56 227.085 35.44 ;
    RECT 362.925 34.56 363.205 35.44 ;
    RECT 223.485 34.56 223.765 35.44 ;
    RECT 359.605 34.56 359.885 35.44 ;
    RECT 220.165 34.56 220.445 35.44 ;
    RECT 356.285 34.56 356.565 35.44 ;
    RECT 352.965 34.56 353.245 35.44 ;
    RECT 216.845 34.56 217.125 35.44 ;
    RECT 349.645 34.56 349.925 35.44 ;
    RECT 213.525 34.56 213.805 35.44 ;
    RECT 346.325 34.56 346.605 35.44 ;
    RECT 210.205 34.56 210.485 35.44 ;
    RECT 343.005 34.56 343.285 35.44 ;
    RECT 206.885 34.56 207.165 35.44 ;
    RECT 339.685 34.56 339.965 35.44 ;
    RECT 203.565 34.56 203.845 35.44 ;
    RECT 336.365 34.56 336.645 35.44 ;
    RECT 266.645 34.56 266.925 35.44 ;
    RECT 263.325 34.56 263.605 35.44 ;
    RECT 260.005 34.56 260.285 35.44 ;
    RECT 256.685 34.56 256.965 35.44 ;
    RECT 253.365 34.56 253.645 35.44 ;
    RECT 250.045 34.56 250.325 35.44 ;
    RECT 246.725 34.56 247.005 35.44 ;
    RECT 243.405 34.56 243.685 35.44 ;
    RECT 240.085 34.56 240.365 35.44 ;
    RECT 236.765 34.56 237.045 35.44 ;
    RECT 333.045 34.56 333.325 35.44 ;
    RECT 329.725 34.56 330.005 35.44 ;
    RECT 326.405 34.56 326.685 35.44 ;
    RECT 323.085 34.56 323.365 35.44 ;
    RECT 319.765 34.56 320.045 35.44 ;
    RECT 316.445 34.56 316.725 35.44 ;
    RECT 313.125 34.56 313.405 35.44 ;
    RECT 309.805 34.56 310.085 35.44 ;
    RECT 306.485 34.56 306.765 35.44 ;
    RECT 303.165 20.16 303.445 21.04 ;
    RECT 372.885 20.16 373.165 21.04 ;
    RECT 369.565 20.16 369.845 21.04 ;
    RECT 299.845 20.16 300.125 21.04 ;
    RECT 296.525 20.16 296.805 21.04 ;
    RECT 293.205 20.16 293.485 21.04 ;
    RECT 289.885 20.16 290.165 21.04 ;
    RECT 286.565 20.16 286.845 21.04 ;
    RECT 283.245 20.16 283.525 21.04 ;
    RECT 279.925 20.16 280.205 21.04 ;
    RECT 276.605 20.16 276.885 21.04 ;
    RECT 273.285 20.16 273.565 21.04 ;
    RECT 269.965 20.16 270.245 21.04 ;
    RECT 233.445 20.16 233.725 21.04 ;
    RECT 230.125 20.16 230.405 21.04 ;
    RECT 366.245 20.16 366.525 21.04 ;
    RECT 226.805 20.16 227.085 21.04 ;
    RECT 362.925 20.16 363.205 21.04 ;
    RECT 223.485 20.16 223.765 21.04 ;
    RECT 359.605 20.16 359.885 21.04 ;
    RECT 220.165 20.16 220.445 21.04 ;
    RECT 356.285 20.16 356.565 21.04 ;
    RECT 352.965 20.16 353.245 21.04 ;
    RECT 216.845 20.16 217.125 21.04 ;
    RECT 349.645 20.16 349.925 21.04 ;
    RECT 213.525 20.16 213.805 21.04 ;
    RECT 346.325 20.16 346.605 21.04 ;
    RECT 210.205 20.16 210.485 21.04 ;
    RECT 343.005 20.16 343.285 21.04 ;
    RECT 206.885 20.16 207.165 21.04 ;
    RECT 339.685 20.16 339.965 21.04 ;
    RECT 203.565 20.16 203.845 21.04 ;
    RECT 336.365 20.16 336.645 21.04 ;
    RECT 266.645 20.16 266.925 21.04 ;
    RECT 263.325 20.16 263.605 21.04 ;
    RECT 260.005 20.16 260.285 21.04 ;
    RECT 256.685 20.16 256.965 21.04 ;
    RECT 253.365 20.16 253.645 21.04 ;
    RECT 250.045 20.16 250.325 21.04 ;
    RECT 246.725 20.16 247.005 21.04 ;
    RECT 243.405 20.16 243.685 21.04 ;
    RECT 240.085 20.16 240.365 21.04 ;
    RECT 236.765 20.16 237.045 21.04 ;
    RECT 333.045 20.16 333.325 21.04 ;
    RECT 329.725 20.16 330.005 21.04 ;
    RECT 326.405 20.16 326.685 21.04 ;
    RECT 323.085 20.16 323.365 21.04 ;
    RECT 319.765 20.16 320.045 21.04 ;
    RECT 316.445 20.16 316.725 21.04 ;
    RECT 313.125 20.16 313.405 21.04 ;
    RECT 309.805 20.16 310.085 21.04 ;
    RECT 306.485 20.16 306.765 21.04 ;
    RECT 303.165 33.84 303.445 34.72 ;
    RECT 372.885 33.84 373.165 34.72 ;
    RECT 369.565 33.84 369.845 34.72 ;
    RECT 299.845 33.84 300.125 34.72 ;
    RECT 296.525 33.84 296.805 34.72 ;
    RECT 293.205 33.84 293.485 34.72 ;
    RECT 289.885 33.84 290.165 34.72 ;
    RECT 286.565 33.84 286.845 34.72 ;
    RECT 283.245 33.84 283.525 34.72 ;
    RECT 279.925 33.84 280.205 34.72 ;
    RECT 276.605 33.84 276.885 34.72 ;
    RECT 273.285 33.84 273.565 34.72 ;
    RECT 269.965 33.84 270.245 34.72 ;
    RECT 233.445 33.84 233.725 34.72 ;
    RECT 230.125 33.84 230.405 34.72 ;
    RECT 366.245 33.84 366.525 34.72 ;
    RECT 226.805 33.84 227.085 34.72 ;
    RECT 362.925 33.84 363.205 34.72 ;
    RECT 223.485 33.84 223.765 34.72 ;
    RECT 359.605 33.84 359.885 34.72 ;
    RECT 220.165 33.84 220.445 34.72 ;
    RECT 356.285 33.84 356.565 34.72 ;
    RECT 352.965 33.84 353.245 34.72 ;
    RECT 216.845 33.84 217.125 34.72 ;
    RECT 349.645 33.84 349.925 34.72 ;
    RECT 213.525 33.84 213.805 34.72 ;
    RECT 346.325 33.84 346.605 34.72 ;
    RECT 210.205 33.84 210.485 34.72 ;
    RECT 343.005 33.84 343.285 34.72 ;
    RECT 206.885 33.84 207.165 34.72 ;
    RECT 339.685 33.84 339.965 34.72 ;
    RECT 203.565 33.84 203.845 34.72 ;
    RECT 336.365 33.84 336.645 34.72 ;
    RECT 266.645 33.84 266.925 34.72 ;
    RECT 263.325 33.84 263.605 34.72 ;
    RECT 260.005 33.84 260.285 34.72 ;
    RECT 256.685 33.84 256.965 34.72 ;
    RECT 253.365 33.84 253.645 34.72 ;
    RECT 250.045 33.84 250.325 34.72 ;
    RECT 246.725 33.84 247.005 34.72 ;
    RECT 243.405 33.84 243.685 34.72 ;
    RECT 240.085 33.84 240.365 34.72 ;
    RECT 236.765 33.84 237.045 34.72 ;
    RECT 333.045 33.84 333.325 34.72 ;
    RECT 329.725 33.84 330.005 34.72 ;
    RECT 326.405 33.84 326.685 34.72 ;
    RECT 323.085 33.84 323.365 34.72 ;
    RECT 319.765 33.84 320.045 34.72 ;
    RECT 316.445 33.84 316.725 34.72 ;
    RECT 313.125 33.84 313.405 34.72 ;
    RECT 309.805 33.84 310.085 34.72 ;
    RECT 306.485 33.84 306.765 34.72 ;
    RECT 303.165 19.44 303.445 20.32 ;
    RECT 372.885 19.44 373.165 20.32 ;
    RECT 369.565 19.44 369.845 20.32 ;
    RECT 299.845 19.44 300.125 20.32 ;
    RECT 296.525 19.44 296.805 20.32 ;
    RECT 293.205 19.44 293.485 20.32 ;
    RECT 289.885 19.44 290.165 20.32 ;
    RECT 286.565 19.44 286.845 20.32 ;
    RECT 283.245 19.44 283.525 20.32 ;
    RECT 279.925 19.44 280.205 20.32 ;
    RECT 276.605 19.44 276.885 20.32 ;
    RECT 273.285 19.44 273.565 20.32 ;
    RECT 269.965 19.44 270.245 20.32 ;
    RECT 233.445 19.44 233.725 20.32 ;
    RECT 230.125 19.44 230.405 20.32 ;
    RECT 366.245 19.44 366.525 20.32 ;
    RECT 226.805 19.44 227.085 20.32 ;
    RECT 362.925 19.44 363.205 20.32 ;
    RECT 223.485 19.44 223.765 20.32 ;
    RECT 359.605 19.44 359.885 20.32 ;
    RECT 220.165 19.44 220.445 20.32 ;
    RECT 356.285 19.44 356.565 20.32 ;
    RECT 352.965 19.44 353.245 20.32 ;
    RECT 216.845 19.44 217.125 20.32 ;
    RECT 349.645 19.44 349.925 20.32 ;
    RECT 213.525 19.44 213.805 20.32 ;
    RECT 346.325 19.44 346.605 20.32 ;
    RECT 210.205 19.44 210.485 20.32 ;
    RECT 343.005 19.44 343.285 20.32 ;
    RECT 206.885 19.44 207.165 20.32 ;
    RECT 339.685 19.44 339.965 20.32 ;
    RECT 203.565 19.44 203.845 20.32 ;
    RECT 336.365 19.44 336.645 20.32 ;
    RECT 266.645 19.44 266.925 20.32 ;
    RECT 263.325 19.44 263.605 20.32 ;
    RECT 260.005 19.44 260.285 20.32 ;
    RECT 256.685 19.44 256.965 20.32 ;
    RECT 253.365 19.44 253.645 20.32 ;
    RECT 250.045 19.44 250.325 20.32 ;
    RECT 246.725 19.44 247.005 20.32 ;
    RECT 243.405 19.44 243.685 20.32 ;
    RECT 240.085 19.44 240.365 20.32 ;
    RECT 236.765 19.44 237.045 20.32 ;
    RECT 333.045 19.44 333.325 20.32 ;
    RECT 329.725 19.44 330.005 20.32 ;
    RECT 326.405 19.44 326.685 20.32 ;
    RECT 323.085 19.44 323.365 20.32 ;
    RECT 319.765 19.44 320.045 20.32 ;
    RECT 316.445 19.44 316.725 20.32 ;
    RECT 313.125 19.44 313.405 20.32 ;
    RECT 309.805 19.44 310.085 20.32 ;
    RECT 306.485 19.44 306.765 20.32 ;
    RECT 303.165 18.72 303.445 19.6 ;
    RECT 372.885 18.72 373.165 19.6 ;
    RECT 369.565 18.72 369.845 19.6 ;
    RECT 299.845 18.72 300.125 19.6 ;
    RECT 296.525 18.72 296.805 19.6 ;
    RECT 293.205 18.72 293.485 19.6 ;
    RECT 289.885 18.72 290.165 19.6 ;
    RECT 286.565 18.72 286.845 19.6 ;
    RECT 283.245 18.72 283.525 19.6 ;
    RECT 279.925 18.72 280.205 19.6 ;
    RECT 276.605 18.72 276.885 19.6 ;
    RECT 273.285 18.72 273.565 19.6 ;
    RECT 269.965 18.72 270.245 19.6 ;
    RECT 233.445 18.72 233.725 19.6 ;
    RECT 230.125 18.72 230.405 19.6 ;
    RECT 366.245 18.72 366.525 19.6 ;
    RECT 226.805 18.72 227.085 19.6 ;
    RECT 362.925 18.72 363.205 19.6 ;
    RECT 223.485 18.72 223.765 19.6 ;
    RECT 359.605 18.72 359.885 19.6 ;
    RECT 220.165 18.72 220.445 19.6 ;
    RECT 356.285 18.72 356.565 19.6 ;
    RECT 352.965 18.72 353.245 19.6 ;
    RECT 216.845 18.72 217.125 19.6 ;
    RECT 349.645 18.72 349.925 19.6 ;
    RECT 213.525 18.72 213.805 19.6 ;
    RECT 346.325 18.72 346.605 19.6 ;
    RECT 210.205 18.72 210.485 19.6 ;
    RECT 343.005 18.72 343.285 19.6 ;
    RECT 206.885 18.72 207.165 19.6 ;
    RECT 339.685 18.72 339.965 19.6 ;
    RECT 203.565 18.72 203.845 19.6 ;
    RECT 336.365 18.72 336.645 19.6 ;
    RECT 266.645 18.72 266.925 19.6 ;
    RECT 263.325 18.72 263.605 19.6 ;
    RECT 260.005 18.72 260.285 19.6 ;
    RECT 256.685 18.72 256.965 19.6 ;
    RECT 253.365 18.72 253.645 19.6 ;
    RECT 250.045 18.72 250.325 19.6 ;
    RECT 246.725 18.72 247.005 19.6 ;
    RECT 243.405 18.72 243.685 19.6 ;
    RECT 240.085 18.72 240.365 19.6 ;
    RECT 236.765 18.72 237.045 19.6 ;
    RECT 333.045 18.72 333.325 19.6 ;
    RECT 329.725 18.72 330.005 19.6 ;
    RECT 326.405 18.72 326.685 19.6 ;
    RECT 323.085 18.72 323.365 19.6 ;
    RECT 319.765 18.72 320.045 19.6 ;
    RECT 316.445 18.72 316.725 19.6 ;
    RECT 313.125 18.72 313.405 19.6 ;
    RECT 309.805 18.72 310.085 19.6 ;
    RECT 306.485 18.72 306.765 19.6 ;
    RECT 233.445 57.68 233.725 58.42 ;
    RECT 230.125 57.68 230.405 58.42 ;
    RECT 226.805 57.68 227.085 58.42 ;
    RECT 223.485 57.68 223.765 58.42 ;
    RECT 220.165 57.68 220.445 58.42 ;
    RECT 216.845 57.68 217.125 58.42 ;
    RECT 213.525 57.68 213.805 58.42 ;
    RECT 210.205 57.68 210.485 58.42 ;
    RECT 206.885 57.68 207.165 58.42 ;
    RECT 203.565 57.68 203.845 58.42 ;
    RECT 372.885 57.68 373.165 58.42 ;
    RECT 369.565 57.68 369.845 58.42 ;
    RECT 366.245 57.68 366.525 58.42 ;
    RECT 362.925 57.68 363.205 58.42 ;
    RECT 359.605 57.68 359.885 58.42 ;
    RECT 356.285 57.68 356.565 58.42 ;
    RECT 352.965 57.68 353.245 58.42 ;
    RECT 349.645 57.68 349.925 58.42 ;
    RECT 346.325 57.68 346.605 58.42 ;
    RECT 343.005 57.68 343.285 58.42 ;
    RECT 339.685 57.68 339.965 58.42 ;
    RECT 336.365 57.68 336.645 58.42 ;
    RECT 333.045 57.68 333.325 58.42 ;
    RECT 329.725 57.68 330.005 58.42 ;
    RECT 326.405 57.68 326.685 58.42 ;
    RECT 323.085 57.68 323.365 58.42 ;
    RECT 319.765 57.68 320.045 58.42 ;
    RECT 316.445 57.68 316.725 58.42 ;
    RECT 313.125 57.68 313.405 58.42 ;
    RECT 309.805 57.68 310.085 58.42 ;
    RECT 306.485 57.68 306.765 58.42 ;
    RECT 303.165 57.68 303.445 58.42 ;
    RECT 299.845 57.68 300.125 58.42 ;
    RECT 296.525 57.68 296.805 58.42 ;
    RECT 293.205 57.68 293.485 58.42 ;
    RECT 289.885 57.68 290.165 58.42 ;
    RECT 286.565 57.68 286.845 58.42 ;
    RECT 283.245 57.68 283.525 58.42 ;
    RECT 279.925 57.68 280.205 58.42 ;
    RECT 276.605 57.68 276.885 58.42 ;
    RECT 273.285 57.68 273.565 58.42 ;
    RECT 269.965 57.68 270.245 58.42 ;
    RECT 266.645 57.68 266.925 58.42 ;
    RECT 263.325 57.68 263.605 58.42 ;
    RECT 260.005 57.68 260.285 58.42 ;
    RECT 256.685 57.68 256.965 58.42 ;
    RECT 253.365 57.68 253.645 58.42 ;
    RECT 250.045 57.68 250.325 58.42 ;
    RECT 246.725 57.68 247.005 58.42 ;
    RECT 243.405 57.68 243.685 58.42 ;
    RECT 240.085 57.68 240.365 58.42 ;
    RECT 236.765 57.68 237.045 58.42 ;
    RECT 303.165 56.88 303.445 57.76 ;
    RECT 372.885 56.88 373.165 57.76 ;
    RECT 369.565 56.88 369.845 57.76 ;
    RECT 299.845 56.88 300.125 57.76 ;
    RECT 296.525 56.88 296.805 57.76 ;
    RECT 293.205 56.88 293.485 57.76 ;
    RECT 289.885 56.88 290.165 57.76 ;
    RECT 286.565 56.88 286.845 57.76 ;
    RECT 283.245 56.88 283.525 57.76 ;
    RECT 279.925 56.88 280.205 57.76 ;
    RECT 276.605 56.88 276.885 57.76 ;
    RECT 273.285 56.88 273.565 57.76 ;
    RECT 269.965 56.88 270.245 57.76 ;
    RECT 233.445 56.88 233.725 57.76 ;
    RECT 230.125 56.88 230.405 57.76 ;
    RECT 366.245 56.88 366.525 57.76 ;
    RECT 226.805 56.88 227.085 57.76 ;
    RECT 362.925 56.88 363.205 57.76 ;
    RECT 223.485 56.88 223.765 57.76 ;
    RECT 359.605 56.88 359.885 57.76 ;
    RECT 220.165 56.88 220.445 57.76 ;
    RECT 356.285 56.88 356.565 57.76 ;
    RECT 352.965 56.88 353.245 57.76 ;
    RECT 216.845 56.88 217.125 57.76 ;
    RECT 349.645 56.88 349.925 57.76 ;
    RECT 213.525 56.88 213.805 57.76 ;
    RECT 346.325 56.88 346.605 57.76 ;
    RECT 210.205 56.88 210.485 57.76 ;
    RECT 343.005 56.88 343.285 57.76 ;
    RECT 206.885 56.88 207.165 57.76 ;
    RECT 339.685 56.88 339.965 57.76 ;
    RECT 203.565 56.88 203.845 57.76 ;
    RECT 336.365 56.88 336.645 57.76 ;
    RECT 266.645 56.88 266.925 57.76 ;
    RECT 263.325 56.88 263.605 57.76 ;
    RECT 260.005 56.88 260.285 57.76 ;
    RECT 256.685 56.88 256.965 57.76 ;
    RECT 253.365 56.88 253.645 57.76 ;
    RECT 250.045 56.88 250.325 57.76 ;
    RECT 246.725 56.88 247.005 57.76 ;
    RECT 243.405 56.88 243.685 57.76 ;
    RECT 240.085 56.88 240.365 57.76 ;
    RECT 236.765 56.88 237.045 57.76 ;
    RECT 333.045 56.88 333.325 57.76 ;
    RECT 329.725 56.88 330.005 57.76 ;
    RECT 326.405 56.88 326.685 57.76 ;
    RECT 323.085 56.88 323.365 57.76 ;
    RECT 319.765 56.88 320.045 57.76 ;
    RECT 316.445 56.88 316.725 57.76 ;
    RECT 313.125 56.88 313.405 57.76 ;
    RECT 309.805 56.88 310.085 57.76 ;
    RECT 306.485 56.88 306.765 57.76 ;
    RECT 303.165 56.16 303.445 57.04 ;
    RECT 372.885 56.16 373.165 57.04 ;
    RECT 369.565 56.16 369.845 57.04 ;
    RECT 299.845 56.16 300.125 57.04 ;
    RECT 296.525 56.16 296.805 57.04 ;
    RECT 293.205 56.16 293.485 57.04 ;
    RECT 289.885 56.16 290.165 57.04 ;
    RECT 286.565 56.16 286.845 57.04 ;
    RECT 283.245 56.16 283.525 57.04 ;
    RECT 279.925 56.16 280.205 57.04 ;
    RECT 276.605 56.16 276.885 57.04 ;
    RECT 273.285 56.16 273.565 57.04 ;
    RECT 269.965 56.16 270.245 57.04 ;
    RECT 233.445 56.16 233.725 57.04 ;
    RECT 230.125 56.16 230.405 57.04 ;
    RECT 366.245 56.16 366.525 57.04 ;
    RECT 226.805 56.16 227.085 57.04 ;
    RECT 362.925 56.16 363.205 57.04 ;
    RECT 223.485 56.16 223.765 57.04 ;
    RECT 359.605 56.16 359.885 57.04 ;
    RECT 220.165 56.16 220.445 57.04 ;
    RECT 356.285 56.16 356.565 57.04 ;
    RECT 352.965 56.16 353.245 57.04 ;
    RECT 216.845 56.16 217.125 57.04 ;
    RECT 349.645 56.16 349.925 57.04 ;
    RECT 213.525 56.16 213.805 57.04 ;
    RECT 346.325 56.16 346.605 57.04 ;
    RECT 210.205 56.16 210.485 57.04 ;
    RECT 343.005 56.16 343.285 57.04 ;
    RECT 206.885 56.16 207.165 57.04 ;
    RECT 339.685 56.16 339.965 57.04 ;
    RECT 203.565 56.16 203.845 57.04 ;
    RECT 336.365 56.16 336.645 57.04 ;
    RECT 266.645 56.16 266.925 57.04 ;
    RECT 263.325 56.16 263.605 57.04 ;
    RECT 260.005 56.16 260.285 57.04 ;
    RECT 256.685 56.16 256.965 57.04 ;
    RECT 253.365 56.16 253.645 57.04 ;
    RECT 250.045 56.16 250.325 57.04 ;
    RECT 246.725 56.16 247.005 57.04 ;
    RECT 243.405 56.16 243.685 57.04 ;
    RECT 240.085 56.16 240.365 57.04 ;
    RECT 236.765 56.16 237.045 57.04 ;
    RECT 333.045 56.16 333.325 57.04 ;
    RECT 329.725 56.16 330.005 57.04 ;
    RECT 326.405 56.16 326.685 57.04 ;
    RECT 323.085 56.16 323.365 57.04 ;
    RECT 319.765 56.16 320.045 57.04 ;
    RECT 316.445 56.16 316.725 57.04 ;
    RECT 313.125 56.16 313.405 57.04 ;
    RECT 309.805 56.16 310.085 57.04 ;
    RECT 306.485 56.16 306.765 57.04 ;
    RECT 303.165 55.44 303.445 56.32 ;
    RECT 372.885 55.44 373.165 56.32 ;
    RECT 369.565 55.44 369.845 56.32 ;
    RECT 299.845 55.44 300.125 56.32 ;
    RECT 296.525 55.44 296.805 56.32 ;
    RECT 293.205 55.44 293.485 56.32 ;
    RECT 289.885 55.44 290.165 56.32 ;
    RECT 286.565 55.44 286.845 56.32 ;
    RECT 283.245 55.44 283.525 56.32 ;
    RECT 279.925 55.44 280.205 56.32 ;
    RECT 276.605 55.44 276.885 56.32 ;
    RECT 273.285 55.44 273.565 56.32 ;
    RECT 269.965 55.44 270.245 56.32 ;
    RECT 233.445 55.44 233.725 56.32 ;
    RECT 230.125 55.44 230.405 56.32 ;
    RECT 366.245 55.44 366.525 56.32 ;
    RECT 226.805 55.44 227.085 56.32 ;
    RECT 362.925 55.44 363.205 56.32 ;
    RECT 223.485 55.44 223.765 56.32 ;
    RECT 359.605 55.44 359.885 56.32 ;
    RECT 220.165 55.44 220.445 56.32 ;
    RECT 356.285 55.44 356.565 56.32 ;
    RECT 352.965 55.44 353.245 56.32 ;
    RECT 216.845 55.44 217.125 56.32 ;
    RECT 349.645 55.44 349.925 56.32 ;
    RECT 213.525 55.44 213.805 56.32 ;
    RECT 346.325 55.44 346.605 56.32 ;
    RECT 210.205 55.44 210.485 56.32 ;
    RECT 343.005 55.44 343.285 56.32 ;
    RECT 206.885 55.44 207.165 56.32 ;
    RECT 339.685 55.44 339.965 56.32 ;
    RECT 203.565 55.44 203.845 56.32 ;
    RECT 336.365 55.44 336.645 56.32 ;
    RECT 266.645 55.44 266.925 56.32 ;
    RECT 263.325 55.44 263.605 56.32 ;
    RECT 260.005 55.44 260.285 56.32 ;
    RECT 256.685 55.44 256.965 56.32 ;
    RECT 253.365 55.44 253.645 56.32 ;
    RECT 250.045 55.44 250.325 56.32 ;
    RECT 246.725 55.44 247.005 56.32 ;
    RECT 243.405 55.44 243.685 56.32 ;
    RECT 240.085 55.44 240.365 56.32 ;
    RECT 236.765 55.44 237.045 56.32 ;
    RECT 333.045 55.44 333.325 56.32 ;
    RECT 329.725 55.44 330.005 56.32 ;
    RECT 326.405 55.44 326.685 56.32 ;
    RECT 323.085 55.44 323.365 56.32 ;
    RECT 319.765 55.44 320.045 56.32 ;
    RECT 316.445 55.44 316.725 56.32 ;
    RECT 313.125 55.44 313.405 56.32 ;
    RECT 309.805 55.44 310.085 56.32 ;
    RECT 306.485 55.44 306.765 56.32 ;
    RECT 303.165 54.72 303.445 55.6 ;
    RECT 372.885 54.72 373.165 55.6 ;
    RECT 369.565 54.72 369.845 55.6 ;
    RECT 299.845 54.72 300.125 55.6 ;
    RECT 296.525 54.72 296.805 55.6 ;
    RECT 293.205 54.72 293.485 55.6 ;
    RECT 289.885 54.72 290.165 55.6 ;
    RECT 286.565 54.72 286.845 55.6 ;
    RECT 283.245 54.72 283.525 55.6 ;
    RECT 279.925 54.72 280.205 55.6 ;
    RECT 276.605 54.72 276.885 55.6 ;
    RECT 273.285 54.72 273.565 55.6 ;
    RECT 269.965 54.72 270.245 55.6 ;
    RECT 233.445 54.72 233.725 55.6 ;
    RECT 230.125 54.72 230.405 55.6 ;
    RECT 366.245 54.72 366.525 55.6 ;
    RECT 226.805 54.72 227.085 55.6 ;
    RECT 362.925 54.72 363.205 55.6 ;
    RECT 223.485 54.72 223.765 55.6 ;
    RECT 359.605 54.72 359.885 55.6 ;
    RECT 220.165 54.72 220.445 55.6 ;
    RECT 356.285 54.72 356.565 55.6 ;
    RECT 352.965 54.72 353.245 55.6 ;
    RECT 216.845 54.72 217.125 55.6 ;
    RECT 349.645 54.72 349.925 55.6 ;
    RECT 213.525 54.72 213.805 55.6 ;
    RECT 346.325 54.72 346.605 55.6 ;
    RECT 210.205 54.72 210.485 55.6 ;
    RECT 343.005 54.72 343.285 55.6 ;
    RECT 206.885 54.72 207.165 55.6 ;
    RECT 339.685 54.72 339.965 55.6 ;
    RECT 203.565 54.72 203.845 55.6 ;
    RECT 336.365 54.72 336.645 55.6 ;
    RECT 266.645 54.72 266.925 55.6 ;
    RECT 263.325 54.72 263.605 55.6 ;
    RECT 260.005 54.72 260.285 55.6 ;
    RECT 256.685 54.72 256.965 55.6 ;
    RECT 253.365 54.72 253.645 55.6 ;
    RECT 250.045 54.72 250.325 55.6 ;
    RECT 246.725 54.72 247.005 55.6 ;
    RECT 243.405 54.72 243.685 55.6 ;
    RECT 240.085 54.72 240.365 55.6 ;
    RECT 236.765 54.72 237.045 55.6 ;
    RECT 333.045 54.72 333.325 55.6 ;
    RECT 329.725 54.72 330.005 55.6 ;
    RECT 326.405 54.72 326.685 55.6 ;
    RECT 323.085 54.72 323.365 55.6 ;
    RECT 319.765 54.72 320.045 55.6 ;
    RECT 316.445 54.72 316.725 55.6 ;
    RECT 313.125 54.72 313.405 55.6 ;
    RECT 309.805 54.72 310.085 55.6 ;
    RECT 306.485 54.72 306.765 55.6 ;
    RECT 303.165 54.0 303.445 54.88 ;
    RECT 372.885 54.0 373.165 54.88 ;
    RECT 369.565 54.0 369.845 54.88 ;
    RECT 299.845 54.0 300.125 54.88 ;
    RECT 296.525 54.0 296.805 54.88 ;
    RECT 293.205 54.0 293.485 54.88 ;
    RECT 289.885 54.0 290.165 54.88 ;
    RECT 286.565 54.0 286.845 54.88 ;
    RECT 283.245 54.0 283.525 54.88 ;
    RECT 279.925 54.0 280.205 54.88 ;
    RECT 276.605 54.0 276.885 54.88 ;
    RECT 273.285 54.0 273.565 54.88 ;
    RECT 269.965 54.0 270.245 54.88 ;
    RECT 233.445 54.0 233.725 54.88 ;
    RECT 230.125 54.0 230.405 54.88 ;
    RECT 366.245 54.0 366.525 54.88 ;
    RECT 226.805 54.0 227.085 54.88 ;
    RECT 362.925 54.0 363.205 54.88 ;
    RECT 223.485 54.0 223.765 54.88 ;
    RECT 359.605 54.0 359.885 54.88 ;
    RECT 220.165 54.0 220.445 54.88 ;
    RECT 356.285 54.0 356.565 54.88 ;
    RECT 352.965 54.0 353.245 54.88 ;
    RECT 216.845 54.0 217.125 54.88 ;
    RECT 349.645 54.0 349.925 54.88 ;
    RECT 213.525 54.0 213.805 54.88 ;
    RECT 346.325 54.0 346.605 54.88 ;
    RECT 210.205 54.0 210.485 54.88 ;
    RECT 343.005 54.0 343.285 54.88 ;
    RECT 206.885 54.0 207.165 54.88 ;
    RECT 339.685 54.0 339.965 54.88 ;
    RECT 203.565 54.0 203.845 54.88 ;
    RECT 336.365 54.0 336.645 54.88 ;
    RECT 266.645 54.0 266.925 54.88 ;
    RECT 263.325 54.0 263.605 54.88 ;
    RECT 260.005 54.0 260.285 54.88 ;
    RECT 256.685 54.0 256.965 54.88 ;
    RECT 253.365 54.0 253.645 54.88 ;
    RECT 250.045 54.0 250.325 54.88 ;
    RECT 246.725 54.0 247.005 54.88 ;
    RECT 243.405 54.0 243.685 54.88 ;
    RECT 240.085 54.0 240.365 54.88 ;
    RECT 236.765 54.0 237.045 54.88 ;
    RECT 333.045 54.0 333.325 54.88 ;
    RECT 329.725 54.0 330.005 54.88 ;
    RECT 326.405 54.0 326.685 54.88 ;
    RECT 323.085 54.0 323.365 54.88 ;
    RECT 319.765 54.0 320.045 54.88 ;
    RECT 316.445 54.0 316.725 54.88 ;
    RECT 313.125 54.0 313.405 54.88 ;
    RECT 309.805 54.0 310.085 54.88 ;
    RECT 306.485 54.0 306.765 54.88 ;
    RECT 303.165 53.28 303.445 54.16 ;
    RECT 372.885 53.28 373.165 54.16 ;
    RECT 369.565 53.28 369.845 54.16 ;
    RECT 299.845 53.28 300.125 54.16 ;
    RECT 296.525 53.28 296.805 54.16 ;
    RECT 293.205 53.28 293.485 54.16 ;
    RECT 289.885 53.28 290.165 54.16 ;
    RECT 286.565 53.28 286.845 54.16 ;
    RECT 283.245 53.28 283.525 54.16 ;
    RECT 279.925 53.28 280.205 54.16 ;
    RECT 276.605 53.28 276.885 54.16 ;
    RECT 273.285 53.28 273.565 54.16 ;
    RECT 269.965 53.28 270.245 54.16 ;
    RECT 233.445 53.28 233.725 54.16 ;
    RECT 230.125 53.28 230.405 54.16 ;
    RECT 366.245 53.28 366.525 54.16 ;
    RECT 226.805 53.28 227.085 54.16 ;
    RECT 362.925 53.28 363.205 54.16 ;
    RECT 223.485 53.28 223.765 54.16 ;
    RECT 359.605 53.28 359.885 54.16 ;
    RECT 220.165 53.28 220.445 54.16 ;
    RECT 356.285 53.28 356.565 54.16 ;
    RECT 352.965 53.28 353.245 54.16 ;
    RECT 216.845 53.28 217.125 54.16 ;
    RECT 349.645 53.28 349.925 54.16 ;
    RECT 213.525 53.28 213.805 54.16 ;
    RECT 346.325 53.28 346.605 54.16 ;
    RECT 210.205 53.28 210.485 54.16 ;
    RECT 343.005 53.28 343.285 54.16 ;
    RECT 206.885 53.28 207.165 54.16 ;
    RECT 339.685 53.28 339.965 54.16 ;
    RECT 203.565 53.28 203.845 54.16 ;
    RECT 336.365 53.28 336.645 54.16 ;
    RECT 266.645 53.28 266.925 54.16 ;
    RECT 263.325 53.28 263.605 54.16 ;
    RECT 260.005 53.28 260.285 54.16 ;
    RECT 256.685 53.28 256.965 54.16 ;
    RECT 253.365 53.28 253.645 54.16 ;
    RECT 250.045 53.28 250.325 54.16 ;
    RECT 246.725 53.28 247.005 54.16 ;
    RECT 243.405 53.28 243.685 54.16 ;
    RECT 240.085 53.28 240.365 54.16 ;
    RECT 236.765 53.28 237.045 54.16 ;
    RECT 333.045 53.28 333.325 54.16 ;
    RECT 329.725 53.28 330.005 54.16 ;
    RECT 326.405 53.28 326.685 54.16 ;
    RECT 323.085 53.28 323.365 54.16 ;
    RECT 319.765 53.28 320.045 54.16 ;
    RECT 316.445 53.28 316.725 54.16 ;
    RECT 313.125 53.28 313.405 54.16 ;
    RECT 309.805 53.28 310.085 54.16 ;
    RECT 306.485 53.28 306.765 54.16 ;
    RECT 303.165 52.56 303.445 53.44 ;
    RECT 372.885 52.56 373.165 53.44 ;
    RECT 369.565 52.56 369.845 53.44 ;
    RECT 299.845 52.56 300.125 53.44 ;
    RECT 296.525 52.56 296.805 53.44 ;
    RECT 293.205 52.56 293.485 53.44 ;
    RECT 289.885 52.56 290.165 53.44 ;
    RECT 286.565 52.56 286.845 53.44 ;
    RECT 283.245 52.56 283.525 53.44 ;
    RECT 279.925 52.56 280.205 53.44 ;
    RECT 276.605 52.56 276.885 53.44 ;
    RECT 273.285 52.56 273.565 53.44 ;
    RECT 269.965 52.56 270.245 53.44 ;
    RECT 233.445 52.56 233.725 53.44 ;
    RECT 230.125 52.56 230.405 53.44 ;
    RECT 366.245 52.56 366.525 53.44 ;
    RECT 226.805 52.56 227.085 53.44 ;
    RECT 362.925 52.56 363.205 53.44 ;
    RECT 223.485 52.56 223.765 53.44 ;
    RECT 359.605 52.56 359.885 53.44 ;
    RECT 220.165 52.56 220.445 53.44 ;
    RECT 356.285 52.56 356.565 53.44 ;
    RECT 352.965 52.56 353.245 53.44 ;
    RECT 216.845 52.56 217.125 53.44 ;
    RECT 349.645 52.56 349.925 53.44 ;
    RECT 213.525 52.56 213.805 53.44 ;
    RECT 346.325 52.56 346.605 53.44 ;
    RECT 210.205 52.56 210.485 53.44 ;
    RECT 343.005 52.56 343.285 53.44 ;
    RECT 206.885 52.56 207.165 53.44 ;
    RECT 339.685 52.56 339.965 53.44 ;
    RECT 203.565 52.56 203.845 53.44 ;
    RECT 336.365 52.56 336.645 53.44 ;
    RECT 266.645 52.56 266.925 53.44 ;
    RECT 263.325 52.56 263.605 53.44 ;
    RECT 260.005 52.56 260.285 53.44 ;
    RECT 256.685 52.56 256.965 53.44 ;
    RECT 253.365 52.56 253.645 53.44 ;
    RECT 250.045 52.56 250.325 53.44 ;
    RECT 246.725 52.56 247.005 53.44 ;
    RECT 243.405 52.56 243.685 53.44 ;
    RECT 240.085 52.56 240.365 53.44 ;
    RECT 236.765 52.56 237.045 53.44 ;
    RECT 333.045 52.56 333.325 53.44 ;
    RECT 329.725 52.56 330.005 53.44 ;
    RECT 326.405 52.56 326.685 53.44 ;
    RECT 323.085 52.56 323.365 53.44 ;
    RECT 319.765 52.56 320.045 53.44 ;
    RECT 316.445 52.56 316.725 53.44 ;
    RECT 313.125 52.56 313.405 53.44 ;
    RECT 309.805 52.56 310.085 53.44 ;
    RECT 306.485 52.56 306.765 53.44 ;
    RECT 303.165 51.84 303.445 52.72 ;
    RECT 372.885 51.84 373.165 52.72 ;
    RECT 369.565 51.84 369.845 52.72 ;
    RECT 299.845 51.84 300.125 52.72 ;
    RECT 296.525 51.84 296.805 52.72 ;
    RECT 293.205 51.84 293.485 52.72 ;
    RECT 289.885 51.84 290.165 52.72 ;
    RECT 286.565 51.84 286.845 52.72 ;
    RECT 283.245 51.84 283.525 52.72 ;
    RECT 279.925 51.84 280.205 52.72 ;
    RECT 276.605 51.84 276.885 52.72 ;
    RECT 273.285 51.84 273.565 52.72 ;
    RECT 269.965 51.84 270.245 52.72 ;
    RECT 233.445 51.84 233.725 52.72 ;
    RECT 230.125 51.84 230.405 52.72 ;
    RECT 366.245 51.84 366.525 52.72 ;
    RECT 226.805 51.84 227.085 52.72 ;
    RECT 362.925 51.84 363.205 52.72 ;
    RECT 223.485 51.84 223.765 52.72 ;
    RECT 359.605 51.84 359.885 52.72 ;
    RECT 220.165 51.84 220.445 52.72 ;
    RECT 356.285 51.84 356.565 52.72 ;
    RECT 352.965 51.84 353.245 52.72 ;
    RECT 216.845 51.84 217.125 52.72 ;
    RECT 349.645 51.84 349.925 52.72 ;
    RECT 213.525 51.84 213.805 52.72 ;
    RECT 346.325 51.84 346.605 52.72 ;
    RECT 210.205 51.84 210.485 52.72 ;
    RECT 343.005 51.84 343.285 52.72 ;
    RECT 206.885 51.84 207.165 52.72 ;
    RECT 339.685 51.84 339.965 52.72 ;
    RECT 203.565 51.84 203.845 52.72 ;
    RECT 336.365 51.84 336.645 52.72 ;
    RECT 266.645 51.84 266.925 52.72 ;
    RECT 263.325 51.84 263.605 52.72 ;
    RECT 260.005 51.84 260.285 52.72 ;
    RECT 256.685 51.84 256.965 52.72 ;
    RECT 253.365 51.84 253.645 52.72 ;
    RECT 250.045 51.84 250.325 52.72 ;
    RECT 246.725 51.84 247.005 52.72 ;
    RECT 243.405 51.84 243.685 52.72 ;
    RECT 240.085 51.84 240.365 52.72 ;
    RECT 236.765 51.84 237.045 52.72 ;
    RECT 333.045 51.84 333.325 52.72 ;
    RECT 329.725 51.84 330.005 52.72 ;
    RECT 326.405 51.84 326.685 52.72 ;
    RECT 323.085 51.84 323.365 52.72 ;
    RECT 319.765 51.84 320.045 52.72 ;
    RECT 316.445 51.84 316.725 52.72 ;
    RECT 313.125 51.84 313.405 52.72 ;
    RECT 309.805 51.84 310.085 52.72 ;
    RECT 306.485 51.84 306.765 52.72 ;
    RECT 303.165 51.12 303.445 52.0 ;
    RECT 372.885 51.12 373.165 52.0 ;
    RECT 369.565 51.12 369.845 52.0 ;
    RECT 299.845 51.12 300.125 52.0 ;
    RECT 296.525 51.12 296.805 52.0 ;
    RECT 293.205 51.12 293.485 52.0 ;
    RECT 289.885 51.12 290.165 52.0 ;
    RECT 286.565 51.12 286.845 52.0 ;
    RECT 283.245 51.12 283.525 52.0 ;
    RECT 279.925 51.12 280.205 52.0 ;
    RECT 276.605 51.12 276.885 52.0 ;
    RECT 273.285 51.12 273.565 52.0 ;
    RECT 269.965 51.12 270.245 52.0 ;
    RECT 233.445 51.12 233.725 52.0 ;
    RECT 230.125 51.12 230.405 52.0 ;
    RECT 366.245 51.12 366.525 52.0 ;
    RECT 226.805 51.12 227.085 52.0 ;
    RECT 362.925 51.12 363.205 52.0 ;
    RECT 223.485 51.12 223.765 52.0 ;
    RECT 359.605 51.12 359.885 52.0 ;
    RECT 220.165 51.12 220.445 52.0 ;
    RECT 356.285 51.12 356.565 52.0 ;
    RECT 352.965 51.12 353.245 52.0 ;
    RECT 216.845 51.12 217.125 52.0 ;
    RECT 349.645 51.12 349.925 52.0 ;
    RECT 213.525 51.12 213.805 52.0 ;
    RECT 346.325 51.12 346.605 52.0 ;
    RECT 210.205 51.12 210.485 52.0 ;
    RECT 343.005 51.12 343.285 52.0 ;
    RECT 206.885 51.12 207.165 52.0 ;
    RECT 339.685 51.12 339.965 52.0 ;
    RECT 203.565 51.12 203.845 52.0 ;
    RECT 336.365 51.12 336.645 52.0 ;
    RECT 266.645 51.12 266.925 52.0 ;
    RECT 263.325 51.12 263.605 52.0 ;
    RECT 260.005 51.12 260.285 52.0 ;
    RECT 256.685 51.12 256.965 52.0 ;
    RECT 253.365 51.12 253.645 52.0 ;
    RECT 250.045 51.12 250.325 52.0 ;
    RECT 246.725 51.12 247.005 52.0 ;
    RECT 243.405 51.12 243.685 52.0 ;
    RECT 240.085 51.12 240.365 52.0 ;
    RECT 236.765 51.12 237.045 52.0 ;
    RECT 333.045 51.12 333.325 52.0 ;
    RECT 329.725 51.12 330.005 52.0 ;
    RECT 326.405 51.12 326.685 52.0 ;
    RECT 323.085 51.12 323.365 52.0 ;
    RECT 319.765 51.12 320.045 52.0 ;
    RECT 316.445 51.12 316.725 52.0 ;
    RECT 313.125 51.12 313.405 52.0 ;
    RECT 309.805 51.12 310.085 52.0 ;
    RECT 306.485 51.12 306.765 52.0 ;
    RECT 303.165 50.4 303.445 51.28 ;
    RECT 372.885 50.4 373.165 51.28 ;
    RECT 369.565 50.4 369.845 51.28 ;
    RECT 299.845 50.4 300.125 51.28 ;
    RECT 296.525 50.4 296.805 51.28 ;
    RECT 293.205 50.4 293.485 51.28 ;
    RECT 289.885 50.4 290.165 51.28 ;
    RECT 286.565 50.4 286.845 51.28 ;
    RECT 283.245 50.4 283.525 51.28 ;
    RECT 279.925 50.4 280.205 51.28 ;
    RECT 276.605 50.4 276.885 51.28 ;
    RECT 273.285 50.4 273.565 51.28 ;
    RECT 269.965 50.4 270.245 51.28 ;
    RECT 233.445 50.4 233.725 51.28 ;
    RECT 230.125 50.4 230.405 51.28 ;
    RECT 366.245 50.4 366.525 51.28 ;
    RECT 226.805 50.4 227.085 51.28 ;
    RECT 362.925 50.4 363.205 51.28 ;
    RECT 223.485 50.4 223.765 51.28 ;
    RECT 359.605 50.4 359.885 51.28 ;
    RECT 220.165 50.4 220.445 51.28 ;
    RECT 356.285 50.4 356.565 51.28 ;
    RECT 352.965 50.4 353.245 51.28 ;
    RECT 216.845 50.4 217.125 51.28 ;
    RECT 349.645 50.4 349.925 51.28 ;
    RECT 213.525 50.4 213.805 51.28 ;
    RECT 346.325 50.4 346.605 51.28 ;
    RECT 210.205 50.4 210.485 51.28 ;
    RECT 343.005 50.4 343.285 51.28 ;
    RECT 206.885 50.4 207.165 51.28 ;
    RECT 339.685 50.4 339.965 51.28 ;
    RECT 203.565 50.4 203.845 51.28 ;
    RECT 336.365 50.4 336.645 51.28 ;
    RECT 266.645 50.4 266.925 51.28 ;
    RECT 263.325 50.4 263.605 51.28 ;
    RECT 260.005 50.4 260.285 51.28 ;
    RECT 256.685 50.4 256.965 51.28 ;
    RECT 253.365 50.4 253.645 51.28 ;
    RECT 250.045 50.4 250.325 51.28 ;
    RECT 246.725 50.4 247.005 51.28 ;
    RECT 243.405 50.4 243.685 51.28 ;
    RECT 240.085 50.4 240.365 51.28 ;
    RECT 236.765 50.4 237.045 51.28 ;
    RECT 333.045 50.4 333.325 51.28 ;
    RECT 329.725 50.4 330.005 51.28 ;
    RECT 326.405 50.4 326.685 51.28 ;
    RECT 323.085 50.4 323.365 51.28 ;
    RECT 319.765 50.4 320.045 51.28 ;
    RECT 316.445 50.4 316.725 51.28 ;
    RECT 313.125 50.4 313.405 51.28 ;
    RECT 309.805 50.4 310.085 51.28 ;
    RECT 306.485 50.4 306.765 51.28 ;
    RECT 303.165 11.52 303.445 12.4 ;
    RECT 369.565 11.52 369.845 12.4 ;
    RECT 299.845 11.52 300.125 12.4 ;
    RECT 296.525 11.52 296.805 12.4 ;
    RECT 293.205 11.52 293.485 12.4 ;
    RECT 289.885 11.52 290.165 12.4 ;
    RECT 286.565 11.52 286.845 12.4 ;
    RECT 283.245 11.52 283.525 12.4 ;
    RECT 279.925 11.52 280.205 12.4 ;
    RECT 276.605 11.52 276.885 12.4 ;
    RECT 273.285 11.52 273.565 12.4 ;
    RECT 269.965 11.52 270.245 12.4 ;
    RECT 233.445 11.52 233.725 12.4 ;
    RECT 230.125 11.52 230.405 12.4 ;
    RECT 366.245 11.52 366.525 12.4 ;
    RECT 226.805 11.52 227.085 12.4 ;
    RECT 362.925 11.52 363.205 12.4 ;
    RECT 223.485 11.52 223.765 12.4 ;
    RECT 359.605 11.52 359.885 12.4 ;
    RECT 220.165 11.52 220.445 12.4 ;
    RECT 356.285 11.52 356.565 12.4 ;
    RECT 352.965 11.52 353.245 12.4 ;
    RECT 216.845 11.52 217.125 12.4 ;
    RECT 349.645 11.52 349.925 12.4 ;
    RECT 213.525 11.52 213.805 12.4 ;
    RECT 346.325 11.52 346.605 12.4 ;
    RECT 210.205 11.52 210.485 12.4 ;
    RECT 343.005 11.52 343.285 12.4 ;
    RECT 206.885 11.52 207.165 12.4 ;
    RECT 339.685 11.52 339.965 12.4 ;
    RECT 336.365 11.52 336.645 12.4 ;
    RECT 266.645 11.52 266.925 12.4 ;
    RECT 263.325 11.52 263.605 12.4 ;
    RECT 372.885 11.52 373.165 12.4 ;
    RECT 260.005 11.52 260.285 12.4 ;
    RECT 256.685 11.52 256.965 12.4 ;
    RECT 253.365 11.52 253.645 12.4 ;
    RECT 250.045 11.52 250.325 12.4 ;
    RECT 246.725 11.52 247.005 12.4 ;
    RECT 243.405 11.52 243.685 12.4 ;
    RECT 203.565 11.52 203.845 12.4 ;
    RECT 240.085 11.52 240.365 12.4 ;
    RECT 236.765 11.52 237.045 12.4 ;
    RECT 333.045 11.52 333.325 12.4 ;
    RECT 329.725 11.52 330.005 12.4 ;
    RECT 326.405 11.52 326.685 12.4 ;
    RECT 323.085 11.52 323.365 12.4 ;
    RECT 319.765 11.52 320.045 12.4 ;
    RECT 316.445 11.52 316.725 12.4 ;
    RECT 313.125 11.52 313.405 12.4 ;
    RECT 309.805 11.52 310.085 12.4 ;
    RECT 306.485 11.52 306.765 12.4 ;
    RECT 303.165 49.68 303.445 50.56 ;
    RECT 372.885 49.68 373.165 50.56 ;
    RECT 369.565 49.68 369.845 50.56 ;
    RECT 299.845 49.68 300.125 50.56 ;
    RECT 296.525 49.68 296.805 50.56 ;
    RECT 293.205 49.68 293.485 50.56 ;
    RECT 289.885 49.68 290.165 50.56 ;
    RECT 286.565 49.68 286.845 50.56 ;
    RECT 283.245 49.68 283.525 50.56 ;
    RECT 279.925 49.68 280.205 50.56 ;
    RECT 276.605 49.68 276.885 50.56 ;
    RECT 273.285 49.68 273.565 50.56 ;
    RECT 269.965 49.68 270.245 50.56 ;
    RECT 233.445 49.68 233.725 50.56 ;
    RECT 230.125 49.68 230.405 50.56 ;
    RECT 366.245 49.68 366.525 50.56 ;
    RECT 226.805 49.68 227.085 50.56 ;
    RECT 362.925 49.68 363.205 50.56 ;
    RECT 223.485 49.68 223.765 50.56 ;
    RECT 359.605 49.68 359.885 50.56 ;
    RECT 220.165 49.68 220.445 50.56 ;
    RECT 356.285 49.68 356.565 50.56 ;
    RECT 352.965 49.68 353.245 50.56 ;
    RECT 216.845 49.68 217.125 50.56 ;
    RECT 349.645 49.68 349.925 50.56 ;
    RECT 213.525 49.68 213.805 50.56 ;
    RECT 346.325 49.68 346.605 50.56 ;
    RECT 210.205 49.68 210.485 50.56 ;
    RECT 343.005 49.68 343.285 50.56 ;
    RECT 206.885 49.68 207.165 50.56 ;
    RECT 339.685 49.68 339.965 50.56 ;
    RECT 203.565 49.68 203.845 50.56 ;
    RECT 336.365 49.68 336.645 50.56 ;
    RECT 266.645 49.68 266.925 50.56 ;
    RECT 263.325 49.68 263.605 50.56 ;
    RECT 260.005 49.68 260.285 50.56 ;
    RECT 256.685 49.68 256.965 50.56 ;
    RECT 253.365 49.68 253.645 50.56 ;
    RECT 250.045 49.68 250.325 50.56 ;
    RECT 246.725 49.68 247.005 50.56 ;
    RECT 243.405 49.68 243.685 50.56 ;
    RECT 240.085 49.68 240.365 50.56 ;
    RECT 236.765 49.68 237.045 50.56 ;
    RECT 333.045 49.68 333.325 50.56 ;
    RECT 329.725 49.68 330.005 50.56 ;
    RECT 326.405 49.68 326.685 50.56 ;
    RECT 323.085 49.68 323.365 50.56 ;
    RECT 319.765 49.68 320.045 50.56 ;
    RECT 316.445 49.68 316.725 50.56 ;
    RECT 313.125 49.68 313.405 50.56 ;
    RECT 309.805 49.68 310.085 50.56 ;
    RECT 306.485 49.68 306.765 50.56 ;
    RECT 303.165 48.96 303.445 49.84 ;
    RECT 372.885 48.96 373.165 49.84 ;
    RECT 369.565 48.96 369.845 49.84 ;
    RECT 299.845 48.96 300.125 49.84 ;
    RECT 296.525 48.96 296.805 49.84 ;
    RECT 293.205 48.96 293.485 49.84 ;
    RECT 289.885 48.96 290.165 49.84 ;
    RECT 286.565 48.96 286.845 49.84 ;
    RECT 283.245 48.96 283.525 49.84 ;
    RECT 279.925 48.96 280.205 49.84 ;
    RECT 276.605 48.96 276.885 49.84 ;
    RECT 273.285 48.96 273.565 49.84 ;
    RECT 269.965 48.96 270.245 49.84 ;
    RECT 233.445 48.96 233.725 49.84 ;
    RECT 230.125 48.96 230.405 49.84 ;
    RECT 366.245 48.96 366.525 49.84 ;
    RECT 226.805 48.96 227.085 49.84 ;
    RECT 362.925 48.96 363.205 49.84 ;
    RECT 223.485 48.96 223.765 49.84 ;
    RECT 359.605 48.96 359.885 49.84 ;
    RECT 220.165 48.96 220.445 49.84 ;
    RECT 356.285 48.96 356.565 49.84 ;
    RECT 352.965 48.96 353.245 49.84 ;
    RECT 216.845 48.96 217.125 49.84 ;
    RECT 349.645 48.96 349.925 49.84 ;
    RECT 213.525 48.96 213.805 49.84 ;
    RECT 346.325 48.96 346.605 49.84 ;
    RECT 210.205 48.96 210.485 49.84 ;
    RECT 343.005 48.96 343.285 49.84 ;
    RECT 206.885 48.96 207.165 49.84 ;
    RECT 339.685 48.96 339.965 49.84 ;
    RECT 203.565 48.96 203.845 49.84 ;
    RECT 336.365 48.96 336.645 49.84 ;
    RECT 266.645 48.96 266.925 49.84 ;
    RECT 263.325 48.96 263.605 49.84 ;
    RECT 260.005 48.96 260.285 49.84 ;
    RECT 256.685 48.96 256.965 49.84 ;
    RECT 253.365 48.96 253.645 49.84 ;
    RECT 250.045 48.96 250.325 49.84 ;
    RECT 246.725 48.96 247.005 49.84 ;
    RECT 243.405 48.96 243.685 49.84 ;
    RECT 240.085 48.96 240.365 49.84 ;
    RECT 236.765 48.96 237.045 49.84 ;
    RECT 333.045 48.96 333.325 49.84 ;
    RECT 329.725 48.96 330.005 49.84 ;
    RECT 326.405 48.96 326.685 49.84 ;
    RECT 323.085 48.96 323.365 49.84 ;
    RECT 319.765 48.96 320.045 49.84 ;
    RECT 316.445 48.96 316.725 49.84 ;
    RECT 313.125 48.96 313.405 49.84 ;
    RECT 309.805 48.96 310.085 49.84 ;
    RECT 306.485 48.96 306.765 49.84 ;
    RECT 303.165 48.24 303.445 49.12 ;
    RECT 372.885 48.24 373.165 49.12 ;
    RECT 369.565 48.24 369.845 49.12 ;
    RECT 299.845 48.24 300.125 49.12 ;
    RECT 296.525 48.24 296.805 49.12 ;
    RECT 293.205 48.24 293.485 49.12 ;
    RECT 289.885 48.24 290.165 49.12 ;
    RECT 286.565 48.24 286.845 49.12 ;
    RECT 283.245 48.24 283.525 49.12 ;
    RECT 279.925 48.24 280.205 49.12 ;
    RECT 276.605 48.24 276.885 49.12 ;
    RECT 273.285 48.24 273.565 49.12 ;
    RECT 269.965 48.24 270.245 49.12 ;
    RECT 233.445 48.24 233.725 49.12 ;
    RECT 230.125 48.24 230.405 49.12 ;
    RECT 366.245 48.24 366.525 49.12 ;
    RECT 226.805 48.24 227.085 49.12 ;
    RECT 362.925 48.24 363.205 49.12 ;
    RECT 223.485 48.24 223.765 49.12 ;
    RECT 359.605 48.24 359.885 49.12 ;
    RECT 220.165 48.24 220.445 49.12 ;
    RECT 356.285 48.24 356.565 49.12 ;
    RECT 352.965 48.24 353.245 49.12 ;
    RECT 216.845 48.24 217.125 49.12 ;
    RECT 349.645 48.24 349.925 49.12 ;
    RECT 213.525 48.24 213.805 49.12 ;
    RECT 346.325 48.24 346.605 49.12 ;
    RECT 210.205 48.24 210.485 49.12 ;
    RECT 343.005 48.24 343.285 49.12 ;
    RECT 206.885 48.24 207.165 49.12 ;
    RECT 339.685 48.24 339.965 49.12 ;
    RECT 203.565 48.24 203.845 49.12 ;
    RECT 336.365 48.24 336.645 49.12 ;
    RECT 266.645 48.24 266.925 49.12 ;
    RECT 263.325 48.24 263.605 49.12 ;
    RECT 260.005 48.24 260.285 49.12 ;
    RECT 256.685 48.24 256.965 49.12 ;
    RECT 253.365 48.24 253.645 49.12 ;
    RECT 250.045 48.24 250.325 49.12 ;
    RECT 246.725 48.24 247.005 49.12 ;
    RECT 243.405 48.24 243.685 49.12 ;
    RECT 240.085 48.24 240.365 49.12 ;
    RECT 236.765 48.24 237.045 49.12 ;
    RECT 333.045 48.24 333.325 49.12 ;
    RECT 329.725 48.24 330.005 49.12 ;
    RECT 326.405 48.24 326.685 49.12 ;
    RECT 323.085 48.24 323.365 49.12 ;
    RECT 319.765 48.24 320.045 49.12 ;
    RECT 316.445 48.24 316.725 49.12 ;
    RECT 313.125 48.24 313.405 49.12 ;
    RECT 309.805 48.24 310.085 49.12 ;
    RECT 306.485 48.24 306.765 49.12 ;
    RECT 303.165 47.52 303.445 48.4 ;
    RECT 372.885 47.52 373.165 48.4 ;
    RECT 369.565 47.52 369.845 48.4 ;
    RECT 299.845 47.52 300.125 48.4 ;
    RECT 296.525 47.52 296.805 48.4 ;
    RECT 293.205 47.52 293.485 48.4 ;
    RECT 289.885 47.52 290.165 48.4 ;
    RECT 286.565 47.52 286.845 48.4 ;
    RECT 283.245 47.52 283.525 48.4 ;
    RECT 279.925 47.52 280.205 48.4 ;
    RECT 276.605 47.52 276.885 48.4 ;
    RECT 273.285 47.52 273.565 48.4 ;
    RECT 269.965 47.52 270.245 48.4 ;
    RECT 233.445 47.52 233.725 48.4 ;
    RECT 230.125 47.52 230.405 48.4 ;
    RECT 366.245 47.52 366.525 48.4 ;
    RECT 226.805 47.52 227.085 48.4 ;
    RECT 362.925 47.52 363.205 48.4 ;
    RECT 223.485 47.52 223.765 48.4 ;
    RECT 359.605 47.52 359.885 48.4 ;
    RECT 220.165 47.52 220.445 48.4 ;
    RECT 356.285 47.52 356.565 48.4 ;
    RECT 352.965 47.52 353.245 48.4 ;
    RECT 216.845 47.52 217.125 48.4 ;
    RECT 349.645 47.52 349.925 48.4 ;
    RECT 213.525 47.52 213.805 48.4 ;
    RECT 346.325 47.52 346.605 48.4 ;
    RECT 210.205 47.52 210.485 48.4 ;
    RECT 343.005 47.52 343.285 48.4 ;
    RECT 206.885 47.52 207.165 48.4 ;
    RECT 339.685 47.52 339.965 48.4 ;
    RECT 203.565 47.52 203.845 48.4 ;
    RECT 336.365 47.52 336.645 48.4 ;
    RECT 266.645 47.52 266.925 48.4 ;
    RECT 263.325 47.52 263.605 48.4 ;
    RECT 260.005 47.52 260.285 48.4 ;
    RECT 256.685 47.52 256.965 48.4 ;
    RECT 253.365 47.52 253.645 48.4 ;
    RECT 250.045 47.52 250.325 48.4 ;
    RECT 246.725 47.52 247.005 48.4 ;
    RECT 243.405 47.52 243.685 48.4 ;
    RECT 240.085 47.52 240.365 48.4 ;
    RECT 236.765 47.52 237.045 48.4 ;
    RECT 333.045 47.52 333.325 48.4 ;
    RECT 329.725 47.52 330.005 48.4 ;
    RECT 326.405 47.52 326.685 48.4 ;
    RECT 323.085 47.52 323.365 48.4 ;
    RECT 319.765 47.52 320.045 48.4 ;
    RECT 316.445 47.52 316.725 48.4 ;
    RECT 313.125 47.52 313.405 48.4 ;
    RECT 309.805 47.52 310.085 48.4 ;
    RECT 306.485 47.52 306.765 48.4 ;
    RECT 303.165 46.8 303.445 47.68 ;
    RECT 372.885 46.8 373.165 47.68 ;
    RECT 369.565 46.8 369.845 47.68 ;
    RECT 299.845 46.8 300.125 47.68 ;
    RECT 296.525 46.8 296.805 47.68 ;
    RECT 293.205 46.8 293.485 47.68 ;
    RECT 289.885 46.8 290.165 47.68 ;
    RECT 286.565 46.8 286.845 47.68 ;
    RECT 283.245 46.8 283.525 47.68 ;
    RECT 279.925 46.8 280.205 47.68 ;
    RECT 276.605 46.8 276.885 47.68 ;
    RECT 273.285 46.8 273.565 47.68 ;
    RECT 269.965 46.8 270.245 47.68 ;
    RECT 233.445 46.8 233.725 47.68 ;
    RECT 230.125 46.8 230.405 47.68 ;
    RECT 366.245 46.8 366.525 47.68 ;
    RECT 226.805 46.8 227.085 47.68 ;
    RECT 362.925 46.8 363.205 47.68 ;
    RECT 223.485 46.8 223.765 47.68 ;
    RECT 359.605 46.8 359.885 47.68 ;
    RECT 220.165 46.8 220.445 47.68 ;
    RECT 356.285 46.8 356.565 47.68 ;
    RECT 352.965 46.8 353.245 47.68 ;
    RECT 216.845 46.8 217.125 47.68 ;
    RECT 349.645 46.8 349.925 47.68 ;
    RECT 213.525 46.8 213.805 47.68 ;
    RECT 346.325 46.8 346.605 47.68 ;
    RECT 210.205 46.8 210.485 47.68 ;
    RECT 343.005 46.8 343.285 47.68 ;
    RECT 206.885 46.8 207.165 47.68 ;
    RECT 339.685 46.8 339.965 47.68 ;
    RECT 203.565 46.8 203.845 47.68 ;
    RECT 336.365 46.8 336.645 47.68 ;
    RECT 266.645 46.8 266.925 47.68 ;
    RECT 263.325 46.8 263.605 47.68 ;
    RECT 260.005 46.8 260.285 47.68 ;
    RECT 256.685 46.8 256.965 47.68 ;
    RECT 253.365 46.8 253.645 47.68 ;
    RECT 250.045 46.8 250.325 47.68 ;
    RECT 246.725 46.8 247.005 47.68 ;
    RECT 243.405 46.8 243.685 47.68 ;
    RECT 240.085 46.8 240.365 47.68 ;
    RECT 236.765 46.8 237.045 47.68 ;
    RECT 333.045 46.8 333.325 47.68 ;
    RECT 329.725 46.8 330.005 47.68 ;
    RECT 326.405 46.8 326.685 47.68 ;
    RECT 323.085 46.8 323.365 47.68 ;
    RECT 319.765 46.8 320.045 47.68 ;
    RECT 316.445 46.8 316.725 47.68 ;
    RECT 313.125 46.8 313.405 47.68 ;
    RECT 309.805 46.8 310.085 47.68 ;
    RECT 306.485 46.8 306.765 47.68 ;
    RECT 303.165 46.08 303.445 46.96 ;
    RECT 372.885 46.08 373.165 46.96 ;
    RECT 369.565 46.08 369.845 46.96 ;
    RECT 299.845 46.08 300.125 46.96 ;
    RECT 296.525 46.08 296.805 46.96 ;
    RECT 293.205 46.08 293.485 46.96 ;
    RECT 289.885 46.08 290.165 46.96 ;
    RECT 286.565 46.08 286.845 46.96 ;
    RECT 283.245 46.08 283.525 46.96 ;
    RECT 279.925 46.08 280.205 46.96 ;
    RECT 276.605 46.08 276.885 46.96 ;
    RECT 273.285 46.08 273.565 46.96 ;
    RECT 269.965 46.08 270.245 46.96 ;
    RECT 233.445 46.08 233.725 46.96 ;
    RECT 230.125 46.08 230.405 46.96 ;
    RECT 366.245 46.08 366.525 46.96 ;
    RECT 226.805 46.08 227.085 46.96 ;
    RECT 362.925 46.08 363.205 46.96 ;
    RECT 223.485 46.08 223.765 46.96 ;
    RECT 359.605 46.08 359.885 46.96 ;
    RECT 220.165 46.08 220.445 46.96 ;
    RECT 356.285 46.08 356.565 46.96 ;
    RECT 352.965 46.08 353.245 46.96 ;
    RECT 216.845 46.08 217.125 46.96 ;
    RECT 349.645 46.08 349.925 46.96 ;
    RECT 213.525 46.08 213.805 46.96 ;
    RECT 346.325 46.08 346.605 46.96 ;
    RECT 210.205 46.08 210.485 46.96 ;
    RECT 343.005 46.08 343.285 46.96 ;
    RECT 206.885 46.08 207.165 46.96 ;
    RECT 339.685 46.08 339.965 46.96 ;
    RECT 203.565 46.08 203.845 46.96 ;
    RECT 336.365 46.08 336.645 46.96 ;
    RECT 266.645 46.08 266.925 46.96 ;
    RECT 263.325 46.08 263.605 46.96 ;
    RECT 260.005 46.08 260.285 46.96 ;
    RECT 256.685 46.08 256.965 46.96 ;
    RECT 253.365 46.08 253.645 46.96 ;
    RECT 250.045 46.08 250.325 46.96 ;
    RECT 246.725 46.08 247.005 46.96 ;
    RECT 243.405 46.08 243.685 46.96 ;
    RECT 240.085 46.08 240.365 46.96 ;
    RECT 236.765 46.08 237.045 46.96 ;
    RECT 333.045 46.08 333.325 46.96 ;
    RECT 329.725 46.08 330.005 46.96 ;
    RECT 326.405 46.08 326.685 46.96 ;
    RECT 323.085 46.08 323.365 46.96 ;
    RECT 319.765 46.08 320.045 46.96 ;
    RECT 316.445 46.08 316.725 46.96 ;
    RECT 313.125 46.08 313.405 46.96 ;
    RECT 309.805 46.08 310.085 46.96 ;
    RECT 306.485 46.08 306.765 46.96 ;
    RECT 303.165 45.36 303.445 46.24 ;
    RECT 372.885 45.36 373.165 46.24 ;
    RECT 369.565 45.36 369.845 46.24 ;
    RECT 299.845 45.36 300.125 46.24 ;
    RECT 296.525 45.36 296.805 46.24 ;
    RECT 293.205 45.36 293.485 46.24 ;
    RECT 289.885 45.36 290.165 46.24 ;
    RECT 286.565 45.36 286.845 46.24 ;
    RECT 283.245 45.36 283.525 46.24 ;
    RECT 279.925 45.36 280.205 46.24 ;
    RECT 276.605 45.36 276.885 46.24 ;
    RECT 273.285 45.36 273.565 46.24 ;
    RECT 269.965 45.36 270.245 46.24 ;
    RECT 233.445 45.36 233.725 46.24 ;
    RECT 230.125 45.36 230.405 46.24 ;
    RECT 366.245 45.36 366.525 46.24 ;
    RECT 226.805 45.36 227.085 46.24 ;
    RECT 362.925 45.36 363.205 46.24 ;
    RECT 223.485 45.36 223.765 46.24 ;
    RECT 359.605 45.36 359.885 46.24 ;
    RECT 220.165 45.36 220.445 46.24 ;
    RECT 356.285 45.36 356.565 46.24 ;
    RECT 352.965 45.36 353.245 46.24 ;
    RECT 216.845 45.36 217.125 46.24 ;
    RECT 349.645 45.36 349.925 46.24 ;
    RECT 213.525 45.36 213.805 46.24 ;
    RECT 346.325 45.36 346.605 46.24 ;
    RECT 210.205 45.36 210.485 46.24 ;
    RECT 343.005 45.36 343.285 46.24 ;
    RECT 206.885 45.36 207.165 46.24 ;
    RECT 339.685 45.36 339.965 46.24 ;
    RECT 203.565 45.36 203.845 46.24 ;
    RECT 336.365 45.36 336.645 46.24 ;
    RECT 266.645 45.36 266.925 46.24 ;
    RECT 263.325 45.36 263.605 46.24 ;
    RECT 260.005 45.36 260.285 46.24 ;
    RECT 256.685 45.36 256.965 46.24 ;
    RECT 253.365 45.36 253.645 46.24 ;
    RECT 250.045 45.36 250.325 46.24 ;
    RECT 246.725 45.36 247.005 46.24 ;
    RECT 243.405 45.36 243.685 46.24 ;
    RECT 240.085 45.36 240.365 46.24 ;
    RECT 236.765 45.36 237.045 46.24 ;
    RECT 333.045 45.36 333.325 46.24 ;
    RECT 329.725 45.36 330.005 46.24 ;
    RECT 326.405 45.36 326.685 46.24 ;
    RECT 323.085 45.36 323.365 46.24 ;
    RECT 319.765 45.36 320.045 46.24 ;
    RECT 316.445 45.36 316.725 46.24 ;
    RECT 313.125 45.36 313.405 46.24 ;
    RECT 309.805 45.36 310.085 46.24 ;
    RECT 306.485 45.36 306.765 46.24 ;
    RECT 303.165 44.64 303.445 45.52 ;
    RECT 372.885 44.64 373.165 45.52 ;
    RECT 369.565 44.64 369.845 45.52 ;
    RECT 299.845 44.64 300.125 45.52 ;
    RECT 296.525 44.64 296.805 45.52 ;
    RECT 293.205 44.64 293.485 45.52 ;
    RECT 289.885 44.64 290.165 45.52 ;
    RECT 286.565 44.64 286.845 45.52 ;
    RECT 283.245 44.64 283.525 45.52 ;
    RECT 279.925 44.64 280.205 45.52 ;
    RECT 276.605 44.64 276.885 45.52 ;
    RECT 273.285 44.64 273.565 45.52 ;
    RECT 269.965 44.64 270.245 45.52 ;
    RECT 233.445 44.64 233.725 45.52 ;
    RECT 230.125 44.64 230.405 45.52 ;
    RECT 366.245 44.64 366.525 45.52 ;
    RECT 226.805 44.64 227.085 45.52 ;
    RECT 362.925 44.64 363.205 45.52 ;
    RECT 223.485 44.64 223.765 45.52 ;
    RECT 359.605 44.64 359.885 45.52 ;
    RECT 220.165 44.64 220.445 45.52 ;
    RECT 356.285 44.64 356.565 45.52 ;
    RECT 352.965 44.64 353.245 45.52 ;
    RECT 216.845 44.64 217.125 45.52 ;
    RECT 349.645 44.64 349.925 45.52 ;
    RECT 213.525 44.64 213.805 45.52 ;
    RECT 346.325 44.64 346.605 45.52 ;
    RECT 210.205 44.64 210.485 45.52 ;
    RECT 343.005 44.64 343.285 45.52 ;
    RECT 206.885 44.64 207.165 45.52 ;
    RECT 339.685 44.64 339.965 45.52 ;
    RECT 203.565 44.64 203.845 45.52 ;
    RECT 336.365 44.64 336.645 45.52 ;
    RECT 266.645 44.64 266.925 45.52 ;
    RECT 263.325 44.64 263.605 45.52 ;
    RECT 260.005 44.64 260.285 45.52 ;
    RECT 256.685 44.64 256.965 45.52 ;
    RECT 253.365 44.64 253.645 45.52 ;
    RECT 250.045 44.64 250.325 45.52 ;
    RECT 246.725 44.64 247.005 45.52 ;
    RECT 243.405 44.64 243.685 45.52 ;
    RECT 240.085 44.64 240.365 45.52 ;
    RECT 236.765 44.64 237.045 45.52 ;
    RECT 333.045 44.64 333.325 45.52 ;
    RECT 329.725 44.64 330.005 45.52 ;
    RECT 326.405 44.64 326.685 45.52 ;
    RECT 323.085 44.64 323.365 45.52 ;
    RECT 319.765 44.64 320.045 45.52 ;
    RECT 316.445 44.64 316.725 45.52 ;
    RECT 313.125 44.64 313.405 45.52 ;
    RECT 309.805 44.64 310.085 45.52 ;
    RECT 306.485 44.64 306.765 45.52 ;
    RECT 303.165 43.92 303.445 44.8 ;
    RECT 372.885 43.92 373.165 44.8 ;
    RECT 369.565 43.92 369.845 44.8 ;
    RECT 299.845 43.92 300.125 44.8 ;
    RECT 296.525 43.92 296.805 44.8 ;
    RECT 293.205 43.92 293.485 44.8 ;
    RECT 289.885 43.92 290.165 44.8 ;
    RECT 286.565 43.92 286.845 44.8 ;
    RECT 283.245 43.92 283.525 44.8 ;
    RECT 279.925 43.92 280.205 44.8 ;
    RECT 276.605 43.92 276.885 44.8 ;
    RECT 273.285 43.92 273.565 44.8 ;
    RECT 269.965 43.92 270.245 44.8 ;
    RECT 233.445 43.92 233.725 44.8 ;
    RECT 230.125 43.92 230.405 44.8 ;
    RECT 366.245 43.92 366.525 44.8 ;
    RECT 226.805 43.92 227.085 44.8 ;
    RECT 362.925 43.92 363.205 44.8 ;
    RECT 223.485 43.92 223.765 44.8 ;
    RECT 359.605 43.92 359.885 44.8 ;
    RECT 220.165 43.92 220.445 44.8 ;
    RECT 356.285 43.92 356.565 44.8 ;
    RECT 352.965 43.92 353.245 44.8 ;
    RECT 216.845 43.92 217.125 44.8 ;
    RECT 349.645 43.92 349.925 44.8 ;
    RECT 213.525 43.92 213.805 44.8 ;
    RECT 346.325 43.92 346.605 44.8 ;
    RECT 210.205 43.92 210.485 44.8 ;
    RECT 343.005 43.92 343.285 44.8 ;
    RECT 206.885 43.92 207.165 44.8 ;
    RECT 339.685 43.92 339.965 44.8 ;
    RECT 203.565 43.92 203.845 44.8 ;
    RECT 336.365 43.92 336.645 44.8 ;
    RECT 266.645 43.92 266.925 44.8 ;
    RECT 263.325 43.92 263.605 44.8 ;
    RECT 260.005 43.92 260.285 44.8 ;
    RECT 256.685 43.92 256.965 44.8 ;
    RECT 253.365 43.92 253.645 44.8 ;
    RECT 250.045 43.92 250.325 44.8 ;
    RECT 246.725 43.92 247.005 44.8 ;
    RECT 243.405 43.92 243.685 44.8 ;
    RECT 240.085 43.92 240.365 44.8 ;
    RECT 236.765 43.92 237.045 44.8 ;
    RECT 333.045 43.92 333.325 44.8 ;
    RECT 329.725 43.92 330.005 44.8 ;
    RECT 326.405 43.92 326.685 44.8 ;
    RECT 323.085 43.92 323.365 44.8 ;
    RECT 319.765 43.92 320.045 44.8 ;
    RECT 316.445 43.92 316.725 44.8 ;
    RECT 313.125 43.92 313.405 44.8 ;
    RECT 309.805 43.92 310.085 44.8 ;
    RECT 306.485 43.92 306.765 44.8 ;
    RECT 303.165 43.2 303.445 44.08 ;
    RECT 372.885 43.2 373.165 44.08 ;
    RECT 369.565 43.2 369.845 44.08 ;
    RECT 299.845 43.2 300.125 44.08 ;
    RECT 296.525 43.2 296.805 44.08 ;
    RECT 293.205 43.2 293.485 44.08 ;
    RECT 289.885 43.2 290.165 44.08 ;
    RECT 286.565 43.2 286.845 44.08 ;
    RECT 283.245 43.2 283.525 44.08 ;
    RECT 279.925 43.2 280.205 44.08 ;
    RECT 276.605 43.2 276.885 44.08 ;
    RECT 273.285 43.2 273.565 44.08 ;
    RECT 269.965 43.2 270.245 44.08 ;
    RECT 233.445 43.2 233.725 44.08 ;
    RECT 230.125 43.2 230.405 44.08 ;
    RECT 366.245 43.2 366.525 44.08 ;
    RECT 226.805 43.2 227.085 44.08 ;
    RECT 362.925 43.2 363.205 44.08 ;
    RECT 223.485 43.2 223.765 44.08 ;
    RECT 359.605 43.2 359.885 44.08 ;
    RECT 220.165 43.2 220.445 44.08 ;
    RECT 356.285 43.2 356.565 44.08 ;
    RECT 352.965 43.2 353.245 44.08 ;
    RECT 216.845 43.2 217.125 44.08 ;
    RECT 349.645 43.2 349.925 44.08 ;
    RECT 213.525 43.2 213.805 44.08 ;
    RECT 346.325 43.2 346.605 44.08 ;
    RECT 210.205 43.2 210.485 44.08 ;
    RECT 343.005 43.2 343.285 44.08 ;
    RECT 206.885 43.2 207.165 44.08 ;
    RECT 339.685 43.2 339.965 44.08 ;
    RECT 203.565 43.2 203.845 44.08 ;
    RECT 336.365 43.2 336.645 44.08 ;
    RECT 266.645 43.2 266.925 44.08 ;
    RECT 263.325 43.2 263.605 44.08 ;
    RECT 260.005 43.2 260.285 44.08 ;
    RECT 256.685 43.2 256.965 44.08 ;
    RECT 253.365 43.2 253.645 44.08 ;
    RECT 250.045 43.2 250.325 44.08 ;
    RECT 246.725 43.2 247.005 44.08 ;
    RECT 243.405 43.2 243.685 44.08 ;
    RECT 240.085 43.2 240.365 44.08 ;
    RECT 236.765 43.2 237.045 44.08 ;
    RECT 333.045 43.2 333.325 44.08 ;
    RECT 329.725 43.2 330.005 44.08 ;
    RECT 326.405 43.2 326.685 44.08 ;
    RECT 323.085 43.2 323.365 44.08 ;
    RECT 319.765 43.2 320.045 44.08 ;
    RECT 316.445 43.2 316.725 44.08 ;
    RECT 313.125 43.2 313.405 44.08 ;
    RECT 309.805 43.2 310.085 44.08 ;
    RECT 306.485 43.2 306.765 44.08 ;
    RECT 303.165 42.48 303.445 43.36 ;
    RECT 372.885 42.48 373.165 43.36 ;
    RECT 369.565 42.48 369.845 43.36 ;
    RECT 299.845 42.48 300.125 43.36 ;
    RECT 296.525 42.48 296.805 43.36 ;
    RECT 293.205 42.48 293.485 43.36 ;
    RECT 289.885 42.48 290.165 43.36 ;
    RECT 286.565 42.48 286.845 43.36 ;
    RECT 283.245 42.48 283.525 43.36 ;
    RECT 279.925 42.48 280.205 43.36 ;
    RECT 276.605 42.48 276.885 43.36 ;
    RECT 273.285 42.48 273.565 43.36 ;
    RECT 269.965 42.48 270.245 43.36 ;
    RECT 233.445 42.48 233.725 43.36 ;
    RECT 230.125 42.48 230.405 43.36 ;
    RECT 366.245 42.48 366.525 43.36 ;
    RECT 226.805 42.48 227.085 43.36 ;
    RECT 362.925 42.48 363.205 43.36 ;
    RECT 223.485 42.48 223.765 43.36 ;
    RECT 359.605 42.48 359.885 43.36 ;
    RECT 220.165 42.48 220.445 43.36 ;
    RECT 356.285 42.48 356.565 43.36 ;
    RECT 352.965 42.48 353.245 43.36 ;
    RECT 216.845 42.48 217.125 43.36 ;
    RECT 349.645 42.48 349.925 43.36 ;
    RECT 213.525 42.48 213.805 43.36 ;
    RECT 346.325 42.48 346.605 43.36 ;
    RECT 210.205 42.48 210.485 43.36 ;
    RECT 343.005 42.48 343.285 43.36 ;
    RECT 206.885 42.48 207.165 43.36 ;
    RECT 339.685 42.48 339.965 43.36 ;
    RECT 203.565 42.48 203.845 43.36 ;
    RECT 336.365 42.48 336.645 43.36 ;
    RECT 266.645 42.48 266.925 43.36 ;
    RECT 263.325 42.48 263.605 43.36 ;
    RECT 260.005 42.48 260.285 43.36 ;
    RECT 256.685 42.48 256.965 43.36 ;
    RECT 253.365 42.48 253.645 43.36 ;
    RECT 250.045 42.48 250.325 43.36 ;
    RECT 246.725 42.48 247.005 43.36 ;
    RECT 243.405 42.48 243.685 43.36 ;
    RECT 240.085 42.48 240.365 43.36 ;
    RECT 236.765 42.48 237.045 43.36 ;
    RECT 333.045 42.48 333.325 43.36 ;
    RECT 329.725 42.48 330.005 43.36 ;
    RECT 326.405 42.48 326.685 43.36 ;
    RECT 323.085 42.48 323.365 43.36 ;
    RECT 319.765 42.48 320.045 43.36 ;
    RECT 316.445 42.48 316.725 43.36 ;
    RECT 313.125 42.48 313.405 43.36 ;
    RECT 309.805 42.48 310.085 43.36 ;
    RECT 306.485 42.48 306.765 43.36 ;
    RECT 303.165 41.76 303.445 42.64 ;
    RECT 372.885 41.76 373.165 42.64 ;
    RECT 369.565 41.76 369.845 42.64 ;
    RECT 299.845 41.76 300.125 42.64 ;
    RECT 296.525 41.76 296.805 42.64 ;
    RECT 293.205 41.76 293.485 42.64 ;
    RECT 289.885 41.76 290.165 42.64 ;
    RECT 286.565 41.76 286.845 42.64 ;
    RECT 283.245 41.76 283.525 42.64 ;
    RECT 279.925 41.76 280.205 42.64 ;
    RECT 276.605 41.76 276.885 42.64 ;
    RECT 273.285 41.76 273.565 42.64 ;
    RECT 269.965 41.76 270.245 42.64 ;
    RECT 233.445 41.76 233.725 42.64 ;
    RECT 230.125 41.76 230.405 42.64 ;
    RECT 366.245 41.76 366.525 42.64 ;
    RECT 226.805 41.76 227.085 42.64 ;
    RECT 362.925 41.76 363.205 42.64 ;
    RECT 223.485 41.76 223.765 42.64 ;
    RECT 359.605 41.76 359.885 42.64 ;
    RECT 220.165 41.76 220.445 42.64 ;
    RECT 356.285 41.76 356.565 42.64 ;
    RECT 352.965 41.76 353.245 42.64 ;
    RECT 216.845 41.76 217.125 42.64 ;
    RECT 349.645 41.76 349.925 42.64 ;
    RECT 213.525 41.76 213.805 42.64 ;
    RECT 346.325 41.76 346.605 42.64 ;
    RECT 210.205 41.76 210.485 42.64 ;
    RECT 343.005 41.76 343.285 42.64 ;
    RECT 206.885 41.76 207.165 42.64 ;
    RECT 339.685 41.76 339.965 42.64 ;
    RECT 203.565 41.76 203.845 42.64 ;
    RECT 336.365 41.76 336.645 42.64 ;
    RECT 266.645 41.76 266.925 42.64 ;
    RECT 263.325 41.76 263.605 42.64 ;
    RECT 260.005 41.76 260.285 42.64 ;
    RECT 256.685 41.76 256.965 42.64 ;
    RECT 253.365 41.76 253.645 42.64 ;
    RECT 250.045 41.76 250.325 42.64 ;
    RECT 246.725 41.76 247.005 42.64 ;
    RECT 243.405 41.76 243.685 42.64 ;
    RECT 240.085 41.76 240.365 42.64 ;
    RECT 236.765 41.76 237.045 42.64 ;
    RECT 333.045 41.76 333.325 42.64 ;
    RECT 329.725 41.76 330.005 42.64 ;
    RECT 326.405 41.76 326.685 42.64 ;
    RECT 323.085 41.76 323.365 42.64 ;
    RECT 319.765 41.76 320.045 42.64 ;
    RECT 316.445 41.76 316.725 42.64 ;
    RECT 313.125 41.76 313.405 42.64 ;
    RECT 309.805 41.76 310.085 42.64 ;
    RECT 306.485 41.76 306.765 42.64 ;
    RECT 303.165 41.04 303.445 41.92 ;
    RECT 372.885 41.04 373.165 41.92 ;
    RECT 369.565 41.04 369.845 41.92 ;
    RECT 299.845 41.04 300.125 41.92 ;
    RECT 296.525 41.04 296.805 41.92 ;
    RECT 293.205 41.04 293.485 41.92 ;
    RECT 289.885 41.04 290.165 41.92 ;
    RECT 286.565 41.04 286.845 41.92 ;
    RECT 283.245 41.04 283.525 41.92 ;
    RECT 279.925 41.04 280.205 41.92 ;
    RECT 276.605 41.04 276.885 41.92 ;
    RECT 273.285 41.04 273.565 41.92 ;
    RECT 269.965 41.04 270.245 41.92 ;
    RECT 233.445 41.04 233.725 41.92 ;
    RECT 230.125 41.04 230.405 41.92 ;
    RECT 366.245 41.04 366.525 41.92 ;
    RECT 226.805 41.04 227.085 41.92 ;
    RECT 362.925 41.04 363.205 41.92 ;
    RECT 223.485 41.04 223.765 41.92 ;
    RECT 359.605 41.04 359.885 41.92 ;
    RECT 220.165 41.04 220.445 41.92 ;
    RECT 356.285 41.04 356.565 41.92 ;
    RECT 352.965 41.04 353.245 41.92 ;
    RECT 216.845 41.04 217.125 41.92 ;
    RECT 349.645 41.04 349.925 41.92 ;
    RECT 213.525 41.04 213.805 41.92 ;
    RECT 346.325 41.04 346.605 41.92 ;
    RECT 210.205 41.04 210.485 41.92 ;
    RECT 343.005 41.04 343.285 41.92 ;
    RECT 206.885 41.04 207.165 41.92 ;
    RECT 339.685 41.04 339.965 41.92 ;
    RECT 203.565 41.04 203.845 41.92 ;
    RECT 336.365 41.04 336.645 41.92 ;
    RECT 266.645 41.04 266.925 41.92 ;
    RECT 263.325 41.04 263.605 41.92 ;
    RECT 260.005 41.04 260.285 41.92 ;
    RECT 256.685 41.04 256.965 41.92 ;
    RECT 253.365 41.04 253.645 41.92 ;
    RECT 250.045 41.04 250.325 41.92 ;
    RECT 246.725 41.04 247.005 41.92 ;
    RECT 243.405 41.04 243.685 41.92 ;
    RECT 240.085 41.04 240.365 41.92 ;
    RECT 236.765 41.04 237.045 41.92 ;
    RECT 333.045 41.04 333.325 41.92 ;
    RECT 329.725 41.04 330.005 41.92 ;
    RECT 326.405 41.04 326.685 41.92 ;
    RECT 323.085 41.04 323.365 41.92 ;
    RECT 319.765 41.04 320.045 41.92 ;
    RECT 316.445 41.04 316.725 41.92 ;
    RECT 313.125 41.04 313.405 41.92 ;
    RECT 309.805 41.04 310.085 41.92 ;
    RECT 306.485 41.04 306.765 41.92 ;
    RECT 303.165 40.32 303.445 41.2 ;
    RECT 372.885 40.32 373.165 41.2 ;
    RECT 369.565 40.32 369.845 41.2 ;
    RECT 299.845 40.32 300.125 41.2 ;
    RECT 296.525 40.32 296.805 41.2 ;
    RECT 293.205 40.32 293.485 41.2 ;
    RECT 289.885 40.32 290.165 41.2 ;
    RECT 286.565 40.32 286.845 41.2 ;
    RECT 283.245 40.32 283.525 41.2 ;
    RECT 279.925 40.32 280.205 41.2 ;
    RECT 276.605 40.32 276.885 41.2 ;
    RECT 273.285 40.32 273.565 41.2 ;
    RECT 269.965 40.32 270.245 41.2 ;
    RECT 233.445 40.32 233.725 41.2 ;
    RECT 230.125 40.32 230.405 41.2 ;
    RECT 366.245 40.32 366.525 41.2 ;
    RECT 226.805 40.32 227.085 41.2 ;
    RECT 362.925 40.32 363.205 41.2 ;
    RECT 223.485 40.32 223.765 41.2 ;
    RECT 359.605 40.32 359.885 41.2 ;
    RECT 220.165 40.32 220.445 41.2 ;
    RECT 356.285 40.32 356.565 41.2 ;
    RECT 352.965 40.32 353.245 41.2 ;
    RECT 216.845 40.32 217.125 41.2 ;
    RECT 349.645 40.32 349.925 41.2 ;
    RECT 213.525 40.32 213.805 41.2 ;
    RECT 346.325 40.32 346.605 41.2 ;
    RECT 210.205 40.32 210.485 41.2 ;
    RECT 343.005 40.32 343.285 41.2 ;
    RECT 206.885 40.32 207.165 41.2 ;
    RECT 339.685 40.32 339.965 41.2 ;
    RECT 203.565 40.32 203.845 41.2 ;
    RECT 336.365 40.32 336.645 41.2 ;
    RECT 266.645 40.32 266.925 41.2 ;
    RECT 263.325 40.32 263.605 41.2 ;
    RECT 260.005 40.32 260.285 41.2 ;
    RECT 256.685 40.32 256.965 41.2 ;
    RECT 253.365 40.32 253.645 41.2 ;
    RECT 250.045 40.32 250.325 41.2 ;
    RECT 246.725 40.32 247.005 41.2 ;
    RECT 243.405 40.32 243.685 41.2 ;
    RECT 240.085 40.32 240.365 41.2 ;
    RECT 236.765 40.32 237.045 41.2 ;
    RECT 333.045 40.32 333.325 41.2 ;
    RECT 329.725 40.32 330.005 41.2 ;
    RECT 326.405 40.32 326.685 41.2 ;
    RECT 323.085 40.32 323.365 41.2 ;
    RECT 319.765 40.32 320.045 41.2 ;
    RECT 316.445 40.32 316.725 41.2 ;
    RECT 313.125 40.32 313.405 41.2 ;
    RECT 309.805 40.32 310.085 41.2 ;
    RECT 306.485 40.32 306.765 41.2 ;
    RECT 303.165 58.34 303.445 59.22 ;
    RECT 369.565 58.34 369.845 59.22 ;
    RECT 299.845 58.34 300.125 59.22 ;
    RECT 296.525 58.34 296.805 59.22 ;
    RECT 293.205 58.34 293.485 59.22 ;
    RECT 289.885 58.34 290.165 59.22 ;
    RECT 286.565 58.34 286.845 59.22 ;
    RECT 283.245 58.34 283.525 59.22 ;
    RECT 279.925 58.34 280.205 59.22 ;
    RECT 276.605 58.34 276.885 59.22 ;
    RECT 273.285 58.34 273.565 59.22 ;
    RECT 269.965 58.34 270.245 59.22 ;
    RECT 233.445 58.34 233.725 59.22 ;
    RECT 230.125 58.34 230.405 59.22 ;
    RECT 366.245 58.34 366.525 59.22 ;
    RECT 226.805 58.34 227.085 59.22 ;
    RECT 362.925 58.34 363.205 59.22 ;
    RECT 223.485 58.34 223.765 59.22 ;
    RECT 359.605 58.34 359.885 59.22 ;
    RECT 220.165 58.34 220.445 59.22 ;
    RECT 356.285 58.34 356.565 59.22 ;
    RECT 352.965 58.34 353.245 59.22 ;
    RECT 216.845 58.34 217.125 59.22 ;
    RECT 349.645 58.34 349.925 59.22 ;
    RECT 213.525 58.34 213.805 59.22 ;
    RECT 346.325 58.34 346.605 59.22 ;
    RECT 210.205 58.34 210.485 59.22 ;
    RECT 343.005 58.34 343.285 59.22 ;
    RECT 206.885 58.34 207.165 59.22 ;
    RECT 339.685 58.34 339.965 59.22 ;
    RECT 336.365 58.34 336.645 59.22 ;
    RECT 266.645 58.34 266.925 59.22 ;
    RECT 263.325 58.34 263.605 59.22 ;
    RECT 260.005 58.34 260.285 59.22 ;
    RECT 256.685 58.34 256.965 59.22 ;
    RECT 253.365 58.34 253.645 59.22 ;
    RECT 250.045 58.34 250.325 59.22 ;
    RECT 246.725 58.34 247.005 59.22 ;
    RECT 243.405 58.34 243.685 59.22 ;
    RECT 240.085 58.34 240.365 59.22 ;
    RECT 236.765 58.34 237.045 59.22 ;
    RECT 372.885 58.34 373.165 59.22 ;
    RECT 333.045 58.34 333.325 59.22 ;
    RECT 329.725 58.34 330.005 59.22 ;
    RECT 326.405 58.34 326.685 59.22 ;
    RECT 203.565 58.34 203.845 59.22 ;
    RECT 323.085 58.34 323.365 59.22 ;
    RECT 319.765 58.34 320.045 59.22 ;
    RECT 316.445 58.34 316.725 59.22 ;
    RECT 313.125 58.34 313.405 59.22 ;
    RECT 309.805 58.34 310.085 59.22 ;
    RECT 306.485 58.34 306.765 59.22 ;
    RECT 303.165 39.6 303.445 40.48 ;
    RECT 372.885 39.6 373.165 40.48 ;
    RECT 369.565 39.6 369.845 40.48 ;
    RECT 299.845 39.6 300.125 40.48 ;
    RECT 296.525 39.6 296.805 40.48 ;
    RECT 293.205 39.6 293.485 40.48 ;
    RECT 289.885 39.6 290.165 40.48 ;
    RECT 286.565 39.6 286.845 40.48 ;
    RECT 283.245 39.6 283.525 40.48 ;
    RECT 279.925 39.6 280.205 40.48 ;
    RECT 276.605 39.6 276.885 40.48 ;
    RECT 273.285 39.6 273.565 40.48 ;
    RECT 269.965 39.6 270.245 40.48 ;
    RECT 233.445 39.6 233.725 40.48 ;
    RECT 230.125 39.6 230.405 40.48 ;
    RECT 366.245 39.6 366.525 40.48 ;
    RECT 226.805 39.6 227.085 40.48 ;
    RECT 362.925 39.6 363.205 40.48 ;
    RECT 223.485 39.6 223.765 40.48 ;
    RECT 359.605 39.6 359.885 40.48 ;
    RECT 220.165 39.6 220.445 40.48 ;
    RECT 356.285 39.6 356.565 40.48 ;
    RECT 352.965 39.6 353.245 40.48 ;
    RECT 216.845 39.6 217.125 40.48 ;
    RECT 349.645 39.6 349.925 40.48 ;
    RECT 213.525 39.6 213.805 40.48 ;
    RECT 346.325 39.6 346.605 40.48 ;
    RECT 210.205 39.6 210.485 40.48 ;
    RECT 343.005 39.6 343.285 40.48 ;
    RECT 206.885 39.6 207.165 40.48 ;
    RECT 339.685 39.6 339.965 40.48 ;
    RECT 203.565 39.6 203.845 40.48 ;
    RECT 336.365 39.6 336.645 40.48 ;
    RECT 266.645 39.6 266.925 40.48 ;
    RECT 263.325 39.6 263.605 40.48 ;
    RECT 260.005 39.6 260.285 40.48 ;
    RECT 256.685 39.6 256.965 40.48 ;
    RECT 253.365 39.6 253.645 40.48 ;
    RECT 250.045 39.6 250.325 40.48 ;
    RECT 246.725 39.6 247.005 40.48 ;
    RECT 243.405 39.6 243.685 40.48 ;
    RECT 240.085 39.6 240.365 40.48 ;
    RECT 236.765 39.6 237.045 40.48 ;
    RECT 333.045 39.6 333.325 40.48 ;
    RECT 329.725 39.6 330.005 40.48 ;
    RECT 326.405 39.6 326.685 40.48 ;
    RECT 323.085 39.6 323.365 40.48 ;
    RECT 319.765 39.6 320.045 40.48 ;
    RECT 316.445 39.6 316.725 40.48 ;
    RECT 313.125 39.6 313.405 40.48 ;
    RECT 309.805 39.6 310.085 40.48 ;
    RECT 306.485 39.6 306.765 40.48 ;
    RECT 303.165 38.88 303.445 39.76 ;
    RECT 372.885 38.88 373.165 39.76 ;
    RECT 369.565 38.88 369.845 39.76 ;
    RECT 299.845 38.88 300.125 39.76 ;
    RECT 296.525 38.88 296.805 39.76 ;
    RECT 293.205 38.88 293.485 39.76 ;
    RECT 289.885 38.88 290.165 39.76 ;
    RECT 286.565 38.88 286.845 39.76 ;
    RECT 283.245 38.88 283.525 39.76 ;
    RECT 279.925 38.88 280.205 39.76 ;
    RECT 276.605 38.88 276.885 39.76 ;
    RECT 273.285 38.88 273.565 39.76 ;
    RECT 269.965 38.88 270.245 39.76 ;
    RECT 233.445 38.88 233.725 39.76 ;
    RECT 230.125 38.88 230.405 39.76 ;
    RECT 366.245 38.88 366.525 39.76 ;
    RECT 226.805 38.88 227.085 39.76 ;
    RECT 362.925 38.88 363.205 39.76 ;
    RECT 223.485 38.88 223.765 39.76 ;
    RECT 359.605 38.88 359.885 39.76 ;
    RECT 220.165 38.88 220.445 39.76 ;
    RECT 356.285 38.88 356.565 39.76 ;
    RECT 352.965 38.88 353.245 39.76 ;
    RECT 216.845 38.88 217.125 39.76 ;
    RECT 349.645 38.88 349.925 39.76 ;
    RECT 213.525 38.88 213.805 39.76 ;
    RECT 346.325 38.88 346.605 39.76 ;
    RECT 210.205 38.88 210.485 39.76 ;
    RECT 343.005 38.88 343.285 39.76 ;
    RECT 206.885 38.88 207.165 39.76 ;
    RECT 339.685 38.88 339.965 39.76 ;
    RECT 203.565 38.88 203.845 39.76 ;
    RECT 336.365 38.88 336.645 39.76 ;
    RECT 266.645 38.88 266.925 39.76 ;
    RECT 263.325 38.88 263.605 39.76 ;
    RECT 260.005 38.88 260.285 39.76 ;
    RECT 256.685 38.88 256.965 39.76 ;
    RECT 253.365 38.88 253.645 39.76 ;
    RECT 250.045 38.88 250.325 39.76 ;
    RECT 246.725 38.88 247.005 39.76 ;
    RECT 243.405 38.88 243.685 39.76 ;
    RECT 240.085 38.88 240.365 39.76 ;
    RECT 236.765 38.88 237.045 39.76 ;
    RECT 333.045 38.88 333.325 39.76 ;
    RECT 329.725 38.88 330.005 39.76 ;
    RECT 326.405 38.88 326.685 39.76 ;
    RECT 323.085 38.88 323.365 39.76 ;
    RECT 319.765 38.88 320.045 39.76 ;
    RECT 316.445 38.88 316.725 39.76 ;
    RECT 313.125 38.88 313.405 39.76 ;
    RECT 309.805 38.88 310.085 39.76 ;
    RECT 306.485 38.88 306.765 39.76 ;
    RECT 303.165 38.16 303.445 39.04 ;
    RECT 372.885 38.16 373.165 39.04 ;
    RECT 369.565 38.16 369.845 39.04 ;
    RECT 299.845 38.16 300.125 39.04 ;
    RECT 296.525 38.16 296.805 39.04 ;
    RECT 293.205 38.16 293.485 39.04 ;
    RECT 289.885 38.16 290.165 39.04 ;
    RECT 286.565 38.16 286.845 39.04 ;
    RECT 283.245 38.16 283.525 39.04 ;
    RECT 279.925 38.16 280.205 39.04 ;
    RECT 276.605 38.16 276.885 39.04 ;
    RECT 273.285 38.16 273.565 39.04 ;
    RECT 269.965 38.16 270.245 39.04 ;
    RECT 233.445 38.16 233.725 39.04 ;
    RECT 230.125 38.16 230.405 39.04 ;
    RECT 366.245 38.16 366.525 39.04 ;
    RECT 226.805 38.16 227.085 39.04 ;
    RECT 362.925 38.16 363.205 39.04 ;
    RECT 223.485 38.16 223.765 39.04 ;
    RECT 359.605 38.16 359.885 39.04 ;
    RECT 220.165 38.16 220.445 39.04 ;
    RECT 356.285 38.16 356.565 39.04 ;
    RECT 352.965 38.16 353.245 39.04 ;
    RECT 216.845 38.16 217.125 39.04 ;
    RECT 349.645 38.16 349.925 39.04 ;
    RECT 213.525 38.16 213.805 39.04 ;
    RECT 346.325 38.16 346.605 39.04 ;
    RECT 210.205 38.16 210.485 39.04 ;
    RECT 343.005 38.16 343.285 39.04 ;
    RECT 206.885 38.16 207.165 39.04 ;
    RECT 339.685 38.16 339.965 39.04 ;
    RECT 203.565 38.16 203.845 39.04 ;
    RECT 336.365 38.16 336.645 39.04 ;
    RECT 266.645 38.16 266.925 39.04 ;
    RECT 263.325 38.16 263.605 39.04 ;
    RECT 260.005 38.16 260.285 39.04 ;
    RECT 256.685 38.16 256.965 39.04 ;
    RECT 253.365 38.16 253.645 39.04 ;
    RECT 250.045 38.16 250.325 39.04 ;
    RECT 246.725 38.16 247.005 39.04 ;
    RECT 243.405 38.16 243.685 39.04 ;
    RECT 240.085 38.16 240.365 39.04 ;
    RECT 236.765 38.16 237.045 39.04 ;
    RECT 333.045 38.16 333.325 39.04 ;
    RECT 329.725 38.16 330.005 39.04 ;
    RECT 326.405 38.16 326.685 39.04 ;
    RECT 323.085 38.16 323.365 39.04 ;
    RECT 319.765 38.16 320.045 39.04 ;
    RECT 316.445 38.16 316.725 39.04 ;
    RECT 313.125 38.16 313.405 39.04 ;
    RECT 309.805 38.16 310.085 39.04 ;
    RECT 306.485 38.16 306.765 39.04 ;
    RECT 303.165 37.44 303.445 38.32 ;
    RECT 372.885 37.44 373.165 38.32 ;
    RECT 369.565 37.44 369.845 38.32 ;
    RECT 299.845 37.44 300.125 38.32 ;
    RECT 296.525 37.44 296.805 38.32 ;
    RECT 293.205 37.44 293.485 38.32 ;
    RECT 289.885 37.44 290.165 38.32 ;
    RECT 286.565 37.44 286.845 38.32 ;
    RECT 283.245 37.44 283.525 38.32 ;
    RECT 279.925 37.44 280.205 38.32 ;
    RECT 276.605 37.44 276.885 38.32 ;
    RECT 273.285 37.44 273.565 38.32 ;
    RECT 269.965 37.44 270.245 38.32 ;
    RECT 233.445 37.44 233.725 38.32 ;
    RECT 230.125 37.44 230.405 38.32 ;
    RECT 366.245 37.44 366.525 38.32 ;
    RECT 226.805 37.44 227.085 38.32 ;
    RECT 362.925 37.44 363.205 38.32 ;
    RECT 223.485 37.44 223.765 38.32 ;
    RECT 359.605 37.44 359.885 38.32 ;
    RECT 220.165 37.44 220.445 38.32 ;
    RECT 356.285 37.44 356.565 38.32 ;
    RECT 352.965 37.44 353.245 38.32 ;
    RECT 216.845 37.44 217.125 38.32 ;
    RECT 349.645 37.44 349.925 38.32 ;
    RECT 213.525 37.44 213.805 38.32 ;
    RECT 346.325 37.44 346.605 38.32 ;
    RECT 210.205 37.44 210.485 38.32 ;
    RECT 343.005 37.44 343.285 38.32 ;
    RECT 206.885 37.44 207.165 38.32 ;
    RECT 339.685 37.44 339.965 38.32 ;
    RECT 203.565 37.44 203.845 38.32 ;
    RECT 336.365 37.44 336.645 38.32 ;
    RECT 266.645 37.44 266.925 38.32 ;
    RECT 263.325 37.44 263.605 38.32 ;
    RECT 260.005 37.44 260.285 38.32 ;
    RECT 256.685 37.44 256.965 38.32 ;
    RECT 253.365 37.44 253.645 38.32 ;
    RECT 250.045 37.44 250.325 38.32 ;
    RECT 246.725 37.44 247.005 38.32 ;
    RECT 243.405 37.44 243.685 38.32 ;
    RECT 240.085 37.44 240.365 38.32 ;
    RECT 236.765 37.44 237.045 38.32 ;
    RECT 333.045 37.44 333.325 38.32 ;
    RECT 329.725 37.44 330.005 38.32 ;
    RECT 326.405 37.44 326.685 38.32 ;
    RECT 323.085 37.44 323.365 38.32 ;
    RECT 319.765 37.44 320.045 38.32 ;
    RECT 316.445 37.44 316.725 38.32 ;
    RECT 313.125 37.44 313.405 38.32 ;
    RECT 309.805 37.44 310.085 38.32 ;
    RECT 306.485 37.44 306.765 38.32 ;
    RECT 303.165 36.72 303.445 37.6 ;
    RECT 372.885 36.72 373.165 37.6 ;
    RECT 369.565 36.72 369.845 37.6 ;
    RECT 299.845 36.72 300.125 37.6 ;
    RECT 296.525 36.72 296.805 37.6 ;
    RECT 293.205 36.72 293.485 37.6 ;
    RECT 289.885 36.72 290.165 37.6 ;
    RECT 286.565 36.72 286.845 37.6 ;
    RECT 283.245 36.72 283.525 37.6 ;
    RECT 279.925 36.72 280.205 37.6 ;
    RECT 276.605 36.72 276.885 37.6 ;
    RECT 273.285 36.72 273.565 37.6 ;
    RECT 269.965 36.72 270.245 37.6 ;
    RECT 233.445 36.72 233.725 37.6 ;
    RECT 230.125 36.72 230.405 37.6 ;
    RECT 366.245 36.72 366.525 37.6 ;
    RECT 226.805 36.72 227.085 37.6 ;
    RECT 362.925 36.72 363.205 37.6 ;
    RECT 223.485 36.72 223.765 37.6 ;
    RECT 359.605 36.72 359.885 37.6 ;
    RECT 220.165 36.72 220.445 37.6 ;
    RECT 356.285 36.72 356.565 37.6 ;
    RECT 352.965 36.72 353.245 37.6 ;
    RECT 216.845 36.72 217.125 37.6 ;
    RECT 349.645 36.72 349.925 37.6 ;
    RECT 213.525 36.72 213.805 37.6 ;
    RECT 346.325 36.72 346.605 37.6 ;
    RECT 210.205 36.72 210.485 37.6 ;
    RECT 343.005 36.72 343.285 37.6 ;
    RECT 206.885 36.72 207.165 37.6 ;
    RECT 339.685 36.72 339.965 37.6 ;
    RECT 203.565 36.72 203.845 37.6 ;
    RECT 336.365 36.72 336.645 37.6 ;
    RECT 266.645 36.72 266.925 37.6 ;
    RECT 263.325 36.72 263.605 37.6 ;
    RECT 260.005 36.72 260.285 37.6 ;
    RECT 256.685 36.72 256.965 37.6 ;
    RECT 253.365 36.72 253.645 37.6 ;
    RECT 250.045 36.72 250.325 37.6 ;
    RECT 246.725 36.72 247.005 37.6 ;
    RECT 243.405 36.72 243.685 37.6 ;
    RECT 240.085 36.72 240.365 37.6 ;
    RECT 236.765 36.72 237.045 37.6 ;
    RECT 333.045 36.72 333.325 37.6 ;
    RECT 329.725 36.72 330.005 37.6 ;
    RECT 326.405 36.72 326.685 37.6 ;
    RECT 323.085 36.72 323.365 37.6 ;
    RECT 319.765 36.72 320.045 37.6 ;
    RECT 316.445 36.72 316.725 37.6 ;
    RECT 313.125 36.72 313.405 37.6 ;
    RECT 309.805 36.72 310.085 37.6 ;
    RECT 306.485 36.72 306.765 37.6 ;
    RECT 303.165 36.0 303.445 36.88 ;
    RECT 372.885 36.0 373.165 36.88 ;
    RECT 369.565 36.0 369.845 36.88 ;
    RECT 299.845 36.0 300.125 36.88 ;
    RECT 296.525 36.0 296.805 36.88 ;
    RECT 293.205 36.0 293.485 36.88 ;
    RECT 289.885 36.0 290.165 36.88 ;
    RECT 286.565 36.0 286.845 36.88 ;
    RECT 283.245 36.0 283.525 36.88 ;
    RECT 279.925 36.0 280.205 36.88 ;
    RECT 276.605 36.0 276.885 36.88 ;
    RECT 273.285 36.0 273.565 36.88 ;
    RECT 269.965 36.0 270.245 36.88 ;
    RECT 233.445 36.0 233.725 36.88 ;
    RECT 230.125 36.0 230.405 36.88 ;
    RECT 366.245 36.0 366.525 36.88 ;
    RECT 226.805 36.0 227.085 36.88 ;
    RECT 362.925 36.0 363.205 36.88 ;
    RECT 223.485 36.0 223.765 36.88 ;
    RECT 359.605 36.0 359.885 36.88 ;
    RECT 220.165 36.0 220.445 36.88 ;
    RECT 356.285 36.0 356.565 36.88 ;
    RECT 352.965 36.0 353.245 36.88 ;
    RECT 216.845 36.0 217.125 36.88 ;
    RECT 349.645 36.0 349.925 36.88 ;
    RECT 213.525 36.0 213.805 36.88 ;
    RECT 346.325 36.0 346.605 36.88 ;
    RECT 210.205 36.0 210.485 36.88 ;
    RECT 343.005 36.0 343.285 36.88 ;
    RECT 206.885 36.0 207.165 36.88 ;
    RECT 339.685 36.0 339.965 36.88 ;
    RECT 203.565 36.0 203.845 36.88 ;
    RECT 336.365 36.0 336.645 36.88 ;
    RECT 266.645 36.0 266.925 36.88 ;
    RECT 263.325 36.0 263.605 36.88 ;
    RECT 260.005 36.0 260.285 36.88 ;
    RECT 256.685 36.0 256.965 36.88 ;
    RECT 253.365 36.0 253.645 36.88 ;
    RECT 250.045 36.0 250.325 36.88 ;
    RECT 246.725 36.0 247.005 36.88 ;
    RECT 243.405 36.0 243.685 36.88 ;
    RECT 240.085 36.0 240.365 36.88 ;
    RECT 236.765 36.0 237.045 36.88 ;
    RECT 333.045 36.0 333.325 36.88 ;
    RECT 329.725 36.0 330.005 36.88 ;
    RECT 326.405 36.0 326.685 36.88 ;
    RECT 323.085 36.0 323.365 36.88 ;
    RECT 319.765 36.0 320.045 36.88 ;
    RECT 316.445 36.0 316.725 36.88 ;
    RECT 313.125 36.0 313.405 36.88 ;
    RECT 309.805 36.0 310.085 36.88 ;
    RECT 306.485 36.0 306.765 36.88 ;
    RECT 61.215 49.68 61.495 50.56 ;
    RECT 57.895 49.68 58.175 50.56 ;
    RECT 54.575 49.68 54.855 50.56 ;
    RECT 51.255 49.68 51.535 50.56 ;
    RECT 47.935 49.68 48.215 50.56 ;
    RECT 44.615 49.68 44.895 50.56 ;
    RECT 41.295 49.68 41.575 50.56 ;
    RECT 37.975 49.68 38.255 50.56 ;
    RECT 34.655 49.68 34.935 50.56 ;
    RECT 130.935 49.68 131.215 50.56 ;
    RECT 127.615 49.68 127.895 50.56 ;
    RECT 124.295 49.68 124.575 50.56 ;
    RECT 120.975 49.68 121.255 50.56 ;
    RECT 117.655 49.68 117.935 50.56 ;
    RECT 114.335 49.68 114.615 50.56 ;
    RECT 111.015 49.68 111.295 50.56 ;
    RECT 107.695 49.68 107.975 50.56 ;
    RECT 104.375 49.68 104.655 50.56 ;
    RECT 101.055 49.68 101.335 50.56 ;
    RECT 170.775 49.68 171.055 50.56 ;
    RECT 167.455 49.68 167.735 50.56 ;
    RECT 97.735 49.68 98.015 50.56 ;
    RECT 94.415 49.68 94.695 50.56 ;
    RECT 91.095 49.68 91.375 50.56 ;
    RECT 87.775 49.68 88.055 50.56 ;
    RECT 84.455 49.68 84.735 50.56 ;
    RECT 81.135 49.68 81.415 50.56 ;
    RECT 77.815 49.68 78.095 50.56 ;
    RECT 74.495 49.68 74.775 50.56 ;
    RECT 71.175 49.68 71.455 50.56 ;
    RECT 31.335 49.68 31.615 50.56 ;
    RECT 67.855 49.68 68.135 50.56 ;
    RECT 28.015 49.68 28.295 50.56 ;
    RECT 24.695 49.68 24.975 50.56 ;
    RECT 21.375 49.68 21.655 50.56 ;
    RECT 18.055 49.68 18.335 50.56 ;
    RECT 14.735 49.68 15.015 50.56 ;
    RECT 11.415 49.68 11.695 50.56 ;
    RECT 8.095 49.68 8.375 50.56 ;
    RECT 4.775 49.68 5.055 50.56 ;
    RECT 164.135 49.68 164.415 50.56 ;
    RECT 1.455 49.68 1.735 50.56 ;
    RECT 160.815 49.68 161.095 50.56 ;
    RECT 157.495 49.68 157.775 50.56 ;
    RECT 154.175 49.68 154.455 50.56 ;
    RECT 150.855 49.68 151.135 50.56 ;
    RECT 147.535 49.68 147.815 50.56 ;
    RECT 144.215 49.68 144.495 50.56 ;
    RECT 140.895 49.68 141.175 50.56 ;
    RECT 137.575 49.68 137.855 50.56 ;
    RECT 134.255 49.68 134.535 50.56 ;
    RECT 64.535 49.68 64.815 50.56 ;
    RECT 61.215 48.96 61.495 49.84 ;
    RECT 57.895 48.96 58.175 49.84 ;
    RECT 54.575 48.96 54.855 49.84 ;
    RECT 51.255 48.96 51.535 49.84 ;
    RECT 47.935 48.96 48.215 49.84 ;
    RECT 44.615 48.96 44.895 49.84 ;
    RECT 41.295 48.96 41.575 49.84 ;
    RECT 37.975 48.96 38.255 49.84 ;
    RECT 34.655 48.96 34.935 49.84 ;
    RECT 130.935 48.96 131.215 49.84 ;
    RECT 127.615 48.96 127.895 49.84 ;
    RECT 124.295 48.96 124.575 49.84 ;
    RECT 120.975 48.96 121.255 49.84 ;
    RECT 117.655 48.96 117.935 49.84 ;
    RECT 114.335 48.96 114.615 49.84 ;
    RECT 111.015 48.96 111.295 49.84 ;
    RECT 107.695 48.96 107.975 49.84 ;
    RECT 104.375 48.96 104.655 49.84 ;
    RECT 101.055 48.96 101.335 49.84 ;
    RECT 170.775 48.96 171.055 49.84 ;
    RECT 167.455 48.96 167.735 49.84 ;
    RECT 97.735 48.96 98.015 49.84 ;
    RECT 94.415 48.96 94.695 49.84 ;
    RECT 91.095 48.96 91.375 49.84 ;
    RECT 87.775 48.96 88.055 49.84 ;
    RECT 84.455 48.96 84.735 49.84 ;
    RECT 81.135 48.96 81.415 49.84 ;
    RECT 77.815 48.96 78.095 49.84 ;
    RECT 74.495 48.96 74.775 49.84 ;
    RECT 71.175 48.96 71.455 49.84 ;
    RECT 31.335 48.96 31.615 49.84 ;
    RECT 67.855 48.96 68.135 49.84 ;
    RECT 28.015 48.96 28.295 49.84 ;
    RECT 24.695 48.96 24.975 49.84 ;
    RECT 21.375 48.96 21.655 49.84 ;
    RECT 18.055 48.96 18.335 49.84 ;
    RECT 14.735 48.96 15.015 49.84 ;
    RECT 11.415 48.96 11.695 49.84 ;
    RECT 8.095 48.96 8.375 49.84 ;
    RECT 4.775 48.96 5.055 49.84 ;
    RECT 164.135 48.96 164.415 49.84 ;
    RECT 1.455 48.96 1.735 49.84 ;
    RECT 160.815 48.96 161.095 49.84 ;
    RECT 157.495 48.96 157.775 49.84 ;
    RECT 154.175 48.96 154.455 49.84 ;
    RECT 150.855 48.96 151.135 49.84 ;
    RECT 147.535 48.96 147.815 49.84 ;
    RECT 144.215 48.96 144.495 49.84 ;
    RECT 140.895 48.96 141.175 49.84 ;
    RECT 137.575 48.96 137.855 49.84 ;
    RECT 134.255 48.96 134.535 49.84 ;
    RECT 64.535 48.96 64.815 49.84 ;
    RECT 61.215 48.24 61.495 49.12 ;
    RECT 57.895 48.24 58.175 49.12 ;
    RECT 54.575 48.24 54.855 49.12 ;
    RECT 51.255 48.24 51.535 49.12 ;
    RECT 47.935 48.24 48.215 49.12 ;
    RECT 44.615 48.24 44.895 49.12 ;
    RECT 41.295 48.24 41.575 49.12 ;
    RECT 37.975 48.24 38.255 49.12 ;
    RECT 34.655 48.24 34.935 49.12 ;
    RECT 130.935 48.24 131.215 49.12 ;
    RECT 127.615 48.24 127.895 49.12 ;
    RECT 124.295 48.24 124.575 49.12 ;
    RECT 120.975 48.24 121.255 49.12 ;
    RECT 117.655 48.24 117.935 49.12 ;
    RECT 114.335 48.24 114.615 49.12 ;
    RECT 111.015 48.24 111.295 49.12 ;
    RECT 107.695 48.24 107.975 49.12 ;
    RECT 104.375 48.24 104.655 49.12 ;
    RECT 101.055 48.24 101.335 49.12 ;
    RECT 170.775 48.24 171.055 49.12 ;
    RECT 167.455 48.24 167.735 49.12 ;
    RECT 97.735 48.24 98.015 49.12 ;
    RECT 94.415 48.24 94.695 49.12 ;
    RECT 91.095 48.24 91.375 49.12 ;
    RECT 87.775 48.24 88.055 49.12 ;
    RECT 84.455 48.24 84.735 49.12 ;
    RECT 81.135 48.24 81.415 49.12 ;
    RECT 77.815 48.24 78.095 49.12 ;
    RECT 74.495 48.24 74.775 49.12 ;
    RECT 71.175 48.24 71.455 49.12 ;
    RECT 31.335 48.24 31.615 49.12 ;
    RECT 67.855 48.24 68.135 49.12 ;
    RECT 28.015 48.24 28.295 49.12 ;
    RECT 24.695 48.24 24.975 49.12 ;
    RECT 21.375 48.24 21.655 49.12 ;
    RECT 18.055 48.24 18.335 49.12 ;
    RECT 14.735 48.24 15.015 49.12 ;
    RECT 11.415 48.24 11.695 49.12 ;
    RECT 8.095 48.24 8.375 49.12 ;
    RECT 4.775 48.24 5.055 49.12 ;
    RECT 164.135 48.24 164.415 49.12 ;
    RECT 1.455 48.24 1.735 49.12 ;
    RECT 160.815 48.24 161.095 49.12 ;
    RECT 157.495 48.24 157.775 49.12 ;
    RECT 154.175 48.24 154.455 49.12 ;
    RECT 150.855 48.24 151.135 49.12 ;
    RECT 147.535 48.24 147.815 49.12 ;
    RECT 144.215 48.24 144.495 49.12 ;
    RECT 140.895 48.24 141.175 49.12 ;
    RECT 137.575 48.24 137.855 49.12 ;
    RECT 134.255 48.24 134.535 49.12 ;
    RECT 64.535 48.24 64.815 49.12 ;
    RECT 61.215 47.52 61.495 48.4 ;
    RECT 57.895 47.52 58.175 48.4 ;
    RECT 54.575 47.52 54.855 48.4 ;
    RECT 51.255 47.52 51.535 48.4 ;
    RECT 47.935 47.52 48.215 48.4 ;
    RECT 44.615 47.52 44.895 48.4 ;
    RECT 41.295 47.52 41.575 48.4 ;
    RECT 37.975 47.52 38.255 48.4 ;
    RECT 34.655 47.52 34.935 48.4 ;
    RECT 130.935 47.52 131.215 48.4 ;
    RECT 127.615 47.52 127.895 48.4 ;
    RECT 124.295 47.52 124.575 48.4 ;
    RECT 120.975 47.52 121.255 48.4 ;
    RECT 117.655 47.52 117.935 48.4 ;
    RECT 114.335 47.52 114.615 48.4 ;
    RECT 111.015 47.52 111.295 48.4 ;
    RECT 107.695 47.52 107.975 48.4 ;
    RECT 104.375 47.52 104.655 48.4 ;
    RECT 101.055 47.52 101.335 48.4 ;
    RECT 170.775 47.52 171.055 48.4 ;
    RECT 167.455 47.52 167.735 48.4 ;
    RECT 97.735 47.52 98.015 48.4 ;
    RECT 94.415 47.52 94.695 48.4 ;
    RECT 91.095 47.52 91.375 48.4 ;
    RECT 87.775 47.52 88.055 48.4 ;
    RECT 84.455 47.52 84.735 48.4 ;
    RECT 81.135 47.52 81.415 48.4 ;
    RECT 77.815 47.52 78.095 48.4 ;
    RECT 74.495 47.52 74.775 48.4 ;
    RECT 71.175 47.52 71.455 48.4 ;
    RECT 31.335 47.52 31.615 48.4 ;
    RECT 67.855 47.52 68.135 48.4 ;
    RECT 28.015 47.52 28.295 48.4 ;
    RECT 24.695 47.52 24.975 48.4 ;
    RECT 21.375 47.52 21.655 48.4 ;
    RECT 18.055 47.52 18.335 48.4 ;
    RECT 14.735 47.52 15.015 48.4 ;
    RECT 11.415 47.52 11.695 48.4 ;
    RECT 8.095 47.52 8.375 48.4 ;
    RECT 4.775 47.52 5.055 48.4 ;
    RECT 164.135 47.52 164.415 48.4 ;
    RECT 1.455 47.52 1.735 48.4 ;
    RECT 160.815 47.52 161.095 48.4 ;
    RECT 157.495 47.52 157.775 48.4 ;
    RECT 154.175 47.52 154.455 48.4 ;
    RECT 150.855 47.52 151.135 48.4 ;
    RECT 147.535 47.52 147.815 48.4 ;
    RECT 144.215 47.52 144.495 48.4 ;
    RECT 140.895 47.52 141.175 48.4 ;
    RECT 137.575 47.52 137.855 48.4 ;
    RECT 134.255 47.52 134.535 48.4 ;
    RECT 64.535 47.52 64.815 48.4 ;
    RECT 61.215 11.52 61.495 12.4 ;
    RECT 57.895 11.52 58.175 12.4 ;
    RECT 54.575 11.52 54.855 12.4 ;
    RECT 51.255 11.52 51.535 12.4 ;
    RECT 47.935 11.52 48.215 12.4 ;
    RECT 44.615 11.52 44.895 12.4 ;
    RECT 41.295 11.52 41.575 12.4 ;
    RECT 37.975 11.52 38.255 12.4 ;
    RECT 34.655 11.52 34.935 12.4 ;
    RECT 130.935 11.52 131.215 12.4 ;
    RECT 127.615 11.52 127.895 12.4 ;
    RECT 124.295 11.52 124.575 12.4 ;
    RECT 120.975 11.52 121.255 12.4 ;
    RECT 117.655 11.52 117.935 12.4 ;
    RECT 114.335 11.52 114.615 12.4 ;
    RECT 111.015 11.52 111.295 12.4 ;
    RECT 107.695 11.52 107.975 12.4 ;
    RECT 104.375 11.52 104.655 12.4 ;
    RECT 101.055 11.52 101.335 12.4 ;
    RECT 167.455 11.52 167.735 12.4 ;
    RECT 97.735 11.52 98.015 12.4 ;
    RECT 94.415 11.52 94.695 12.4 ;
    RECT 91.095 11.52 91.375 12.4 ;
    RECT 87.775 11.52 88.055 12.4 ;
    RECT 84.455 11.52 84.735 12.4 ;
    RECT 81.135 11.52 81.415 12.4 ;
    RECT 77.815 11.52 78.095 12.4 ;
    RECT 74.495 11.52 74.775 12.4 ;
    RECT 71.175 11.52 71.455 12.4 ;
    RECT 31.335 11.52 31.615 12.4 ;
    RECT 67.855 11.52 68.135 12.4 ;
    RECT 28.015 11.52 28.295 12.4 ;
    RECT 24.695 11.52 24.975 12.4 ;
    RECT 21.375 11.52 21.655 12.4 ;
    RECT 18.055 11.52 18.335 12.4 ;
    RECT 14.735 11.52 15.015 12.4 ;
    RECT 11.415 11.52 11.695 12.4 ;
    RECT 8.095 11.52 8.375 12.4 ;
    RECT 4.775 11.52 5.055 12.4 ;
    RECT 164.135 11.52 164.415 12.4 ;
    RECT 160.815 11.52 161.095 12.4 ;
    RECT 157.495 11.52 157.775 12.4 ;
    RECT 154.175 11.52 154.455 12.4 ;
    RECT 150.855 11.52 151.135 12.4 ;
    RECT 170.775 11.52 171.055 12.4 ;
    RECT 147.535 11.52 147.815 12.4 ;
    RECT 144.215 11.52 144.495 12.4 ;
    RECT 140.895 11.52 141.175 12.4 ;
    RECT 137.575 11.52 137.855 12.4 ;
    RECT 134.255 11.52 134.535 12.4 ;
    RECT 1.455 11.52 1.735 12.4 ;
    RECT 64.535 11.52 64.815 12.4 ;
    RECT 61.215 18.0 61.495 18.88 ;
    RECT 57.895 18.0 58.175 18.88 ;
    RECT 54.575 18.0 54.855 18.88 ;
    RECT 51.255 18.0 51.535 18.88 ;
    RECT 47.935 18.0 48.215 18.88 ;
    RECT 44.615 18.0 44.895 18.88 ;
    RECT 41.295 18.0 41.575 18.88 ;
    RECT 37.975 18.0 38.255 18.88 ;
    RECT 34.655 18.0 34.935 18.88 ;
    RECT 130.935 18.0 131.215 18.88 ;
    RECT 127.615 18.0 127.895 18.88 ;
    RECT 124.295 18.0 124.575 18.88 ;
    RECT 120.975 18.0 121.255 18.88 ;
    RECT 117.655 18.0 117.935 18.88 ;
    RECT 114.335 18.0 114.615 18.88 ;
    RECT 111.015 18.0 111.295 18.88 ;
    RECT 107.695 18.0 107.975 18.88 ;
    RECT 104.375 18.0 104.655 18.88 ;
    RECT 101.055 18.0 101.335 18.88 ;
    RECT 170.775 18.0 171.055 18.88 ;
    RECT 167.455 18.0 167.735 18.88 ;
    RECT 97.735 18.0 98.015 18.88 ;
    RECT 94.415 18.0 94.695 18.88 ;
    RECT 91.095 18.0 91.375 18.88 ;
    RECT 87.775 18.0 88.055 18.88 ;
    RECT 84.455 18.0 84.735 18.88 ;
    RECT 81.135 18.0 81.415 18.88 ;
    RECT 77.815 18.0 78.095 18.88 ;
    RECT 74.495 18.0 74.775 18.88 ;
    RECT 71.175 18.0 71.455 18.88 ;
    RECT 31.335 18.0 31.615 18.88 ;
    RECT 67.855 18.0 68.135 18.88 ;
    RECT 28.015 18.0 28.295 18.88 ;
    RECT 24.695 18.0 24.975 18.88 ;
    RECT 21.375 18.0 21.655 18.88 ;
    RECT 18.055 18.0 18.335 18.88 ;
    RECT 14.735 18.0 15.015 18.88 ;
    RECT 11.415 18.0 11.695 18.88 ;
    RECT 8.095 18.0 8.375 18.88 ;
    RECT 4.775 18.0 5.055 18.88 ;
    RECT 164.135 18.0 164.415 18.88 ;
    RECT 1.455 18.0 1.735 18.88 ;
    RECT 160.815 18.0 161.095 18.88 ;
    RECT 157.495 18.0 157.775 18.88 ;
    RECT 154.175 18.0 154.455 18.88 ;
    RECT 150.855 18.0 151.135 18.88 ;
    RECT 147.535 18.0 147.815 18.88 ;
    RECT 144.215 18.0 144.495 18.88 ;
    RECT 140.895 18.0 141.175 18.88 ;
    RECT 137.575 18.0 137.855 18.88 ;
    RECT 134.255 18.0 134.535 18.88 ;
    RECT 64.535 18.0 64.815 18.88 ;
    RECT 61.215 17.28 61.495 18.16 ;
    RECT 57.895 17.28 58.175 18.16 ;
    RECT 54.575 17.28 54.855 18.16 ;
    RECT 51.255 17.28 51.535 18.16 ;
    RECT 47.935 17.28 48.215 18.16 ;
    RECT 44.615 17.28 44.895 18.16 ;
    RECT 41.295 17.28 41.575 18.16 ;
    RECT 37.975 17.28 38.255 18.16 ;
    RECT 34.655 17.28 34.935 18.16 ;
    RECT 130.935 17.28 131.215 18.16 ;
    RECT 127.615 17.28 127.895 18.16 ;
    RECT 124.295 17.28 124.575 18.16 ;
    RECT 120.975 17.28 121.255 18.16 ;
    RECT 117.655 17.28 117.935 18.16 ;
    RECT 114.335 17.28 114.615 18.16 ;
    RECT 111.015 17.28 111.295 18.16 ;
    RECT 107.695 17.28 107.975 18.16 ;
    RECT 104.375 17.28 104.655 18.16 ;
    RECT 101.055 17.28 101.335 18.16 ;
    RECT 170.775 17.28 171.055 18.16 ;
    RECT 167.455 17.28 167.735 18.16 ;
    RECT 97.735 17.28 98.015 18.16 ;
    RECT 94.415 17.28 94.695 18.16 ;
    RECT 91.095 17.28 91.375 18.16 ;
    RECT 87.775 17.28 88.055 18.16 ;
    RECT 84.455 17.28 84.735 18.16 ;
    RECT 81.135 17.28 81.415 18.16 ;
    RECT 77.815 17.28 78.095 18.16 ;
    RECT 74.495 17.28 74.775 18.16 ;
    RECT 71.175 17.28 71.455 18.16 ;
    RECT 31.335 17.28 31.615 18.16 ;
    RECT 67.855 17.28 68.135 18.16 ;
    RECT 28.015 17.28 28.295 18.16 ;
    RECT 24.695 17.28 24.975 18.16 ;
    RECT 21.375 17.28 21.655 18.16 ;
    RECT 18.055 17.28 18.335 18.16 ;
    RECT 14.735 17.28 15.015 18.16 ;
    RECT 11.415 17.28 11.695 18.16 ;
    RECT 8.095 17.28 8.375 18.16 ;
    RECT 4.775 17.28 5.055 18.16 ;
    RECT 164.135 17.28 164.415 18.16 ;
    RECT 1.455 17.28 1.735 18.16 ;
    RECT 160.815 17.28 161.095 18.16 ;
    RECT 157.495 17.28 157.775 18.16 ;
    RECT 154.175 17.28 154.455 18.16 ;
    RECT 150.855 17.28 151.135 18.16 ;
    RECT 147.535 17.28 147.815 18.16 ;
    RECT 144.215 17.28 144.495 18.16 ;
    RECT 140.895 17.28 141.175 18.16 ;
    RECT 137.575 17.28 137.855 18.16 ;
    RECT 134.255 17.28 134.535 18.16 ;
    RECT 64.535 17.28 64.815 18.16 ;
    RECT 61.215 16.56 61.495 17.44 ;
    RECT 57.895 16.56 58.175 17.44 ;
    RECT 54.575 16.56 54.855 17.44 ;
    RECT 51.255 16.56 51.535 17.44 ;
    RECT 47.935 16.56 48.215 17.44 ;
    RECT 44.615 16.56 44.895 17.44 ;
    RECT 41.295 16.56 41.575 17.44 ;
    RECT 37.975 16.56 38.255 17.44 ;
    RECT 34.655 16.56 34.935 17.44 ;
    RECT 130.935 16.56 131.215 17.44 ;
    RECT 127.615 16.56 127.895 17.44 ;
    RECT 124.295 16.56 124.575 17.44 ;
    RECT 120.975 16.56 121.255 17.44 ;
    RECT 117.655 16.56 117.935 17.44 ;
    RECT 114.335 16.56 114.615 17.44 ;
    RECT 111.015 16.56 111.295 17.44 ;
    RECT 107.695 16.56 107.975 17.44 ;
    RECT 104.375 16.56 104.655 17.44 ;
    RECT 101.055 16.56 101.335 17.44 ;
    RECT 170.775 16.56 171.055 17.44 ;
    RECT 167.455 16.56 167.735 17.44 ;
    RECT 97.735 16.56 98.015 17.44 ;
    RECT 94.415 16.56 94.695 17.44 ;
    RECT 91.095 16.56 91.375 17.44 ;
    RECT 87.775 16.56 88.055 17.44 ;
    RECT 84.455 16.56 84.735 17.44 ;
    RECT 81.135 16.56 81.415 17.44 ;
    RECT 77.815 16.56 78.095 17.44 ;
    RECT 74.495 16.56 74.775 17.44 ;
    RECT 71.175 16.56 71.455 17.44 ;
    RECT 31.335 16.56 31.615 17.44 ;
    RECT 67.855 16.56 68.135 17.44 ;
    RECT 28.015 16.56 28.295 17.44 ;
    RECT 24.695 16.56 24.975 17.44 ;
    RECT 21.375 16.56 21.655 17.44 ;
    RECT 18.055 16.56 18.335 17.44 ;
    RECT 14.735 16.56 15.015 17.44 ;
    RECT 11.415 16.56 11.695 17.44 ;
    RECT 8.095 16.56 8.375 17.44 ;
    RECT 4.775 16.56 5.055 17.44 ;
    RECT 164.135 16.56 164.415 17.44 ;
    RECT 1.455 16.56 1.735 17.44 ;
    RECT 160.815 16.56 161.095 17.44 ;
    RECT 157.495 16.56 157.775 17.44 ;
    RECT 154.175 16.56 154.455 17.44 ;
    RECT 150.855 16.56 151.135 17.44 ;
    RECT 147.535 16.56 147.815 17.44 ;
    RECT 144.215 16.56 144.495 17.44 ;
    RECT 140.895 16.56 141.175 17.44 ;
    RECT 137.575 16.56 137.855 17.44 ;
    RECT 134.255 16.56 134.535 17.44 ;
    RECT 64.535 16.56 64.815 17.44 ;
    RECT 61.215 15.84 61.495 16.72 ;
    RECT 57.895 15.84 58.175 16.72 ;
    RECT 54.575 15.84 54.855 16.72 ;
    RECT 51.255 15.84 51.535 16.72 ;
    RECT 47.935 15.84 48.215 16.72 ;
    RECT 44.615 15.84 44.895 16.72 ;
    RECT 41.295 15.84 41.575 16.72 ;
    RECT 37.975 15.84 38.255 16.72 ;
    RECT 34.655 15.84 34.935 16.72 ;
    RECT 130.935 15.84 131.215 16.72 ;
    RECT 127.615 15.84 127.895 16.72 ;
    RECT 124.295 15.84 124.575 16.72 ;
    RECT 120.975 15.84 121.255 16.72 ;
    RECT 117.655 15.84 117.935 16.72 ;
    RECT 114.335 15.84 114.615 16.72 ;
    RECT 111.015 15.84 111.295 16.72 ;
    RECT 107.695 15.84 107.975 16.72 ;
    RECT 104.375 15.84 104.655 16.72 ;
    RECT 101.055 15.84 101.335 16.72 ;
    RECT 170.775 15.84 171.055 16.72 ;
    RECT 167.455 15.84 167.735 16.72 ;
    RECT 97.735 15.84 98.015 16.72 ;
    RECT 94.415 15.84 94.695 16.72 ;
    RECT 91.095 15.84 91.375 16.72 ;
    RECT 87.775 15.84 88.055 16.72 ;
    RECT 84.455 15.84 84.735 16.72 ;
    RECT 81.135 15.84 81.415 16.72 ;
    RECT 77.815 15.84 78.095 16.72 ;
    RECT 74.495 15.84 74.775 16.72 ;
    RECT 71.175 15.84 71.455 16.72 ;
    RECT 31.335 15.84 31.615 16.72 ;
    RECT 67.855 15.84 68.135 16.72 ;
    RECT 28.015 15.84 28.295 16.72 ;
    RECT 24.695 15.84 24.975 16.72 ;
    RECT 21.375 15.84 21.655 16.72 ;
    RECT 18.055 15.84 18.335 16.72 ;
    RECT 14.735 15.84 15.015 16.72 ;
    RECT 11.415 15.84 11.695 16.72 ;
    RECT 8.095 15.84 8.375 16.72 ;
    RECT 4.775 15.84 5.055 16.72 ;
    RECT 164.135 15.84 164.415 16.72 ;
    RECT 1.455 15.84 1.735 16.72 ;
    RECT 160.815 15.84 161.095 16.72 ;
    RECT 157.495 15.84 157.775 16.72 ;
    RECT 154.175 15.84 154.455 16.72 ;
    RECT 150.855 15.84 151.135 16.72 ;
    RECT 147.535 15.84 147.815 16.72 ;
    RECT 144.215 15.84 144.495 16.72 ;
    RECT 140.895 15.84 141.175 16.72 ;
    RECT 137.575 15.84 137.855 16.72 ;
    RECT 134.255 15.84 134.535 16.72 ;
    RECT 64.535 15.84 64.815 16.72 ;
    RECT 61.215 46.8 61.495 47.68 ;
    RECT 57.895 46.8 58.175 47.68 ;
    RECT 54.575 46.8 54.855 47.68 ;
    RECT 51.255 46.8 51.535 47.68 ;
    RECT 47.935 46.8 48.215 47.68 ;
    RECT 44.615 46.8 44.895 47.68 ;
    RECT 41.295 46.8 41.575 47.68 ;
    RECT 37.975 46.8 38.255 47.68 ;
    RECT 34.655 46.8 34.935 47.68 ;
    RECT 130.935 46.8 131.215 47.68 ;
    RECT 127.615 46.8 127.895 47.68 ;
    RECT 124.295 46.8 124.575 47.68 ;
    RECT 120.975 46.8 121.255 47.68 ;
    RECT 117.655 46.8 117.935 47.68 ;
    RECT 114.335 46.8 114.615 47.68 ;
    RECT 111.015 46.8 111.295 47.68 ;
    RECT 107.695 46.8 107.975 47.68 ;
    RECT 104.375 46.8 104.655 47.68 ;
    RECT 101.055 46.8 101.335 47.68 ;
    RECT 170.775 46.8 171.055 47.68 ;
    RECT 167.455 46.8 167.735 47.68 ;
    RECT 97.735 46.8 98.015 47.68 ;
    RECT 94.415 46.8 94.695 47.68 ;
    RECT 91.095 46.8 91.375 47.68 ;
    RECT 87.775 46.8 88.055 47.68 ;
    RECT 84.455 46.8 84.735 47.68 ;
    RECT 81.135 46.8 81.415 47.68 ;
    RECT 77.815 46.8 78.095 47.68 ;
    RECT 74.495 46.8 74.775 47.68 ;
    RECT 71.175 46.8 71.455 47.68 ;
    RECT 31.335 46.8 31.615 47.68 ;
    RECT 67.855 46.8 68.135 47.68 ;
    RECT 28.015 46.8 28.295 47.68 ;
    RECT 24.695 46.8 24.975 47.68 ;
    RECT 21.375 46.8 21.655 47.68 ;
    RECT 18.055 46.8 18.335 47.68 ;
    RECT 14.735 46.8 15.015 47.68 ;
    RECT 11.415 46.8 11.695 47.68 ;
    RECT 8.095 46.8 8.375 47.68 ;
    RECT 4.775 46.8 5.055 47.68 ;
    RECT 164.135 46.8 164.415 47.68 ;
    RECT 1.455 46.8 1.735 47.68 ;
    RECT 160.815 46.8 161.095 47.68 ;
    RECT 157.495 46.8 157.775 47.68 ;
    RECT 154.175 46.8 154.455 47.68 ;
    RECT 150.855 46.8 151.135 47.68 ;
    RECT 147.535 46.8 147.815 47.68 ;
    RECT 144.215 46.8 144.495 47.68 ;
    RECT 140.895 46.8 141.175 47.68 ;
    RECT 137.575 46.8 137.855 47.68 ;
    RECT 134.255 46.8 134.535 47.68 ;
    RECT 64.535 46.8 64.815 47.68 ;
    RECT 61.215 15.12 61.495 16.0 ;
    RECT 57.895 15.12 58.175 16.0 ;
    RECT 54.575 15.12 54.855 16.0 ;
    RECT 51.255 15.12 51.535 16.0 ;
    RECT 47.935 15.12 48.215 16.0 ;
    RECT 44.615 15.12 44.895 16.0 ;
    RECT 41.295 15.12 41.575 16.0 ;
    RECT 37.975 15.12 38.255 16.0 ;
    RECT 34.655 15.12 34.935 16.0 ;
    RECT 130.935 15.12 131.215 16.0 ;
    RECT 127.615 15.12 127.895 16.0 ;
    RECT 124.295 15.12 124.575 16.0 ;
    RECT 120.975 15.12 121.255 16.0 ;
    RECT 117.655 15.12 117.935 16.0 ;
    RECT 114.335 15.12 114.615 16.0 ;
    RECT 111.015 15.12 111.295 16.0 ;
    RECT 107.695 15.12 107.975 16.0 ;
    RECT 104.375 15.12 104.655 16.0 ;
    RECT 101.055 15.12 101.335 16.0 ;
    RECT 170.775 15.12 171.055 16.0 ;
    RECT 167.455 15.12 167.735 16.0 ;
    RECT 97.735 15.12 98.015 16.0 ;
    RECT 94.415 15.12 94.695 16.0 ;
    RECT 91.095 15.12 91.375 16.0 ;
    RECT 87.775 15.12 88.055 16.0 ;
    RECT 84.455 15.12 84.735 16.0 ;
    RECT 81.135 15.12 81.415 16.0 ;
    RECT 77.815 15.12 78.095 16.0 ;
    RECT 74.495 15.12 74.775 16.0 ;
    RECT 71.175 15.12 71.455 16.0 ;
    RECT 31.335 15.12 31.615 16.0 ;
    RECT 67.855 15.12 68.135 16.0 ;
    RECT 28.015 15.12 28.295 16.0 ;
    RECT 24.695 15.12 24.975 16.0 ;
    RECT 21.375 15.12 21.655 16.0 ;
    RECT 18.055 15.12 18.335 16.0 ;
    RECT 14.735 15.12 15.015 16.0 ;
    RECT 11.415 15.12 11.695 16.0 ;
    RECT 8.095 15.12 8.375 16.0 ;
    RECT 4.775 15.12 5.055 16.0 ;
    RECT 164.135 15.12 164.415 16.0 ;
    RECT 1.455 15.12 1.735 16.0 ;
    RECT 160.815 15.12 161.095 16.0 ;
    RECT 157.495 15.12 157.775 16.0 ;
    RECT 154.175 15.12 154.455 16.0 ;
    RECT 150.855 15.12 151.135 16.0 ;
    RECT 147.535 15.12 147.815 16.0 ;
    RECT 144.215 15.12 144.495 16.0 ;
    RECT 140.895 15.12 141.175 16.0 ;
    RECT 137.575 15.12 137.855 16.0 ;
    RECT 134.255 15.12 134.535 16.0 ;
    RECT 64.535 15.12 64.815 16.0 ;
    RECT 61.215 46.08 61.495 46.96 ;
    RECT 57.895 46.08 58.175 46.96 ;
    RECT 54.575 46.08 54.855 46.96 ;
    RECT 51.255 46.08 51.535 46.96 ;
    RECT 47.935 46.08 48.215 46.96 ;
    RECT 44.615 46.08 44.895 46.96 ;
    RECT 41.295 46.08 41.575 46.96 ;
    RECT 37.975 46.08 38.255 46.96 ;
    RECT 34.655 46.08 34.935 46.96 ;
    RECT 130.935 46.08 131.215 46.96 ;
    RECT 127.615 46.08 127.895 46.96 ;
    RECT 124.295 46.08 124.575 46.96 ;
    RECT 120.975 46.08 121.255 46.96 ;
    RECT 117.655 46.08 117.935 46.96 ;
    RECT 114.335 46.08 114.615 46.96 ;
    RECT 111.015 46.08 111.295 46.96 ;
    RECT 107.695 46.08 107.975 46.96 ;
    RECT 104.375 46.08 104.655 46.96 ;
    RECT 101.055 46.08 101.335 46.96 ;
    RECT 170.775 46.08 171.055 46.96 ;
    RECT 167.455 46.08 167.735 46.96 ;
    RECT 97.735 46.08 98.015 46.96 ;
    RECT 94.415 46.08 94.695 46.96 ;
    RECT 91.095 46.08 91.375 46.96 ;
    RECT 87.775 46.08 88.055 46.96 ;
    RECT 84.455 46.08 84.735 46.96 ;
    RECT 81.135 46.08 81.415 46.96 ;
    RECT 77.815 46.08 78.095 46.96 ;
    RECT 74.495 46.08 74.775 46.96 ;
    RECT 71.175 46.08 71.455 46.96 ;
    RECT 31.335 46.08 31.615 46.96 ;
    RECT 67.855 46.08 68.135 46.96 ;
    RECT 28.015 46.08 28.295 46.96 ;
    RECT 24.695 46.08 24.975 46.96 ;
    RECT 21.375 46.08 21.655 46.96 ;
    RECT 18.055 46.08 18.335 46.96 ;
    RECT 14.735 46.08 15.015 46.96 ;
    RECT 11.415 46.08 11.695 46.96 ;
    RECT 8.095 46.08 8.375 46.96 ;
    RECT 4.775 46.08 5.055 46.96 ;
    RECT 164.135 46.08 164.415 46.96 ;
    RECT 1.455 46.08 1.735 46.96 ;
    RECT 160.815 46.08 161.095 46.96 ;
    RECT 157.495 46.08 157.775 46.96 ;
    RECT 154.175 46.08 154.455 46.96 ;
    RECT 150.855 46.08 151.135 46.96 ;
    RECT 147.535 46.08 147.815 46.96 ;
    RECT 144.215 46.08 144.495 46.96 ;
    RECT 140.895 46.08 141.175 46.96 ;
    RECT 137.575 46.08 137.855 46.96 ;
    RECT 134.255 46.08 134.535 46.96 ;
    RECT 64.535 46.08 64.815 46.96 ;
    RECT 61.215 14.4 61.495 15.28 ;
    RECT 57.895 14.4 58.175 15.28 ;
    RECT 54.575 14.4 54.855 15.28 ;
    RECT 51.255 14.4 51.535 15.28 ;
    RECT 47.935 14.4 48.215 15.28 ;
    RECT 44.615 14.4 44.895 15.28 ;
    RECT 41.295 14.4 41.575 15.28 ;
    RECT 37.975 14.4 38.255 15.28 ;
    RECT 34.655 14.4 34.935 15.28 ;
    RECT 130.935 14.4 131.215 15.28 ;
    RECT 127.615 14.4 127.895 15.28 ;
    RECT 124.295 14.4 124.575 15.28 ;
    RECT 120.975 14.4 121.255 15.28 ;
    RECT 117.655 14.4 117.935 15.28 ;
    RECT 114.335 14.4 114.615 15.28 ;
    RECT 111.015 14.4 111.295 15.28 ;
    RECT 107.695 14.4 107.975 15.28 ;
    RECT 104.375 14.4 104.655 15.28 ;
    RECT 101.055 14.4 101.335 15.28 ;
    RECT 170.775 14.4 171.055 15.28 ;
    RECT 167.455 14.4 167.735 15.28 ;
    RECT 97.735 14.4 98.015 15.28 ;
    RECT 94.415 14.4 94.695 15.28 ;
    RECT 91.095 14.4 91.375 15.28 ;
    RECT 87.775 14.4 88.055 15.28 ;
    RECT 84.455 14.4 84.735 15.28 ;
    RECT 81.135 14.4 81.415 15.28 ;
    RECT 77.815 14.4 78.095 15.28 ;
    RECT 74.495 14.4 74.775 15.28 ;
    RECT 71.175 14.4 71.455 15.28 ;
    RECT 31.335 14.4 31.615 15.28 ;
    RECT 67.855 14.4 68.135 15.28 ;
    RECT 28.015 14.4 28.295 15.28 ;
    RECT 24.695 14.4 24.975 15.28 ;
    RECT 21.375 14.4 21.655 15.28 ;
    RECT 18.055 14.4 18.335 15.28 ;
    RECT 14.735 14.4 15.015 15.28 ;
    RECT 11.415 14.4 11.695 15.28 ;
    RECT 8.095 14.4 8.375 15.28 ;
    RECT 4.775 14.4 5.055 15.28 ;
    RECT 164.135 14.4 164.415 15.28 ;
    RECT 1.455 14.4 1.735 15.28 ;
    RECT 160.815 14.4 161.095 15.28 ;
    RECT 157.495 14.4 157.775 15.28 ;
    RECT 154.175 14.4 154.455 15.28 ;
    RECT 150.855 14.4 151.135 15.28 ;
    RECT 147.535 14.4 147.815 15.28 ;
    RECT 144.215 14.4 144.495 15.28 ;
    RECT 140.895 14.4 141.175 15.28 ;
    RECT 137.575 14.4 137.855 15.28 ;
    RECT 134.255 14.4 134.535 15.28 ;
    RECT 64.535 14.4 64.815 15.28 ;
    RECT 61.215 45.36 61.495 46.24 ;
    RECT 57.895 45.36 58.175 46.24 ;
    RECT 54.575 45.36 54.855 46.24 ;
    RECT 51.255 45.36 51.535 46.24 ;
    RECT 47.935 45.36 48.215 46.24 ;
    RECT 44.615 45.36 44.895 46.24 ;
    RECT 41.295 45.36 41.575 46.24 ;
    RECT 37.975 45.36 38.255 46.24 ;
    RECT 34.655 45.36 34.935 46.24 ;
    RECT 130.935 45.36 131.215 46.24 ;
    RECT 127.615 45.36 127.895 46.24 ;
    RECT 124.295 45.36 124.575 46.24 ;
    RECT 120.975 45.36 121.255 46.24 ;
    RECT 117.655 45.36 117.935 46.24 ;
    RECT 114.335 45.36 114.615 46.24 ;
    RECT 111.015 45.36 111.295 46.24 ;
    RECT 107.695 45.36 107.975 46.24 ;
    RECT 104.375 45.36 104.655 46.24 ;
    RECT 101.055 45.36 101.335 46.24 ;
    RECT 170.775 45.36 171.055 46.24 ;
    RECT 167.455 45.36 167.735 46.24 ;
    RECT 97.735 45.36 98.015 46.24 ;
    RECT 94.415 45.36 94.695 46.24 ;
    RECT 91.095 45.36 91.375 46.24 ;
    RECT 87.775 45.36 88.055 46.24 ;
    RECT 84.455 45.36 84.735 46.24 ;
    RECT 81.135 45.36 81.415 46.24 ;
    RECT 77.815 45.36 78.095 46.24 ;
    RECT 74.495 45.36 74.775 46.24 ;
    RECT 71.175 45.36 71.455 46.24 ;
    RECT 31.335 45.36 31.615 46.24 ;
    RECT 67.855 45.36 68.135 46.24 ;
    RECT 28.015 45.36 28.295 46.24 ;
    RECT 24.695 45.36 24.975 46.24 ;
    RECT 21.375 45.36 21.655 46.24 ;
    RECT 18.055 45.36 18.335 46.24 ;
    RECT 14.735 45.36 15.015 46.24 ;
    RECT 11.415 45.36 11.695 46.24 ;
    RECT 8.095 45.36 8.375 46.24 ;
    RECT 4.775 45.36 5.055 46.24 ;
    RECT 164.135 45.36 164.415 46.24 ;
    RECT 1.455 45.36 1.735 46.24 ;
    RECT 160.815 45.36 161.095 46.24 ;
    RECT 157.495 45.36 157.775 46.24 ;
    RECT 154.175 45.36 154.455 46.24 ;
    RECT 150.855 45.36 151.135 46.24 ;
    RECT 147.535 45.36 147.815 46.24 ;
    RECT 144.215 45.36 144.495 46.24 ;
    RECT 140.895 45.36 141.175 46.24 ;
    RECT 137.575 45.36 137.855 46.24 ;
    RECT 134.255 45.36 134.535 46.24 ;
    RECT 64.535 45.36 64.815 46.24 ;
    RECT 61.215 13.68 61.495 14.56 ;
    RECT 57.895 13.68 58.175 14.56 ;
    RECT 54.575 13.68 54.855 14.56 ;
    RECT 51.255 13.68 51.535 14.56 ;
    RECT 47.935 13.68 48.215 14.56 ;
    RECT 44.615 13.68 44.895 14.56 ;
    RECT 41.295 13.68 41.575 14.56 ;
    RECT 37.975 13.68 38.255 14.56 ;
    RECT 34.655 13.68 34.935 14.56 ;
    RECT 130.935 13.68 131.215 14.56 ;
    RECT 127.615 13.68 127.895 14.56 ;
    RECT 124.295 13.68 124.575 14.56 ;
    RECT 120.975 13.68 121.255 14.56 ;
    RECT 117.655 13.68 117.935 14.56 ;
    RECT 114.335 13.68 114.615 14.56 ;
    RECT 111.015 13.68 111.295 14.56 ;
    RECT 107.695 13.68 107.975 14.56 ;
    RECT 104.375 13.68 104.655 14.56 ;
    RECT 101.055 13.68 101.335 14.56 ;
    RECT 170.775 13.68 171.055 14.56 ;
    RECT 167.455 13.68 167.735 14.56 ;
    RECT 97.735 13.68 98.015 14.56 ;
    RECT 94.415 13.68 94.695 14.56 ;
    RECT 91.095 13.68 91.375 14.56 ;
    RECT 87.775 13.68 88.055 14.56 ;
    RECT 84.455 13.68 84.735 14.56 ;
    RECT 81.135 13.68 81.415 14.56 ;
    RECT 77.815 13.68 78.095 14.56 ;
    RECT 74.495 13.68 74.775 14.56 ;
    RECT 71.175 13.68 71.455 14.56 ;
    RECT 31.335 13.68 31.615 14.56 ;
    RECT 67.855 13.68 68.135 14.56 ;
    RECT 28.015 13.68 28.295 14.56 ;
    RECT 24.695 13.68 24.975 14.56 ;
    RECT 21.375 13.68 21.655 14.56 ;
    RECT 18.055 13.68 18.335 14.56 ;
    RECT 14.735 13.68 15.015 14.56 ;
    RECT 11.415 13.68 11.695 14.56 ;
    RECT 8.095 13.68 8.375 14.56 ;
    RECT 4.775 13.68 5.055 14.56 ;
    RECT 164.135 13.68 164.415 14.56 ;
    RECT 1.455 13.68 1.735 14.56 ;
    RECT 160.815 13.68 161.095 14.56 ;
    RECT 157.495 13.68 157.775 14.56 ;
    RECT 154.175 13.68 154.455 14.56 ;
    RECT 150.855 13.68 151.135 14.56 ;
    RECT 147.535 13.68 147.815 14.56 ;
    RECT 144.215 13.68 144.495 14.56 ;
    RECT 140.895 13.68 141.175 14.56 ;
    RECT 137.575 13.68 137.855 14.56 ;
    RECT 134.255 13.68 134.535 14.56 ;
    RECT 64.535 13.68 64.815 14.56 ;
    RECT 61.215 44.64 61.495 45.52 ;
    RECT 57.895 44.64 58.175 45.52 ;
    RECT 54.575 44.64 54.855 45.52 ;
    RECT 51.255 44.64 51.535 45.52 ;
    RECT 47.935 44.64 48.215 45.52 ;
    RECT 44.615 44.64 44.895 45.52 ;
    RECT 41.295 44.64 41.575 45.52 ;
    RECT 37.975 44.64 38.255 45.52 ;
    RECT 34.655 44.64 34.935 45.52 ;
    RECT 130.935 44.64 131.215 45.52 ;
    RECT 127.615 44.64 127.895 45.52 ;
    RECT 124.295 44.64 124.575 45.52 ;
    RECT 120.975 44.64 121.255 45.52 ;
    RECT 117.655 44.64 117.935 45.52 ;
    RECT 114.335 44.64 114.615 45.52 ;
    RECT 111.015 44.64 111.295 45.52 ;
    RECT 107.695 44.64 107.975 45.52 ;
    RECT 104.375 44.64 104.655 45.52 ;
    RECT 101.055 44.64 101.335 45.52 ;
    RECT 170.775 44.64 171.055 45.52 ;
    RECT 167.455 44.64 167.735 45.52 ;
    RECT 97.735 44.64 98.015 45.52 ;
    RECT 94.415 44.64 94.695 45.52 ;
    RECT 91.095 44.64 91.375 45.52 ;
    RECT 87.775 44.64 88.055 45.52 ;
    RECT 84.455 44.64 84.735 45.52 ;
    RECT 81.135 44.64 81.415 45.52 ;
    RECT 77.815 44.64 78.095 45.52 ;
    RECT 74.495 44.64 74.775 45.52 ;
    RECT 71.175 44.64 71.455 45.52 ;
    RECT 31.335 44.64 31.615 45.52 ;
    RECT 67.855 44.64 68.135 45.52 ;
    RECT 28.015 44.64 28.295 45.52 ;
    RECT 24.695 44.64 24.975 45.52 ;
    RECT 21.375 44.64 21.655 45.52 ;
    RECT 18.055 44.64 18.335 45.52 ;
    RECT 14.735 44.64 15.015 45.52 ;
    RECT 11.415 44.64 11.695 45.52 ;
    RECT 8.095 44.64 8.375 45.52 ;
    RECT 4.775 44.64 5.055 45.52 ;
    RECT 164.135 44.64 164.415 45.52 ;
    RECT 1.455 44.64 1.735 45.52 ;
    RECT 160.815 44.64 161.095 45.52 ;
    RECT 157.495 44.64 157.775 45.52 ;
    RECT 154.175 44.64 154.455 45.52 ;
    RECT 150.855 44.64 151.135 45.52 ;
    RECT 147.535 44.64 147.815 45.52 ;
    RECT 144.215 44.64 144.495 45.52 ;
    RECT 140.895 44.64 141.175 45.52 ;
    RECT 137.575 44.64 137.855 45.52 ;
    RECT 134.255 44.64 134.535 45.52 ;
    RECT 64.535 44.64 64.815 45.52 ;
    RECT 61.215 12.96 61.495 13.84 ;
    RECT 57.895 12.96 58.175 13.84 ;
    RECT 54.575 12.96 54.855 13.84 ;
    RECT 51.255 12.96 51.535 13.84 ;
    RECT 47.935 12.96 48.215 13.84 ;
    RECT 44.615 12.96 44.895 13.84 ;
    RECT 41.295 12.96 41.575 13.84 ;
    RECT 37.975 12.96 38.255 13.84 ;
    RECT 34.655 12.96 34.935 13.84 ;
    RECT 130.935 12.96 131.215 13.84 ;
    RECT 127.615 12.96 127.895 13.84 ;
    RECT 124.295 12.96 124.575 13.84 ;
    RECT 120.975 12.96 121.255 13.84 ;
    RECT 117.655 12.96 117.935 13.84 ;
    RECT 114.335 12.96 114.615 13.84 ;
    RECT 111.015 12.96 111.295 13.84 ;
    RECT 107.695 12.96 107.975 13.84 ;
    RECT 104.375 12.96 104.655 13.84 ;
    RECT 101.055 12.96 101.335 13.84 ;
    RECT 170.775 12.96 171.055 13.84 ;
    RECT 167.455 12.96 167.735 13.84 ;
    RECT 97.735 12.96 98.015 13.84 ;
    RECT 94.415 12.96 94.695 13.84 ;
    RECT 91.095 12.96 91.375 13.84 ;
    RECT 87.775 12.96 88.055 13.84 ;
    RECT 84.455 12.96 84.735 13.84 ;
    RECT 81.135 12.96 81.415 13.84 ;
    RECT 77.815 12.96 78.095 13.84 ;
    RECT 74.495 12.96 74.775 13.84 ;
    RECT 71.175 12.96 71.455 13.84 ;
    RECT 31.335 12.96 31.615 13.84 ;
    RECT 67.855 12.96 68.135 13.84 ;
    RECT 28.015 12.96 28.295 13.84 ;
    RECT 24.695 12.96 24.975 13.84 ;
    RECT 21.375 12.96 21.655 13.84 ;
    RECT 18.055 12.96 18.335 13.84 ;
    RECT 14.735 12.96 15.015 13.84 ;
    RECT 11.415 12.96 11.695 13.84 ;
    RECT 8.095 12.96 8.375 13.84 ;
    RECT 4.775 12.96 5.055 13.84 ;
    RECT 164.135 12.96 164.415 13.84 ;
    RECT 1.455 12.96 1.735 13.84 ;
    RECT 160.815 12.96 161.095 13.84 ;
    RECT 157.495 12.96 157.775 13.84 ;
    RECT 154.175 12.96 154.455 13.84 ;
    RECT 150.855 12.96 151.135 13.84 ;
    RECT 147.535 12.96 147.815 13.84 ;
    RECT 144.215 12.96 144.495 13.84 ;
    RECT 140.895 12.96 141.175 13.84 ;
    RECT 137.575 12.96 137.855 13.84 ;
    RECT 134.255 12.96 134.535 13.84 ;
    RECT 64.535 12.96 64.815 13.84 ;
    RECT 61.215 43.92 61.495 44.8 ;
    RECT 57.895 43.92 58.175 44.8 ;
    RECT 54.575 43.92 54.855 44.8 ;
    RECT 51.255 43.92 51.535 44.8 ;
    RECT 47.935 43.92 48.215 44.8 ;
    RECT 44.615 43.92 44.895 44.8 ;
    RECT 41.295 43.92 41.575 44.8 ;
    RECT 37.975 43.92 38.255 44.8 ;
    RECT 34.655 43.92 34.935 44.8 ;
    RECT 130.935 43.92 131.215 44.8 ;
    RECT 127.615 43.92 127.895 44.8 ;
    RECT 124.295 43.92 124.575 44.8 ;
    RECT 120.975 43.92 121.255 44.8 ;
    RECT 117.655 43.92 117.935 44.8 ;
    RECT 114.335 43.92 114.615 44.8 ;
    RECT 111.015 43.92 111.295 44.8 ;
    RECT 107.695 43.92 107.975 44.8 ;
    RECT 104.375 43.92 104.655 44.8 ;
    RECT 101.055 43.92 101.335 44.8 ;
    RECT 170.775 43.92 171.055 44.8 ;
    RECT 167.455 43.92 167.735 44.8 ;
    RECT 97.735 43.92 98.015 44.8 ;
    RECT 94.415 43.92 94.695 44.8 ;
    RECT 91.095 43.92 91.375 44.8 ;
    RECT 87.775 43.92 88.055 44.8 ;
    RECT 84.455 43.92 84.735 44.8 ;
    RECT 81.135 43.92 81.415 44.8 ;
    RECT 77.815 43.92 78.095 44.8 ;
    RECT 74.495 43.92 74.775 44.8 ;
    RECT 71.175 43.92 71.455 44.8 ;
    RECT 31.335 43.92 31.615 44.8 ;
    RECT 67.855 43.92 68.135 44.8 ;
    RECT 28.015 43.92 28.295 44.8 ;
    RECT 24.695 43.92 24.975 44.8 ;
    RECT 21.375 43.92 21.655 44.8 ;
    RECT 18.055 43.92 18.335 44.8 ;
    RECT 14.735 43.92 15.015 44.8 ;
    RECT 11.415 43.92 11.695 44.8 ;
    RECT 8.095 43.92 8.375 44.8 ;
    RECT 4.775 43.92 5.055 44.8 ;
    RECT 164.135 43.92 164.415 44.8 ;
    RECT 1.455 43.92 1.735 44.8 ;
    RECT 160.815 43.92 161.095 44.8 ;
    RECT 157.495 43.92 157.775 44.8 ;
    RECT 154.175 43.92 154.455 44.8 ;
    RECT 150.855 43.92 151.135 44.8 ;
    RECT 147.535 43.92 147.815 44.8 ;
    RECT 144.215 43.92 144.495 44.8 ;
    RECT 140.895 43.92 141.175 44.8 ;
    RECT 137.575 43.92 137.855 44.8 ;
    RECT 134.255 43.92 134.535 44.8 ;
    RECT 64.535 43.92 64.815 44.8 ;
    RECT 61.215 12.24 61.495 13.12 ;
    RECT 57.895 12.24 58.175 13.12 ;
    RECT 54.575 12.24 54.855 13.12 ;
    RECT 51.255 12.24 51.535 13.12 ;
    RECT 47.935 12.24 48.215 13.12 ;
    RECT 44.615 12.24 44.895 13.12 ;
    RECT 41.295 12.24 41.575 13.12 ;
    RECT 37.975 12.24 38.255 13.12 ;
    RECT 34.655 12.24 34.935 13.12 ;
    RECT 130.935 12.24 131.215 13.12 ;
    RECT 127.615 12.24 127.895 13.12 ;
    RECT 124.295 12.24 124.575 13.12 ;
    RECT 120.975 12.24 121.255 13.12 ;
    RECT 117.655 12.24 117.935 13.12 ;
    RECT 114.335 12.24 114.615 13.12 ;
    RECT 111.015 12.24 111.295 13.12 ;
    RECT 107.695 12.24 107.975 13.12 ;
    RECT 104.375 12.24 104.655 13.12 ;
    RECT 101.055 12.24 101.335 13.12 ;
    RECT 170.775 12.24 171.055 13.12 ;
    RECT 167.455 12.24 167.735 13.12 ;
    RECT 97.735 12.24 98.015 13.12 ;
    RECT 94.415 12.24 94.695 13.12 ;
    RECT 91.095 12.24 91.375 13.12 ;
    RECT 87.775 12.24 88.055 13.12 ;
    RECT 84.455 12.24 84.735 13.12 ;
    RECT 81.135 12.24 81.415 13.12 ;
    RECT 77.815 12.24 78.095 13.12 ;
    RECT 74.495 12.24 74.775 13.12 ;
    RECT 71.175 12.24 71.455 13.12 ;
    RECT 31.335 12.24 31.615 13.12 ;
    RECT 67.855 12.24 68.135 13.12 ;
    RECT 28.015 12.24 28.295 13.12 ;
    RECT 24.695 12.24 24.975 13.12 ;
    RECT 21.375 12.24 21.655 13.12 ;
    RECT 18.055 12.24 18.335 13.12 ;
    RECT 14.735 12.24 15.015 13.12 ;
    RECT 11.415 12.24 11.695 13.12 ;
    RECT 8.095 12.24 8.375 13.12 ;
    RECT 4.775 12.24 5.055 13.12 ;
    RECT 164.135 12.24 164.415 13.12 ;
    RECT 1.455 12.24 1.735 13.12 ;
    RECT 160.815 12.24 161.095 13.12 ;
    RECT 157.495 12.24 157.775 13.12 ;
    RECT 154.175 12.24 154.455 13.12 ;
    RECT 150.855 12.24 151.135 13.12 ;
    RECT 147.535 12.24 147.815 13.12 ;
    RECT 144.215 12.24 144.495 13.12 ;
    RECT 140.895 12.24 141.175 13.12 ;
    RECT 137.575 12.24 137.855 13.12 ;
    RECT 134.255 12.24 134.535 13.12 ;
    RECT 64.535 12.24 64.815 13.12 ;
    RECT 61.215 43.2 61.495 44.08 ;
    RECT 57.895 43.2 58.175 44.08 ;
    RECT 54.575 43.2 54.855 44.08 ;
    RECT 51.255 43.2 51.535 44.08 ;
    RECT 47.935 43.2 48.215 44.08 ;
    RECT 44.615 43.2 44.895 44.08 ;
    RECT 41.295 43.2 41.575 44.08 ;
    RECT 37.975 43.2 38.255 44.08 ;
    RECT 34.655 43.2 34.935 44.08 ;
    RECT 130.935 43.2 131.215 44.08 ;
    RECT 127.615 43.2 127.895 44.08 ;
    RECT 124.295 43.2 124.575 44.08 ;
    RECT 120.975 43.2 121.255 44.08 ;
    RECT 117.655 43.2 117.935 44.08 ;
    RECT 114.335 43.2 114.615 44.08 ;
    RECT 111.015 43.2 111.295 44.08 ;
    RECT 107.695 43.2 107.975 44.08 ;
    RECT 104.375 43.2 104.655 44.08 ;
    RECT 101.055 43.2 101.335 44.08 ;
    RECT 170.775 43.2 171.055 44.08 ;
    RECT 167.455 43.2 167.735 44.08 ;
    RECT 97.735 43.2 98.015 44.08 ;
    RECT 94.415 43.2 94.695 44.08 ;
    RECT 91.095 43.2 91.375 44.08 ;
    RECT 87.775 43.2 88.055 44.08 ;
    RECT 84.455 43.2 84.735 44.08 ;
    RECT 81.135 43.2 81.415 44.08 ;
    RECT 77.815 43.2 78.095 44.08 ;
    RECT 74.495 43.2 74.775 44.08 ;
    RECT 71.175 43.2 71.455 44.08 ;
    RECT 31.335 43.2 31.615 44.08 ;
    RECT 67.855 43.2 68.135 44.08 ;
    RECT 28.015 43.2 28.295 44.08 ;
    RECT 24.695 43.2 24.975 44.08 ;
    RECT 21.375 43.2 21.655 44.08 ;
    RECT 18.055 43.2 18.335 44.08 ;
    RECT 14.735 43.2 15.015 44.08 ;
    RECT 11.415 43.2 11.695 44.08 ;
    RECT 8.095 43.2 8.375 44.08 ;
    RECT 4.775 43.2 5.055 44.08 ;
    RECT 164.135 43.2 164.415 44.08 ;
    RECT 1.455 43.2 1.735 44.08 ;
    RECT 160.815 43.2 161.095 44.08 ;
    RECT 157.495 43.2 157.775 44.08 ;
    RECT 154.175 43.2 154.455 44.08 ;
    RECT 150.855 43.2 151.135 44.08 ;
    RECT 147.535 43.2 147.815 44.08 ;
    RECT 144.215 43.2 144.495 44.08 ;
    RECT 140.895 43.2 141.175 44.08 ;
    RECT 137.575 43.2 137.855 44.08 ;
    RECT 134.255 43.2 134.535 44.08 ;
    RECT 64.535 43.2 64.815 44.08 ;
    RECT 61.215 42.48 61.495 43.36 ;
    RECT 57.895 42.48 58.175 43.36 ;
    RECT 54.575 42.48 54.855 43.36 ;
    RECT 51.255 42.48 51.535 43.36 ;
    RECT 47.935 42.48 48.215 43.36 ;
    RECT 44.615 42.48 44.895 43.36 ;
    RECT 41.295 42.48 41.575 43.36 ;
    RECT 37.975 42.48 38.255 43.36 ;
    RECT 34.655 42.48 34.935 43.36 ;
    RECT 130.935 42.48 131.215 43.36 ;
    RECT 127.615 42.48 127.895 43.36 ;
    RECT 124.295 42.48 124.575 43.36 ;
    RECT 120.975 42.48 121.255 43.36 ;
    RECT 117.655 42.48 117.935 43.36 ;
    RECT 114.335 42.48 114.615 43.36 ;
    RECT 111.015 42.48 111.295 43.36 ;
    RECT 107.695 42.48 107.975 43.36 ;
    RECT 104.375 42.48 104.655 43.36 ;
    RECT 101.055 42.48 101.335 43.36 ;
    RECT 170.775 42.48 171.055 43.36 ;
    RECT 167.455 42.48 167.735 43.36 ;
    RECT 97.735 42.48 98.015 43.36 ;
    RECT 94.415 42.48 94.695 43.36 ;
    RECT 91.095 42.48 91.375 43.36 ;
    RECT 87.775 42.48 88.055 43.36 ;
    RECT 84.455 42.48 84.735 43.36 ;
    RECT 81.135 42.48 81.415 43.36 ;
    RECT 77.815 42.48 78.095 43.36 ;
    RECT 74.495 42.48 74.775 43.36 ;
    RECT 71.175 42.48 71.455 43.36 ;
    RECT 31.335 42.48 31.615 43.36 ;
    RECT 67.855 42.48 68.135 43.36 ;
    RECT 28.015 42.48 28.295 43.36 ;
    RECT 24.695 42.48 24.975 43.36 ;
    RECT 21.375 42.48 21.655 43.36 ;
    RECT 18.055 42.48 18.335 43.36 ;
    RECT 14.735 42.48 15.015 43.36 ;
    RECT 11.415 42.48 11.695 43.36 ;
    RECT 8.095 42.48 8.375 43.36 ;
    RECT 4.775 42.48 5.055 43.36 ;
    RECT 164.135 42.48 164.415 43.36 ;
    RECT 1.455 42.48 1.735 43.36 ;
    RECT 160.815 42.48 161.095 43.36 ;
    RECT 157.495 42.48 157.775 43.36 ;
    RECT 154.175 42.48 154.455 43.36 ;
    RECT 150.855 42.48 151.135 43.36 ;
    RECT 147.535 42.48 147.815 43.36 ;
    RECT 144.215 42.48 144.495 43.36 ;
    RECT 140.895 42.48 141.175 43.36 ;
    RECT 137.575 42.48 137.855 43.36 ;
    RECT 134.255 42.48 134.535 43.36 ;
    RECT 64.535 42.48 64.815 43.36 ;
    RECT 61.215 41.76 61.495 42.64 ;
    RECT 57.895 41.76 58.175 42.64 ;
    RECT 54.575 41.76 54.855 42.64 ;
    RECT 51.255 41.76 51.535 42.64 ;
    RECT 47.935 41.76 48.215 42.64 ;
    RECT 44.615 41.76 44.895 42.64 ;
    RECT 41.295 41.76 41.575 42.64 ;
    RECT 37.975 41.76 38.255 42.64 ;
    RECT 34.655 41.76 34.935 42.64 ;
    RECT 130.935 41.76 131.215 42.64 ;
    RECT 127.615 41.76 127.895 42.64 ;
    RECT 124.295 41.76 124.575 42.64 ;
    RECT 120.975 41.76 121.255 42.64 ;
    RECT 117.655 41.76 117.935 42.64 ;
    RECT 114.335 41.76 114.615 42.64 ;
    RECT 111.015 41.76 111.295 42.64 ;
    RECT 107.695 41.76 107.975 42.64 ;
    RECT 104.375 41.76 104.655 42.64 ;
    RECT 101.055 41.76 101.335 42.64 ;
    RECT 170.775 41.76 171.055 42.64 ;
    RECT 167.455 41.76 167.735 42.64 ;
    RECT 97.735 41.76 98.015 42.64 ;
    RECT 94.415 41.76 94.695 42.64 ;
    RECT 91.095 41.76 91.375 42.64 ;
    RECT 87.775 41.76 88.055 42.64 ;
    RECT 84.455 41.76 84.735 42.64 ;
    RECT 81.135 41.76 81.415 42.64 ;
    RECT 77.815 41.76 78.095 42.64 ;
    RECT 74.495 41.76 74.775 42.64 ;
    RECT 71.175 41.76 71.455 42.64 ;
    RECT 31.335 41.76 31.615 42.64 ;
    RECT 67.855 41.76 68.135 42.64 ;
    RECT 28.015 41.76 28.295 42.64 ;
    RECT 24.695 41.76 24.975 42.64 ;
    RECT 21.375 41.76 21.655 42.64 ;
    RECT 18.055 41.76 18.335 42.64 ;
    RECT 14.735 41.76 15.015 42.64 ;
    RECT 11.415 41.76 11.695 42.64 ;
    RECT 8.095 41.76 8.375 42.64 ;
    RECT 4.775 41.76 5.055 42.64 ;
    RECT 164.135 41.76 164.415 42.64 ;
    RECT 1.455 41.76 1.735 42.64 ;
    RECT 160.815 41.76 161.095 42.64 ;
    RECT 157.495 41.76 157.775 42.64 ;
    RECT 154.175 41.76 154.455 42.64 ;
    RECT 150.855 41.76 151.135 42.64 ;
    RECT 147.535 41.76 147.815 42.64 ;
    RECT 144.215 41.76 144.495 42.64 ;
    RECT 140.895 41.76 141.175 42.64 ;
    RECT 137.575 41.76 137.855 42.64 ;
    RECT 134.255 41.76 134.535 42.64 ;
    RECT 64.535 41.76 64.815 42.64 ;
    RECT 61.215 41.04 61.495 41.92 ;
    RECT 57.895 41.04 58.175 41.92 ;
    RECT 54.575 41.04 54.855 41.92 ;
    RECT 51.255 41.04 51.535 41.92 ;
    RECT 47.935 41.04 48.215 41.92 ;
    RECT 44.615 41.04 44.895 41.92 ;
    RECT 41.295 41.04 41.575 41.92 ;
    RECT 37.975 41.04 38.255 41.92 ;
    RECT 34.655 41.04 34.935 41.92 ;
    RECT 130.935 41.04 131.215 41.92 ;
    RECT 127.615 41.04 127.895 41.92 ;
    RECT 124.295 41.04 124.575 41.92 ;
    RECT 120.975 41.04 121.255 41.92 ;
    RECT 117.655 41.04 117.935 41.92 ;
    RECT 114.335 41.04 114.615 41.92 ;
    RECT 111.015 41.04 111.295 41.92 ;
    RECT 107.695 41.04 107.975 41.92 ;
    RECT 104.375 41.04 104.655 41.92 ;
    RECT 101.055 41.04 101.335 41.92 ;
    RECT 170.775 41.04 171.055 41.92 ;
    RECT 167.455 41.04 167.735 41.92 ;
    RECT 97.735 41.04 98.015 41.92 ;
    RECT 94.415 41.04 94.695 41.92 ;
    RECT 91.095 41.04 91.375 41.92 ;
    RECT 87.775 41.04 88.055 41.92 ;
    RECT 84.455 41.04 84.735 41.92 ;
    RECT 81.135 41.04 81.415 41.92 ;
    RECT 77.815 41.04 78.095 41.92 ;
    RECT 74.495 41.04 74.775 41.92 ;
    RECT 71.175 41.04 71.455 41.92 ;
    RECT 31.335 41.04 31.615 41.92 ;
    RECT 67.855 41.04 68.135 41.92 ;
    RECT 28.015 41.04 28.295 41.92 ;
    RECT 24.695 41.04 24.975 41.92 ;
    RECT 21.375 41.04 21.655 41.92 ;
    RECT 18.055 41.04 18.335 41.92 ;
    RECT 14.735 41.04 15.015 41.92 ;
    RECT 11.415 41.04 11.695 41.92 ;
    RECT 8.095 41.04 8.375 41.92 ;
    RECT 4.775 41.04 5.055 41.92 ;
    RECT 164.135 41.04 164.415 41.92 ;
    RECT 1.455 41.04 1.735 41.92 ;
    RECT 160.815 41.04 161.095 41.92 ;
    RECT 157.495 41.04 157.775 41.92 ;
    RECT 154.175 41.04 154.455 41.92 ;
    RECT 150.855 41.04 151.135 41.92 ;
    RECT 147.535 41.04 147.815 41.92 ;
    RECT 144.215 41.04 144.495 41.92 ;
    RECT 140.895 41.04 141.175 41.92 ;
    RECT 137.575 41.04 137.855 41.92 ;
    RECT 134.255 41.04 134.535 41.92 ;
    RECT 64.535 41.04 64.815 41.92 ;
    RECT 61.215 40.32 61.495 41.2 ;
    RECT 57.895 40.32 58.175 41.2 ;
    RECT 54.575 40.32 54.855 41.2 ;
    RECT 51.255 40.32 51.535 41.2 ;
    RECT 47.935 40.32 48.215 41.2 ;
    RECT 44.615 40.32 44.895 41.2 ;
    RECT 41.295 40.32 41.575 41.2 ;
    RECT 37.975 40.32 38.255 41.2 ;
    RECT 34.655 40.32 34.935 41.2 ;
    RECT 130.935 40.32 131.215 41.2 ;
    RECT 127.615 40.32 127.895 41.2 ;
    RECT 124.295 40.32 124.575 41.2 ;
    RECT 120.975 40.32 121.255 41.2 ;
    RECT 117.655 40.32 117.935 41.2 ;
    RECT 114.335 40.32 114.615 41.2 ;
    RECT 111.015 40.32 111.295 41.2 ;
    RECT 107.695 40.32 107.975 41.2 ;
    RECT 104.375 40.32 104.655 41.2 ;
    RECT 101.055 40.32 101.335 41.2 ;
    RECT 170.775 40.32 171.055 41.2 ;
    RECT 167.455 40.32 167.735 41.2 ;
    RECT 97.735 40.32 98.015 41.2 ;
    RECT 94.415 40.32 94.695 41.2 ;
    RECT 91.095 40.32 91.375 41.2 ;
    RECT 87.775 40.32 88.055 41.2 ;
    RECT 84.455 40.32 84.735 41.2 ;
    RECT 81.135 40.32 81.415 41.2 ;
    RECT 77.815 40.32 78.095 41.2 ;
    RECT 74.495 40.32 74.775 41.2 ;
    RECT 71.175 40.32 71.455 41.2 ;
    RECT 31.335 40.32 31.615 41.2 ;
    RECT 67.855 40.32 68.135 41.2 ;
    RECT 28.015 40.32 28.295 41.2 ;
    RECT 24.695 40.32 24.975 41.2 ;
    RECT 21.375 40.32 21.655 41.2 ;
    RECT 18.055 40.32 18.335 41.2 ;
    RECT 14.735 40.32 15.015 41.2 ;
    RECT 11.415 40.32 11.695 41.2 ;
    RECT 8.095 40.32 8.375 41.2 ;
    RECT 4.775 40.32 5.055 41.2 ;
    RECT 164.135 40.32 164.415 41.2 ;
    RECT 1.455 40.32 1.735 41.2 ;
    RECT 160.815 40.32 161.095 41.2 ;
    RECT 157.495 40.32 157.775 41.2 ;
    RECT 154.175 40.32 154.455 41.2 ;
    RECT 150.855 40.32 151.135 41.2 ;
    RECT 147.535 40.32 147.815 41.2 ;
    RECT 144.215 40.32 144.495 41.2 ;
    RECT 140.895 40.32 141.175 41.2 ;
    RECT 137.575 40.32 137.855 41.2 ;
    RECT 134.255 40.32 134.535 41.2 ;
    RECT 64.535 40.32 64.815 41.2 ;
    RECT 61.215 39.6 61.495 40.48 ;
    RECT 57.895 39.6 58.175 40.48 ;
    RECT 54.575 39.6 54.855 40.48 ;
    RECT 51.255 39.6 51.535 40.48 ;
    RECT 47.935 39.6 48.215 40.48 ;
    RECT 44.615 39.6 44.895 40.48 ;
    RECT 41.295 39.6 41.575 40.48 ;
    RECT 37.975 39.6 38.255 40.48 ;
    RECT 34.655 39.6 34.935 40.48 ;
    RECT 130.935 39.6 131.215 40.48 ;
    RECT 127.615 39.6 127.895 40.48 ;
    RECT 124.295 39.6 124.575 40.48 ;
    RECT 120.975 39.6 121.255 40.48 ;
    RECT 117.655 39.6 117.935 40.48 ;
    RECT 114.335 39.6 114.615 40.48 ;
    RECT 111.015 39.6 111.295 40.48 ;
    RECT 107.695 39.6 107.975 40.48 ;
    RECT 104.375 39.6 104.655 40.48 ;
    RECT 101.055 39.6 101.335 40.48 ;
    RECT 170.775 39.6 171.055 40.48 ;
    RECT 167.455 39.6 167.735 40.48 ;
    RECT 97.735 39.6 98.015 40.48 ;
    RECT 94.415 39.6 94.695 40.48 ;
    RECT 91.095 39.6 91.375 40.48 ;
    RECT 87.775 39.6 88.055 40.48 ;
    RECT 84.455 39.6 84.735 40.48 ;
    RECT 81.135 39.6 81.415 40.48 ;
    RECT 77.815 39.6 78.095 40.48 ;
    RECT 74.495 39.6 74.775 40.48 ;
    RECT 71.175 39.6 71.455 40.48 ;
    RECT 31.335 39.6 31.615 40.48 ;
    RECT 67.855 39.6 68.135 40.48 ;
    RECT 28.015 39.6 28.295 40.48 ;
    RECT 24.695 39.6 24.975 40.48 ;
    RECT 21.375 39.6 21.655 40.48 ;
    RECT 18.055 39.6 18.335 40.48 ;
    RECT 14.735 39.6 15.015 40.48 ;
    RECT 11.415 39.6 11.695 40.48 ;
    RECT 8.095 39.6 8.375 40.48 ;
    RECT 4.775 39.6 5.055 40.48 ;
    RECT 164.135 39.6 164.415 40.48 ;
    RECT 1.455 39.6 1.735 40.48 ;
    RECT 160.815 39.6 161.095 40.48 ;
    RECT 157.495 39.6 157.775 40.48 ;
    RECT 154.175 39.6 154.455 40.48 ;
    RECT 150.855 39.6 151.135 40.48 ;
    RECT 147.535 39.6 147.815 40.48 ;
    RECT 144.215 39.6 144.495 40.48 ;
    RECT 140.895 39.6 141.175 40.48 ;
    RECT 137.575 39.6 137.855 40.48 ;
    RECT 134.255 39.6 134.535 40.48 ;
    RECT 64.535 39.6 64.815 40.48 ;
    RECT 61.215 58.34 61.495 59.22 ;
    RECT 57.895 58.34 58.175 59.22 ;
    RECT 54.575 58.34 54.855 59.22 ;
    RECT 170.775 58.34 171.055 59.22 ;
    RECT 51.255 58.34 51.535 59.22 ;
    RECT 47.935 58.34 48.215 59.22 ;
    RECT 44.615 58.34 44.895 59.22 ;
    RECT 41.295 58.34 41.575 59.22 ;
    RECT 37.975 58.34 38.255 59.22 ;
    RECT 34.655 58.34 34.935 59.22 ;
    RECT 1.455 58.34 1.735 59.22 ;
    RECT 130.935 58.34 131.215 59.22 ;
    RECT 127.615 58.34 127.895 59.22 ;
    RECT 124.295 58.34 124.575 59.22 ;
    RECT 120.975 58.34 121.255 59.22 ;
    RECT 117.655 58.34 117.935 59.22 ;
    RECT 114.335 58.34 114.615 59.22 ;
    RECT 111.015 58.34 111.295 59.22 ;
    RECT 107.695 58.34 107.975 59.22 ;
    RECT 104.375 58.34 104.655 59.22 ;
    RECT 101.055 58.34 101.335 59.22 ;
    RECT 167.455 58.34 167.735 59.22 ;
    RECT 97.735 58.34 98.015 59.22 ;
    RECT 94.415 58.34 94.695 59.22 ;
    RECT 91.095 58.34 91.375 59.22 ;
    RECT 87.775 58.34 88.055 59.22 ;
    RECT 84.455 58.34 84.735 59.22 ;
    RECT 81.135 58.34 81.415 59.22 ;
    RECT 77.815 58.34 78.095 59.22 ;
    RECT 74.495 58.34 74.775 59.22 ;
    RECT 71.175 58.34 71.455 59.22 ;
    RECT 31.335 58.34 31.615 59.22 ;
    RECT 67.855 58.34 68.135 59.22 ;
    RECT 28.015 58.34 28.295 59.22 ;
    RECT 24.695 58.34 24.975 59.22 ;
    RECT 21.375 58.34 21.655 59.22 ;
    RECT 18.055 58.34 18.335 59.22 ;
    RECT 14.735 58.34 15.015 59.22 ;
    RECT 11.415 58.34 11.695 59.22 ;
    RECT 8.095 58.34 8.375 59.22 ;
    RECT 4.775 58.34 5.055 59.22 ;
    RECT 164.135 58.34 164.415 59.22 ;
    RECT 160.815 58.34 161.095 59.22 ;
    RECT 157.495 58.34 157.775 59.22 ;
    RECT 154.175 58.34 154.455 59.22 ;
    RECT 150.855 58.34 151.135 59.22 ;
    RECT 147.535 58.34 147.815 59.22 ;
    RECT 144.215 58.34 144.495 59.22 ;
    RECT 140.895 58.34 141.175 59.22 ;
    RECT 137.575 58.34 137.855 59.22 ;
    RECT 134.255 58.34 134.535 59.22 ;
    RECT 64.535 58.34 64.815 59.22 ;
    RECT 61.215 38.88 61.495 39.76 ;
    RECT 57.895 38.88 58.175 39.76 ;
    RECT 54.575 38.88 54.855 39.76 ;
    RECT 51.255 38.88 51.535 39.76 ;
    RECT 47.935 38.88 48.215 39.76 ;
    RECT 44.615 38.88 44.895 39.76 ;
    RECT 41.295 38.88 41.575 39.76 ;
    RECT 37.975 38.88 38.255 39.76 ;
    RECT 34.655 38.88 34.935 39.76 ;
    RECT 130.935 38.88 131.215 39.76 ;
    RECT 127.615 38.88 127.895 39.76 ;
    RECT 124.295 38.88 124.575 39.76 ;
    RECT 120.975 38.88 121.255 39.76 ;
    RECT 117.655 38.88 117.935 39.76 ;
    RECT 114.335 38.88 114.615 39.76 ;
    RECT 111.015 38.88 111.295 39.76 ;
    RECT 107.695 38.88 107.975 39.76 ;
    RECT 104.375 38.88 104.655 39.76 ;
    RECT 101.055 38.88 101.335 39.76 ;
    RECT 170.775 38.88 171.055 39.76 ;
    RECT 167.455 38.88 167.735 39.76 ;
    RECT 97.735 38.88 98.015 39.76 ;
    RECT 94.415 38.88 94.695 39.76 ;
    RECT 91.095 38.88 91.375 39.76 ;
    RECT 87.775 38.88 88.055 39.76 ;
    RECT 84.455 38.88 84.735 39.76 ;
    RECT 81.135 38.88 81.415 39.76 ;
    RECT 77.815 38.88 78.095 39.76 ;
    RECT 74.495 38.88 74.775 39.76 ;
    RECT 71.175 38.88 71.455 39.76 ;
    RECT 31.335 38.88 31.615 39.76 ;
    RECT 67.855 38.88 68.135 39.76 ;
    RECT 28.015 38.88 28.295 39.76 ;
    RECT 24.695 38.88 24.975 39.76 ;
    RECT 21.375 38.88 21.655 39.76 ;
    RECT 18.055 38.88 18.335 39.76 ;
    RECT 14.735 38.88 15.015 39.76 ;
    RECT 11.415 38.88 11.695 39.76 ;
    RECT 8.095 38.88 8.375 39.76 ;
    RECT 4.775 38.88 5.055 39.76 ;
    RECT 164.135 38.88 164.415 39.76 ;
    RECT 1.455 38.88 1.735 39.76 ;
    RECT 160.815 38.88 161.095 39.76 ;
    RECT 157.495 38.88 157.775 39.76 ;
    RECT 154.175 38.88 154.455 39.76 ;
    RECT 150.855 38.88 151.135 39.76 ;
    RECT 147.535 38.88 147.815 39.76 ;
    RECT 144.215 38.88 144.495 39.76 ;
    RECT 140.895 38.88 141.175 39.76 ;
    RECT 137.575 38.88 137.855 39.76 ;
    RECT 134.255 38.88 134.535 39.76 ;
    RECT 64.535 38.88 64.815 39.76 ;
    RECT 61.215 38.16 61.495 39.04 ;
    RECT 57.895 38.16 58.175 39.04 ;
    RECT 54.575 38.16 54.855 39.04 ;
    RECT 51.255 38.16 51.535 39.04 ;
    RECT 47.935 38.16 48.215 39.04 ;
    RECT 44.615 38.16 44.895 39.04 ;
    RECT 41.295 38.16 41.575 39.04 ;
    RECT 37.975 38.16 38.255 39.04 ;
    RECT 34.655 38.16 34.935 39.04 ;
    RECT 130.935 38.16 131.215 39.04 ;
    RECT 127.615 38.16 127.895 39.04 ;
    RECT 124.295 38.16 124.575 39.04 ;
    RECT 120.975 38.16 121.255 39.04 ;
    RECT 117.655 38.16 117.935 39.04 ;
    RECT 114.335 38.16 114.615 39.04 ;
    RECT 111.015 38.16 111.295 39.04 ;
    RECT 107.695 38.16 107.975 39.04 ;
    RECT 104.375 38.16 104.655 39.04 ;
    RECT 101.055 38.16 101.335 39.04 ;
    RECT 170.775 38.16 171.055 39.04 ;
    RECT 167.455 38.16 167.735 39.04 ;
    RECT 97.735 38.16 98.015 39.04 ;
    RECT 94.415 38.16 94.695 39.04 ;
    RECT 91.095 38.16 91.375 39.04 ;
    RECT 87.775 38.16 88.055 39.04 ;
    RECT 84.455 38.16 84.735 39.04 ;
    RECT 81.135 38.16 81.415 39.04 ;
    RECT 77.815 38.16 78.095 39.04 ;
    RECT 74.495 38.16 74.775 39.04 ;
    RECT 71.175 38.16 71.455 39.04 ;
    RECT 31.335 38.16 31.615 39.04 ;
    RECT 67.855 38.16 68.135 39.04 ;
    RECT 28.015 38.16 28.295 39.04 ;
    RECT 24.695 38.16 24.975 39.04 ;
    RECT 21.375 38.16 21.655 39.04 ;
    RECT 18.055 38.16 18.335 39.04 ;
    RECT 14.735 38.16 15.015 39.04 ;
    RECT 11.415 38.16 11.695 39.04 ;
    RECT 8.095 38.16 8.375 39.04 ;
    RECT 4.775 38.16 5.055 39.04 ;
    RECT 164.135 38.16 164.415 39.04 ;
    RECT 1.455 38.16 1.735 39.04 ;
    RECT 160.815 38.16 161.095 39.04 ;
    RECT 157.495 38.16 157.775 39.04 ;
    RECT 154.175 38.16 154.455 39.04 ;
    RECT 150.855 38.16 151.135 39.04 ;
    RECT 147.535 38.16 147.815 39.04 ;
    RECT 144.215 38.16 144.495 39.04 ;
    RECT 140.895 38.16 141.175 39.04 ;
    RECT 137.575 38.16 137.855 39.04 ;
    RECT 134.255 38.16 134.535 39.04 ;
    RECT 64.535 38.16 64.815 39.04 ;
    RECT 61.215 37.44 61.495 38.32 ;
    RECT 57.895 37.44 58.175 38.32 ;
    RECT 54.575 37.44 54.855 38.32 ;
    RECT 51.255 37.44 51.535 38.32 ;
    RECT 47.935 37.44 48.215 38.32 ;
    RECT 44.615 37.44 44.895 38.32 ;
    RECT 41.295 37.44 41.575 38.32 ;
    RECT 37.975 37.44 38.255 38.32 ;
    RECT 34.655 37.44 34.935 38.32 ;
    RECT 130.935 37.44 131.215 38.32 ;
    RECT 127.615 37.44 127.895 38.32 ;
    RECT 124.295 37.44 124.575 38.32 ;
    RECT 120.975 37.44 121.255 38.32 ;
    RECT 117.655 37.44 117.935 38.32 ;
    RECT 114.335 37.44 114.615 38.32 ;
    RECT 111.015 37.44 111.295 38.32 ;
    RECT 107.695 37.44 107.975 38.32 ;
    RECT 104.375 37.44 104.655 38.32 ;
    RECT 101.055 37.44 101.335 38.32 ;
    RECT 170.775 37.44 171.055 38.32 ;
    RECT 167.455 37.44 167.735 38.32 ;
    RECT 97.735 37.44 98.015 38.32 ;
    RECT 94.415 37.44 94.695 38.32 ;
    RECT 91.095 37.44 91.375 38.32 ;
    RECT 87.775 37.44 88.055 38.32 ;
    RECT 84.455 37.44 84.735 38.32 ;
    RECT 81.135 37.44 81.415 38.32 ;
    RECT 77.815 37.44 78.095 38.32 ;
    RECT 74.495 37.44 74.775 38.32 ;
    RECT 71.175 37.44 71.455 38.32 ;
    RECT 31.335 37.44 31.615 38.32 ;
    RECT 67.855 37.44 68.135 38.32 ;
    RECT 28.015 37.44 28.295 38.32 ;
    RECT 24.695 37.44 24.975 38.32 ;
    RECT 21.375 37.44 21.655 38.32 ;
    RECT 18.055 37.44 18.335 38.32 ;
    RECT 14.735 37.44 15.015 38.32 ;
    RECT 11.415 37.44 11.695 38.32 ;
    RECT 8.095 37.44 8.375 38.32 ;
    RECT 4.775 37.44 5.055 38.32 ;
    RECT 164.135 37.44 164.415 38.32 ;
    RECT 1.455 37.44 1.735 38.32 ;
    RECT 160.815 37.44 161.095 38.32 ;
    RECT 157.495 37.44 157.775 38.32 ;
    RECT 154.175 37.44 154.455 38.32 ;
    RECT 150.855 37.44 151.135 38.32 ;
    RECT 147.535 37.44 147.815 38.32 ;
    RECT 144.215 37.44 144.495 38.32 ;
    RECT 140.895 37.44 141.175 38.32 ;
    RECT 137.575 37.44 137.855 38.32 ;
    RECT 134.255 37.44 134.535 38.32 ;
    RECT 64.535 37.44 64.815 38.32 ;
    RECT 61.215 36.72 61.495 37.6 ;
    RECT 57.895 36.72 58.175 37.6 ;
    RECT 54.575 36.72 54.855 37.6 ;
    RECT 51.255 36.72 51.535 37.6 ;
    RECT 47.935 36.72 48.215 37.6 ;
    RECT 44.615 36.72 44.895 37.6 ;
    RECT 41.295 36.72 41.575 37.6 ;
    RECT 37.975 36.72 38.255 37.6 ;
    RECT 34.655 36.72 34.935 37.6 ;
    RECT 130.935 36.72 131.215 37.6 ;
    RECT 127.615 36.72 127.895 37.6 ;
    RECT 124.295 36.72 124.575 37.6 ;
    RECT 120.975 36.72 121.255 37.6 ;
    RECT 117.655 36.72 117.935 37.6 ;
    RECT 114.335 36.72 114.615 37.6 ;
    RECT 111.015 36.72 111.295 37.6 ;
    RECT 107.695 36.72 107.975 37.6 ;
    RECT 104.375 36.72 104.655 37.6 ;
    RECT 101.055 36.72 101.335 37.6 ;
    RECT 170.775 36.72 171.055 37.6 ;
    RECT 167.455 36.72 167.735 37.6 ;
    RECT 97.735 36.72 98.015 37.6 ;
    RECT 94.415 36.72 94.695 37.6 ;
    RECT 91.095 36.72 91.375 37.6 ;
    RECT 87.775 36.72 88.055 37.6 ;
    RECT 84.455 36.72 84.735 37.6 ;
    RECT 81.135 36.72 81.415 37.6 ;
    RECT 77.815 36.72 78.095 37.6 ;
    RECT 74.495 36.72 74.775 37.6 ;
    RECT 71.175 36.72 71.455 37.6 ;
    RECT 31.335 36.72 31.615 37.6 ;
    RECT 67.855 36.72 68.135 37.6 ;
    RECT 28.015 36.72 28.295 37.6 ;
    RECT 24.695 36.72 24.975 37.6 ;
    RECT 21.375 36.72 21.655 37.6 ;
    RECT 18.055 36.72 18.335 37.6 ;
    RECT 14.735 36.72 15.015 37.6 ;
    RECT 11.415 36.72 11.695 37.6 ;
    RECT 8.095 36.72 8.375 37.6 ;
    RECT 4.775 36.72 5.055 37.6 ;
    RECT 164.135 36.72 164.415 37.6 ;
    RECT 1.455 36.72 1.735 37.6 ;
    RECT 160.815 36.72 161.095 37.6 ;
    RECT 157.495 36.72 157.775 37.6 ;
    RECT 154.175 36.72 154.455 37.6 ;
    RECT 150.855 36.72 151.135 37.6 ;
    RECT 147.535 36.72 147.815 37.6 ;
    RECT 144.215 36.72 144.495 37.6 ;
    RECT 140.895 36.72 141.175 37.6 ;
    RECT 137.575 36.72 137.855 37.6 ;
    RECT 134.255 36.72 134.535 37.6 ;
    RECT 64.535 36.72 64.815 37.6 ;
    RECT 61.215 36.0 61.495 36.88 ;
    RECT 57.895 36.0 58.175 36.88 ;
    RECT 54.575 36.0 54.855 36.88 ;
    RECT 51.255 36.0 51.535 36.88 ;
    RECT 47.935 36.0 48.215 36.88 ;
    RECT 44.615 36.0 44.895 36.88 ;
    RECT 41.295 36.0 41.575 36.88 ;
    RECT 37.975 36.0 38.255 36.88 ;
    RECT 34.655 36.0 34.935 36.88 ;
    RECT 130.935 36.0 131.215 36.88 ;
    RECT 127.615 36.0 127.895 36.88 ;
    RECT 124.295 36.0 124.575 36.88 ;
    RECT 120.975 36.0 121.255 36.88 ;
    RECT 117.655 36.0 117.935 36.88 ;
    RECT 114.335 36.0 114.615 36.88 ;
    RECT 111.015 36.0 111.295 36.88 ;
    RECT 107.695 36.0 107.975 36.88 ;
    RECT 104.375 36.0 104.655 36.88 ;
    RECT 101.055 36.0 101.335 36.88 ;
    RECT 170.775 36.0 171.055 36.88 ;
    RECT 167.455 36.0 167.735 36.88 ;
    RECT 97.735 36.0 98.015 36.88 ;
    RECT 94.415 36.0 94.695 36.88 ;
    RECT 91.095 36.0 91.375 36.88 ;
    RECT 87.775 36.0 88.055 36.88 ;
    RECT 84.455 36.0 84.735 36.88 ;
    RECT 81.135 36.0 81.415 36.88 ;
    RECT 77.815 36.0 78.095 36.88 ;
    RECT 74.495 36.0 74.775 36.88 ;
    RECT 71.175 36.0 71.455 36.88 ;
    RECT 31.335 36.0 31.615 36.88 ;
    RECT 67.855 36.0 68.135 36.88 ;
    RECT 28.015 36.0 28.295 36.88 ;
    RECT 24.695 36.0 24.975 36.88 ;
    RECT 21.375 36.0 21.655 36.88 ;
    RECT 18.055 36.0 18.335 36.88 ;
    RECT 14.735 36.0 15.015 36.88 ;
    RECT 11.415 36.0 11.695 36.88 ;
    RECT 8.095 36.0 8.375 36.88 ;
    RECT 4.775 36.0 5.055 36.88 ;
    RECT 164.135 36.0 164.415 36.88 ;
    RECT 1.455 36.0 1.735 36.88 ;
    RECT 160.815 36.0 161.095 36.88 ;
    RECT 157.495 36.0 157.775 36.88 ;
    RECT 154.175 36.0 154.455 36.88 ;
    RECT 150.855 36.0 151.135 36.88 ;
    RECT 147.535 36.0 147.815 36.88 ;
    RECT 144.215 36.0 144.495 36.88 ;
    RECT 140.895 36.0 141.175 36.88 ;
    RECT 137.575 36.0 137.855 36.88 ;
    RECT 134.255 36.0 134.535 36.88 ;
    RECT 64.535 36.0 64.815 36.88 ;
    RECT 61.215 33.12 61.495 34.0 ;
    RECT 57.895 33.12 58.175 34.0 ;
    RECT 54.575 33.12 54.855 34.0 ;
    RECT 51.255 33.12 51.535 34.0 ;
    RECT 47.935 33.12 48.215 34.0 ;
    RECT 44.615 33.12 44.895 34.0 ;
    RECT 41.295 33.12 41.575 34.0 ;
    RECT 37.975 33.12 38.255 34.0 ;
    RECT 34.655 33.12 34.935 34.0 ;
    RECT 130.935 33.12 131.215 34.0 ;
    RECT 127.615 33.12 127.895 34.0 ;
    RECT 124.295 33.12 124.575 34.0 ;
    RECT 120.975 33.12 121.255 34.0 ;
    RECT 117.655 33.12 117.935 34.0 ;
    RECT 114.335 33.12 114.615 34.0 ;
    RECT 111.015 33.12 111.295 34.0 ;
    RECT 107.695 33.12 107.975 34.0 ;
    RECT 104.375 33.12 104.655 34.0 ;
    RECT 101.055 33.12 101.335 34.0 ;
    RECT 170.775 33.12 171.055 34.0 ;
    RECT 167.455 33.12 167.735 34.0 ;
    RECT 97.735 33.12 98.015 34.0 ;
    RECT 94.415 33.12 94.695 34.0 ;
    RECT 91.095 33.12 91.375 34.0 ;
    RECT 87.775 33.12 88.055 34.0 ;
    RECT 84.455 33.12 84.735 34.0 ;
    RECT 81.135 33.12 81.415 34.0 ;
    RECT 77.815 33.12 78.095 34.0 ;
    RECT 74.495 33.12 74.775 34.0 ;
    RECT 71.175 33.12 71.455 34.0 ;
    RECT 31.335 33.12 31.615 34.0 ;
    RECT 67.855 33.12 68.135 34.0 ;
    RECT 28.015 33.12 28.295 34.0 ;
    RECT 24.695 33.12 24.975 34.0 ;
    RECT 21.375 33.12 21.655 34.0 ;
    RECT 18.055 33.12 18.335 34.0 ;
    RECT 14.735 33.12 15.015 34.0 ;
    RECT 11.415 33.12 11.695 34.0 ;
    RECT 8.095 33.12 8.375 34.0 ;
    RECT 4.775 33.12 5.055 34.0 ;
    RECT 164.135 33.12 164.415 34.0 ;
    RECT 1.455 33.12 1.735 34.0 ;
    RECT 160.815 33.12 161.095 34.0 ;
    RECT 157.495 33.12 157.775 34.0 ;
    RECT 154.175 33.12 154.455 34.0 ;
    RECT 150.855 33.12 151.135 34.0 ;
    RECT 147.535 33.12 147.815 34.0 ;
    RECT 144.215 33.12 144.495 34.0 ;
    RECT 140.895 33.12 141.175 34.0 ;
    RECT 137.575 33.12 137.855 34.0 ;
    RECT 134.255 33.12 134.535 34.0 ;
    RECT 64.535 33.12 64.815 34.0 ;
    RECT 61.215 32.4 61.495 33.28 ;
    RECT 57.895 32.4 58.175 33.28 ;
    RECT 54.575 32.4 54.855 33.28 ;
    RECT 51.255 32.4 51.535 33.28 ;
    RECT 47.935 32.4 48.215 33.28 ;
    RECT 44.615 32.4 44.895 33.28 ;
    RECT 41.295 32.4 41.575 33.28 ;
    RECT 37.975 32.4 38.255 33.28 ;
    RECT 34.655 32.4 34.935 33.28 ;
    RECT 130.935 32.4 131.215 33.28 ;
    RECT 127.615 32.4 127.895 33.28 ;
    RECT 124.295 32.4 124.575 33.28 ;
    RECT 120.975 32.4 121.255 33.28 ;
    RECT 117.655 32.4 117.935 33.28 ;
    RECT 114.335 32.4 114.615 33.28 ;
    RECT 111.015 32.4 111.295 33.28 ;
    RECT 107.695 32.4 107.975 33.28 ;
    RECT 104.375 32.4 104.655 33.28 ;
    RECT 101.055 32.4 101.335 33.28 ;
    RECT 170.775 32.4 171.055 33.28 ;
    RECT 167.455 32.4 167.735 33.28 ;
    RECT 97.735 32.4 98.015 33.28 ;
    RECT 94.415 32.4 94.695 33.28 ;
    RECT 91.095 32.4 91.375 33.28 ;
    RECT 87.775 32.4 88.055 33.28 ;
    RECT 84.455 32.4 84.735 33.28 ;
    RECT 81.135 32.4 81.415 33.28 ;
    RECT 77.815 32.4 78.095 33.28 ;
    RECT 74.495 32.4 74.775 33.28 ;
    RECT 71.175 32.4 71.455 33.28 ;
    RECT 31.335 32.4 31.615 33.28 ;
    RECT 67.855 32.4 68.135 33.28 ;
    RECT 28.015 32.4 28.295 33.28 ;
    RECT 24.695 32.4 24.975 33.28 ;
    RECT 21.375 32.4 21.655 33.28 ;
    RECT 18.055 32.4 18.335 33.28 ;
    RECT 14.735 32.4 15.015 33.28 ;
    RECT 11.415 32.4 11.695 33.28 ;
    RECT 8.095 32.4 8.375 33.28 ;
    RECT 4.775 32.4 5.055 33.28 ;
    RECT 164.135 32.4 164.415 33.28 ;
    RECT 1.455 32.4 1.735 33.28 ;
    RECT 160.815 32.4 161.095 33.28 ;
    RECT 157.495 32.4 157.775 33.28 ;
    RECT 154.175 32.4 154.455 33.28 ;
    RECT 150.855 32.4 151.135 33.28 ;
    RECT 147.535 32.4 147.815 33.28 ;
    RECT 144.215 32.4 144.495 33.28 ;
    RECT 140.895 32.4 141.175 33.28 ;
    RECT 137.575 32.4 137.855 33.28 ;
    RECT 134.255 32.4 134.535 33.28 ;
    RECT 64.535 32.4 64.815 33.28 ;
    RECT 61.215 31.68 61.495 32.56 ;
    RECT 57.895 31.68 58.175 32.56 ;
    RECT 54.575 31.68 54.855 32.56 ;
    RECT 51.255 31.68 51.535 32.56 ;
    RECT 47.935 31.68 48.215 32.56 ;
    RECT 44.615 31.68 44.895 32.56 ;
    RECT 41.295 31.68 41.575 32.56 ;
    RECT 37.975 31.68 38.255 32.56 ;
    RECT 34.655 31.68 34.935 32.56 ;
    RECT 130.935 31.68 131.215 32.56 ;
    RECT 127.615 31.68 127.895 32.56 ;
    RECT 124.295 31.68 124.575 32.56 ;
    RECT 120.975 31.68 121.255 32.56 ;
    RECT 117.655 31.68 117.935 32.56 ;
    RECT 114.335 31.68 114.615 32.56 ;
    RECT 111.015 31.68 111.295 32.56 ;
    RECT 107.695 31.68 107.975 32.56 ;
    RECT 104.375 31.68 104.655 32.56 ;
    RECT 101.055 31.68 101.335 32.56 ;
    RECT 170.775 31.68 171.055 32.56 ;
    RECT 167.455 31.68 167.735 32.56 ;
    RECT 97.735 31.68 98.015 32.56 ;
    RECT 94.415 31.68 94.695 32.56 ;
    RECT 91.095 31.68 91.375 32.56 ;
    RECT 87.775 31.68 88.055 32.56 ;
    RECT 84.455 31.68 84.735 32.56 ;
    RECT 81.135 31.68 81.415 32.56 ;
    RECT 77.815 31.68 78.095 32.56 ;
    RECT 74.495 31.68 74.775 32.56 ;
    RECT 71.175 31.68 71.455 32.56 ;
    RECT 31.335 31.68 31.615 32.56 ;
    RECT 67.855 31.68 68.135 32.56 ;
    RECT 28.015 31.68 28.295 32.56 ;
    RECT 24.695 31.68 24.975 32.56 ;
    RECT 21.375 31.68 21.655 32.56 ;
    RECT 18.055 31.68 18.335 32.56 ;
    RECT 14.735 31.68 15.015 32.56 ;
    RECT 11.415 31.68 11.695 32.56 ;
    RECT 8.095 31.68 8.375 32.56 ;
    RECT 4.775 31.68 5.055 32.56 ;
    RECT 164.135 31.68 164.415 32.56 ;
    RECT 1.455 31.68 1.735 32.56 ;
    RECT 160.815 31.68 161.095 32.56 ;
    RECT 157.495 31.68 157.775 32.56 ;
    RECT 154.175 31.68 154.455 32.56 ;
    RECT 150.855 31.68 151.135 32.56 ;
    RECT 147.535 31.68 147.815 32.56 ;
    RECT 144.215 31.68 144.495 32.56 ;
    RECT 140.895 31.68 141.175 32.56 ;
    RECT 137.575 31.68 137.855 32.56 ;
    RECT 134.255 31.68 134.535 32.56 ;
    RECT 64.535 31.68 64.815 32.56 ;
    RECT 61.215 30.96 61.495 31.84 ;
    RECT 57.895 30.96 58.175 31.84 ;
    RECT 54.575 30.96 54.855 31.84 ;
    RECT 51.255 30.96 51.535 31.84 ;
    RECT 47.935 30.96 48.215 31.84 ;
    RECT 44.615 30.96 44.895 31.84 ;
    RECT 41.295 30.96 41.575 31.84 ;
    RECT 37.975 30.96 38.255 31.84 ;
    RECT 34.655 30.96 34.935 31.84 ;
    RECT 130.935 30.96 131.215 31.84 ;
    RECT 127.615 30.96 127.895 31.84 ;
    RECT 124.295 30.96 124.575 31.84 ;
    RECT 120.975 30.96 121.255 31.84 ;
    RECT 117.655 30.96 117.935 31.84 ;
    RECT 114.335 30.96 114.615 31.84 ;
    RECT 111.015 30.96 111.295 31.84 ;
    RECT 107.695 30.96 107.975 31.84 ;
    RECT 104.375 30.96 104.655 31.84 ;
    RECT 101.055 30.96 101.335 31.84 ;
    RECT 170.775 30.96 171.055 31.84 ;
    RECT 167.455 30.96 167.735 31.84 ;
    RECT 97.735 30.96 98.015 31.84 ;
    RECT 94.415 30.96 94.695 31.84 ;
    RECT 91.095 30.96 91.375 31.84 ;
    RECT 87.775 30.96 88.055 31.84 ;
    RECT 84.455 30.96 84.735 31.84 ;
    RECT 81.135 30.96 81.415 31.84 ;
    RECT 77.815 30.96 78.095 31.84 ;
    RECT 74.495 30.96 74.775 31.84 ;
    RECT 71.175 30.96 71.455 31.84 ;
    RECT 31.335 30.96 31.615 31.84 ;
    RECT 67.855 30.96 68.135 31.84 ;
    RECT 28.015 30.96 28.295 31.84 ;
    RECT 24.695 30.96 24.975 31.84 ;
    RECT 21.375 30.96 21.655 31.84 ;
    RECT 18.055 30.96 18.335 31.84 ;
    RECT 14.735 30.96 15.015 31.84 ;
    RECT 11.415 30.96 11.695 31.84 ;
    RECT 8.095 30.96 8.375 31.84 ;
    RECT 4.775 30.96 5.055 31.84 ;
    RECT 164.135 30.96 164.415 31.84 ;
    RECT 1.455 30.96 1.735 31.84 ;
    RECT 160.815 30.96 161.095 31.84 ;
    RECT 157.495 30.96 157.775 31.84 ;
    RECT 154.175 30.96 154.455 31.84 ;
    RECT 150.855 30.96 151.135 31.84 ;
    RECT 147.535 30.96 147.815 31.84 ;
    RECT 144.215 30.96 144.495 31.84 ;
    RECT 140.895 30.96 141.175 31.84 ;
    RECT 137.575 30.96 137.855 31.84 ;
    RECT 134.255 30.96 134.535 31.84 ;
    RECT 64.535 30.96 64.815 31.84 ;
    RECT 61.215 30.24 61.495 31.12 ;
    RECT 57.895 30.24 58.175 31.12 ;
    RECT 54.575 30.24 54.855 31.12 ;
    RECT 51.255 30.24 51.535 31.12 ;
    RECT 47.935 30.24 48.215 31.12 ;
    RECT 44.615 30.24 44.895 31.12 ;
    RECT 41.295 30.24 41.575 31.12 ;
    RECT 37.975 30.24 38.255 31.12 ;
    RECT 34.655 30.24 34.935 31.12 ;
    RECT 130.935 30.24 131.215 31.12 ;
    RECT 127.615 30.24 127.895 31.12 ;
    RECT 124.295 30.24 124.575 31.12 ;
    RECT 120.975 30.24 121.255 31.12 ;
    RECT 117.655 30.24 117.935 31.12 ;
    RECT 114.335 30.24 114.615 31.12 ;
    RECT 111.015 30.24 111.295 31.12 ;
    RECT 107.695 30.24 107.975 31.12 ;
    RECT 104.375 30.24 104.655 31.12 ;
    RECT 101.055 30.24 101.335 31.12 ;
    RECT 170.775 30.24 171.055 31.12 ;
    RECT 167.455 30.24 167.735 31.12 ;
    RECT 97.735 30.24 98.015 31.12 ;
    RECT 94.415 30.24 94.695 31.12 ;
    RECT 91.095 30.24 91.375 31.12 ;
    RECT 87.775 30.24 88.055 31.12 ;
    RECT 84.455 30.24 84.735 31.12 ;
    RECT 81.135 30.24 81.415 31.12 ;
    RECT 77.815 30.24 78.095 31.12 ;
    RECT 74.495 30.24 74.775 31.12 ;
    RECT 71.175 30.24 71.455 31.12 ;
    RECT 31.335 30.24 31.615 31.12 ;
    RECT 67.855 30.24 68.135 31.12 ;
    RECT 28.015 30.24 28.295 31.12 ;
    RECT 24.695 30.24 24.975 31.12 ;
    RECT 21.375 30.24 21.655 31.12 ;
    RECT 18.055 30.24 18.335 31.12 ;
    RECT 14.735 30.24 15.015 31.12 ;
    RECT 11.415 30.24 11.695 31.12 ;
    RECT 8.095 30.24 8.375 31.12 ;
    RECT 4.775 30.24 5.055 31.12 ;
    RECT 164.135 30.24 164.415 31.12 ;
    RECT 1.455 30.24 1.735 31.12 ;
    RECT 160.815 30.24 161.095 31.12 ;
    RECT 157.495 30.24 157.775 31.12 ;
    RECT 154.175 30.24 154.455 31.12 ;
    RECT 150.855 30.24 151.135 31.12 ;
    RECT 147.535 30.24 147.815 31.12 ;
    RECT 144.215 30.24 144.495 31.12 ;
    RECT 140.895 30.24 141.175 31.12 ;
    RECT 137.575 30.24 137.855 31.12 ;
    RECT 134.255 30.24 134.535 31.12 ;
    RECT 64.535 30.24 64.815 31.12 ;
    RECT 61.215 29.52 61.495 30.4 ;
    RECT 57.895 29.52 58.175 30.4 ;
    RECT 54.575 29.52 54.855 30.4 ;
    RECT 51.255 29.52 51.535 30.4 ;
    RECT 47.935 29.52 48.215 30.4 ;
    RECT 44.615 29.52 44.895 30.4 ;
    RECT 41.295 29.52 41.575 30.4 ;
    RECT 37.975 29.52 38.255 30.4 ;
    RECT 34.655 29.52 34.935 30.4 ;
    RECT 130.935 29.52 131.215 30.4 ;
    RECT 127.615 29.52 127.895 30.4 ;
    RECT 124.295 29.52 124.575 30.4 ;
    RECT 120.975 29.52 121.255 30.4 ;
    RECT 117.655 29.52 117.935 30.4 ;
    RECT 114.335 29.52 114.615 30.4 ;
    RECT 111.015 29.52 111.295 30.4 ;
    RECT 107.695 29.52 107.975 30.4 ;
    RECT 104.375 29.52 104.655 30.4 ;
    RECT 101.055 29.52 101.335 30.4 ;
    RECT 170.775 29.52 171.055 30.4 ;
    RECT 167.455 29.52 167.735 30.4 ;
    RECT 97.735 29.52 98.015 30.4 ;
    RECT 94.415 29.52 94.695 30.4 ;
    RECT 91.095 29.52 91.375 30.4 ;
    RECT 87.775 29.52 88.055 30.4 ;
    RECT 84.455 29.52 84.735 30.4 ;
    RECT 81.135 29.52 81.415 30.4 ;
    RECT 77.815 29.52 78.095 30.4 ;
    RECT 74.495 29.52 74.775 30.4 ;
    RECT 71.175 29.52 71.455 30.4 ;
    RECT 31.335 29.52 31.615 30.4 ;
    RECT 67.855 29.52 68.135 30.4 ;
    RECT 28.015 29.52 28.295 30.4 ;
    RECT 24.695 29.52 24.975 30.4 ;
    RECT 21.375 29.52 21.655 30.4 ;
    RECT 18.055 29.52 18.335 30.4 ;
    RECT 14.735 29.52 15.015 30.4 ;
    RECT 11.415 29.52 11.695 30.4 ;
    RECT 8.095 29.52 8.375 30.4 ;
    RECT 4.775 29.52 5.055 30.4 ;
    RECT 164.135 29.52 164.415 30.4 ;
    RECT 1.455 29.52 1.735 30.4 ;
    RECT 160.815 29.52 161.095 30.4 ;
    RECT 157.495 29.52 157.775 30.4 ;
    RECT 154.175 29.52 154.455 30.4 ;
    RECT 150.855 29.52 151.135 30.4 ;
    RECT 147.535 29.52 147.815 30.4 ;
    RECT 144.215 29.52 144.495 30.4 ;
    RECT 140.895 29.52 141.175 30.4 ;
    RECT 137.575 29.52 137.855 30.4 ;
    RECT 134.255 29.52 134.535 30.4 ;
    RECT 64.535 29.52 64.815 30.4 ;
    RECT 61.215 28.8 61.495 29.68 ;
    RECT 57.895 28.8 58.175 29.68 ;
    RECT 54.575 28.8 54.855 29.68 ;
    RECT 51.255 28.8 51.535 29.68 ;
    RECT 47.935 28.8 48.215 29.68 ;
    RECT 44.615 28.8 44.895 29.68 ;
    RECT 41.295 28.8 41.575 29.68 ;
    RECT 37.975 28.8 38.255 29.68 ;
    RECT 34.655 28.8 34.935 29.68 ;
    RECT 130.935 28.8 131.215 29.68 ;
    RECT 127.615 28.8 127.895 29.68 ;
    RECT 124.295 28.8 124.575 29.68 ;
    RECT 120.975 28.8 121.255 29.68 ;
    RECT 117.655 28.8 117.935 29.68 ;
    RECT 114.335 28.8 114.615 29.68 ;
    RECT 111.015 28.8 111.295 29.68 ;
    RECT 107.695 28.8 107.975 29.68 ;
    RECT 104.375 28.8 104.655 29.68 ;
    RECT 101.055 28.8 101.335 29.68 ;
    RECT 170.775 28.8 171.055 29.68 ;
    RECT 167.455 28.8 167.735 29.68 ;
    RECT 97.735 28.8 98.015 29.68 ;
    RECT 94.415 28.8 94.695 29.68 ;
    RECT 91.095 28.8 91.375 29.68 ;
    RECT 87.775 28.8 88.055 29.68 ;
    RECT 84.455 28.8 84.735 29.68 ;
    RECT 81.135 28.8 81.415 29.68 ;
    RECT 77.815 28.8 78.095 29.68 ;
    RECT 74.495 28.8 74.775 29.68 ;
    RECT 71.175 28.8 71.455 29.68 ;
    RECT 31.335 28.8 31.615 29.68 ;
    RECT 67.855 28.8 68.135 29.68 ;
    RECT 28.015 28.8 28.295 29.68 ;
    RECT 24.695 28.8 24.975 29.68 ;
    RECT 21.375 28.8 21.655 29.68 ;
    RECT 18.055 28.8 18.335 29.68 ;
    RECT 14.735 28.8 15.015 29.68 ;
    RECT 11.415 28.8 11.695 29.68 ;
    RECT 8.095 28.8 8.375 29.68 ;
    RECT 4.775 28.8 5.055 29.68 ;
    RECT 164.135 28.8 164.415 29.68 ;
    RECT 1.455 28.8 1.735 29.68 ;
    RECT 160.815 28.8 161.095 29.68 ;
    RECT 157.495 28.8 157.775 29.68 ;
    RECT 154.175 28.8 154.455 29.68 ;
    RECT 150.855 28.8 151.135 29.68 ;
    RECT 147.535 28.8 147.815 29.68 ;
    RECT 144.215 28.8 144.495 29.68 ;
    RECT 140.895 28.8 141.175 29.68 ;
    RECT 137.575 28.8 137.855 29.68 ;
    RECT 134.255 28.8 134.535 29.68 ;
    RECT 64.535 28.8 64.815 29.68 ;
    RECT 61.215 28.08 61.495 28.96 ;
    RECT 57.895 28.08 58.175 28.96 ;
    RECT 54.575 28.08 54.855 28.96 ;
    RECT 51.255 28.08 51.535 28.96 ;
    RECT 47.935 28.08 48.215 28.96 ;
    RECT 44.615 28.08 44.895 28.96 ;
    RECT 41.295 28.08 41.575 28.96 ;
    RECT 37.975 28.08 38.255 28.96 ;
    RECT 34.655 28.08 34.935 28.96 ;
    RECT 130.935 28.08 131.215 28.96 ;
    RECT 127.615 28.08 127.895 28.96 ;
    RECT 124.295 28.08 124.575 28.96 ;
    RECT 120.975 28.08 121.255 28.96 ;
    RECT 117.655 28.08 117.935 28.96 ;
    RECT 114.335 28.08 114.615 28.96 ;
    RECT 111.015 28.08 111.295 28.96 ;
    RECT 107.695 28.08 107.975 28.96 ;
    RECT 104.375 28.08 104.655 28.96 ;
    RECT 101.055 28.08 101.335 28.96 ;
    RECT 170.775 28.08 171.055 28.96 ;
    RECT 167.455 28.08 167.735 28.96 ;
    RECT 97.735 28.08 98.015 28.96 ;
    RECT 94.415 28.08 94.695 28.96 ;
    RECT 91.095 28.08 91.375 28.96 ;
    RECT 87.775 28.08 88.055 28.96 ;
    RECT 84.455 28.08 84.735 28.96 ;
    RECT 81.135 28.08 81.415 28.96 ;
    RECT 77.815 28.08 78.095 28.96 ;
    RECT 74.495 28.08 74.775 28.96 ;
    RECT 71.175 28.08 71.455 28.96 ;
    RECT 31.335 28.08 31.615 28.96 ;
    RECT 67.855 28.08 68.135 28.96 ;
    RECT 28.015 28.08 28.295 28.96 ;
    RECT 24.695 28.08 24.975 28.96 ;
    RECT 21.375 28.08 21.655 28.96 ;
    RECT 18.055 28.08 18.335 28.96 ;
    RECT 14.735 28.08 15.015 28.96 ;
    RECT 11.415 28.08 11.695 28.96 ;
    RECT 8.095 28.08 8.375 28.96 ;
    RECT 4.775 28.08 5.055 28.96 ;
    RECT 164.135 28.08 164.415 28.96 ;
    RECT 1.455 28.08 1.735 28.96 ;
    RECT 160.815 28.08 161.095 28.96 ;
    RECT 157.495 28.08 157.775 28.96 ;
    RECT 154.175 28.08 154.455 28.96 ;
    RECT 150.855 28.08 151.135 28.96 ;
    RECT 147.535 28.08 147.815 28.96 ;
    RECT 144.215 28.08 144.495 28.96 ;
    RECT 140.895 28.08 141.175 28.96 ;
    RECT 137.575 28.08 137.855 28.96 ;
    RECT 134.255 28.08 134.535 28.96 ;
    RECT 64.535 28.08 64.815 28.96 ;
    RECT 61.215 27.36 61.495 28.24 ;
    RECT 57.895 27.36 58.175 28.24 ;
    RECT 54.575 27.36 54.855 28.24 ;
    RECT 51.255 27.36 51.535 28.24 ;
    RECT 47.935 27.36 48.215 28.24 ;
    RECT 44.615 27.36 44.895 28.24 ;
    RECT 41.295 27.36 41.575 28.24 ;
    RECT 37.975 27.36 38.255 28.24 ;
    RECT 34.655 27.36 34.935 28.24 ;
    RECT 130.935 27.36 131.215 28.24 ;
    RECT 127.615 27.36 127.895 28.24 ;
    RECT 124.295 27.36 124.575 28.24 ;
    RECT 120.975 27.36 121.255 28.24 ;
    RECT 117.655 27.36 117.935 28.24 ;
    RECT 114.335 27.36 114.615 28.24 ;
    RECT 111.015 27.36 111.295 28.24 ;
    RECT 107.695 27.36 107.975 28.24 ;
    RECT 104.375 27.36 104.655 28.24 ;
    RECT 101.055 27.36 101.335 28.24 ;
    RECT 170.775 27.36 171.055 28.24 ;
    RECT 167.455 27.36 167.735 28.24 ;
    RECT 97.735 27.36 98.015 28.24 ;
    RECT 94.415 27.36 94.695 28.24 ;
    RECT 91.095 27.36 91.375 28.24 ;
    RECT 87.775 27.36 88.055 28.24 ;
    RECT 84.455 27.36 84.735 28.24 ;
    RECT 81.135 27.36 81.415 28.24 ;
    RECT 77.815 27.36 78.095 28.24 ;
    RECT 74.495 27.36 74.775 28.24 ;
    RECT 71.175 27.36 71.455 28.24 ;
    RECT 31.335 27.36 31.615 28.24 ;
    RECT 67.855 27.36 68.135 28.24 ;
    RECT 28.015 27.36 28.295 28.24 ;
    RECT 24.695 27.36 24.975 28.24 ;
    RECT 21.375 27.36 21.655 28.24 ;
    RECT 18.055 27.36 18.335 28.24 ;
    RECT 14.735 27.36 15.015 28.24 ;
    RECT 11.415 27.36 11.695 28.24 ;
    RECT 8.095 27.36 8.375 28.24 ;
    RECT 4.775 27.36 5.055 28.24 ;
    RECT 164.135 27.36 164.415 28.24 ;
    RECT 1.455 27.36 1.735 28.24 ;
    RECT 160.815 27.36 161.095 28.24 ;
    RECT 157.495 27.36 157.775 28.24 ;
    RECT 154.175 27.36 154.455 28.24 ;
    RECT 150.855 27.36 151.135 28.24 ;
    RECT 147.535 27.36 147.815 28.24 ;
    RECT 144.215 27.36 144.495 28.24 ;
    RECT 140.895 27.36 141.175 28.24 ;
    RECT 137.575 27.36 137.855 28.24 ;
    RECT 134.255 27.36 134.535 28.24 ;
    RECT 64.535 27.36 64.815 28.24 ;
    RECT 61.215 26.64 61.495 27.52 ;
    RECT 57.895 26.64 58.175 27.52 ;
    RECT 54.575 26.64 54.855 27.52 ;
    RECT 51.255 26.64 51.535 27.52 ;
    RECT 47.935 26.64 48.215 27.52 ;
    RECT 44.615 26.64 44.895 27.52 ;
    RECT 41.295 26.64 41.575 27.52 ;
    RECT 37.975 26.64 38.255 27.52 ;
    RECT 34.655 26.64 34.935 27.52 ;
    RECT 130.935 26.64 131.215 27.52 ;
    RECT 127.615 26.64 127.895 27.52 ;
    RECT 124.295 26.64 124.575 27.52 ;
    RECT 120.975 26.64 121.255 27.52 ;
    RECT 117.655 26.64 117.935 27.52 ;
    RECT 114.335 26.64 114.615 27.52 ;
    RECT 111.015 26.64 111.295 27.52 ;
    RECT 107.695 26.64 107.975 27.52 ;
    RECT 104.375 26.64 104.655 27.52 ;
    RECT 101.055 26.64 101.335 27.52 ;
    RECT 170.775 26.64 171.055 27.52 ;
    RECT 167.455 26.64 167.735 27.52 ;
    RECT 97.735 26.64 98.015 27.52 ;
    RECT 94.415 26.64 94.695 27.52 ;
    RECT 91.095 26.64 91.375 27.52 ;
    RECT 87.775 26.64 88.055 27.52 ;
    RECT 84.455 26.64 84.735 27.52 ;
    RECT 81.135 26.64 81.415 27.52 ;
    RECT 77.815 26.64 78.095 27.52 ;
    RECT 74.495 26.64 74.775 27.52 ;
    RECT 71.175 26.64 71.455 27.52 ;
    RECT 31.335 26.64 31.615 27.52 ;
    RECT 67.855 26.64 68.135 27.52 ;
    RECT 28.015 26.64 28.295 27.52 ;
    RECT 24.695 26.64 24.975 27.52 ;
    RECT 21.375 26.64 21.655 27.52 ;
    RECT 18.055 26.64 18.335 27.52 ;
    RECT 14.735 26.64 15.015 27.52 ;
    RECT 11.415 26.64 11.695 27.52 ;
    RECT 8.095 26.64 8.375 27.52 ;
    RECT 4.775 26.64 5.055 27.52 ;
    RECT 164.135 26.64 164.415 27.52 ;
    RECT 1.455 26.64 1.735 27.52 ;
    RECT 160.815 26.64 161.095 27.52 ;
    RECT 157.495 26.64 157.775 27.52 ;
    RECT 154.175 26.64 154.455 27.52 ;
    RECT 150.855 26.64 151.135 27.52 ;
    RECT 147.535 26.64 147.815 27.52 ;
    RECT 144.215 26.64 144.495 27.52 ;
    RECT 140.895 26.64 141.175 27.52 ;
    RECT 137.575 26.64 137.855 27.52 ;
    RECT 134.255 26.64 134.535 27.52 ;
    RECT 64.535 26.64 64.815 27.52 ;
    RECT 61.215 25.92 61.495 26.8 ;
    RECT 57.895 25.92 58.175 26.8 ;
    RECT 54.575 25.92 54.855 26.8 ;
    RECT 51.255 25.92 51.535 26.8 ;
    RECT 47.935 25.92 48.215 26.8 ;
    RECT 44.615 25.92 44.895 26.8 ;
    RECT 41.295 25.92 41.575 26.8 ;
    RECT 37.975 25.92 38.255 26.8 ;
    RECT 34.655 25.92 34.935 26.8 ;
    RECT 130.935 25.92 131.215 26.8 ;
    RECT 127.615 25.92 127.895 26.8 ;
    RECT 124.295 25.92 124.575 26.8 ;
    RECT 120.975 25.92 121.255 26.8 ;
    RECT 117.655 25.92 117.935 26.8 ;
    RECT 114.335 25.92 114.615 26.8 ;
    RECT 111.015 25.92 111.295 26.8 ;
    RECT 107.695 25.92 107.975 26.8 ;
    RECT 104.375 25.92 104.655 26.8 ;
    RECT 101.055 25.92 101.335 26.8 ;
    RECT 170.775 25.92 171.055 26.8 ;
    RECT 167.455 25.92 167.735 26.8 ;
    RECT 97.735 25.92 98.015 26.8 ;
    RECT 94.415 25.92 94.695 26.8 ;
    RECT 91.095 25.92 91.375 26.8 ;
    RECT 87.775 25.92 88.055 26.8 ;
    RECT 84.455 25.92 84.735 26.8 ;
    RECT 81.135 25.92 81.415 26.8 ;
    RECT 77.815 25.92 78.095 26.8 ;
    RECT 74.495 25.92 74.775 26.8 ;
    RECT 71.175 25.92 71.455 26.8 ;
    RECT 31.335 25.92 31.615 26.8 ;
    RECT 67.855 25.92 68.135 26.8 ;
    RECT 28.015 25.92 28.295 26.8 ;
    RECT 24.695 25.92 24.975 26.8 ;
    RECT 21.375 25.92 21.655 26.8 ;
    RECT 18.055 25.92 18.335 26.8 ;
    RECT 14.735 25.92 15.015 26.8 ;
    RECT 11.415 25.92 11.695 26.8 ;
    RECT 8.095 25.92 8.375 26.8 ;
    RECT 4.775 25.92 5.055 26.8 ;
    RECT 164.135 25.92 164.415 26.8 ;
    RECT 1.455 25.92 1.735 26.8 ;
    RECT 160.815 25.92 161.095 26.8 ;
    RECT 157.495 25.92 157.775 26.8 ;
    RECT 154.175 25.92 154.455 26.8 ;
    RECT 150.855 25.92 151.135 26.8 ;
    RECT 147.535 25.92 147.815 26.8 ;
    RECT 144.215 25.92 144.495 26.8 ;
    RECT 140.895 25.92 141.175 26.8 ;
    RECT 137.575 25.92 137.855 26.8 ;
    RECT 134.255 25.92 134.535 26.8 ;
    RECT 64.535 25.92 64.815 26.8 ;
    RECT 61.215 25.2 61.495 26.08 ;
    RECT 57.895 25.2 58.175 26.08 ;
    RECT 54.575 25.2 54.855 26.08 ;
    RECT 51.255 25.2 51.535 26.08 ;
    RECT 47.935 25.2 48.215 26.08 ;
    RECT 44.615 25.2 44.895 26.08 ;
    RECT 41.295 25.2 41.575 26.08 ;
    RECT 37.975 25.2 38.255 26.08 ;
    RECT 34.655 25.2 34.935 26.08 ;
    RECT 130.935 25.2 131.215 26.08 ;
    RECT 127.615 25.2 127.895 26.08 ;
    RECT 124.295 25.2 124.575 26.08 ;
    RECT 120.975 25.2 121.255 26.08 ;
    RECT 117.655 25.2 117.935 26.08 ;
    RECT 114.335 25.2 114.615 26.08 ;
    RECT 111.015 25.2 111.295 26.08 ;
    RECT 107.695 25.2 107.975 26.08 ;
    RECT 104.375 25.2 104.655 26.08 ;
    RECT 101.055 25.2 101.335 26.08 ;
    RECT 170.775 25.2 171.055 26.08 ;
    RECT 167.455 25.2 167.735 26.08 ;
    RECT 97.735 25.2 98.015 26.08 ;
    RECT 94.415 25.2 94.695 26.08 ;
    RECT 91.095 25.2 91.375 26.08 ;
    RECT 87.775 25.2 88.055 26.08 ;
    RECT 84.455 25.2 84.735 26.08 ;
    RECT 81.135 25.2 81.415 26.08 ;
    RECT 77.815 25.2 78.095 26.08 ;
    RECT 74.495 25.2 74.775 26.08 ;
    RECT 71.175 25.2 71.455 26.08 ;
    RECT 31.335 25.2 31.615 26.08 ;
    RECT 67.855 25.2 68.135 26.08 ;
    RECT 28.015 25.2 28.295 26.08 ;
    RECT 24.695 25.2 24.975 26.08 ;
    RECT 21.375 25.2 21.655 26.08 ;
    RECT 18.055 25.2 18.335 26.08 ;
    RECT 14.735 25.2 15.015 26.08 ;
    RECT 11.415 25.2 11.695 26.08 ;
    RECT 8.095 25.2 8.375 26.08 ;
    RECT 4.775 25.2 5.055 26.08 ;
    RECT 164.135 25.2 164.415 26.08 ;
    RECT 1.455 25.2 1.735 26.08 ;
    RECT 160.815 25.2 161.095 26.08 ;
    RECT 157.495 25.2 157.775 26.08 ;
    RECT 154.175 25.2 154.455 26.08 ;
    RECT 150.855 25.2 151.135 26.08 ;
    RECT 147.535 25.2 147.815 26.08 ;
    RECT 144.215 25.2 144.495 26.08 ;
    RECT 140.895 25.2 141.175 26.08 ;
    RECT 137.575 25.2 137.855 26.08 ;
    RECT 134.255 25.2 134.535 26.08 ;
    RECT 64.535 25.2 64.815 26.08 ;
    RECT 61.215 24.48 61.495 25.36 ;
    RECT 57.895 24.48 58.175 25.36 ;
    RECT 54.575 24.48 54.855 25.36 ;
    RECT 51.255 24.48 51.535 25.36 ;
    RECT 47.935 24.48 48.215 25.36 ;
    RECT 44.615 24.48 44.895 25.36 ;
    RECT 41.295 24.48 41.575 25.36 ;
    RECT 37.975 24.48 38.255 25.36 ;
    RECT 34.655 24.48 34.935 25.36 ;
    RECT 130.935 24.48 131.215 25.36 ;
    RECT 127.615 24.48 127.895 25.36 ;
    RECT 124.295 24.48 124.575 25.36 ;
    RECT 120.975 24.48 121.255 25.36 ;
    RECT 117.655 24.48 117.935 25.36 ;
    RECT 114.335 24.48 114.615 25.36 ;
    RECT 111.015 24.48 111.295 25.36 ;
    RECT 107.695 24.48 107.975 25.36 ;
    RECT 104.375 24.48 104.655 25.36 ;
    RECT 101.055 24.48 101.335 25.36 ;
    RECT 170.775 24.48 171.055 25.36 ;
    RECT 167.455 24.48 167.735 25.36 ;
    RECT 97.735 24.48 98.015 25.36 ;
    RECT 94.415 24.48 94.695 25.36 ;
    RECT 91.095 24.48 91.375 25.36 ;
    RECT 87.775 24.48 88.055 25.36 ;
    RECT 84.455 24.48 84.735 25.36 ;
    RECT 81.135 24.48 81.415 25.36 ;
    RECT 77.815 24.48 78.095 25.36 ;
    RECT 74.495 24.48 74.775 25.36 ;
    RECT 71.175 24.48 71.455 25.36 ;
    RECT 31.335 24.48 31.615 25.36 ;
    RECT 67.855 24.48 68.135 25.36 ;
    RECT 28.015 24.48 28.295 25.36 ;
    RECT 24.695 24.48 24.975 25.36 ;
    RECT 21.375 24.48 21.655 25.36 ;
    RECT 18.055 24.48 18.335 25.36 ;
    RECT 14.735 24.48 15.015 25.36 ;
    RECT 11.415 24.48 11.695 25.36 ;
    RECT 8.095 24.48 8.375 25.36 ;
    RECT 4.775 24.48 5.055 25.36 ;
    RECT 164.135 24.48 164.415 25.36 ;
    RECT 1.455 24.48 1.735 25.36 ;
    RECT 160.815 24.48 161.095 25.36 ;
    RECT 157.495 24.48 157.775 25.36 ;
    RECT 154.175 24.48 154.455 25.36 ;
    RECT 150.855 24.48 151.135 25.36 ;
    RECT 147.535 24.48 147.815 25.36 ;
    RECT 144.215 24.48 144.495 25.36 ;
    RECT 140.895 24.48 141.175 25.36 ;
    RECT 137.575 24.48 137.855 25.36 ;
    RECT 134.255 24.48 134.535 25.36 ;
    RECT 64.535 24.48 64.815 25.36 ;
    RECT 61.215 23.76 61.495 24.64 ;
    RECT 57.895 23.76 58.175 24.64 ;
    RECT 54.575 23.76 54.855 24.64 ;
    RECT 51.255 23.76 51.535 24.64 ;
    RECT 47.935 23.76 48.215 24.64 ;
    RECT 44.615 23.76 44.895 24.64 ;
    RECT 41.295 23.76 41.575 24.64 ;
    RECT 37.975 23.76 38.255 24.64 ;
    RECT 34.655 23.76 34.935 24.64 ;
    RECT 130.935 23.76 131.215 24.64 ;
    RECT 127.615 23.76 127.895 24.64 ;
    RECT 124.295 23.76 124.575 24.64 ;
    RECT 120.975 23.76 121.255 24.64 ;
    RECT 117.655 23.76 117.935 24.64 ;
    RECT 114.335 23.76 114.615 24.64 ;
    RECT 111.015 23.76 111.295 24.64 ;
    RECT 107.695 23.76 107.975 24.64 ;
    RECT 104.375 23.76 104.655 24.64 ;
    RECT 101.055 23.76 101.335 24.64 ;
    RECT 170.775 23.76 171.055 24.64 ;
    RECT 167.455 23.76 167.735 24.64 ;
    RECT 97.735 23.76 98.015 24.64 ;
    RECT 94.415 23.76 94.695 24.64 ;
    RECT 91.095 23.76 91.375 24.64 ;
    RECT 87.775 23.76 88.055 24.64 ;
    RECT 84.455 23.76 84.735 24.64 ;
    RECT 81.135 23.76 81.415 24.64 ;
    RECT 77.815 23.76 78.095 24.64 ;
    RECT 74.495 23.76 74.775 24.64 ;
    RECT 71.175 23.76 71.455 24.64 ;
    RECT 31.335 23.76 31.615 24.64 ;
    RECT 67.855 23.76 68.135 24.64 ;
    RECT 28.015 23.76 28.295 24.64 ;
    RECT 24.695 23.76 24.975 24.64 ;
    RECT 21.375 23.76 21.655 24.64 ;
    RECT 18.055 23.76 18.335 24.64 ;
    RECT 14.735 23.76 15.015 24.64 ;
    RECT 11.415 23.76 11.695 24.64 ;
    RECT 8.095 23.76 8.375 24.64 ;
    RECT 4.775 23.76 5.055 24.64 ;
    RECT 164.135 23.76 164.415 24.64 ;
    RECT 1.455 23.76 1.735 24.64 ;
    RECT 160.815 23.76 161.095 24.64 ;
    RECT 157.495 23.76 157.775 24.64 ;
    RECT 154.175 23.76 154.455 24.64 ;
    RECT 150.855 23.76 151.135 24.64 ;
    RECT 147.535 23.76 147.815 24.64 ;
    RECT 144.215 23.76 144.495 24.64 ;
    RECT 140.895 23.76 141.175 24.64 ;
    RECT 137.575 23.76 137.855 24.64 ;
    RECT 134.255 23.76 134.535 24.64 ;
    RECT 64.535 23.76 64.815 24.64 ;
    RECT 61.215 23.04 61.495 23.92 ;
    RECT 57.895 23.04 58.175 23.92 ;
    RECT 54.575 23.04 54.855 23.92 ;
    RECT 51.255 23.04 51.535 23.92 ;
    RECT 47.935 23.04 48.215 23.92 ;
    RECT 44.615 23.04 44.895 23.92 ;
    RECT 41.295 23.04 41.575 23.92 ;
    RECT 37.975 23.04 38.255 23.92 ;
    RECT 34.655 23.04 34.935 23.92 ;
    RECT 130.935 23.04 131.215 23.92 ;
    RECT 127.615 23.04 127.895 23.92 ;
    RECT 124.295 23.04 124.575 23.92 ;
    RECT 120.975 23.04 121.255 23.92 ;
    RECT 117.655 23.04 117.935 23.92 ;
    RECT 114.335 23.04 114.615 23.92 ;
    RECT 111.015 23.04 111.295 23.92 ;
    RECT 107.695 23.04 107.975 23.92 ;
    RECT 104.375 23.04 104.655 23.92 ;
    RECT 101.055 23.04 101.335 23.92 ;
    RECT 170.775 23.04 171.055 23.92 ;
    RECT 167.455 23.04 167.735 23.92 ;
    RECT 97.735 23.04 98.015 23.92 ;
    RECT 94.415 23.04 94.695 23.92 ;
    RECT 91.095 23.04 91.375 23.92 ;
    RECT 87.775 23.04 88.055 23.92 ;
    RECT 84.455 23.04 84.735 23.92 ;
    RECT 81.135 23.04 81.415 23.92 ;
    RECT 77.815 23.04 78.095 23.92 ;
    RECT 74.495 23.04 74.775 23.92 ;
    RECT 71.175 23.04 71.455 23.92 ;
    RECT 31.335 23.04 31.615 23.92 ;
    RECT 67.855 23.04 68.135 23.92 ;
    RECT 28.015 23.04 28.295 23.92 ;
    RECT 24.695 23.04 24.975 23.92 ;
    RECT 21.375 23.04 21.655 23.92 ;
    RECT 18.055 23.04 18.335 23.92 ;
    RECT 14.735 23.04 15.015 23.92 ;
    RECT 11.415 23.04 11.695 23.92 ;
    RECT 8.095 23.04 8.375 23.92 ;
    RECT 4.775 23.04 5.055 23.92 ;
    RECT 164.135 23.04 164.415 23.92 ;
    RECT 1.455 23.04 1.735 23.92 ;
    RECT 160.815 23.04 161.095 23.92 ;
    RECT 157.495 23.04 157.775 23.92 ;
    RECT 154.175 23.04 154.455 23.92 ;
    RECT 150.855 23.04 151.135 23.92 ;
    RECT 147.535 23.04 147.815 23.92 ;
    RECT 144.215 23.04 144.495 23.92 ;
    RECT 140.895 23.04 141.175 23.92 ;
    RECT 137.575 23.04 137.855 23.92 ;
    RECT 134.255 23.04 134.535 23.92 ;
    RECT 64.535 23.04 64.815 23.92 ;
    RECT 61.215 22.32 61.495 23.2 ;
    RECT 57.895 22.32 58.175 23.2 ;
    RECT 54.575 22.32 54.855 23.2 ;
    RECT 51.255 22.32 51.535 23.2 ;
    RECT 47.935 22.32 48.215 23.2 ;
    RECT 44.615 22.32 44.895 23.2 ;
    RECT 41.295 22.32 41.575 23.2 ;
    RECT 37.975 22.32 38.255 23.2 ;
    RECT 34.655 22.32 34.935 23.2 ;
    RECT 130.935 22.32 131.215 23.2 ;
    RECT 127.615 22.32 127.895 23.2 ;
    RECT 124.295 22.32 124.575 23.2 ;
    RECT 120.975 22.32 121.255 23.2 ;
    RECT 117.655 22.32 117.935 23.2 ;
    RECT 114.335 22.32 114.615 23.2 ;
    RECT 111.015 22.32 111.295 23.2 ;
    RECT 107.695 22.32 107.975 23.2 ;
    RECT 104.375 22.32 104.655 23.2 ;
    RECT 101.055 22.32 101.335 23.2 ;
    RECT 170.775 22.32 171.055 23.2 ;
    RECT 167.455 22.32 167.735 23.2 ;
    RECT 97.735 22.32 98.015 23.2 ;
    RECT 94.415 22.32 94.695 23.2 ;
    RECT 91.095 22.32 91.375 23.2 ;
    RECT 87.775 22.32 88.055 23.2 ;
    RECT 84.455 22.32 84.735 23.2 ;
    RECT 81.135 22.32 81.415 23.2 ;
    RECT 77.815 22.32 78.095 23.2 ;
    RECT 74.495 22.32 74.775 23.2 ;
    RECT 71.175 22.32 71.455 23.2 ;
    RECT 31.335 22.32 31.615 23.2 ;
    RECT 67.855 22.32 68.135 23.2 ;
    RECT 28.015 22.32 28.295 23.2 ;
    RECT 24.695 22.32 24.975 23.2 ;
    RECT 21.375 22.32 21.655 23.2 ;
    RECT 18.055 22.32 18.335 23.2 ;
    RECT 14.735 22.32 15.015 23.2 ;
    RECT 11.415 22.32 11.695 23.2 ;
    RECT 8.095 22.32 8.375 23.2 ;
    RECT 4.775 22.32 5.055 23.2 ;
    RECT 164.135 22.32 164.415 23.2 ;
    RECT 1.455 22.32 1.735 23.2 ;
    RECT 160.815 22.32 161.095 23.2 ;
    RECT 157.495 22.32 157.775 23.2 ;
    RECT 154.175 22.32 154.455 23.2 ;
    RECT 150.855 22.32 151.135 23.2 ;
    RECT 147.535 22.32 147.815 23.2 ;
    RECT 144.215 22.32 144.495 23.2 ;
    RECT 140.895 22.32 141.175 23.2 ;
    RECT 137.575 22.32 137.855 23.2 ;
    RECT 134.255 22.32 134.535 23.2 ;
    RECT 64.535 22.32 64.815 23.2 ;
    RECT 61.215 35.28 61.495 36.16 ;
    RECT 57.895 35.28 58.175 36.16 ;
    RECT 54.575 35.28 54.855 36.16 ;
    RECT 51.255 35.28 51.535 36.16 ;
    RECT 47.935 35.28 48.215 36.16 ;
    RECT 44.615 35.28 44.895 36.16 ;
    RECT 41.295 35.28 41.575 36.16 ;
    RECT 37.975 35.28 38.255 36.16 ;
    RECT 34.655 35.28 34.935 36.16 ;
    RECT 130.935 35.28 131.215 36.16 ;
    RECT 127.615 35.28 127.895 36.16 ;
    RECT 124.295 35.28 124.575 36.16 ;
    RECT 120.975 35.28 121.255 36.16 ;
    RECT 117.655 35.28 117.935 36.16 ;
    RECT 114.335 35.28 114.615 36.16 ;
    RECT 111.015 35.28 111.295 36.16 ;
    RECT 107.695 35.28 107.975 36.16 ;
    RECT 104.375 35.28 104.655 36.16 ;
    RECT 101.055 35.28 101.335 36.16 ;
    RECT 170.775 35.28 171.055 36.16 ;
    RECT 167.455 35.28 167.735 36.16 ;
    RECT 97.735 35.28 98.015 36.16 ;
    RECT 94.415 35.28 94.695 36.16 ;
    RECT 91.095 35.28 91.375 36.16 ;
    RECT 87.775 35.28 88.055 36.16 ;
    RECT 84.455 35.28 84.735 36.16 ;
    RECT 81.135 35.28 81.415 36.16 ;
    RECT 77.815 35.28 78.095 36.16 ;
    RECT 74.495 35.28 74.775 36.16 ;
    RECT 71.175 35.28 71.455 36.16 ;
    RECT 31.335 35.28 31.615 36.16 ;
    RECT 67.855 35.28 68.135 36.16 ;
    RECT 28.015 35.28 28.295 36.16 ;
    RECT 24.695 35.28 24.975 36.16 ;
    RECT 21.375 35.28 21.655 36.16 ;
    RECT 18.055 35.28 18.335 36.16 ;
    RECT 14.735 35.28 15.015 36.16 ;
    RECT 11.415 35.28 11.695 36.16 ;
    RECT 8.095 35.28 8.375 36.16 ;
    RECT 4.775 35.28 5.055 36.16 ;
    RECT 164.135 35.28 164.415 36.16 ;
    RECT 1.455 35.28 1.735 36.16 ;
    RECT 160.815 35.28 161.095 36.16 ;
    RECT 157.495 35.28 157.775 36.16 ;
    RECT 154.175 35.28 154.455 36.16 ;
    RECT 150.855 35.28 151.135 36.16 ;
    RECT 147.535 35.28 147.815 36.16 ;
    RECT 144.215 35.28 144.495 36.16 ;
    RECT 140.895 35.28 141.175 36.16 ;
    RECT 137.575 35.28 137.855 36.16 ;
    RECT 134.255 35.28 134.535 36.16 ;
    RECT 64.535 35.28 64.815 36.16 ;
    RECT 61.215 21.6 61.495 22.48 ;
    RECT 57.895 21.6 58.175 22.48 ;
    RECT 54.575 21.6 54.855 22.48 ;
    RECT 51.255 21.6 51.535 22.48 ;
    RECT 47.935 21.6 48.215 22.48 ;
    RECT 44.615 21.6 44.895 22.48 ;
    RECT 41.295 21.6 41.575 22.48 ;
    RECT 37.975 21.6 38.255 22.48 ;
    RECT 34.655 21.6 34.935 22.48 ;
    RECT 130.935 21.6 131.215 22.48 ;
    RECT 127.615 21.6 127.895 22.48 ;
    RECT 124.295 21.6 124.575 22.48 ;
    RECT 120.975 21.6 121.255 22.48 ;
    RECT 117.655 21.6 117.935 22.48 ;
    RECT 114.335 21.6 114.615 22.48 ;
    RECT 111.015 21.6 111.295 22.48 ;
    RECT 107.695 21.6 107.975 22.48 ;
    RECT 104.375 21.6 104.655 22.48 ;
    RECT 101.055 21.6 101.335 22.48 ;
    RECT 170.775 21.6 171.055 22.48 ;
    RECT 167.455 21.6 167.735 22.48 ;
    RECT 97.735 21.6 98.015 22.48 ;
    RECT 94.415 21.6 94.695 22.48 ;
    RECT 91.095 21.6 91.375 22.48 ;
    RECT 87.775 21.6 88.055 22.48 ;
    RECT 84.455 21.6 84.735 22.48 ;
    RECT 81.135 21.6 81.415 22.48 ;
    RECT 77.815 21.6 78.095 22.48 ;
    RECT 74.495 21.6 74.775 22.48 ;
    RECT 71.175 21.6 71.455 22.48 ;
    RECT 31.335 21.6 31.615 22.48 ;
    RECT 67.855 21.6 68.135 22.48 ;
    RECT 28.015 21.6 28.295 22.48 ;
    RECT 24.695 21.6 24.975 22.48 ;
    RECT 21.375 21.6 21.655 22.48 ;
    RECT 18.055 21.6 18.335 22.48 ;
    RECT 14.735 21.6 15.015 22.48 ;
    RECT 11.415 21.6 11.695 22.48 ;
    RECT 8.095 21.6 8.375 22.48 ;
    RECT 4.775 21.6 5.055 22.48 ;
    RECT 164.135 21.6 164.415 22.48 ;
    RECT 1.455 21.6 1.735 22.48 ;
    RECT 160.815 21.6 161.095 22.48 ;
    RECT 157.495 21.6 157.775 22.48 ;
    RECT 154.175 21.6 154.455 22.48 ;
    RECT 150.855 21.6 151.135 22.48 ;
    RECT 147.535 21.6 147.815 22.48 ;
    RECT 144.215 21.6 144.495 22.48 ;
    RECT 140.895 21.6 141.175 22.48 ;
    RECT 137.575 21.6 137.855 22.48 ;
    RECT 134.255 21.6 134.535 22.48 ;
    RECT 64.535 21.6 64.815 22.48 ;
    RECT 61.215 20.88 61.495 21.76 ;
    RECT 57.895 20.88 58.175 21.76 ;
    RECT 54.575 20.88 54.855 21.76 ;
    RECT 51.255 20.88 51.535 21.76 ;
    RECT 47.935 20.88 48.215 21.76 ;
    RECT 44.615 20.88 44.895 21.76 ;
    RECT 41.295 20.88 41.575 21.76 ;
    RECT 37.975 20.88 38.255 21.76 ;
    RECT 34.655 20.88 34.935 21.76 ;
    RECT 130.935 20.88 131.215 21.76 ;
    RECT 127.615 20.88 127.895 21.76 ;
    RECT 124.295 20.88 124.575 21.76 ;
    RECT 120.975 20.88 121.255 21.76 ;
    RECT 117.655 20.88 117.935 21.76 ;
    RECT 114.335 20.88 114.615 21.76 ;
    RECT 111.015 20.88 111.295 21.76 ;
    RECT 107.695 20.88 107.975 21.76 ;
    RECT 104.375 20.88 104.655 21.76 ;
    RECT 101.055 20.88 101.335 21.76 ;
    RECT 170.775 20.88 171.055 21.76 ;
    RECT 167.455 20.88 167.735 21.76 ;
    RECT 97.735 20.88 98.015 21.76 ;
    RECT 94.415 20.88 94.695 21.76 ;
    RECT 91.095 20.88 91.375 21.76 ;
    RECT 87.775 20.88 88.055 21.76 ;
    RECT 84.455 20.88 84.735 21.76 ;
    RECT 81.135 20.88 81.415 21.76 ;
    RECT 77.815 20.88 78.095 21.76 ;
    RECT 74.495 20.88 74.775 21.76 ;
    RECT 71.175 20.88 71.455 21.76 ;
    RECT 31.335 20.88 31.615 21.76 ;
    RECT 67.855 20.88 68.135 21.76 ;
    RECT 28.015 20.88 28.295 21.76 ;
    RECT 24.695 20.88 24.975 21.76 ;
    RECT 21.375 20.88 21.655 21.76 ;
    RECT 18.055 20.88 18.335 21.76 ;
    RECT 14.735 20.88 15.015 21.76 ;
    RECT 11.415 20.88 11.695 21.76 ;
    RECT 8.095 20.88 8.375 21.76 ;
    RECT 4.775 20.88 5.055 21.76 ;
    RECT 164.135 20.88 164.415 21.76 ;
    RECT 1.455 20.88 1.735 21.76 ;
    RECT 160.815 20.88 161.095 21.76 ;
    RECT 157.495 20.88 157.775 21.76 ;
    RECT 154.175 20.88 154.455 21.76 ;
    RECT 150.855 20.88 151.135 21.76 ;
    RECT 147.535 20.88 147.815 21.76 ;
    RECT 144.215 20.88 144.495 21.76 ;
    RECT 140.895 20.88 141.175 21.76 ;
    RECT 137.575 20.88 137.855 21.76 ;
    RECT 134.255 20.88 134.535 21.76 ;
    RECT 64.535 20.88 64.815 21.76 ;
    RECT 61.215 20.16 61.495 21.04 ;
    RECT 57.895 20.16 58.175 21.04 ;
    RECT 54.575 20.16 54.855 21.04 ;
    RECT 51.255 20.16 51.535 21.04 ;
    RECT 47.935 20.16 48.215 21.04 ;
    RECT 44.615 20.16 44.895 21.04 ;
    RECT 41.295 20.16 41.575 21.04 ;
    RECT 37.975 20.16 38.255 21.04 ;
    RECT 34.655 20.16 34.935 21.04 ;
    RECT 130.935 20.16 131.215 21.04 ;
    RECT 127.615 20.16 127.895 21.04 ;
    RECT 124.295 20.16 124.575 21.04 ;
    RECT 120.975 20.16 121.255 21.04 ;
    RECT 117.655 20.16 117.935 21.04 ;
    RECT 114.335 20.16 114.615 21.04 ;
    RECT 111.015 20.16 111.295 21.04 ;
    RECT 107.695 20.16 107.975 21.04 ;
    RECT 104.375 20.16 104.655 21.04 ;
    RECT 101.055 20.16 101.335 21.04 ;
    RECT 170.775 20.16 171.055 21.04 ;
    RECT 167.455 20.16 167.735 21.04 ;
    RECT 97.735 20.16 98.015 21.04 ;
    RECT 94.415 20.16 94.695 21.04 ;
    RECT 91.095 20.16 91.375 21.04 ;
    RECT 87.775 20.16 88.055 21.04 ;
    RECT 84.455 20.16 84.735 21.04 ;
    RECT 81.135 20.16 81.415 21.04 ;
    RECT 77.815 20.16 78.095 21.04 ;
    RECT 74.495 20.16 74.775 21.04 ;
    RECT 71.175 20.16 71.455 21.04 ;
    RECT 31.335 20.16 31.615 21.04 ;
    RECT 67.855 20.16 68.135 21.04 ;
    RECT 28.015 20.16 28.295 21.04 ;
    RECT 24.695 20.16 24.975 21.04 ;
    RECT 21.375 20.16 21.655 21.04 ;
    RECT 18.055 20.16 18.335 21.04 ;
    RECT 14.735 20.16 15.015 21.04 ;
    RECT 11.415 20.16 11.695 21.04 ;
    RECT 8.095 20.16 8.375 21.04 ;
    RECT 4.775 20.16 5.055 21.04 ;
    RECT 164.135 20.16 164.415 21.04 ;
    RECT 1.455 20.16 1.735 21.04 ;
    RECT 160.815 20.16 161.095 21.04 ;
    RECT 157.495 20.16 157.775 21.04 ;
    RECT 154.175 20.16 154.455 21.04 ;
    RECT 150.855 20.16 151.135 21.04 ;
    RECT 147.535 20.16 147.815 21.04 ;
    RECT 144.215 20.16 144.495 21.04 ;
    RECT 140.895 20.16 141.175 21.04 ;
    RECT 137.575 20.16 137.855 21.04 ;
    RECT 134.255 20.16 134.535 21.04 ;
    RECT 64.535 20.16 64.815 21.04 ;
    RECT 61.215 19.44 61.495 20.32 ;
    RECT 57.895 19.44 58.175 20.32 ;
    RECT 54.575 19.44 54.855 20.32 ;
    RECT 51.255 19.44 51.535 20.32 ;
    RECT 47.935 19.44 48.215 20.32 ;
    RECT 44.615 19.44 44.895 20.32 ;
    RECT 41.295 19.44 41.575 20.32 ;
    RECT 37.975 19.44 38.255 20.32 ;
    RECT 34.655 19.44 34.935 20.32 ;
    RECT 130.935 19.44 131.215 20.32 ;
    RECT 127.615 19.44 127.895 20.32 ;
    RECT 124.295 19.44 124.575 20.32 ;
    RECT 120.975 19.44 121.255 20.32 ;
    RECT 117.655 19.44 117.935 20.32 ;
    RECT 114.335 19.44 114.615 20.32 ;
    RECT 111.015 19.44 111.295 20.32 ;
    RECT 107.695 19.44 107.975 20.32 ;
    RECT 104.375 19.44 104.655 20.32 ;
    RECT 101.055 19.44 101.335 20.32 ;
    RECT 170.775 19.44 171.055 20.32 ;
    RECT 167.455 19.44 167.735 20.32 ;
    RECT 97.735 19.44 98.015 20.32 ;
    RECT 94.415 19.44 94.695 20.32 ;
    RECT 91.095 19.44 91.375 20.32 ;
    RECT 87.775 19.44 88.055 20.32 ;
    RECT 84.455 19.44 84.735 20.32 ;
    RECT 81.135 19.44 81.415 20.32 ;
    RECT 77.815 19.44 78.095 20.32 ;
    RECT 74.495 19.44 74.775 20.32 ;
    RECT 71.175 19.44 71.455 20.32 ;
    RECT 31.335 19.44 31.615 20.32 ;
    RECT 67.855 19.44 68.135 20.32 ;
    RECT 28.015 19.44 28.295 20.32 ;
    RECT 24.695 19.44 24.975 20.32 ;
    RECT 21.375 19.44 21.655 20.32 ;
    RECT 18.055 19.44 18.335 20.32 ;
    RECT 14.735 19.44 15.015 20.32 ;
    RECT 11.415 19.44 11.695 20.32 ;
    RECT 8.095 19.44 8.375 20.32 ;
    RECT 4.775 19.44 5.055 20.32 ;
    RECT 164.135 19.44 164.415 20.32 ;
    RECT 1.455 19.44 1.735 20.32 ;
    RECT 160.815 19.44 161.095 20.32 ;
    RECT 157.495 19.44 157.775 20.32 ;
    RECT 154.175 19.44 154.455 20.32 ;
    RECT 150.855 19.44 151.135 20.32 ;
    RECT 147.535 19.44 147.815 20.32 ;
    RECT 144.215 19.44 144.495 20.32 ;
    RECT 140.895 19.44 141.175 20.32 ;
    RECT 137.575 19.44 137.855 20.32 ;
    RECT 134.255 19.44 134.535 20.32 ;
    RECT 64.535 19.44 64.815 20.32 ;
    RECT 61.215 18.72 61.495 19.6 ;
    RECT 57.895 18.72 58.175 19.6 ;
    RECT 54.575 18.72 54.855 19.6 ;
    RECT 51.255 18.72 51.535 19.6 ;
    RECT 47.935 18.72 48.215 19.6 ;
    RECT 44.615 18.72 44.895 19.6 ;
    RECT 41.295 18.72 41.575 19.6 ;
    RECT 37.975 18.72 38.255 19.6 ;
    RECT 34.655 18.72 34.935 19.6 ;
    RECT 130.935 18.72 131.215 19.6 ;
    RECT 127.615 18.72 127.895 19.6 ;
    RECT 124.295 18.72 124.575 19.6 ;
    RECT 120.975 18.72 121.255 19.6 ;
    RECT 117.655 18.72 117.935 19.6 ;
    RECT 114.335 18.72 114.615 19.6 ;
    RECT 111.015 18.72 111.295 19.6 ;
    RECT 107.695 18.72 107.975 19.6 ;
    RECT 104.375 18.72 104.655 19.6 ;
    RECT 101.055 18.72 101.335 19.6 ;
    RECT 170.775 18.72 171.055 19.6 ;
    RECT 167.455 18.72 167.735 19.6 ;
    RECT 97.735 18.72 98.015 19.6 ;
    RECT 94.415 18.72 94.695 19.6 ;
    RECT 91.095 18.72 91.375 19.6 ;
    RECT 87.775 18.72 88.055 19.6 ;
    RECT 84.455 18.72 84.735 19.6 ;
    RECT 81.135 18.72 81.415 19.6 ;
    RECT 77.815 18.72 78.095 19.6 ;
    RECT 74.495 18.72 74.775 19.6 ;
    RECT 71.175 18.72 71.455 19.6 ;
    RECT 31.335 18.72 31.615 19.6 ;
    RECT 67.855 18.72 68.135 19.6 ;
    RECT 28.015 18.72 28.295 19.6 ;
    RECT 24.695 18.72 24.975 19.6 ;
    RECT 21.375 18.72 21.655 19.6 ;
    RECT 18.055 18.72 18.335 19.6 ;
    RECT 14.735 18.72 15.015 19.6 ;
    RECT 11.415 18.72 11.695 19.6 ;
    RECT 8.095 18.72 8.375 19.6 ;
    RECT 4.775 18.72 5.055 19.6 ;
    RECT 164.135 18.72 164.415 19.6 ;
    RECT 1.455 18.72 1.735 19.6 ;
    RECT 160.815 18.72 161.095 19.6 ;
    RECT 157.495 18.72 157.775 19.6 ;
    RECT 154.175 18.72 154.455 19.6 ;
    RECT 150.855 18.72 151.135 19.6 ;
    RECT 147.535 18.72 147.815 19.6 ;
    RECT 144.215 18.72 144.495 19.6 ;
    RECT 140.895 18.72 141.175 19.6 ;
    RECT 137.575 18.72 137.855 19.6 ;
    RECT 134.255 18.72 134.535 19.6 ;
    RECT 64.535 18.72 64.815 19.6 ;
    RECT 31.335 57.68 31.615 58.42 ;
    RECT 28.015 57.68 28.295 58.42 ;
    RECT 24.695 57.68 24.975 58.42 ;
    RECT 21.375 57.68 21.655 58.42 ;
    RECT 18.055 57.68 18.335 58.42 ;
    RECT 14.735 57.68 15.015 58.42 ;
    RECT 11.415 57.68 11.695 58.42 ;
    RECT 8.095 57.68 8.375 58.42 ;
    RECT 4.775 57.68 5.055 58.42 ;
    RECT 1.455 57.68 1.735 58.42 ;
    RECT 170.775 57.68 171.055 58.42 ;
    RECT 167.455 57.68 167.735 58.42 ;
    RECT 164.135 57.68 164.415 58.42 ;
    RECT 160.815 57.68 161.095 58.42 ;
    RECT 157.495 57.68 157.775 58.42 ;
    RECT 154.175 57.68 154.455 58.42 ;
    RECT 150.855 57.68 151.135 58.42 ;
    RECT 147.535 57.68 147.815 58.42 ;
    RECT 144.215 57.68 144.495 58.42 ;
    RECT 140.895 57.68 141.175 58.42 ;
    RECT 137.575 57.68 137.855 58.42 ;
    RECT 134.255 57.68 134.535 58.42 ;
    RECT 130.935 57.68 131.215 58.42 ;
    RECT 127.615 57.68 127.895 58.42 ;
    RECT 124.295 57.68 124.575 58.42 ;
    RECT 120.975 57.68 121.255 58.42 ;
    RECT 117.655 57.68 117.935 58.42 ;
    RECT 114.335 57.68 114.615 58.42 ;
    RECT 111.015 57.68 111.295 58.42 ;
    RECT 107.695 57.68 107.975 58.42 ;
    RECT 104.375 57.68 104.655 58.42 ;
    RECT 101.055 57.68 101.335 58.42 ;
    RECT 97.735 57.68 98.015 58.42 ;
    RECT 94.415 57.68 94.695 58.42 ;
    RECT 91.095 57.68 91.375 58.42 ;
    RECT 87.775 57.68 88.055 58.42 ;
    RECT 84.455 57.68 84.735 58.42 ;
    RECT 81.135 57.68 81.415 58.42 ;
    RECT 77.815 57.68 78.095 58.42 ;
    RECT 74.495 57.68 74.775 58.42 ;
    RECT 71.175 57.68 71.455 58.42 ;
    RECT 67.855 57.68 68.135 58.42 ;
    RECT 64.535 57.68 64.815 58.42 ;
    RECT 61.215 57.68 61.495 58.42 ;
    RECT 57.895 57.68 58.175 58.42 ;
    RECT 54.575 57.68 54.855 58.42 ;
    RECT 51.255 57.68 51.535 58.42 ;
    RECT 47.935 57.68 48.215 58.42 ;
    RECT 44.615 57.68 44.895 58.42 ;
    RECT 41.295 57.68 41.575 58.42 ;
    RECT 37.975 57.68 38.255 58.42 ;
    RECT 34.655 57.68 34.935 58.42 ;
    RECT 61.215 56.88 61.495 57.76 ;
    RECT 57.895 56.88 58.175 57.76 ;
    RECT 54.575 56.88 54.855 57.76 ;
    RECT 51.255 56.88 51.535 57.76 ;
    RECT 47.935 56.88 48.215 57.76 ;
    RECT 44.615 56.88 44.895 57.76 ;
    RECT 41.295 56.88 41.575 57.76 ;
    RECT 37.975 56.88 38.255 57.76 ;
    RECT 34.655 56.88 34.935 57.76 ;
    RECT 130.935 56.88 131.215 57.76 ;
    RECT 127.615 56.88 127.895 57.76 ;
    RECT 124.295 56.88 124.575 57.76 ;
    RECT 120.975 56.88 121.255 57.76 ;
    RECT 117.655 56.88 117.935 57.76 ;
    RECT 114.335 56.88 114.615 57.76 ;
    RECT 111.015 56.88 111.295 57.76 ;
    RECT 107.695 56.88 107.975 57.76 ;
    RECT 104.375 56.88 104.655 57.76 ;
    RECT 101.055 56.88 101.335 57.76 ;
    RECT 170.775 56.88 171.055 57.76 ;
    RECT 167.455 56.88 167.735 57.76 ;
    RECT 97.735 56.88 98.015 57.76 ;
    RECT 94.415 56.88 94.695 57.76 ;
    RECT 91.095 56.88 91.375 57.76 ;
    RECT 87.775 56.88 88.055 57.76 ;
    RECT 84.455 56.88 84.735 57.76 ;
    RECT 81.135 56.88 81.415 57.76 ;
    RECT 77.815 56.88 78.095 57.76 ;
    RECT 74.495 56.88 74.775 57.76 ;
    RECT 71.175 56.88 71.455 57.76 ;
    RECT 31.335 56.88 31.615 57.76 ;
    RECT 67.855 56.88 68.135 57.76 ;
    RECT 28.015 56.88 28.295 57.76 ;
    RECT 24.695 56.88 24.975 57.76 ;
    RECT 21.375 56.88 21.655 57.76 ;
    RECT 18.055 56.88 18.335 57.76 ;
    RECT 14.735 56.88 15.015 57.76 ;
    RECT 11.415 56.88 11.695 57.76 ;
    RECT 8.095 56.88 8.375 57.76 ;
    RECT 4.775 56.88 5.055 57.76 ;
    RECT 164.135 56.88 164.415 57.76 ;
    RECT 1.455 56.88 1.735 57.76 ;
    RECT 160.815 56.88 161.095 57.76 ;
    RECT 157.495 56.88 157.775 57.76 ;
    RECT 154.175 56.88 154.455 57.76 ;
    RECT 150.855 56.88 151.135 57.76 ;
    RECT 147.535 56.88 147.815 57.76 ;
    RECT 144.215 56.88 144.495 57.76 ;
    RECT 140.895 56.88 141.175 57.76 ;
    RECT 137.575 56.88 137.855 57.76 ;
    RECT 134.255 56.88 134.535 57.76 ;
    RECT 64.535 56.88 64.815 57.76 ;
    RECT 61.215 56.16 61.495 57.04 ;
    RECT 57.895 56.16 58.175 57.04 ;
    RECT 54.575 56.16 54.855 57.04 ;
    RECT 51.255 56.16 51.535 57.04 ;
    RECT 47.935 56.16 48.215 57.04 ;
    RECT 44.615 56.16 44.895 57.04 ;
    RECT 41.295 56.16 41.575 57.04 ;
    RECT 37.975 56.16 38.255 57.04 ;
    RECT 34.655 56.16 34.935 57.04 ;
    RECT 130.935 56.16 131.215 57.04 ;
    RECT 127.615 56.16 127.895 57.04 ;
    RECT 124.295 56.16 124.575 57.04 ;
    RECT 120.975 56.16 121.255 57.04 ;
    RECT 117.655 56.16 117.935 57.04 ;
    RECT 114.335 56.16 114.615 57.04 ;
    RECT 111.015 56.16 111.295 57.04 ;
    RECT 107.695 56.16 107.975 57.04 ;
    RECT 104.375 56.16 104.655 57.04 ;
    RECT 101.055 56.16 101.335 57.04 ;
    RECT 170.775 56.16 171.055 57.04 ;
    RECT 167.455 56.16 167.735 57.04 ;
    RECT 97.735 56.16 98.015 57.04 ;
    RECT 94.415 56.16 94.695 57.04 ;
    RECT 91.095 56.16 91.375 57.04 ;
    RECT 87.775 56.16 88.055 57.04 ;
    RECT 84.455 56.16 84.735 57.04 ;
    RECT 81.135 56.16 81.415 57.04 ;
    RECT 77.815 56.16 78.095 57.04 ;
    RECT 74.495 56.16 74.775 57.04 ;
    RECT 71.175 56.16 71.455 57.04 ;
    RECT 31.335 56.16 31.615 57.04 ;
    RECT 67.855 56.16 68.135 57.04 ;
    RECT 28.015 56.16 28.295 57.04 ;
    RECT 24.695 56.16 24.975 57.04 ;
    RECT 21.375 56.16 21.655 57.04 ;
    RECT 18.055 56.16 18.335 57.04 ;
    RECT 14.735 56.16 15.015 57.04 ;
    RECT 11.415 56.16 11.695 57.04 ;
    RECT 8.095 56.16 8.375 57.04 ;
    RECT 4.775 56.16 5.055 57.04 ;
    RECT 164.135 56.16 164.415 57.04 ;
    RECT 1.455 56.16 1.735 57.04 ;
    RECT 160.815 56.16 161.095 57.04 ;
    RECT 157.495 56.16 157.775 57.04 ;
    RECT 154.175 56.16 154.455 57.04 ;
    RECT 150.855 56.16 151.135 57.04 ;
    RECT 147.535 56.16 147.815 57.04 ;
    RECT 144.215 56.16 144.495 57.04 ;
    RECT 140.895 56.16 141.175 57.04 ;
    RECT 137.575 56.16 137.855 57.04 ;
    RECT 134.255 56.16 134.535 57.04 ;
    RECT 64.535 56.16 64.815 57.04 ;
    RECT 61.215 55.44 61.495 56.32 ;
    RECT 57.895 55.44 58.175 56.32 ;
    RECT 54.575 55.44 54.855 56.32 ;
    RECT 51.255 55.44 51.535 56.32 ;
    RECT 47.935 55.44 48.215 56.32 ;
    RECT 44.615 55.44 44.895 56.32 ;
    RECT 41.295 55.44 41.575 56.32 ;
    RECT 37.975 55.44 38.255 56.32 ;
    RECT 34.655 55.44 34.935 56.32 ;
    RECT 130.935 55.44 131.215 56.32 ;
    RECT 127.615 55.44 127.895 56.32 ;
    RECT 124.295 55.44 124.575 56.32 ;
    RECT 120.975 55.44 121.255 56.32 ;
    RECT 117.655 55.44 117.935 56.32 ;
    RECT 114.335 55.44 114.615 56.32 ;
    RECT 111.015 55.44 111.295 56.32 ;
    RECT 107.695 55.44 107.975 56.32 ;
    RECT 104.375 55.44 104.655 56.32 ;
    RECT 101.055 55.44 101.335 56.32 ;
    RECT 170.775 55.44 171.055 56.32 ;
    RECT 167.455 55.44 167.735 56.32 ;
    RECT 97.735 55.44 98.015 56.32 ;
    RECT 94.415 55.44 94.695 56.32 ;
    RECT 91.095 55.44 91.375 56.32 ;
    RECT 87.775 55.44 88.055 56.32 ;
    RECT 84.455 55.44 84.735 56.32 ;
    RECT 81.135 55.44 81.415 56.32 ;
    RECT 77.815 55.44 78.095 56.32 ;
    RECT 74.495 55.44 74.775 56.32 ;
    RECT 71.175 55.44 71.455 56.32 ;
    RECT 31.335 55.44 31.615 56.32 ;
    RECT 67.855 55.44 68.135 56.32 ;
    RECT 28.015 55.44 28.295 56.32 ;
    RECT 24.695 55.44 24.975 56.32 ;
    RECT 21.375 55.44 21.655 56.32 ;
    RECT 18.055 55.44 18.335 56.32 ;
    RECT 14.735 55.44 15.015 56.32 ;
    RECT 11.415 55.44 11.695 56.32 ;
    RECT 8.095 55.44 8.375 56.32 ;
    RECT 4.775 55.44 5.055 56.32 ;
    RECT 164.135 55.44 164.415 56.32 ;
    RECT 1.455 55.44 1.735 56.32 ;
    RECT 160.815 55.44 161.095 56.32 ;
    RECT 157.495 55.44 157.775 56.32 ;
    RECT 154.175 55.44 154.455 56.32 ;
    RECT 150.855 55.44 151.135 56.32 ;
    RECT 147.535 55.44 147.815 56.32 ;
    RECT 144.215 55.44 144.495 56.32 ;
    RECT 140.895 55.44 141.175 56.32 ;
    RECT 137.575 55.44 137.855 56.32 ;
    RECT 134.255 55.44 134.535 56.32 ;
    RECT 64.535 55.44 64.815 56.32 ;
    RECT 61.215 54.72 61.495 55.6 ;
    RECT 57.895 54.72 58.175 55.6 ;
    RECT 54.575 54.72 54.855 55.6 ;
    RECT 51.255 54.72 51.535 55.6 ;
    RECT 47.935 54.72 48.215 55.6 ;
    RECT 44.615 54.72 44.895 55.6 ;
    RECT 41.295 54.72 41.575 55.6 ;
    RECT 37.975 54.72 38.255 55.6 ;
    RECT 34.655 54.72 34.935 55.6 ;
    RECT 130.935 54.72 131.215 55.6 ;
    RECT 127.615 54.72 127.895 55.6 ;
    RECT 124.295 54.72 124.575 55.6 ;
    RECT 120.975 54.72 121.255 55.6 ;
    RECT 117.655 54.72 117.935 55.6 ;
    RECT 114.335 54.72 114.615 55.6 ;
    RECT 111.015 54.72 111.295 55.6 ;
    RECT 107.695 54.72 107.975 55.6 ;
    RECT 104.375 54.72 104.655 55.6 ;
    RECT 101.055 54.72 101.335 55.6 ;
    RECT 170.775 54.72 171.055 55.6 ;
    RECT 167.455 54.72 167.735 55.6 ;
    RECT 97.735 54.72 98.015 55.6 ;
    RECT 94.415 54.72 94.695 55.6 ;
    RECT 91.095 54.72 91.375 55.6 ;
    RECT 87.775 54.72 88.055 55.6 ;
    RECT 84.455 54.72 84.735 55.6 ;
    RECT 81.135 54.72 81.415 55.6 ;
    RECT 77.815 54.72 78.095 55.6 ;
    RECT 74.495 54.72 74.775 55.6 ;
    RECT 71.175 54.72 71.455 55.6 ;
    RECT 31.335 54.72 31.615 55.6 ;
    RECT 67.855 54.72 68.135 55.6 ;
    RECT 28.015 54.72 28.295 55.6 ;
    RECT 24.695 54.72 24.975 55.6 ;
    RECT 21.375 54.72 21.655 55.6 ;
    RECT 18.055 54.72 18.335 55.6 ;
    RECT 14.735 54.72 15.015 55.6 ;
    RECT 11.415 54.72 11.695 55.6 ;
    RECT 8.095 54.72 8.375 55.6 ;
    RECT 4.775 54.72 5.055 55.6 ;
    RECT 164.135 54.72 164.415 55.6 ;
    RECT 1.455 54.72 1.735 55.6 ;
    RECT 160.815 54.72 161.095 55.6 ;
    RECT 157.495 54.72 157.775 55.6 ;
    RECT 154.175 54.72 154.455 55.6 ;
    RECT 150.855 54.72 151.135 55.6 ;
    RECT 147.535 54.72 147.815 55.6 ;
    RECT 144.215 54.72 144.495 55.6 ;
    RECT 140.895 54.72 141.175 55.6 ;
    RECT 137.575 54.72 137.855 55.6 ;
    RECT 134.255 54.72 134.535 55.6 ;
    RECT 64.535 54.72 64.815 55.6 ;
    RECT 31.335 59.14 31.615 60.67 ;
    RECT 28.015 59.14 28.295 60.67 ;
    RECT 24.695 59.14 24.975 60.67 ;
    RECT 21.375 59.14 21.655 60.67 ;
    RECT 18.055 59.14 18.335 60.67 ;
    RECT 14.735 59.14 15.015 60.67 ;
    RECT 11.415 59.14 11.695 60.67 ;
    RECT 8.095 59.14 8.375 60.67 ;
    RECT 4.775 59.14 5.055 60.67 ;
    RECT 1.455 59.14 1.735 60.67 ;
    RECT 170.775 59.14 171.055 60.67 ;
    RECT 167.455 59.14 167.735 60.67 ;
    RECT 164.135 59.14 164.415 60.67 ;
    RECT 160.815 59.14 161.095 60.67 ;
    RECT 157.495 59.14 157.775 60.67 ;
    RECT 154.175 59.14 154.455 60.67 ;
    RECT 150.855 59.14 151.135 60.67 ;
    RECT 147.535 59.14 147.815 60.67 ;
    RECT 144.215 59.14 144.495 60.67 ;
    RECT 140.895 59.14 141.175 60.67 ;
    RECT 137.575 59.14 137.855 60.67 ;
    RECT 134.255 59.14 134.535 60.67 ;
    RECT 130.935 59.14 131.215 60.67 ;
    RECT 127.615 59.14 127.895 60.67 ;
    RECT 124.295 59.14 124.575 60.67 ;
    RECT 120.975 59.14 121.255 60.67 ;
    RECT 117.655 59.14 117.935 60.67 ;
    RECT 114.335 59.14 114.615 60.67 ;
    RECT 111.015 59.14 111.295 60.67 ;
    RECT 107.695 59.14 107.975 60.67 ;
    RECT 104.375 59.14 104.655 60.67 ;
    RECT 101.055 59.14 101.335 60.67 ;
    RECT 97.735 59.14 98.015 60.67 ;
    RECT 94.415 59.14 94.695 60.67 ;
    RECT 91.095 59.14 91.375 60.67 ;
    RECT 87.775 59.14 88.055 60.67 ;
    RECT 84.455 59.14 84.735 60.67 ;
    RECT 81.135 59.14 81.415 60.67 ;
    RECT 77.815 59.14 78.095 60.67 ;
    RECT 74.495 59.14 74.775 60.67 ;
    RECT 71.175 59.14 71.455 60.67 ;
    RECT 67.855 59.14 68.135 60.67 ;
    RECT 64.535 59.14 64.815 60.67 ;
    RECT 61.215 59.14 61.495 60.67 ;
    RECT 57.895 59.14 58.175 60.67 ;
    RECT 54.575 59.14 54.855 60.67 ;
    RECT 51.255 59.14 51.535 60.67 ;
    RECT 47.935 59.14 48.215 60.67 ;
    RECT 44.615 59.14 44.895 60.67 ;
    RECT 41.295 59.14 41.575 60.67 ;
    RECT 37.975 59.14 38.255 60.67 ;
    RECT 34.655 59.14 34.935 60.67 ;
    RECT 61.215 33.84 61.495 34.72 ;
    RECT 57.895 33.84 58.175 34.72 ;
    RECT 54.575 33.84 54.855 34.72 ;
    RECT 51.255 33.84 51.535 34.72 ;
    RECT 47.935 33.84 48.215 34.72 ;
    RECT 44.615 33.84 44.895 34.72 ;
    RECT 41.295 33.84 41.575 34.72 ;
    RECT 37.975 33.84 38.255 34.72 ;
    RECT 34.655 33.84 34.935 34.72 ;
    RECT 130.935 33.84 131.215 34.72 ;
    RECT 127.615 33.84 127.895 34.72 ;
    RECT 124.295 33.84 124.575 34.72 ;
    RECT 120.975 33.84 121.255 34.72 ;
    RECT 117.655 33.84 117.935 34.72 ;
    RECT 114.335 33.84 114.615 34.72 ;
    RECT 111.015 33.84 111.295 34.72 ;
    RECT 107.695 33.84 107.975 34.72 ;
    RECT 104.375 33.84 104.655 34.72 ;
    RECT 101.055 33.84 101.335 34.72 ;
    RECT 170.775 33.84 171.055 34.72 ;
    RECT 167.455 33.84 167.735 34.72 ;
    RECT 97.735 33.84 98.015 34.72 ;
    RECT 94.415 33.84 94.695 34.72 ;
    RECT 91.095 33.84 91.375 34.72 ;
    RECT 87.775 33.84 88.055 34.72 ;
    RECT 84.455 33.84 84.735 34.72 ;
    RECT 81.135 33.84 81.415 34.72 ;
    RECT 77.815 33.84 78.095 34.72 ;
    RECT 74.495 33.84 74.775 34.72 ;
    RECT 71.175 33.84 71.455 34.72 ;
    RECT 31.335 33.84 31.615 34.72 ;
    RECT 67.855 33.84 68.135 34.72 ;
    RECT 28.015 33.84 28.295 34.72 ;
    RECT 24.695 33.84 24.975 34.72 ;
    RECT 21.375 33.84 21.655 34.72 ;
    RECT 18.055 33.84 18.335 34.72 ;
    RECT 14.735 33.84 15.015 34.72 ;
    RECT 11.415 33.84 11.695 34.72 ;
    RECT 8.095 33.84 8.375 34.72 ;
    RECT 4.775 33.84 5.055 34.72 ;
    RECT 164.135 33.84 164.415 34.72 ;
    RECT 1.455 33.84 1.735 34.72 ;
    RECT 160.815 33.84 161.095 34.72 ;
    RECT 157.495 33.84 157.775 34.72 ;
    RECT 154.175 33.84 154.455 34.72 ;
    RECT 150.855 33.84 151.135 34.72 ;
    RECT 147.535 33.84 147.815 34.72 ;
    RECT 144.215 33.84 144.495 34.72 ;
    RECT 140.895 33.84 141.175 34.72 ;
    RECT 137.575 33.84 137.855 34.72 ;
    RECT 134.255 33.84 134.535 34.72 ;
    RECT 64.535 33.84 64.815 34.72 ;
    RECT 61.215 34.56 61.495 35.44 ;
    RECT 57.895 34.56 58.175 35.44 ;
    RECT 54.575 34.56 54.855 35.44 ;
    RECT 51.255 34.56 51.535 35.44 ;
    RECT 47.935 34.56 48.215 35.44 ;
    RECT 44.615 34.56 44.895 35.44 ;
    RECT 41.295 34.56 41.575 35.44 ;
    RECT 37.975 34.56 38.255 35.44 ;
    RECT 34.655 34.56 34.935 35.44 ;
    RECT 130.935 34.56 131.215 35.44 ;
    RECT 127.615 34.56 127.895 35.44 ;
    RECT 124.295 34.56 124.575 35.44 ;
    RECT 120.975 34.56 121.255 35.44 ;
    RECT 117.655 34.56 117.935 35.44 ;
    RECT 114.335 34.56 114.615 35.44 ;
    RECT 111.015 34.56 111.295 35.44 ;
    RECT 107.695 34.56 107.975 35.44 ;
    RECT 104.375 34.56 104.655 35.44 ;
    RECT 101.055 34.56 101.335 35.44 ;
    RECT 170.775 34.56 171.055 35.44 ;
    RECT 167.455 34.56 167.735 35.44 ;
    RECT 97.735 34.56 98.015 35.44 ;
    RECT 94.415 34.56 94.695 35.44 ;
    RECT 91.095 34.56 91.375 35.44 ;
    RECT 87.775 34.56 88.055 35.44 ;
    RECT 84.455 34.56 84.735 35.44 ;
    RECT 81.135 34.56 81.415 35.44 ;
    RECT 77.815 34.56 78.095 35.44 ;
    RECT 74.495 34.56 74.775 35.44 ;
    RECT 71.175 34.56 71.455 35.44 ;
    RECT 31.335 34.56 31.615 35.44 ;
    RECT 67.855 34.56 68.135 35.44 ;
    RECT 28.015 34.56 28.295 35.44 ;
    RECT 24.695 34.56 24.975 35.44 ;
    RECT 21.375 34.56 21.655 35.44 ;
    RECT 18.055 34.56 18.335 35.44 ;
    RECT 14.735 34.56 15.015 35.44 ;
    RECT 11.415 34.56 11.695 35.44 ;
    RECT 8.095 34.56 8.375 35.44 ;
    RECT 4.775 34.56 5.055 35.44 ;
    RECT 164.135 34.56 164.415 35.44 ;
    RECT 1.455 34.56 1.735 35.44 ;
    RECT 160.815 34.56 161.095 35.44 ;
    RECT 157.495 34.56 157.775 35.44 ;
    RECT 154.175 34.56 154.455 35.44 ;
    RECT 150.855 34.56 151.135 35.44 ;
    RECT 147.535 34.56 147.815 35.44 ;
    RECT 144.215 34.56 144.495 35.44 ;
    RECT 140.895 34.56 141.175 35.44 ;
    RECT 137.575 34.56 137.855 35.44 ;
    RECT 134.255 34.56 134.535 35.44 ;
    RECT 64.535 34.56 64.815 35.44 ;
    RECT 61.215 54.0 61.495 54.88 ;
    RECT 57.895 54.0 58.175 54.88 ;
    RECT 54.575 54.0 54.855 54.88 ;
    RECT 51.255 54.0 51.535 54.88 ;
    RECT 47.935 54.0 48.215 54.88 ;
    RECT 44.615 54.0 44.895 54.88 ;
    RECT 41.295 54.0 41.575 54.88 ;
    RECT 37.975 54.0 38.255 54.88 ;
    RECT 34.655 54.0 34.935 54.88 ;
    RECT 130.935 54.0 131.215 54.88 ;
    RECT 127.615 54.0 127.895 54.88 ;
    RECT 124.295 54.0 124.575 54.88 ;
    RECT 120.975 54.0 121.255 54.88 ;
    RECT 117.655 54.0 117.935 54.88 ;
    RECT 114.335 54.0 114.615 54.88 ;
    RECT 111.015 54.0 111.295 54.88 ;
    RECT 107.695 54.0 107.975 54.88 ;
    RECT 104.375 54.0 104.655 54.88 ;
    RECT 101.055 54.0 101.335 54.88 ;
    RECT 170.775 54.0 171.055 54.88 ;
    RECT 167.455 54.0 167.735 54.88 ;
    RECT 97.735 54.0 98.015 54.88 ;
    RECT 94.415 54.0 94.695 54.88 ;
    RECT 91.095 54.0 91.375 54.88 ;
    RECT 87.775 54.0 88.055 54.88 ;
    RECT 84.455 54.0 84.735 54.88 ;
    RECT 81.135 54.0 81.415 54.88 ;
    RECT 77.815 54.0 78.095 54.88 ;
    RECT 74.495 54.0 74.775 54.88 ;
    RECT 71.175 54.0 71.455 54.88 ;
    RECT 31.335 54.0 31.615 54.88 ;
    RECT 67.855 54.0 68.135 54.88 ;
    RECT 28.015 54.0 28.295 54.88 ;
    RECT 24.695 54.0 24.975 54.88 ;
    RECT 21.375 54.0 21.655 54.88 ;
    RECT 18.055 54.0 18.335 54.88 ;
    RECT 14.735 54.0 15.015 54.88 ;
    RECT 11.415 54.0 11.695 54.88 ;
    RECT 8.095 54.0 8.375 54.88 ;
    RECT 4.775 54.0 5.055 54.88 ;
    RECT 164.135 54.0 164.415 54.88 ;
    RECT 1.455 54.0 1.735 54.88 ;
    RECT 160.815 54.0 161.095 54.88 ;
    RECT 157.495 54.0 157.775 54.88 ;
    RECT 154.175 54.0 154.455 54.88 ;
    RECT 150.855 54.0 151.135 54.88 ;
    RECT 147.535 54.0 147.815 54.88 ;
    RECT 144.215 54.0 144.495 54.88 ;
    RECT 140.895 54.0 141.175 54.88 ;
    RECT 137.575 54.0 137.855 54.88 ;
    RECT 134.255 54.0 134.535 54.88 ;
    RECT 64.535 54.0 64.815 54.88 ;
    RECT 61.215 53.28 61.495 54.16 ;
    RECT 57.895 53.28 58.175 54.16 ;
    RECT 54.575 53.28 54.855 54.16 ;
    RECT 51.255 53.28 51.535 54.16 ;
    RECT 47.935 53.28 48.215 54.16 ;
    RECT 44.615 53.28 44.895 54.16 ;
    RECT 41.295 53.28 41.575 54.16 ;
    RECT 37.975 53.28 38.255 54.16 ;
    RECT 34.655 53.28 34.935 54.16 ;
    RECT 130.935 53.28 131.215 54.16 ;
    RECT 127.615 53.28 127.895 54.16 ;
    RECT 124.295 53.28 124.575 54.16 ;
    RECT 120.975 53.28 121.255 54.16 ;
    RECT 117.655 53.28 117.935 54.16 ;
    RECT 114.335 53.28 114.615 54.16 ;
    RECT 111.015 53.28 111.295 54.16 ;
    RECT 107.695 53.28 107.975 54.16 ;
    RECT 104.375 53.28 104.655 54.16 ;
    RECT 101.055 53.28 101.335 54.16 ;
    RECT 170.775 53.28 171.055 54.16 ;
    RECT 167.455 53.28 167.735 54.16 ;
    RECT 97.735 53.28 98.015 54.16 ;
    RECT 94.415 53.28 94.695 54.16 ;
    RECT 91.095 53.28 91.375 54.16 ;
    RECT 87.775 53.28 88.055 54.16 ;
    RECT 84.455 53.28 84.735 54.16 ;
    RECT 81.135 53.28 81.415 54.16 ;
    RECT 77.815 53.28 78.095 54.16 ;
    RECT 74.495 53.28 74.775 54.16 ;
    RECT 71.175 53.28 71.455 54.16 ;
    RECT 31.335 53.28 31.615 54.16 ;
    RECT 67.855 53.28 68.135 54.16 ;
    RECT 28.015 53.28 28.295 54.16 ;
    RECT 24.695 53.28 24.975 54.16 ;
    RECT 21.375 53.28 21.655 54.16 ;
    RECT 18.055 53.28 18.335 54.16 ;
    RECT 14.735 53.28 15.015 54.16 ;
    RECT 11.415 53.28 11.695 54.16 ;
    RECT 8.095 53.28 8.375 54.16 ;
    RECT 4.775 53.28 5.055 54.16 ;
    RECT 164.135 53.28 164.415 54.16 ;
    RECT 1.455 53.28 1.735 54.16 ;
    RECT 160.815 53.28 161.095 54.16 ;
    RECT 157.495 53.28 157.775 54.16 ;
    RECT 154.175 53.28 154.455 54.16 ;
    RECT 150.855 53.28 151.135 54.16 ;
    RECT 147.535 53.28 147.815 54.16 ;
    RECT 144.215 53.28 144.495 54.16 ;
    RECT 140.895 53.28 141.175 54.16 ;
    RECT 137.575 53.28 137.855 54.16 ;
    RECT 134.255 53.28 134.535 54.16 ;
    RECT 64.535 53.28 64.815 54.16 ;
    RECT 61.215 52.56 61.495 53.44 ;
    RECT 57.895 52.56 58.175 53.44 ;
    RECT 54.575 52.56 54.855 53.44 ;
    RECT 51.255 52.56 51.535 53.44 ;
    RECT 47.935 52.56 48.215 53.44 ;
    RECT 44.615 52.56 44.895 53.44 ;
    RECT 41.295 52.56 41.575 53.44 ;
    RECT 37.975 52.56 38.255 53.44 ;
    RECT 34.655 52.56 34.935 53.44 ;
    RECT 130.935 52.56 131.215 53.44 ;
    RECT 127.615 52.56 127.895 53.44 ;
    RECT 124.295 52.56 124.575 53.44 ;
    RECT 120.975 52.56 121.255 53.44 ;
    RECT 117.655 52.56 117.935 53.44 ;
    RECT 114.335 52.56 114.615 53.44 ;
    RECT 111.015 52.56 111.295 53.44 ;
    RECT 107.695 52.56 107.975 53.44 ;
    RECT 104.375 52.56 104.655 53.44 ;
    RECT 101.055 52.56 101.335 53.44 ;
    RECT 170.775 52.56 171.055 53.44 ;
    RECT 167.455 52.56 167.735 53.44 ;
    RECT 97.735 52.56 98.015 53.44 ;
    RECT 94.415 52.56 94.695 53.44 ;
    RECT 91.095 52.56 91.375 53.44 ;
    RECT 87.775 52.56 88.055 53.44 ;
    RECT 84.455 52.56 84.735 53.44 ;
    RECT 81.135 52.56 81.415 53.44 ;
    RECT 77.815 52.56 78.095 53.44 ;
    RECT 74.495 52.56 74.775 53.44 ;
    RECT 71.175 52.56 71.455 53.44 ;
    RECT 31.335 52.56 31.615 53.44 ;
    RECT 67.855 52.56 68.135 53.44 ;
    RECT 28.015 52.56 28.295 53.44 ;
    RECT 24.695 52.56 24.975 53.44 ;
    RECT 21.375 52.56 21.655 53.44 ;
    RECT 18.055 52.56 18.335 53.44 ;
    RECT 14.735 52.56 15.015 53.44 ;
    RECT 11.415 52.56 11.695 53.44 ;
    RECT 8.095 52.56 8.375 53.44 ;
    RECT 4.775 52.56 5.055 53.44 ;
    RECT 164.135 52.56 164.415 53.44 ;
    RECT 1.455 52.56 1.735 53.44 ;
    RECT 160.815 52.56 161.095 53.44 ;
    RECT 157.495 52.56 157.775 53.44 ;
    RECT 154.175 52.56 154.455 53.44 ;
    RECT 150.855 52.56 151.135 53.44 ;
    RECT 147.535 52.56 147.815 53.44 ;
    RECT 144.215 52.56 144.495 53.44 ;
    RECT 140.895 52.56 141.175 53.44 ;
    RECT 137.575 52.56 137.855 53.44 ;
    RECT 134.255 52.56 134.535 53.44 ;
    RECT 64.535 52.56 64.815 53.44 ;
    RECT 61.215 51.84 61.495 52.72 ;
    RECT 57.895 51.84 58.175 52.72 ;
    RECT 54.575 51.84 54.855 52.72 ;
    RECT 51.255 51.84 51.535 52.72 ;
    RECT 47.935 51.84 48.215 52.72 ;
    RECT 44.615 51.84 44.895 52.72 ;
    RECT 41.295 51.84 41.575 52.72 ;
    RECT 37.975 51.84 38.255 52.72 ;
    RECT 34.655 51.84 34.935 52.72 ;
    RECT 130.935 51.84 131.215 52.72 ;
    RECT 127.615 51.84 127.895 52.72 ;
    RECT 124.295 51.84 124.575 52.72 ;
    RECT 120.975 51.84 121.255 52.72 ;
    RECT 117.655 51.84 117.935 52.72 ;
    RECT 114.335 51.84 114.615 52.72 ;
    RECT 111.015 51.84 111.295 52.72 ;
    RECT 107.695 51.84 107.975 52.72 ;
    RECT 104.375 51.84 104.655 52.72 ;
    RECT 101.055 51.84 101.335 52.72 ;
    RECT 170.775 51.84 171.055 52.72 ;
    RECT 167.455 51.84 167.735 52.72 ;
    RECT 97.735 51.84 98.015 52.72 ;
    RECT 94.415 51.84 94.695 52.72 ;
    RECT 91.095 51.84 91.375 52.72 ;
    RECT 87.775 51.84 88.055 52.72 ;
    RECT 84.455 51.84 84.735 52.72 ;
    RECT 81.135 51.84 81.415 52.72 ;
    RECT 77.815 51.84 78.095 52.72 ;
    RECT 74.495 51.84 74.775 52.72 ;
    RECT 71.175 51.84 71.455 52.72 ;
    RECT 31.335 51.84 31.615 52.72 ;
    RECT 67.855 51.84 68.135 52.72 ;
    RECT 28.015 51.84 28.295 52.72 ;
    RECT 24.695 51.84 24.975 52.72 ;
    RECT 21.375 51.84 21.655 52.72 ;
    RECT 18.055 51.84 18.335 52.72 ;
    RECT 14.735 51.84 15.015 52.72 ;
    RECT 11.415 51.84 11.695 52.72 ;
    RECT 8.095 51.84 8.375 52.72 ;
    RECT 4.775 51.84 5.055 52.72 ;
    RECT 164.135 51.84 164.415 52.72 ;
    RECT 1.455 51.84 1.735 52.72 ;
    RECT 160.815 51.84 161.095 52.72 ;
    RECT 157.495 51.84 157.775 52.72 ;
    RECT 154.175 51.84 154.455 52.72 ;
    RECT 150.855 51.84 151.135 52.72 ;
    RECT 147.535 51.84 147.815 52.72 ;
    RECT 144.215 51.84 144.495 52.72 ;
    RECT 140.895 51.84 141.175 52.72 ;
    RECT 137.575 51.84 137.855 52.72 ;
    RECT 134.255 51.84 134.535 52.72 ;
    RECT 64.535 51.84 64.815 52.72 ;
    RECT 61.215 51.12 61.495 52.0 ;
    RECT 57.895 51.12 58.175 52.0 ;
    RECT 54.575 51.12 54.855 52.0 ;
    RECT 51.255 51.12 51.535 52.0 ;
    RECT 47.935 51.12 48.215 52.0 ;
    RECT 44.615 51.12 44.895 52.0 ;
    RECT 41.295 51.12 41.575 52.0 ;
    RECT 37.975 51.12 38.255 52.0 ;
    RECT 34.655 51.12 34.935 52.0 ;
    RECT 130.935 51.12 131.215 52.0 ;
    RECT 127.615 51.12 127.895 52.0 ;
    RECT 124.295 51.12 124.575 52.0 ;
    RECT 120.975 51.12 121.255 52.0 ;
    RECT 117.655 51.12 117.935 52.0 ;
    RECT 114.335 51.12 114.615 52.0 ;
    RECT 111.015 51.12 111.295 52.0 ;
    RECT 107.695 51.12 107.975 52.0 ;
    RECT 104.375 51.12 104.655 52.0 ;
    RECT 101.055 51.12 101.335 52.0 ;
    RECT 170.775 51.12 171.055 52.0 ;
    RECT 167.455 51.12 167.735 52.0 ;
    RECT 97.735 51.12 98.015 52.0 ;
    RECT 94.415 51.12 94.695 52.0 ;
    RECT 91.095 51.12 91.375 52.0 ;
    RECT 87.775 51.12 88.055 52.0 ;
    RECT 84.455 51.12 84.735 52.0 ;
    RECT 81.135 51.12 81.415 52.0 ;
    RECT 77.815 51.12 78.095 52.0 ;
    RECT 74.495 51.12 74.775 52.0 ;
    RECT 71.175 51.12 71.455 52.0 ;
    RECT 31.335 51.12 31.615 52.0 ;
    RECT 67.855 51.12 68.135 52.0 ;
    RECT 28.015 51.12 28.295 52.0 ;
    RECT 24.695 51.12 24.975 52.0 ;
    RECT 21.375 51.12 21.655 52.0 ;
    RECT 18.055 51.12 18.335 52.0 ;
    RECT 14.735 51.12 15.015 52.0 ;
    RECT 11.415 51.12 11.695 52.0 ;
    RECT 8.095 51.12 8.375 52.0 ;
    RECT 4.775 51.12 5.055 52.0 ;
    RECT 164.135 51.12 164.415 52.0 ;
    RECT 1.455 51.12 1.735 52.0 ;
    RECT 160.815 51.12 161.095 52.0 ;
    RECT 157.495 51.12 157.775 52.0 ;
    RECT 154.175 51.12 154.455 52.0 ;
    RECT 150.855 51.12 151.135 52.0 ;
    RECT 147.535 51.12 147.815 52.0 ;
    RECT 144.215 51.12 144.495 52.0 ;
    RECT 140.895 51.12 141.175 52.0 ;
    RECT 137.575 51.12 137.855 52.0 ;
    RECT 134.255 51.12 134.535 52.0 ;
    RECT 64.535 51.12 64.815 52.0 ;
    RECT 61.215 50.4 61.495 51.28 ;
    RECT 57.895 50.4 58.175 51.28 ;
    RECT 54.575 50.4 54.855 51.28 ;
    RECT 51.255 50.4 51.535 51.28 ;
    RECT 47.935 50.4 48.215 51.28 ;
    RECT 44.615 50.4 44.895 51.28 ;
    RECT 41.295 50.4 41.575 51.28 ;
    RECT 37.975 50.4 38.255 51.28 ;
    RECT 34.655 50.4 34.935 51.28 ;
    RECT 130.935 50.4 131.215 51.28 ;
    RECT 127.615 50.4 127.895 51.28 ;
    RECT 124.295 50.4 124.575 51.28 ;
    RECT 120.975 50.4 121.255 51.28 ;
    RECT 117.655 50.4 117.935 51.28 ;
    RECT 114.335 50.4 114.615 51.28 ;
    RECT 111.015 50.4 111.295 51.28 ;
    RECT 107.695 50.4 107.975 51.28 ;
    RECT 104.375 50.4 104.655 51.28 ;
    RECT 101.055 50.4 101.335 51.28 ;
    RECT 170.775 50.4 171.055 51.28 ;
    RECT 167.455 50.4 167.735 51.28 ;
    RECT 97.735 50.4 98.015 51.28 ;
    RECT 94.415 50.4 94.695 51.28 ;
    RECT 91.095 50.4 91.375 51.28 ;
    RECT 87.775 50.4 88.055 51.28 ;
    RECT 84.455 50.4 84.735 51.28 ;
    RECT 81.135 50.4 81.415 51.28 ;
    RECT 77.815 50.4 78.095 51.28 ;
    RECT 74.495 50.4 74.775 51.28 ;
    RECT 71.175 50.4 71.455 51.28 ;
    RECT 31.335 50.4 31.615 51.28 ;
    RECT 67.855 50.4 68.135 51.28 ;
    RECT 28.015 50.4 28.295 51.28 ;
    RECT 24.695 50.4 24.975 51.28 ;
    RECT 21.375 50.4 21.655 51.28 ;
    RECT 18.055 50.4 18.335 51.28 ;
    RECT 14.735 50.4 15.015 51.28 ;
    RECT 11.415 50.4 11.695 51.28 ;
    RECT 8.095 50.4 8.375 51.28 ;
    RECT 4.775 50.4 5.055 51.28 ;
    RECT 164.135 50.4 164.415 51.28 ;
    RECT 1.455 50.4 1.735 51.28 ;
    RECT 160.815 50.4 161.095 51.28 ;
    RECT 157.495 50.4 157.775 51.28 ;
    RECT 154.175 50.4 154.455 51.28 ;
    RECT 150.855 50.4 151.135 51.28 ;
    RECT 147.535 50.4 147.815 51.28 ;
    RECT 144.215 50.4 144.495 51.28 ;
    RECT 140.895 50.4 141.175 51.28 ;
    RECT 137.575 50.4 137.855 51.28 ;
    RECT 134.255 50.4 134.535 51.28 ;
    RECT 64.535 50.4 64.815 51.28 ;
    RECT 187.83 56.96 187.91 57.68 ;
    RECT 192.82 56.96 193.09 57.68 ;
    RECT 187.83 56.24 187.91 56.96 ;
    RECT 192.82 56.24 193.09 56.96 ;
    RECT 187.83 55.52 187.91 56.24 ;
    RECT 192.82 55.52 193.09 56.24 ;
    RECT 187.83 54.8 187.91 55.52 ;
    RECT 192.82 54.8 193.09 55.52 ;
    RECT 187.83 54.08 187.91 54.8 ;
    RECT 192.82 54.08 193.09 54.8 ;
    RECT 187.83 53.36 187.91 54.08 ;
    RECT 192.82 53.36 193.09 54.08 ;
    RECT 187.83 52.64 187.91 53.36 ;
    RECT 192.82 52.64 193.09 53.36 ;
    RECT 187.83 51.92 187.91 52.64 ;
    RECT 192.82 51.92 193.09 52.64 ;
    RECT 187.83 51.2 187.91 51.92 ;
    RECT 192.82 51.2 193.09 51.92 ;
    RECT 187.83 50.48 187.91 51.2 ;
    RECT 192.82 50.48 193.09 51.2 ;
    RECT 187.83 49.76 187.91 50.48 ;
    RECT 192.82 49.76 193.09 50.48 ;
    RECT 187.83 49.04 187.91 49.76 ;
    RECT 192.82 49.04 193.09 49.76 ;
    RECT 187.83 58.42 187.91 59.14 ;
    RECT 192.82 58.42 193.09 59.14 ;
    RECT 187.83 48.32 187.91 49.04 ;
    RECT 192.82 48.32 193.09 49.04 ;
    RECT 187.83 47.6 187.91 48.32 ;
    RECT 192.82 47.6 193.09 48.32 ;
    RECT 187.83 46.88 187.91 47.6 ;
    RECT 192.82 46.88 193.09 47.6 ;
    RECT 187.83 46.16 187.91 46.88 ;
    RECT 192.82 46.16 193.09 46.88 ;
    RECT 187.83 45.44 187.91 46.16 ;
    RECT 192.82 45.44 193.09 46.16 ;
    RECT 187.83 44.72 187.91 45.44 ;
    RECT 192.82 44.72 193.09 45.44 ;
    RECT 187.83 44.0 187.91 44.72 ;
    RECT 192.82 44.0 193.09 44.72 ;
    RECT 187.83 43.28 187.91 44.0 ;
    RECT 192.82 43.28 193.09 44.0 ;
    RECT 187.83 42.56 187.91 43.28 ;
    RECT 192.82 42.56 193.09 43.28 ;
    RECT 187.83 41.84 187.91 42.56 ;
    RECT 192.82 41.84 193.09 42.56 ;
    RECT 187.83 57.68 187.91 58.42 ;
    RECT 192.82 57.68 193.09 58.42 ;
    RECT 187.83 41.12 187.91 41.84 ;
    RECT 192.82 41.12 193.09 41.84 ;
    RECT 187.83 40.4 187.91 41.12 ;
    RECT 192.82 40.4 193.09 41.12 ;
    RECT 187.83 39.68 187.91 40.4 ;
    RECT 192.82 39.68 193.09 40.4 ;
    RECT 187.83 38.96 187.91 39.68 ;
    RECT 192.82 38.96 193.09 39.68 ;
    RECT 187.83 38.24 187.91 38.96 ;
    RECT 192.82 38.24 193.09 38.96 ;
    RECT 187.83 37.52 187.91 38.24 ;
    RECT 192.82 37.52 193.09 38.24 ;
    RECT 187.83 36.8 187.91 37.52 ;
    RECT 192.82 36.8 193.09 37.52 ;
    RECT 187.83 36.08 187.91 36.8 ;
    RECT 192.82 36.08 193.09 36.8 ;
    RECT 187.83 35.36 187.91 36.08 ;
    RECT 192.82 35.36 193.09 36.08 ;
    RECT 187.83 34.64 187.91 35.36 ;
    RECT 192.82 34.64 193.09 35.36 ;
    RECT 181.455 11.6 181.665 29.24 ;
    RECT 187.83 11.645 187.91 34.785 ;
    RECT 192.82 11.435 193.09 34.64 ;
    RECT 174.79 60.175 174.98 60.67 ;
    RECT 187.83 59.14 187.91 60.6 ;
    RECT 192.82 59.14 193.09 60.67 ;
    RECT 366.245 9.705 366.525 10.07 ;
    RECT 362.925 9.705 363.205 10.07 ;
    RECT 359.605 9.705 359.885 10.07 ;
    RECT 356.285 9.705 356.565 10.07 ;
    RECT 352.965 9.705 353.245 10.07 ;
    RECT 349.645 9.705 349.925 10.07 ;
    RECT 346.325 9.705 346.605 10.07 ;
    RECT 343.005 9.705 343.285 10.07 ;
    RECT 339.685 9.705 339.965 10.07 ;
    RECT 336.365 9.705 336.645 10.07 ;
    RECT 333.045 9.705 333.325 10.07 ;
    RECT 329.725 9.705 330.005 10.07 ;
    RECT 326.405 9.705 326.685 10.07 ;
    RECT 323.085 9.705 323.365 10.07 ;
    RECT 319.765 9.705 320.045 10.07 ;
    RECT 316.445 9.705 316.725 10.07 ;
    RECT 313.125 9.705 313.405 10.07 ;
    RECT 309.805 9.705 310.085 10.07 ;
    RECT 306.485 9.705 306.765 10.07 ;
    RECT 303.165 9.705 303.445 10.07 ;
    RECT 233.445 9.705 233.725 10.07 ;
    RECT 230.125 9.705 230.405 10.07 ;
    RECT 226.805 9.705 227.085 10.07 ;
    RECT 223.485 9.705 223.765 10.07 ;
    RECT 220.165 9.705 220.445 10.07 ;
    RECT 299.845 9.705 300.125 10.07 ;
    RECT 216.845 9.705 217.125 10.07 ;
    RECT 296.525 9.705 296.805 10.07 ;
    RECT 213.525 9.705 213.805 10.07 ;
    RECT 293.205 9.705 293.485 10.07 ;
    RECT 210.205 9.705 210.485 10.07 ;
    RECT 289.885 9.705 290.165 10.07 ;
    RECT 206.885 9.705 207.165 10.07 ;
    RECT 286.565 9.705 286.845 10.07 ;
    RECT 283.245 9.705 283.525 10.07 ;
    RECT 279.925 9.705 280.205 10.07 ;
    RECT 276.605 9.705 276.885 10.07 ;
    RECT 273.285 9.705 273.565 10.07 ;
    RECT 269.965 9.705 270.245 10.07 ;
    RECT 266.645 9.705 266.925 10.07 ;
    RECT 263.325 9.705 263.605 10.07 ;
    RECT 260.005 9.705 260.285 10.07 ;
    RECT 256.685 9.705 256.965 10.07 ;
    RECT 253.365 9.705 253.645 10.07 ;
    RECT 250.045 9.705 250.325 10.07 ;
    RECT 246.725 9.705 247.005 10.07 ;
    RECT 243.405 9.705 243.685 10.07 ;
    RECT 240.085 9.705 240.365 10.07 ;
    RECT 236.765 9.705 237.045 10.07 ;
    RECT 372.885 9.705 373.165 10.07 ;
    RECT 203.565 9.705 203.845 10.07 ;
    RECT 369.565 9.705 369.845 10.07 ;
    RECT 372.885 10.07 373.165 11.6 ;
    RECT 369.565 10.07 369.845 11.6 ;
    RECT 366.245 10.07 366.525 11.6 ;
    RECT 362.925 10.07 363.205 11.6 ;
    RECT 359.605 10.07 359.885 11.6 ;
    RECT 356.285 10.07 356.565 11.6 ;
    RECT 352.965 10.07 353.245 11.6 ;
    RECT 349.645 10.07 349.925 11.6 ;
    RECT 346.325 10.07 346.605 11.6 ;
    RECT 343.005 10.07 343.285 11.6 ;
    RECT 339.685 10.07 339.965 11.6 ;
    RECT 336.365 10.07 336.645 11.6 ;
    RECT 333.045 10.07 333.325 11.6 ;
    RECT 329.725 10.07 330.005 11.6 ;
    RECT 326.405 10.07 326.685 11.6 ;
    RECT 323.085 10.07 323.365 11.6 ;
    RECT 319.765 10.07 320.045 11.6 ;
    RECT 316.445 10.07 316.725 11.6 ;
    RECT 313.125 10.07 313.405 11.6 ;
    RECT 309.805 10.07 310.085 11.6 ;
    RECT 306.485 10.07 306.765 11.6 ;
    RECT 303.165 10.07 303.445 11.6 ;
    RECT 299.845 10.07 300.125 11.6 ;
    RECT 296.525 10.07 296.805 11.6 ;
    RECT 293.205 10.07 293.485 11.6 ;
    RECT 289.885 10.07 290.165 11.6 ;
    RECT 286.565 10.07 286.845 11.6 ;
    RECT 283.245 10.07 283.525 11.6 ;
    RECT 279.925 10.07 280.205 11.6 ;
    RECT 276.605 10.07 276.885 11.6 ;
    RECT 273.285 10.07 273.565 11.6 ;
    RECT 269.965 10.07 270.245 11.6 ;
    RECT 266.645 10.07 266.925 11.6 ;
    RECT 263.325 10.07 263.605 11.6 ;
    RECT 260.005 10.07 260.285 11.6 ;
    RECT 256.685 10.07 256.965 11.6 ;
    RECT 253.365 10.07 253.645 11.6 ;
    RECT 250.045 10.07 250.325 11.6 ;
    RECT 246.725 10.07 247.005 11.6 ;
    RECT 243.405 10.07 243.685 11.6 ;
    RECT 240.085 10.07 240.365 11.6 ;
    RECT 236.765 10.07 237.045 11.6 ;
    RECT 233.445 10.07 233.725 11.6 ;
    RECT 230.125 10.07 230.405 11.6 ;
    RECT 226.805 10.07 227.085 11.6 ;
    RECT 223.485 10.07 223.765 11.6 ;
    RECT 220.165 10.07 220.445 11.6 ;
    RECT 216.845 10.07 217.125 11.6 ;
    RECT 213.525 10.07 213.805 11.6 ;
    RECT 210.205 10.07 210.485 11.6 ;
    RECT 206.885 10.07 207.165 11.6 ;
    RECT 203.565 10.07 203.845 11.6 ;
    RECT 181.455 0.815 181.665 11.6 ;
    RECT 192.82 1.72 193.09 11.635 ;
    RECT 197.215 3.255 197.3 5.305 ;
    RECT 170.775 10.07 171.055 11.6 ;
    RECT 167.455 10.07 167.735 11.6 ;
    RECT 164.135 10.07 164.415 11.6 ;
    RECT 160.815 10.07 161.095 11.6 ;
    RECT 157.495 10.07 157.775 11.6 ;
    RECT 154.175 10.07 154.455 11.6 ;
    RECT 150.855 10.07 151.135 11.6 ;
    RECT 147.535 10.07 147.815 11.6 ;
    RECT 144.215 10.07 144.495 11.6 ;
    RECT 140.895 10.07 141.175 11.6 ;
    RECT 137.575 10.07 137.855 11.6 ;
    RECT 134.255 10.07 134.535 11.6 ;
    RECT 130.935 10.07 131.215 11.6 ;
    RECT 127.615 10.07 127.895 11.6 ;
    RECT 124.295 10.07 124.575 11.6 ;
    RECT 120.975 10.07 121.255 11.6 ;
    RECT 117.655 10.07 117.935 11.6 ;
    RECT 114.335 10.07 114.615 11.6 ;
    RECT 111.015 10.07 111.295 11.6 ;
    RECT 107.695 10.07 107.975 11.6 ;
    RECT 104.375 10.07 104.655 11.6 ;
    RECT 101.055 10.07 101.335 11.6 ;
    RECT 97.735 10.07 98.015 11.6 ;
    RECT 94.415 10.07 94.695 11.6 ;
    RECT 91.095 10.07 91.375 11.6 ;
    RECT 87.775 10.07 88.055 11.6 ;
    RECT 84.455 10.07 84.735 11.6 ;
    RECT 81.135 10.07 81.415 11.6 ;
    RECT 77.815 10.07 78.095 11.6 ;
    RECT 74.495 10.07 74.775 11.6 ;
    RECT 71.175 10.07 71.455 11.6 ;
    RECT 67.855 10.07 68.135 11.6 ;
    RECT 64.535 10.07 64.815 11.6 ;
    RECT 61.215 10.07 61.495 11.6 ;
    RECT 57.895 10.07 58.175 11.6 ;
    RECT 54.575 10.07 54.855 11.6 ;
    RECT 51.255 10.07 51.535 11.6 ;
    RECT 47.935 10.07 48.215 11.6 ;
    RECT 44.615 10.07 44.895 11.6 ;
    RECT 41.295 10.07 41.575 11.6 ;
    RECT 37.975 10.07 38.255 11.6 ;
    RECT 34.655 10.07 34.935 11.6 ;
    RECT 31.335 10.07 31.615 11.6 ;
    RECT 28.015 10.07 28.295 11.6 ;
    RECT 24.695 10.07 24.975 11.6 ;
    RECT 21.375 10.07 21.655 11.6 ;
    RECT 18.055 10.07 18.335 11.6 ;
    RECT 14.735 10.07 15.015 11.6 ;
    RECT 11.415 10.07 11.695 11.6 ;
    RECT 8.095 10.07 8.375 11.6 ;
    RECT 4.775 10.07 5.055 11.6 ;
    RECT 1.455 10.07 1.735 11.6 ;
    RECT 64.535 9.705 64.815 10.07 ;
    RECT 61.215 9.705 61.495 10.07 ;
    RECT 57.895 9.705 58.175 10.07 ;
    RECT 54.575 9.705 54.855 10.07 ;
    RECT 51.255 9.705 51.535 10.07 ;
    RECT 47.935 9.705 48.215 10.07 ;
    RECT 44.615 9.705 44.895 10.07 ;
    RECT 41.295 9.705 41.575 10.07 ;
    RECT 37.975 9.705 38.255 10.07 ;
    RECT 34.655 9.705 34.935 10.07 ;
    RECT 31.335 9.705 31.615 10.07 ;
    RECT 28.015 9.705 28.295 10.07 ;
    RECT 24.695 9.705 24.975 10.07 ;
    RECT 21.375 9.705 21.655 10.07 ;
    RECT 18.055 9.705 18.335 10.07 ;
    RECT 14.735 9.705 15.015 10.07 ;
    RECT 11.415 9.705 11.695 10.07 ;
    RECT 8.095 9.705 8.375 10.07 ;
    RECT 4.775 9.705 5.055 10.07 ;
    RECT 170.775 9.705 171.055 10.07 ;
    RECT 1.455 9.705 1.735 10.07 ;
    RECT 167.455 9.705 167.735 10.07 ;
    RECT 164.135 9.705 164.415 10.07 ;
    RECT 160.815 9.705 161.095 10.07 ;
    RECT 157.495 9.705 157.775 10.07 ;
    RECT 154.175 9.705 154.455 10.07 ;
    RECT 150.855 9.705 151.135 10.07 ;
    RECT 147.535 9.705 147.815 10.07 ;
    RECT 144.215 9.705 144.495 10.07 ;
    RECT 140.895 9.705 141.175 10.07 ;
    RECT 137.575 9.705 137.855 10.07 ;
    RECT 134.255 9.705 134.535 10.07 ;
    RECT 130.935 9.705 131.215 10.07 ;
    RECT 127.615 9.705 127.895 10.07 ;
    RECT 124.295 9.705 124.575 10.07 ;
    RECT 120.975 9.705 121.255 10.07 ;
    RECT 117.655 9.705 117.935 10.07 ;
    RECT 114.335 9.705 114.615 10.07 ;
    RECT 111.015 9.705 111.295 10.07 ;
    RECT 107.695 9.705 107.975 10.07 ;
    RECT 104.375 9.705 104.655 10.07 ;
    RECT 101.055 9.705 101.335 10.07 ;
    RECT 97.735 9.705 98.015 10.07 ;
    RECT 94.415 9.705 94.695 10.07 ;
    RECT 91.095 9.705 91.375 10.07 ;
    RECT 87.775 9.705 88.055 10.07 ;
    RECT 84.455 9.705 84.735 10.07 ;
    RECT 81.135 9.705 81.415 10.07 ;
    RECT 77.815 9.705 78.095 10.07 ;
    RECT 74.495 9.705 74.775 10.07 ;
    RECT 71.175 9.705 71.455 10.07 ;
    RECT 67.855 9.705 68.135 10.07 ;
    RECT 266.645 60.67 266.925 61.185 ;
    RECT 263.325 60.67 263.605 61.185 ;
    RECT 260.005 60.67 260.285 61.185 ;
    RECT 256.685 60.67 256.965 61.185 ;
    RECT 253.365 60.67 253.645 61.185 ;
    RECT 250.045 60.67 250.325 61.185 ;
    RECT 246.725 60.67 247.005 61.185 ;
    RECT 243.405 60.67 243.685 61.185 ;
    RECT 240.085 60.67 240.365 61.185 ;
    RECT 236.765 60.67 237.045 61.185 ;
    RECT 170.775 60.67 171.055 61.185 ;
    RECT 167.455 60.67 167.735 61.185 ;
    RECT 164.135 60.67 164.415 61.185 ;
    RECT 160.815 60.67 161.095 61.185 ;
    RECT 157.495 60.67 157.775 61.185 ;
    RECT 154.175 60.67 154.455 61.185 ;
    RECT 150.855 60.67 151.135 61.185 ;
    RECT 147.535 60.67 147.815 61.185 ;
    RECT 144.215 60.67 144.495 61.185 ;
    RECT 140.895 60.67 141.175 61.185 ;
    RECT 137.575 60.67 137.855 61.185 ;
    RECT 134.255 60.67 134.535 61.185 ;
    RECT 130.935 60.67 131.215 61.185 ;
    RECT 127.615 60.67 127.895 61.185 ;
    RECT 124.295 60.67 124.575 61.185 ;
    RECT 120.975 60.67 121.255 61.185 ;
    RECT 117.655 60.67 117.935 61.185 ;
    RECT 114.335 60.67 114.615 61.185 ;
    RECT 111.015 60.67 111.295 61.185 ;
    RECT 107.695 60.67 107.975 61.185 ;
    RECT 233.445 60.67 233.725 61.185 ;
    RECT 104.375 60.67 104.655 61.185 ;
    RECT 230.125 60.67 230.405 61.185 ;
    RECT 101.055 60.67 101.335 61.185 ;
    RECT 226.805 60.67 227.085 61.185 ;
    RECT 223.485 60.67 223.765 61.185 ;
    RECT 220.165 60.67 220.445 61.185 ;
    RECT 216.845 60.67 217.125 61.185 ;
    RECT 213.525 60.67 213.805 61.185 ;
    RECT 210.205 60.67 210.485 61.185 ;
    RECT 206.885 60.67 207.165 61.185 ;
    RECT 203.565 60.67 203.845 61.185 ;
    RECT 97.735 60.67 98.015 61.185 ;
    RECT 94.415 60.67 94.695 61.185 ;
    RECT 91.095 60.67 91.375 61.185 ;
    RECT 87.775 60.67 88.055 61.185 ;
    RECT 84.455 60.67 84.735 61.185 ;
    RECT 81.135 60.67 81.415 61.185 ;
    RECT 77.815 60.67 78.095 61.185 ;
    RECT 74.495 60.67 74.775 61.185 ;
    RECT 71.175 60.67 71.455 61.185 ;
    RECT 67.855 60.67 68.135 61.185 ;
    RECT 64.535 60.67 64.815 61.185 ;
    RECT 61.215 60.67 61.495 61.185 ;
    RECT 57.895 60.67 58.175 61.185 ;
    RECT 54.575 60.67 54.855 61.185 ;
    RECT 51.255 60.67 51.535 61.185 ;
    RECT 47.935 60.67 48.215 61.185 ;
    RECT 44.615 60.67 44.895 61.185 ;
    RECT 41.295 60.67 41.575 61.185 ;
    RECT 37.975 60.67 38.255 61.185 ;
    RECT 34.655 60.67 34.935 61.185 ;
    RECT 372.885 60.67 373.165 61.185 ;
    RECT 369.565 60.67 369.845 61.185 ;
    RECT 366.245 60.67 366.525 61.185 ;
    RECT 362.925 60.67 363.205 61.185 ;
    RECT 359.605 60.67 359.885 61.185 ;
    RECT 31.335 60.67 31.615 61.185 ;
    RECT 356.285 60.67 356.565 61.185 ;
    RECT 28.015 60.67 28.295 61.185 ;
    RECT 352.965 60.67 353.245 61.185 ;
    RECT 24.695 60.67 24.975 61.185 ;
    RECT 349.645 60.67 349.925 61.185 ;
    RECT 21.375 60.67 21.655 61.185 ;
    RECT 346.325 60.67 346.605 61.185 ;
    RECT 18.055 60.67 18.335 61.185 ;
    RECT 343.005 60.67 343.285 61.185 ;
    RECT 14.735 60.67 15.015 61.185 ;
    RECT 339.685 60.67 339.965 61.185 ;
    RECT 11.415 60.67 11.695 61.185 ;
    RECT 336.365 60.67 336.645 61.185 ;
    RECT 8.095 60.67 8.375 61.185 ;
    RECT 4.775 60.67 5.055 61.185 ;
    RECT 1.455 60.67 1.735 61.185 ;
    RECT 174.79 60.67 174.98 60.99 ;
    RECT 192.82 60.67 193.09 61.185 ;
    RECT 333.045 60.67 333.325 61.185 ;
    RECT 329.725 60.67 330.005 61.185 ;
    RECT 326.405 60.67 326.685 61.185 ;
    RECT 323.085 60.67 323.365 61.185 ;
    RECT 319.765 60.67 320.045 61.185 ;
    RECT 316.445 60.67 316.725 61.185 ;
    RECT 313.125 60.67 313.405 61.185 ;
    RECT 309.805 60.67 310.085 61.185 ;
    RECT 306.485 60.67 306.765 61.185 ;
    RECT 303.165 60.67 303.445 61.185 ;
    RECT 299.845 60.67 300.125 61.185 ;
    RECT 296.525 60.67 296.805 61.185 ;
    RECT 293.205 60.67 293.485 61.185 ;
    RECT 289.885 60.67 290.165 61.185 ;
    RECT 286.565 60.67 286.845 61.185 ;
    RECT 283.245 60.67 283.525 61.185 ;
    RECT 279.925 60.67 280.205 61.185 ;
    RECT 276.605 60.67 276.885 61.185 ;
    RECT 273.285 60.67 273.565 61.185 ;
    RECT 269.965 60.67 270.245 61.185 ;
    END
  END sram520x104

END LIBRARY

